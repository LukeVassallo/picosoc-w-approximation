* NGSPICE file created from pcpi_div.ext - technology: gf180mcuD

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_1 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_1 D CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_64 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_64 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__antenna abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__antenna I VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_2 I0 I1 S Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_1 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_1 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_1 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_2 D CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_1 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_2 A1 A2 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_2 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_8 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_1 A1 A2 A3 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_4 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_1 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_2 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or3_1 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_2 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_1 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_2 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_1 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_1 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_2 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_2 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_1 A1 A2 A3 A4 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_2 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_2 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_1 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_2 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_2 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_1 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_2 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_2 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_2 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_1 A1 A2 A3 B1 B2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_1 A1 A2 A3 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_1 A1 A2 B1 B2 C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_4 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_2 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_2 A1 A2 A3 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_4 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_1 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

.subckt pcpi_div clk pcpi_div_rd[0] pcpi_div_rd[10] pcpi_div_rd[11] pcpi_div_rd[12]
+ pcpi_div_rd[13] pcpi_div_rd[14] pcpi_div_rd[15] pcpi_div_rd[16] pcpi_div_rd[17]
+ pcpi_div_rd[18] pcpi_div_rd[19] pcpi_div_rd[1] pcpi_div_rd[20] pcpi_div_rd[21] pcpi_div_rd[22]
+ pcpi_div_rd[23] pcpi_div_rd[24] pcpi_div_rd[25] pcpi_div_rd[26] pcpi_div_rd[27]
+ pcpi_div_rd[28] pcpi_div_rd[29] pcpi_div_rd[2] pcpi_div_rd[30] pcpi_div_rd[31] pcpi_div_rd[3]
+ pcpi_div_rd[4] pcpi_div_rd[5] pcpi_div_rd[6] pcpi_div_rd[7] pcpi_div_rd[8] pcpi_div_rd[9]
+ pcpi_div_ready pcpi_div_valid pcpi_div_wait pcpi_div_wr pcpi_insn[0] pcpi_insn[10]
+ pcpi_insn[11] pcpi_insn[12] pcpi_insn[13] pcpi_insn[14] pcpi_insn[15] pcpi_insn[16]
+ pcpi_insn[17] pcpi_insn[18] pcpi_insn[19] pcpi_insn[1] pcpi_insn[20] pcpi_insn[21]
+ pcpi_insn[22] pcpi_insn[23] pcpi_insn[24] pcpi_insn[25] pcpi_insn[26] pcpi_insn[27]
+ pcpi_insn[28] pcpi_insn[29] pcpi_insn[2] pcpi_insn[30] pcpi_insn[31] pcpi_insn[3]
+ pcpi_insn[4] pcpi_insn[5] pcpi_insn[6] pcpi_insn[7] pcpi_insn[8] pcpi_insn[9] pcpi_rs1[0]
+ pcpi_rs1[10] pcpi_rs1[11] pcpi_rs1[12] pcpi_rs1[13] pcpi_rs1[14] pcpi_rs1[15] pcpi_rs1[16]
+ pcpi_rs1[17] pcpi_rs1[18] pcpi_rs1[19] pcpi_rs1[1] pcpi_rs1[20] pcpi_rs1[21] pcpi_rs1[22]
+ pcpi_rs1[23] pcpi_rs1[24] pcpi_rs1[25] pcpi_rs1[26] pcpi_rs1[27] pcpi_rs1[28] pcpi_rs1[29]
+ pcpi_rs1[2] pcpi_rs1[30] pcpi_rs1[31] pcpi_rs1[3] pcpi_rs1[4] pcpi_rs1[5] pcpi_rs1[6]
+ pcpi_rs1[7] pcpi_rs1[8] pcpi_rs1[9] pcpi_rs2[0] pcpi_rs2[10] pcpi_rs2[11] pcpi_rs2[12]
+ pcpi_rs2[13] pcpi_rs2[14] pcpi_rs2[15] pcpi_rs2[16] pcpi_rs2[17] pcpi_rs2[18] pcpi_rs2[19]
+ pcpi_rs2[1] pcpi_rs2[20] pcpi_rs2[21] pcpi_rs2[22] pcpi_rs2[23] pcpi_rs2[24] pcpi_rs2[25]
+ pcpi_rs2[26] pcpi_rs2[27] pcpi_rs2[28] pcpi_rs2[29] pcpi_rs2[2] pcpi_rs2[30] pcpi_rs2[31]
+ pcpi_rs2[3] pcpi_rs2[4] pcpi_rs2[5] pcpi_rs2[6] pcpi_rs2[7] pcpi_rs2[8] pcpi_rs2[9]
+ resetn vdd vss
X_2106_ picorv32_pcpi_div_inst_0.quotient_msk\[15\] _0317_ picorv32_pcpi_div_inst_0.quotient\[15\]
+ _0319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2037_ picorv32_pcpi_div_inst_0.divisor\[29\] _0265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_64_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2939_ _0093_ clknet_4_12_0_clk picorv32_pcpi_div_inst_0.quotient\[24\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_9_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_17_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input73_I pcpi_rs2[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2706__A1 _0405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2349__B _0406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1445__A1 _0952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_43_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1996__A2 _1095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_58_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1606_ _1110_ _1111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3005__CLK clknet_4_10_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2655_ picorv32_pcpi_div_inst_0.divisor\[36\] _0753_ _0778_ _0779_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2724_ _0768_ _0839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_14_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1468_ _0954_ _0985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1537_ _0954_ _1048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2586_ picorv32_pcpi_div_inst_0.dividend\[31\] _0717_ _0401_ _0718_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_10_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_49_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_40_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1978__A2 picorv32_pcpi_div_inst_0.dividend\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_56_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_5_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3028__CLK clknet_4_1_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2440_ _0580_ _0583_ _0585_ _0586_ _0587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_2371_ _0206_ _0524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__1657__A1 _1153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_4_12_0_clk clknet_0_clk clknet_4_12_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_46_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1847__I _1320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_42_353 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2638_ net73 _0763_ _0764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2569_ _1233_ _0702_ _0678_ _0703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2707_ _0824_ picorv32_pcpi_div_inst_0.divisor\[41\] _0395_ _0825_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_input36_I pcpi_rs1[25] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1639__A1 _1116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1940_ _1346_ _1188_ _1391_ _1392_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_28_147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1871_ picorv32_pcpi_div_inst_0.divisor\[17\] _1336_ _1334_ picorv32_pcpi_div_inst_0.divisor\[18\]
+ _1337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_16_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_353 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2423_ net24 _0558_ _0434_ _0571_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_10_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_67_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_67_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2285_ _0417_ _0445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2354_ _0427_ _0508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_19_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_456 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2358__A2 _1041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_13_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2860__CLK clknet_4_12_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2070_ picorv32_pcpi_div_inst_0.quotient_msk\[2\] _0294_ picorv32_pcpi_div_inst_0.quotient\[2\]
+ _0296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_56_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2972_ _0126_ clknet_4_13_0_clk picorv32_pcpi_div_inst_0.quotient_msk\[25\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_48_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_28_Left_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_8_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1785_ net4 net3 _1255_ _1267_ _1270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_0_29_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1923_ _1372_ picorv32_pcpi_div_inst_0.dividend\[17\] picorv32_pcpi_div_inst_0.dividend\[16\]
+ _1374_ _1375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_0_21_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1854_ _1324_ _1321_ _1317_ picorv32_pcpi_div_inst_0.divisor\[12\] _1326_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_12_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2406_ _0433_ _0552_ _0555_ _0556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_12_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2199_ picorv32_pcpi_div_inst_0.quotient_msk\[19\] _0375_ _0372_ picorv32_pcpi_div_inst_0.quotient_msk\[20\]
+ _0376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2337_ _1309_ _1025_ _0483_ _0493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1860__I _1320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2268_ _0427_ _0429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_47_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_50_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_10_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1570_ _0988_ _1073_ _1077_ _0002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_21_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2122_ _0326_ _0328_ _0090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_49_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2053_ picorv32_pcpi_div_inst_0.divisor\[43\] picorv32_pcpi_div_inst_0.divisor\[42\]
+ picorv32_pcpi_div_inst_0.divisor\[41\] picorv32_pcpi_div_inst_0.divisor\[40\] _0281_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
X_2955_ _0109_ clknet_4_7_0_clk picorv32_pcpi_div_inst_0.quotient_msk\[8\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_29_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1768_ net5 _1255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1906_ _1352_ _1360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_40_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2886_ _0040_ clknet_4_3_0_clk picorv32_pcpi_div_inst_0.divisor\[2\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2430__A1 net22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1837_ picorv32_pcpi_div_inst_0.divisor\[8\] _1313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1699_ _0983_ _1193_ _1194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1590__I _0957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2497__A1 _0414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2249__A1 _0402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_23_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput86 net86 pcpi_div_rd[11] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput97 net97 pcpi_div_rd[21] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_46_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1622_ _1123_ _1124_ _1125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2671_ picorv32_pcpi_div_inst_0.divisor\[38\] _0783_ _0792_ _0793_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_26_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2412__A1 _0459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2740_ picorv32_pcpi_div_inst_0.divisor\[45\] _0853_ _0854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1484_ picorv32_pcpi_div_inst_0.quotient\[4\] _0999_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1553_ _1029_ _1062_ _1063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2479__A1 net26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2105_ _0314_ _0318_ _0083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_49_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_37_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2036_ _0250_ _0260_ _0263_ _0264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_27_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2938_ _0092_ clknet_4_14_0_clk picorv32_pcpi_div_inst_0.quotient\[23\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_43_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2869_ _0009_ clknet_4_11_0_clk net93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_32_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input66_I pcpi_rs2[23] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_15_Left_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_55_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_43_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2642__A1 _0747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1495__I _0955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1709__B _1202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_59_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_54_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2723_ _0795_ _0837_ _0838_ _0181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1605_ _1030_ _1108_ _1107_ _0985_ _1110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_1536_ _0968_ _1044_ _1047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2654_ _0775_ _0777_ _0778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2585_ _0586_ _0713_ _0716_ _0717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_1_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1467_ _0962_ _0951_ _0983_ _0984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_37_318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2019_ picorv32_pcpi_div_inst_0.divisor\[24\] picorv32_pcpi_div_inst_0.dividend\[24\]
+ _0247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_9_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_45_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_9_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_0_Left_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_56_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2967__CLK clknet_4_15_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2370_ net20 _0522_ _0523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_19_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_62_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2706_ _0405_ _0822_ _0823_ _0824_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1519_ picorv32_pcpi_div_inst_0.quotient\[4\] picorv32_pcpi_div_inst_0.quotient\[5\]
+ picorv32_pcpi_div_inst_0.quotient\[6\] _0998_ _1031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_49_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2637_ net62 _0748_ _0762_ _0763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2499_ _0455_ _0639_ _0640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2568_ _0698_ _0701_ _0404_ _0702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_2_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_12_Right_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2845__A1 _0469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input29_I pcpi_rs1[19] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_21_Right_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_65_468 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_52_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_36_Left_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_33_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_30_Right_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_45_Left_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_56_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_16_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_54_Left_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_43_118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2553__B _0490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1870_ _1320_ _1336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_24_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_63_Left_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1575__A1 _1078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2353_ _1041_ _0429_ _0507_ _0142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_12_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2422_ _0459_ _0569_ _0570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_67_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_67_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2284_ _0413_ _0444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_59_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1999_ _0224_ _0225_ _0226_ _0227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3018__CLK clknet_4_4_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_13_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1557__A1 picorv32_pcpi_div_inst_0.dividend\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_21_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_4_11_0_clk clknet_0_clk clknet_4_11_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XPHY_EDGE_ROW_3_Left_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2971_ _0125_ clknet_4_13_0_clk picorv32_pcpi_div_inst_0.quotient_msk\[24\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_56_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1922_ picorv32_pcpi_div_inst_0.divisor\[16\] _1374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__1796__A1 picorv32_pcpi_div_inst_0.running vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1784_ net3 _1255_ _1269_ _0035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_1853_ _1325_ _0048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_12_324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2336_ net48 _0491_ _0492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2405_ _0439_ _0554_ _0555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_67_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2198_ _0362_ _0375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2267_ _0428_ _0135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_62_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_10_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_26_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_21_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2121_ picorv32_pcpi_div_inst_0.quotient_msk\[21\] _0323_ picorv32_pcpi_div_inst_0.quotient\[21\]
+ _0328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_49_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_49_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2052_ _0276_ _0277_ _0278_ _0279_ _0280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_2954_ _0108_ clknet_4_7_0_clk picorv32_pcpi_div_inst_0.quotient_msk\[7\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_44_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1905_ _1359_ _0066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_29_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2885_ _0039_ clknet_4_3_0_clk picorv32_pcpi_div_inst_0.divisor\[1\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2430__A2 net23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1767_ net3 _1254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1698_ picorv32_pcpi_div_inst_0.dividend\[23\] picorv32_pcpi_div_inst_0.dividend\[22\]
+ _1178_ _1193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_32_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_6_Right_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1836_ _1312_ _0044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_4_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_12_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2319_ _1016_ _0476_ _0427_ _0477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_input11_I pcpi_insn[29] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2850__CLK clknet_4_4_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput98 net98 pcpi_div_rd[22] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput87 net87 pcpi_div_rd[12] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_31_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_59_Right_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_58_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_46_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1621_ _1113_ _1100_ _1102_ _1124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_1552_ _1060_ _1061_ _1062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2670_ _0775_ _0791_ _0792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_14_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2104_ picorv32_pcpi_div_inst_0.quotient_msk\[14\] _0317_ _1108_ _0318_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1483_ picorv32_pcpi_div_inst_0.quotient\[0\] picorv32_pcpi_div_inst_0.quotient\[1\]
+ picorv32_pcpi_div_inst_0.quotient\[2\] picorv32_pcpi_div_inst_0.quotient\[3\] _0998_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or4_2
XANTENNA__2873__CLK clknet_4_11_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input3_I pcpi_insn[12] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2479__A2 net27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_37_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2035_ _0261_ _0262_ _0263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_27_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2937_ _0091_ clknet_4_14_0_clk picorv32_pcpi_div_inst_0.quotient\[22\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2868_ _0008_ clknet_4_11_0_clk net92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_17_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1819_ picorv32_pcpi_div_inst_0.divisor\[1\] _1299_ _1295_ _1300_ _1301_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_7_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input59_I pcpi_rs2[17] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2799_ _0878_ _0903_ _0904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_63_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2896__CLK clknet_4_9_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2330__A1 _0405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_59_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_503 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2722_ picorv32_pcpi_div_inst_0.divisor\[43\] _0819_ _0838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_14_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1604_ _1030_ _1107_ _1108_ _1109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2653_ net77 _0776_ _0777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2584_ _0714_ _0398_ _0715_ _0716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_22_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1535_ picorv32_pcpi_div_inst_0.dividend\[8\] _1046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_1466_ _0982_ _0983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_38_83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_49_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2018_ picorv32_pcpi_div_inst_0.divisor\[25\] picorv32_pcpi_div_inst_0.dividend\[25\]
+ _0246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_9_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_45_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2615__A2 _1291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2303__A1 _0459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_62_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2911__CLK clknet_4_6_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_19_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2705_ picorv32_pcpi_div_inst_0.divisor\[42\] _0581_ _0823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2636_ _0754_ _0762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_6_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1518_ _0972_ _1030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_1449_ _0957_ _0967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2567_ net40 _0700_ _0701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_2498_ net31 net32 _0577_ _0622_ _0639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_0_52_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2533__A1 net35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2934__CLK clknet_4_14_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_16_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1575__A2 _1042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_355 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2283_ _0981_ _0429_ _0443_ _0136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_10_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2352_ _0431_ _0506_ _0507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2421_ _1422_ _0223_ _0567_ _0569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_19_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_67_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1802__A3 _1285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2463__C _0342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2957__CLK clknet_4_13_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2619_ _1298_ _0747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_30_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1998_ _1328_ _1095_ _0226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2515__A1 net35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input41_I pcpi_rs1[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_491 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_13_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_29_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2970_ _0124_ clknet_4_13_0_clk picorv32_pcpi_div_inst_0.quotient_msk\[23\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_56_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1921_ _1372_ _1134_ _1373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1852_ _1322_ _1321_ _1317_ _1324_ _1325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1783_ net4 _1266_ _1269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_24_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2266_ _0962_ _0426_ _0427_ _0428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2335_ net47 _0478_ _0490_ _0491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2404_ _0201_ _0553_ _0554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2197_ _0374_ _0119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_62_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_26_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2120_ _0326_ _0327_ _0089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_49_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2051_ picorv32_pcpi_div_inst_0.divisor\[59\] picorv32_pcpi_div_inst_0.divisor\[58\]
+ picorv32_pcpi_div_inst_0.divisor\[57\] picorv32_pcpi_div_inst_0.divisor\[56\] _0279_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_16_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2953_ _0107_ clknet_4_7_0_clk picorv32_pcpi_div_inst_0.quotient_msk\[6\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_44_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3008__CLK clknet_4_6_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1904_ _1356_ _1353_ _1358_ picorv32_pcpi_div_inst_0.divisor\[29\] _1359_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_32_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_32_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2884_ _0038_ clknet_4_3_0_clk picorv32_pcpi_div_inst_0.divisor\[0\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_4_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1835_ _1309_ _1308_ _1306_ _1311_ _1312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_17_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1766_ _1091_ _1248_ _1253_ _0024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1697_ picorv32_pcpi_div_inst_0.dividend\[24\] _1192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2469__B _0612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_12_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2249_ _0402_ _0410_ _0411_ _0134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2318_ _0469_ _0471_ _0475_ _0476_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_67_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_4_10_0_clk clknet_0_clk clknet_4_10_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_7_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput99 net99 pcpi_div_rd[23] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput88 net88 pcpi_div_rd[13] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__1696__A1 _1091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1482_ _0959_ _0997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1620_ _1096_ _1123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1551_ _1046_ _1044_ _0967_ _1061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_1_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2103_ _0301_ _0317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_37_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2034_ picorv32_pcpi_div_inst_0.divisor\[28\] picorv32_pcpi_div_inst_0.dividend\[28\]
+ _0262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_9_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2936_ _0090_ clknet_4_14_0_clk picorv32_pcpi_div_inst_0.quotient\[21\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1611__A1 _1113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2867_ _0007_ clknet_4_11_0_clk net91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_32_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1818_ picorv32_pcpi_div_inst_0.divisor\[2\] _1300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2798_ net66 _0902_ _0903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__1678__A1 _1091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1749_ _1116_ _1235_ _1238_ _0021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2218__I _1297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_59_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_42_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2652_ _0720_ _0756_ _0776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2721_ picorv32_pcpi_div_inst_0.divisor\[44\] _0826_ _0836_ _0837_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1603_ picorv32_pcpi_div_inst_0.quotient\[14\] _1108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1465_ _0957_ _0982_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1534_ _1041_ _1042_ _1044_ _1045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_2583_ net40 net42 _0699_ _0416_ _0715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_22_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_10_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_10_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2990__CLK clknet_4_8_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1651__B _1135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2017_ _0243_ _0244_ _0245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_65_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2919_ _0073_ clknet_4_7_0_clk picorv32_pcpi_div_inst_0.quotient\[4\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1877__I _1316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input71_I pcpi_rs2[28] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2863__CLK clknet_4_11_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_62_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_19_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2635_ _0747_ _0760_ _0761_ _0170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2704_ net52 _0821_ _0822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_6_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_49_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1448_ _0965_ _0966_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1517_ _0964_ _1029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2497_ _0414_ _0637_ _0638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2566_ _0612_ _0699_ _0700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_10_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2886__CLK clknet_4_3_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_2_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2533__A2 net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_16_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2420_ _0223_ _0567_ _1422_ _0568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__3041__CLK clknet_4_1_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_67_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2282_ _0431_ _0442_ _0443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2351_ _0489_ _0500_ _0505_ _0506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_19_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_429 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_47_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1997_ picorv32_pcpi_div_inst_0.divisor\[12\] _1078_ _0225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_19_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__1890__I _1315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2549_ _0398_ _0684_ _0685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2618_ _0744_ _0746_ _0168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input34_I pcpi_rs1[23] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2901__CLK clknet_4_9_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1493__A2 _1007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_29_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1920_ picorv32_pcpi_div_inst_0.divisor\[17\] _1372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1851_ picorv32_pcpi_div_inst_0.divisor\[11\] _1324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1782_ _1268_ _0034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_24_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2403_ _0225_ _0546_ _0553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2196_ picorv32_pcpi_div_inst_0.quotient_msk\[18\] _0369_ _0372_ picorv32_pcpi_div_inst_0.quotient_msk\[19\]
+ _0374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2265_ _0329_ _0427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2334_ _0418_ _0490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_47_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2924__CLK clknet_4_13_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2424__A1 net25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1744__B _1202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2575__B _0641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2050_ picorv32_pcpi_div_inst_0.divisor\[61\] picorv32_pcpi_div_inst_0.divisor\[60\]
+ picorv32_pcpi_div_inst_0.divisor\[62\] _0278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_2952_ _0106_ clknet_4_7_0_clk picorv32_pcpi_div_inst_0.quotient_msk\[5\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_32_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1903_ _1349_ _1358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2883_ _0037_ clknet_4_5_0_clk net116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1765_ _1037_ _1252_ _1253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_44_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_32_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1834_ picorv32_pcpi_div_inst_0.divisor\[7\] _1311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_4_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1696_ _1091_ _1187_ _1191_ _0015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2179_ picorv32_pcpi_div_inst_0.quotient_msk\[11\] _0363_ _0359_ picorv32_pcpi_div_inst_0.quotient_msk\[12\]
+ _0364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_57_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2248_ _0952_ _0305_ _0411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2317_ _1409_ _0473_ _0474_ _0475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_35_248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2406__A1 _0433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput89 net89 pcpi_div_rd[14] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_58_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1481_ _0988_ _0990_ _0996_ _0025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_22_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1550_ _1059_ _1060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2102_ _0314_ _0316_ _0082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_37_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2033_ picorv32_pcpi_div_inst_0.divisor\[29\] picorv32_pcpi_div_inst_0.dividend\[29\]
+ _0261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_27_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2479__A4 net29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2935_ _0089_ clknet_4_15_0_clk picorv32_pcpi_div_inst_0.quotient\[20\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_49_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_45_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1748_ _1153_ _1237_ _1238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2866_ _0006_ clknet_4_11_0_clk net90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_13_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2797_ net65 _0891_ _0898_ _0902_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1817_ _1298_ _1299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_40_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1679_ picorv32_pcpi_div_inst_0.dividend\[22\] _1176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_0_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_48_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_42_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1469__B _0985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1602_ _1106_ _1107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2144__I _0290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2582_ net43 _0714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2651_ _0432_ _0775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2720_ _0811_ _0835_ _0836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_59_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1533_ _1043_ _1044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1464_ _0980_ _0981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_10_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_65_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2085__A2 _0305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2016_ picorv32_pcpi_div_inst_0.divisor\[26\] picorv32_pcpi_div_inst_0.dividend\[26\]
+ _0244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XPHY_EDGE_ROW_19_Left_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_64_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2918_ _0072_ clknet_4_7_0_clk picorv32_pcpi_div_inst_0.quotient\[3\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_9_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2849_ _0035_ clknet_4_4_0_clk picorv32_pcpi_div_inst_0.instr_rem vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_13_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input64_I pcpi_rs2[21] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_19_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1578__A1 picorv32_pcpi_div_inst_0.dividend\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_27_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1516_ _0988_ _1023_ _1028_ _0028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_42_357 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2634_ picorv32_pcpi_div_inst_0.divisor\[32\] _0751_ _0761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2565_ net38 net39 _0682_ _0699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_2703_ net82 _0814_ _0812_ _0821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_10_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1447_ _0964_ _0965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2496_ _0237_ _0636_ _0637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_53_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3048_ net116 net118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_2_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2980__CLK clknet_4_3_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_4_6_0_clk_I clknet_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_10_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_10_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_67_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_32_Left_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2281_ _0433_ _0436_ _0438_ _0441_ _0442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__2288__A2 _0981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2350_ _0502_ _0503_ _0504_ _0505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_35_20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_51_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1996_ _1328_ _1095_ _0224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_15_324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2548_ net38 _0460_ _0682_ _0684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_2617_ _0737_ _0297_ _0745_ _0746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_23_390 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2853__CLK clknet_4_12_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2479_ net26 net27 net28 net29 _0622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XANTENNA_input27_I pcpi_rs1[17] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2242__I _0404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_21_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_29_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1781_ net4 _1254_ _1255_ _1267_ _1268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_0_24_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1850_ _1323_ _0047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_4_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_12_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2876__CLK clknet_4_12_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2402_ net23 _0551_ _0552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_20_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2333_ _0432_ _0489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2195_ _0373_ _0118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2264_ _0414_ _0421_ _0422_ _0425_ _0426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_47_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_35_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1979_ picorv32_pcpi_div_inst_0.divisor\[9\] picorv32_pcpi_div_inst_0.dividend\[9\]
+ _0207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_15_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3031__CLK clknet_4_0_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_7_Left_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2700__I _0387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2899__CLK clknet_4_9_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2951_ _0105_ clknet_4_7_0_clk picorv32_pcpi_div_inst_0.quotient_msk\[4\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1902_ _1357_ _0065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_29_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2882_ _0024_ clknet_4_12_0_clk net108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1764_ _1249_ _1251_ _1252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_32_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1833_ _1310_ _0043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_12_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1695_ _1037_ _1190_ _1191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2316_ _1409_ _0473_ _0449_ _0474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2178_ _0362_ _0363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_48_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2247_ _0403_ _0405_ _0409_ _0410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_clkbuf_4_14_0_clk_I clknet_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_499 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_19_Right_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_22_433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1480_ _0992_ _0994_ _0995_ _0996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_28_Right_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_1_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2101_ picorv32_pcpi_div_inst_0.quotient_msk\[13\] _0310_ picorv32_pcpi_div_inst_0.quotient\[13\]
+ _0316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2914__CLK clknet_4_4_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_37_Right_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_37_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2032_ _0252_ _0259_ _0260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_27_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2934_ _0088_ clknet_4_14_0_clk picorv32_pcpi_div_inst_0.quotient\[19\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_57_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2865_ _0005_ clknet_4_14_0_clk net89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_45_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1747_ picorv32_pcpi_div_inst_0.quotient\[29\] _1236_ _1237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_1678_ _1091_ _1171_ _1175_ _0013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_46_Right_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1816_ _1297_ _1298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_40_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2572__A1 net42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_7_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2796_ _0897_ _0396_ _0900_ _0901_ _0191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_13_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_13_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_55_Right_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_67_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_64_Right_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2937__CLK clknet_4_14_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2250__I _1364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_42_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1601_ _1051_ _1031_ _1087_ _1105_ _1106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_0_54_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1532_ _1035_ _1034_ _1043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_2650_ _0769_ _0773_ _0774_ _0172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2581_ _0269_ _0712_ _0713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__2554__A1 net39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_425 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input1_I pcpi_div_valid vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1463_ picorv32_pcpi_div_inst_0.dividend\[2\] _0980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_2015_ _0242_ _0243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_9_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2917_ _0071_ clknet_4_5_0_clk picorv32_pcpi_div_inst_0.quotient\[2\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_45_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2848_ _0034_ clknet_4_4_0_clk picorv32_pcpi_div_inst_0.instr_divu vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1596__A2 _1078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input57_I pcpi_rs2[15] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2779_ net63 _0886_ _0887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__1520__A2 _1031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_5_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_4_2_0_clk_I clknet_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_20_Left_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2224__B1 _1294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_42_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2702_ _0795_ _0818_ _0820_ _0178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_24_77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1515_ _1025_ _1026_ _1027_ _1028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2633_ picorv32_pcpi_div_inst_0.divisor\[33\] _0753_ _0759_ _0760_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2564_ _0261_ _0697_ _0698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2495_ _0231_ _0620_ _1389_ _0636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2527__A1 _0424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1446_ picorv32_pcpi_div_inst_0.instr_divu picorv32_pcpi_div_inst_0.instr_div _0964_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_2_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_61_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_53_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3047_ _0199_ clknet_4_3_0_clk picorv32_pcpi_div_inst_0.divisor\[61\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_18_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2766__A1 _0405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2206__B1 _0378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1980__A2 _1046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_67_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2280_ _0439_ _0440_ _0441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_19_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_15_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2616_ _0416_ _0736_ _0745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_2_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1995_ _0222_ picorv32_pcpi_div_inst_0.dividend\[14\] _0223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1429_ _0949_ _0032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2478_ _0618_ _0620_ _0621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2547_ _0456_ _0682_ net38 _0683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_46_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1780_ _1266_ _1267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_24_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_12_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2401_ net22 _0540_ _0445_ _0551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2332_ _0454_ _0487_ _0488_ _0140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2194_ picorv32_pcpi_div_inst_0.quotient_msk\[17\] _0369_ _0372_ picorv32_pcpi_div_inst_0.quotient_msk\[18\]
+ _0373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__1469__A1 _0981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2263_ _0424_ _1401_ _0425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_47_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_35_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_23_Left_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_1_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1978_ picorv32_pcpi_div_inst_0.divisor\[10\] picorv32_pcpi_div_inst_0.dividend\[10\]
+ _0206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_15_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2970__CLK clknet_4_13_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_4_10_0_clk_I clknet_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_51_Left_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_61_250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_60_Left_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1699__A1 _0983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2950_ _0104_ clknet_4_5_0_clk picorv32_pcpi_div_inst_0.quotient_msk\[3\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2881_ _0023_ clknet_4_6_0_clk net107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1901_ picorv32_pcpi_div_inst_0.divisor\[27\] _1353_ _1350_ _1356_ _1357_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_32_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1832_ picorv32_pcpi_div_inst_0.divisor\[5\] _1308_ _1306_ _1309_ _1310_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_8_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1694_ _1188_ _1189_ _1190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1763_ _0967_ _1250_ _1251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_4_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1507__I picorv32_pcpi_div_inst_0.outsign vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2246_ _0407_ _0408_ _0409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2315_ _0463_ _0464_ _0472_ _0473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2993__CLK clknet_4_8_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2177_ _1297_ _0362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_48_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_23_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2073__I _0297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2866__CLK clknet_4_11_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2100_ _0314_ _0315_ _0081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_45_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_37_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2031_ _0241_ picorv32_pcpi_div_inst_0.dividend\[27\] _0245_ _0258_ _0259_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_27_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2933_ _0087_ clknet_4_15_0_clk picorv32_pcpi_div_inst_0.quotient\[18\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2864_ _0004_ clknet_4_14_0_clk net88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_45_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1815_ _1289_ _1297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2795_ picorv32_pcpi_div_inst_0.divisor\[54\] _0808_ _0809_ _0901_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1746_ _1224_ _1223_ _0958_ _1236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1677_ _1037_ _1174_ _1175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3021__CLK clknet_4_4_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2229_ _0393_ _0132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2889__CLK clknet_4_2_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2012__A1 _0211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_42_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3044__CLK clknet_4_2_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1600_ picorv32_pcpi_div_inst_0.quotient\[12\] picorv32_pcpi_div_inst_0.quotient\[13\]
+ _1105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1462_ picorv32_pcpi_div_inst_0.quotient\[2\] _0978_ _0979_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1531_ _0983_ _1042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2580_ _0706_ _0271_ _0711_ _0712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_1_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2014_ _0241_ picorv32_pcpi_div_inst_0.dividend\[27\] _0242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_9_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2916_ _0070_ clknet_4_7_0_clk picorv32_pcpi_div_inst_0.quotient\[1\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_45_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2847_ _0944_ _0199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_5_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2778_ _0728_ _0804_ _0886_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1729_ picorv32_pcpi_div_inst_0.quotient\[27\] _1220_ _1221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_TAPCELL_ROW_56_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_5_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1586__B _1021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2904__CLK clknet_4_10_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2261__I _1364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2472__A1 _0586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2171__I _1315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_40_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2632_ _0519_ _0758_ _0759_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_27_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2701_ picorv32_pcpi_div_inst_0.divisor\[40\] _0819_ _0820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_6_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1445_ _0952_ _0960_ _0962_ _0963_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1514_ _1025_ _1026_ _0985_ _1027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2494_ _0635_ _0155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2563_ _0696_ _1228_ _0691_ _0697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_2_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3046_ _0198_ clknet_4_3_0_clk picorv32_pcpi_div_inst_0.divisor\[60\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2927__CLK clknet_4_15_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_61_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_53_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_37_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2463__A1 _0598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_18_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_359 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1425__I _0945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2206__B2 picorv32_pcpi_div_inst_0.quotient_msk\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_32_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_67_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2166__I _1352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2445__A1 _0211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_15_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1994_ picorv32_pcpi_div_inst_0.divisor\[14\] _0222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_42_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2615_ picorv32_pcpi_div_inst_0.divisor\[62\] _1291_ _0744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1428_ picorv32_pcpi_div_inst_0.instr_remu picorv32_pcpi_div_inst_0.instr_rem _0947_
+ _0948_ _0949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_2477_ _1376_ _1381_ _0619_ _0620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_2546_ net37 _0670_ _0682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__2436__A1 _0581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3029_ _0181_ clknet_4_1_0_clk picorv32_pcpi_div_inst_0.divisor\[43\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_46_495 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_12_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2400_ _1078_ _0508_ _0550_ _0146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_46_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2262_ _0423_ _0424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_20_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_351 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2331_ _1024_ _0292_ _0488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2193_ _0358_ _0372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_46_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2418__A1 _0454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1977_ picorv32_pcpi_div_inst_0.divisor\[11\] picorv32_pcpi_div_inst_0.dividend\[11\]
+ _0205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_2529_ net36 _0666_ _0667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_11_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input32_I pcpi_rs1[21] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2409__A1 net22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2709__I _0782_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2880_ _0021_ clknet_4_12_0_clk net105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_37_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1900_ picorv32_pcpi_div_inst_0.divisor\[28\] _1356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_29_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1831_ picorv32_pcpi_div_inst_0.divisor\[6\] _1309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_52_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1693_ picorv32_pcpi_div_inst_0.dividend\[22\] _1178_ _1096_ _1189_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1762_ _1239_ _1233_ _1228_ _1230_ _1250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_0_12_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2176_ _0361_ _0111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2619__I _1298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2639__A1 _0519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2245_ _1399_ picorv32_pcpi_div_inst_0.dividend\[0\] _0408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2314_ _1418_ _1005_ _0472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_48_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_23_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_31_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_1_Right_1 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_66_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1608__I _0955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2030_ _0254_ _0256_ _0257_ _0258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2439__I _0449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2932_ _0086_ clknet_4_14_0_clk picorv32_pcpi_div_inst_0.quotient\[17\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_45_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_37_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2960__CLK clknet_4_13_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1745_ _1233_ _1234_ _1235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2863_ _0003_ clknet_4_11_0_clk net87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_40_210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1814_ _1296_ _0038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_25_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2794_ _0399_ _0899_ _0900_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_40_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1676_ _1172_ _1173_ _1174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2159_ picorv32_pcpi_div_inst_0.quotient_msk\[4\] _0349_ _0346_ picorv32_pcpi_div_inst_0.quotient_msk\[5\]
+ _0351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2228_ picorv32_pcpi_div_inst_0.quotient_msk\[31\] _1291_ _0297_ _0393_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__1532__A1 _1035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1599__A1 _1100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_8_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2983__CLK clknet_4_3_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1461_ _0953_ _0971_ _0977_ _0978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_22_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1530_ _1040_ _1041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__1514__A1 _1025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2013_ picorv32_pcpi_div_inst_0.divisor\[27\] _0241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2915_ _0069_ clknet_4_6_0_clk picorv32_pcpi_div_inst_0.quotient\[0\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1728_ _1209_ _1208_ _0958_ _1220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2846_ _0943_ picorv32_pcpi_div_inst_0.divisor\[61\] _0395_ _0944_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2777_ picorv32_pcpi_div_inst_0.divisor\[51\] _0885_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2856__CLK clknet_4_6_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1659_ picorv32_pcpi_div_inst_0.dividend\[20\] _1158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__1505__A1 _1016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output101_I net101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_56_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_64_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3011__CLK clknet_4_3_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2562_ _1356_ _0696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2631_ net62 _0757_ _0758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2700_ _0387_ _0819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_2_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_15_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2879__CLK clknet_4_12_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1513_ _1016_ _1017_ _0959_ _1026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2493_ picorv32_pcpi_div_inst_0.dividend\[21\] _0633_ _0634_ _0635_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1444_ _0961_ _0962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_4_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_53_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1531__I _0983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3045_ _0197_ clknet_4_2_0_clk picorv32_pcpi_div_inst_0.divisor\[59\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_61_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_18_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input62_I pcpi_rs2[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2829_ _0912_ _0928_ _0929_ _0196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3034__CLK clknet_4_0_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_1_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2272__I _0432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_15_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1993_ _0220_ picorv32_pcpi_div_inst_0.dividend\[15\] _0221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2614_ _1254_ _1255_ _1269_ _0167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_42_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2545_ _0242_ _0680_ _0681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_23_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1427_ net83 _0948_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2476_ _0591_ _0235_ _0619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1892__B1 _1350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3028_ _0180_ clknet_4_1_0_clk picorv32_pcpi_div_inst_0.divisor\[42\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_61_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_12_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2192_ _0371_ _0117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2177__I _1297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2261_ _1364_ _0423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2330_ _0405_ _0480_ _0483_ _0486_ _0487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_55_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1976_ _0200_ _0203_ _0204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2528_ net35 _0652_ _0612_ _0666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_11_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2087__I _0297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2459_ _0603_ _0604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2409__A2 net23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input25_I pcpi_rs1[15] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_26_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1761_ picorv32_pcpi_div_inst_0.dividend\[31\] _1249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_1830_ _1298_ _1308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_40_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1692_ picorv32_pcpi_div_inst_0.dividend\[23\] _1188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_25_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2313_ net46 _0470_ _0471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2175_ picorv32_pcpi_div_inst_0.quotient_msk\[10\] _0355_ _0359_ picorv32_pcpi_div_inst_0.quotient_msk\[11\]
+ _0361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2244_ _0406_ _0407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_48_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_23_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_31_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1959_ _1409_ _1410_ _1411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_16_433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_499 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2566__A1 _0612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2318__A1 _0469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1541__A2 _1031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2931_ _0085_ clknet_4_14_0_clk picorv32_pcpi_div_inst_0.quotient\[16\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_45_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_0_clk clk clknet_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_2862_ _0002_ clknet_4_13_0_clk net86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1744_ _1229_ _1230_ _1202_ _1234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_40_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1813_ picorv32_pcpi_div_inst_0.divisor\[0\] _1291_ _1295_ picorv32_pcpi_div_inst_0.divisor\[1\]
+ _1296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_7_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2793_ net65 _0898_ _0899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1675_ picorv32_pcpi_div_inst_0.dividend\[20\] _1160_ _1096_ _1173_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1532__A2 _1034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2309__A1 _1005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_15_Right_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2158_ _0350_ _0104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2089_ _0307_ _0308_ _0077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2227_ _0392_ _0131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_48_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_24_Right_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2365__I _1364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_39_Left_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_33_Right_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2548__A1 net38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_16_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_59_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_48_Left_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_42_Right_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_57_Left_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_54_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_51_Right_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2539__A1 _0658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1460_ _0972_ _0977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_38_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_66_Left_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_60_Right_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_54_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2012_ _0211_ _0230_ _0239_ _0240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_2914_ _0068_ clknet_4_4_0_clk picorv32_pcpi_div_inst_0.divisor\[30\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2845_ _0469_ _0941_ _0942_ _0943_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_5_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1658_ _1112_ _1152_ _1157_ _0010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1727_ _1217_ _1218_ _1219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2776_ _0867_ _0882_ _0884_ _0188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_13_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1589_ _1094_ _1095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_64_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_56_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1439__I picorv32_pcpi_div_inst_0.outsign vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_67_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2209__B1 _0378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2561_ _0695_ _0162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2492_ _0430_ _0634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_2630_ _0748_ _0756_ _0757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1512_ _1024_ _1025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_1443_ picorv32_pcpi_div_inst_0.dividend\[1\] _0961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_10_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1812__I _1294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_53_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1671__B2 _1169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3044_ _0196_ clknet_4_2_0_clk picorv32_pcpi_div_inst_0.divisor\[58\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_18_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_61_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2828_ picorv32_pcpi_div_inst_0.divisor\[58\] _0923_ _0929_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1974__A2 picorv32_pcpi_div_inst_0.dividend\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2759_ _0846_ _0869_ _0870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_input55_I pcpi_rs2[13] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_1_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1965__A2 _1016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_35_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_15_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1992_ picorv32_pcpi_div_inst_0.divisor\[15\] _0220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2613_ _0743_ _0166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2475_ _1383_ _1384_ _0618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2544_ _0251_ _1213_ _0674_ _0680_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__1807__I _1289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2996__CLK clknet_4_9_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_66_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1426_ _0946_ _0947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_3027_ _0179_ clknet_4_1_0_clk picorv32_pcpi_div_inst_0.divisor\[41\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_61_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3001__CLK clknet_4_11_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2869__CLK clknet_4_11_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1635__A1 _1134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_353 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2191_ picorv32_pcpi_div_inst_0.quotient_msk\[16\] _0369_ _0366_ picorv32_pcpi_div_inst_0.quotient_msk\[17\]
+ _0371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_46_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2260_ _1399_ _0951_ _1400_ _0422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_47_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3024__CLK clknet_4_1_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1975_ _0201_ _0202_ _0203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_2527_ _0424_ _0664_ _0665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2458_ _0579_ net27 _0577_ _0603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA_input18_I pcpi_insn[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_26_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2389_ net47 net48 _0478_ _0539_ _0540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XTAP_TAPCELL_ROW_34_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1447__I _0964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2281__A1 _0433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3047__CLK clknet_4_3_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1691_ picorv32_pcpi_div_inst_0.quotient\[23\] _1186_ _1187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1760_ picorv32_pcpi_div_inst_0.quotient\[31\] _1247_ _1248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__2584__A2 _0398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2188__I _0362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_27_Left_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2312_ net45 _0457_ _0419_ _0470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2174_ _0360_ _0110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_57_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_48_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2243_ _0397_ _0406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_11_Left_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2651__I _0432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_23_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1889_ _1348_ _0061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_31_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_31_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1958_ picorv32_pcpi_div_inst_0.divisor\[4\] picorv32_pcpi_div_inst_0.dividend\[4\]
+ _1410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_16_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2098__I _0313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2263__A1 _0424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2907__CLK clknet_4_10_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2930_ _0084_ clknet_4_15_0_clk picorv32_pcpi_div_inst_0.quotient\[15\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_57_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2861_ _0001_ clknet_4_12_0_clk net85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1674_ picorv32_pcpi_div_inst_0.dividend\[21\] _1172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_1743_ picorv32_pcpi_div_inst_0.dividend\[29\] _1233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2309__A2 _0305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2792_ _0728_ _0729_ _0803_ _0898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1812_ _1294_ _1295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2226_ picorv32_pcpi_div_inst_0.quotient_msk\[30\] _0388_ _1294_ picorv32_pcpi_div_inst_0.quotient_msk\[31\]
+ _0392_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__1815__I _1289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2157_ picorv32_pcpi_div_inst_0.quotient_msk\[3\] _0349_ _0346_ picorv32_pcpi_div_inst_0.quotient_msk\[4\]
+ _0350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2088_ picorv32_pcpi_div_inst_0.quotient_msk\[8\] _0302_ _1050_ _0308_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_48_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_59_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2484__A1 _0598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2236__A1 picorv32_pcpi_div_inst_0.running vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_429 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_54_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2011_ _0231_ _0235_ _0237_ _0238_ _0239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_57_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2913_ _0067_ clknet_4_4_0_clk picorv32_pcpi_div_inst_0.divisor\[29\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2844_ picorv32_pcpi_div_inst_0.divisor\[62\] _0424_ _0942_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1986__B1 _1041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1657_ _1153_ _1156_ _1157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1726_ _1213_ _1214_ _1202_ _1218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1588_ picorv32_pcpi_div_inst_0.dividend\[13\] _1094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2775_ picorv32_pcpi_div_inst_0.divisor\[50\] _0883_ _0884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_0_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_13_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2209_ picorv32_pcpi_div_inst_0.quotient_msk\[23\] _0381_ _0378_ picorv32_pcpi_div_inst_0.quotient_msk\[24\]
+ _0382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_56_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_64_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_14_Left_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_63_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1901__B1 _1350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2209__A1 picorv32_pcpi_div_inst_0.quotient_msk\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_4_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_315 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1442_ _0959_ _0960_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_49_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2560_ _1229_ _0694_ _0678_ _0695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_35_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2491_ _0414_ _0629_ _0632_ _0633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1511_ picorv32_pcpi_div_inst_0.dividend\[6\] _1024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_65_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3043_ _0195_ clknet_4_2_0_clk picorv32_pcpi_div_inst_0.divisor\[57\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_53_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_18_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_61_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2758_ net59 _0868_ _0869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2827_ picorv32_pcpi_div_inst_0.divisor\[59\] _0466_ _0927_ _0928_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1709_ _1192_ _1193_ _1202_ _1203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2689_ _1290_ _0809_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_1_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_input48_I pcpi_rs1[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_1_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1662__A2 _0997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_55_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2612_ _1042_ _0742_ _1366_ _0743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1991_ _0215_ _0218_ _0200_ _0203_ _0219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_TAPCELL_ROW_15_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1425_ _0945_ _0946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2543_ _0679_ _0160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2474_ _0617_ _0153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_66_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1892__A2 _1343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3026_ _0178_ clknet_4_1_0_clk picorv32_pcpi_div_inst_0.divisor\[40\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_58_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1644__A2 _1042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2841__A1 _1291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2940__CLK clknet_4_13_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1883__A2 _1343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_29_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2190_ _0370_ _0116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2963__CLK clknet_4_15_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1974_ picorv32_pcpi_div_inst_0.divisor\[12\] picorv32_pcpi_div_inst_0.dividend\[12\]
+ _0202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_30_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_39_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2526_ _0246_ _0256_ _0659_ _0664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_2457_ _0599_ _0601_ _0602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_11_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2388_ net49 net50 net20 net21 _0539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_0_66_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3009_ _0163_ clknet_4_3_0_clk picorv32_pcpi_div_inst_0.dividend\[29\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_26_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_34_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2508__B _0612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2986__CLK clknet_4_2_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1690_ picorv32_pcpi_div_inst_0.quotient\[22\] _1183_ _1135_ _1186_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_25_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_2_Left_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_0_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_57_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2242_ _0404_ _0405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2311_ _0413_ _0469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2173_ picorv32_pcpi_div_inst_0.quotient_msk\[9\] _0355_ _0359_ picorv32_pcpi_div_inst_0.quotient_msk\[10\]
+ _0360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_48_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_31_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_23_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1957_ picorv32_pcpi_div_inst_0.divisor\[5\] picorv32_pcpi_div_inst_0.dividend\[5\]
+ _1409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_16_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2859__CLK clknet_4_12_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1888_ _1346_ _1343_ _1340_ picorv32_pcpi_div_inst_0.divisor\[24\] _1348_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2509_ net34 _0648_ _0649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA_input30_I pcpi_rs1[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1526__A1 _1035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3014__CLK clknet_4_4_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_57_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2860_ _0031_ clknet_4_12_0_clk net115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_45_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1811_ _1293_ _1294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_43_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2791_ picorv32_pcpi_div_inst_0.divisor\[53\] _0897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1673_ picorv32_pcpi_div_inst_0.quotient\[21\] _1170_ _1171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__1765__A1 _1037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1742_ _1225_ _1227_ _1232_ _1010_ _0020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_40_213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_0_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2225_ _0391_ _0130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_0_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2156_ _1352_ _0349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2087_ _0297_ _0307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_36_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_36_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_5_Right_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_17_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1756__A1 _0977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input78_I pcpi_rs2[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2989_ _0143_ clknet_4_8_0_clk picorv32_pcpi_div_inst_0.dividend\[9\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3037__CLK clknet_4_0_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_59_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2010_ picorv32_pcpi_div_inst_0.divisor\[23\] picorv32_pcpi_div_inst_0.dividend\[23\]
+ _0238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2912_ _0066_ clknet_4_4_0_clk picorv32_pcpi_div_inst_0.divisor\[28\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_18_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1725_ picorv32_pcpi_div_inst_0.dividend\[27\] _1217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2843_ _0719_ _0940_ _0941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2774_ _0394_ _0883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1587_ picorv32_pcpi_div_inst_0.quotient\[13\] _1092_ _1093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1656_ picorv32_pcpi_div_inst_0.quotient\[19\] _1155_ _1156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_13_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2208_ _0362_ _0381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_56_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2139_ _1366_ _0339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_64_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_4_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1510_ picorv32_pcpi_div_inst_0.quotient\[6\] _1022_ _1023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1441_ _0958_ _0959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_50_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2490_ _1382_ _0630_ _0631_ _0632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3042_ _0194_ clknet_4_2_0_clk picorv32_pcpi_div_inst_0.divisor\[56\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_4_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_61_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_18_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1708_ _1020_ _1202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_41_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2688_ _0641_ _0808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_5_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2757_ net58 _0861_ _0840_ _0868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2826_ _0918_ _0926_ _0927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1639_ _1116_ _1140_ _1141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_41_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_1_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2127__A1 picorv32_pcpi_div_inst_0.quotient_msk\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_59_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1990_ _0216_ _0217_ _0218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_42_149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2542_ _1213_ _0677_ _0678_ _0679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2611_ _0738_ _0740_ _0741_ _0742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_27_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1424_ picorv32_pcpi_div_inst_0.instr_divu picorv32_pcpi_div_inst_0.instr_div _0945_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_2473_ _1150_ _0616_ _0574_ _0617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__2892__CLK clknet_4_8_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3025_ _0177_ clknet_4_1_0_clk picorv32_pcpi_div_inst_0.divisor\[39\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_41_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_input60_I pcpi_rs2[18] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2809_ _1298_ _0912_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_1_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_29_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1973_ picorv32_pcpi_div_inst_0.divisor\[13\] picorv32_pcpi_div_inst_0.dividend\[13\]
+ _0201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2525_ _0256_ _0659_ _0246_ _0663_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_11_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2456_ _0584_ _0234_ _0600_ _0601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2387_ _0454_ _0537_ _0538_ _0145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3008_ _0162_ clknet_4_6_0_clk picorv32_pcpi_div_inst_0.dividend\[28\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_26_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_34_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2502__A1 net33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2172_ _0358_ _0359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_57_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2241_ _0397_ _0404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2310_ _0454_ _0467_ _0468_ _0138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2930__CLK clknet_4_15_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_23_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1887_ _1347_ _0060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_31_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1956_ _1406_ _1407_ _1408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2508_ net33 _0639_ _0612_ _0648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_3_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_39_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2439_ _0449_ _0586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA_input23_I pcpi_rs1[13] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_22_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_57_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1741_ _1229_ _1231_ _1232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1810_ _1292_ _1289_ _1293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2790_ _0867_ _0895_ _0896_ _0190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1672_ picorv32_pcpi_div_inst_0.quotient\[20\] _1166_ _1135_ _1170_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2155_ _0348_ _0103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2224_ picorv32_pcpi_div_inst_0.quotient_msk\[29\] _0388_ _1294_ picorv32_pcpi_div_inst_0.quotient_msk\[30\]
+ _0391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_36_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2086_ _1051_ _0306_ _1367_ _0076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_48_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1939_ picorv32_pcpi_div_inst_0.divisor\[22\] _1176_ _1391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_31_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2988_ _0142_ clknet_4_8_0_clk picorv32_pcpi_div_inst_0.dividend\[8\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_7_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_59_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_54_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_42_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_11_Right_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_62_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_20_Right_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_54_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_7_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2849__CLK clknet_4_4_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2911_ _0065_ clknet_4_6_0_clk picorv32_pcpi_div_inst_0.divisor\[27\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_35_Left_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1986__A2 _1060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_394 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1724_ _1210_ _1212_ _1216_ _1010_ _0018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XPHY_EDGE_ROW_44_Left_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2999__CLK clknet_4_9_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2842_ _0735_ _0804_ _0940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2773_ picorv32_pcpi_div_inst_0.divisor\[51\] _0855_ _0881_ _0882_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1586_ picorv32_pcpi_div_inst_0.quotient\[12\] _1088_ _1021_ _1092_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1655_ _0982_ _1154_ _1155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1910__A2 _1360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1842__I _1316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2207_ _0380_ _0123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2069_ _1367_ _0295_ _0070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2138_ _0333_ _0338_ _0096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_EDGE_ROW_53_Left_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_64_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_62_Left_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_48_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_36_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3004__CLK clknet_4_12_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2154__A2 _1360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_4_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1440_ _0957_ _0958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2145__A2 _0342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3041_ _0193_ clknet_4_1_0_clk picorv32_pcpi_div_inst_0.divisor\[55\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_61_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_45_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3027__CLK clknet_4_1_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2825_ net70 _0925_ _0926_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_18_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_18_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1638_ _1138_ _1139_ _1140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_1707_ picorv32_pcpi_div_inst_0.dividend\[25\] _1201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2687_ _0399_ _0806_ _0807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2756_ _0768_ _0867_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1569_ _1029_ _1076_ _1077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1572__I picorv32_pcpi_div_inst_0.dividend\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_52_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_1_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_64_423 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_9_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2541_ _0291_ _0678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_2610_ picorv32_pcpi_div_inst_0.instr_rem _0714_ _0741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2472_ _0586_ _0611_ _0615_ _0616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_2_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3024_ _0176_ clknet_4_1_0_clk picorv32_pcpi_div_inst_0.divisor\[38\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_46_423 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2808_ _0907_ _0747_ _0910_ _0911_ _0193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_41_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2739_ _0394_ _0853_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_14_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input53_I pcpi_rs2[11] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_29_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1972_ _1422_ _1423_ _0200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_51_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_49_Right_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2524_ _0662_ _0158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2455_ _1373_ _1375_ _0600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_11_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_58_Right_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2386_ picorv32_pcpi_div_inst_0.dividend\[11\] _0292_ _0538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_34_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3007_ _0161_ clknet_4_3_0_clk picorv32_pcpi_div_inst_0.dividend\[27\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2275__A1 net41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_26_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_67_Right_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_61_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_61_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2882__CLK clknet_4_12_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2171_ _1315_ _0358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2240_ net19 _0403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_7_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_43_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1886_ _1344_ _1343_ _1340_ _1346_ _1347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_31_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1955_ picorv32_pcpi_div_inst_0.divisor\[6\] picorv32_pcpi_div_inst_0.dividend\[6\]
+ _1407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_16_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2507_ _0238_ _0646_ _0647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2438_ _0584_ _0233_ _0585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_11_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input16_I pcpi_insn[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_39_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2248__A1 _0952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2369_ _0520_ _0521_ _0522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_34_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1526__A3 _1034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2487__A1 net32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1671_ _1161_ _1163_ _1168_ _1169_ _0012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1740_ _1006_ _1230_ _1231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_25_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_13_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input8_I pcpi_insn[26] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2154_ picorv32_pcpi_div_inst_0.quotient_msk\[2\] _1360_ _0346_ picorv32_pcpi_div_inst_0.quotient_msk\[3\]
+ _0348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2085_ picorv32_pcpi_div_inst_0.quotient_msk\[7\] _0305_ _0306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2223_ _0390_ _0129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_17_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_48_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2987_ _0141_ clknet_4_8_0_clk picorv32_pcpi_div_inst_0.dividend\[7\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_8_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1938_ _1344_ _1177_ _1386_ _1389_ _1390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_31_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput80 pcpi_rs2[7] net80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2705__A2 _0581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2402__A1 net23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1869_ _1335_ _0054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__1524__B _1035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_50_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_42_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_7_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2910_ _0064_ clknet_4_11_0_clk picorv32_pcpi_div_inst_0.divisor\[26\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2632__A1 _0519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2841_ _1291_ _0938_ _0939_ _0198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1654_ picorv32_pcpi_div_inst_0.quotient\[16\] _1138_ picorv32_pcpi_div_inst_0.quotient\[18\]
+ _1131_ _1154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or4_1
X_1723_ _1213_ _1215_ _1216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_0_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2772_ _0878_ _0880_ _0881_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_13_248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2206_ picorv32_pcpi_div_inst_0.quotient_msk\[22\] _0375_ _0378_ picorv32_pcpi_div_inst_0.quotient_msk\[23\]
+ _0380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1585_ _0966_ _1091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_28_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2137_ picorv32_pcpi_div_inst_0.quotient_msk\[27\] _0336_ picorv32_pcpi_div_inst_0.quotient\[27\]
+ _0338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2068_ picorv32_pcpi_div_inst_0.quotient_msk\[1\] _0294_ _0971_ _0295_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_48_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_64_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_input83_I resetn vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_4_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_55_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3040_ _0192_ clknet_4_0_0_clk picorv32_pcpi_div_inst_0.divisor\[54\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2966__CLK clknet_4_15_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_14_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2824_ _0733_ _0848_ _0925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1637_ _1129_ _1131_ _0982_ _1139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1706_ _1195_ _1197_ _1200_ _1169_ _0016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__1592__A1 _1095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2686_ net81 _0805_ _0806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2755_ _0839_ _0865_ _0866_ _0185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_18_Left_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1499_ _0960_ _1011_ _1012_ _1013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1568_ _1074_ _1075_ _1076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_52_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_1_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_44_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1886__A2 _1343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_9_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2989__CLK clknet_4_8_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1810__A2 _1289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2540_ _0444_ _0672_ _0674_ _0676_ _0677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_2471_ _0581_ _0614_ _0615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_23_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3023_ _0175_ clknet_4_1_0_clk picorv32_pcpi_div_inst_0.divisor\[37\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_58_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2807_ picorv32_pcpi_div_inst_0.divisor\[56\] _0808_ _0809_ _0911_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2738_ picorv32_pcpi_div_inst_0.divisor\[46\] _0826_ _0851_ _0852_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2669_ net79 _0790_ _0791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA_input46_I pcpi_rs1[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_29_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_12_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1556__A1 _0993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3017__CLK clknet_4_4_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_55_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1971_ picorv32_pcpi_div_inst_0.divisor\[14\] picorv32_pcpi_div_inst_0.dividend\[14\]
+ _1423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2523_ _1192_ _0661_ _0634_ _0662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2454_ _1370_ _0599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2385_ _0534_ _0536_ _0459_ _0537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xinput1 pcpi_div_valid net1 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3006_ _0160_ clknet_4_6_0_clk picorv32_pcpi_div_inst_0.dividend\[26\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_52_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_34_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1538__A1 _1046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_0_clk_I clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_4_9_0_clk_I clknet_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2170_ _0357_ _0109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_28_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1954_ picorv32_pcpi_div_inst_0.divisor\[7\] picorv32_pcpi_div_inst_0.dividend\[7\]
+ _1406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_51_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1885_ picorv32_pcpi_div_inst_0.divisor\[23\] _1346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_31_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2506_ _0236_ _0636_ _0645_ _0646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2437_ _0211_ _0230_ _0584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_11_176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2368_ net49 net50 _0498_ _0521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_39_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_39_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2248__A2 _0305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2692__I _0432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2299_ net45 _0456_ _0457_ _0458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_TAPCELL_ROW_22_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_6_Left_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_45_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1670_ _1048_ _1169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_7_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2222_ picorv32_pcpi_div_inst_0.quotient_msk\[28\] _0388_ _0384_ picorv32_pcpi_div_inst_0.quotient_msk\[29\]
+ _0390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2153_ _0347_ _0102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2084_ _0291_ _0305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1937_ _1387_ _1388_ _1389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_8_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2986_ _0140_ clknet_4_2_0_clk picorv32_pcpi_div_inst_0.dividend\[6\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1856__I _1316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1799_ picorv32_pcpi_div_inst_0.quotient_msk\[18\] picorv32_pcpi_div_inst_0.quotient_msk\[17\]
+ picorv32_pcpi_div_inst_0.quotient_msk\[16\] picorv32_pcpi_div_inst_0.quotient_msk\[15\]
+ _1283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_31_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput81 pcpi_rs2[8] net81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1868_ picorv32_pcpi_div_inst_0.divisor\[16\] _1330_ _1334_ picorv32_pcpi_div_inst_0.divisor\[17\]
+ _1335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xinput70 pcpi_rs2[27] net70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2872__CLK clknet_4_11_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_42_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_50_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_58_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_7_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2771_ net61 _0879_ _0880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2840_ picorv32_pcpi_div_inst_0.divisor\[60\] _0923_ _0939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2396__A1 _0404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1653_ _0946_ _1153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1584_ _1082_ _1085_ _1090_ _1055_ _0003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1722_ _1006_ _1214_ _1215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_21_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_0_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2895__CLK clknet_4_8_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_9_Right_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_13_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2205_ _0379_ _0122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_28_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_0_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_64_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2067_ _0291_ _0294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2136_ _0333_ _0337_ _0095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_48_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2969_ _0123_ clknet_4_15_0_clk picorv32_pcpi_div_inst_0.quotient_msk\[22\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_44_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input76_I pcpi_rs2[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2387__A1 _0454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1898__B1 _1350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_55_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_4_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_50_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2378__A1 _0519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2550__A1 _0586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1705_ picorv32_pcpi_div_inst_0.quotient\[24\] _1199_ _1200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_45_116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2823_ _0912_ _0922_ _0924_ _0195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2754_ picorv32_pcpi_div_inst_0.divisor\[47\] _0853_ _0866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_18_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1636_ picorv32_pcpi_div_inst_0.quotient\[17\] _1138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1567_ picorv32_pcpi_div_inst_0.dividend\[10\] _1064_ _0967_ _1075_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2685_ _0802_ _0804_ _0805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2119_ picorv32_pcpi_div_inst_0.quotient_msk\[20\] _0323_ picorv32_pcpi_div_inst_0.quotient\[20\]
+ _0327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1498_ picorv32_pcpi_div_inst_0.quotient\[5\] _1012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2844__A2 _0424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_1_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_52_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2910__CLK clknet_4_11_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_9_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2220__B1 _0384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1574__A2 _1080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2470_ net29 _0613_ _0614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__2933__CLK clknet_4_15_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3022_ _0174_ clknet_4_1_0_clk picorv32_pcpi_div_inst_0.divisor\[36\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_58_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2211__B1 _0378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2668_ _0789_ _0756_ _0790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2737_ _0846_ _0850_ _0851_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2806_ _0598_ _0909_ _0910_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_67_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1619_ _1121_ _1122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_input39_I pcpi_rs1[28] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2599_ net66 net65 _0730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_49_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_12_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2956__CLK clknet_4_13_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_20_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2808__A2 _0747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_4_5_0_clk_I clknet_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1970_ picorv32_pcpi_div_inst_0.divisor\[15\] picorv32_pcpi_div_inst_0.dividend\[15\]
+ _1422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2522_ _0414_ _0654_ _0657_ _0660_ _0661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_11_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2453_ _0404_ _0598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_2384_ _0205_ _0535_ _0536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_11_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput2 pcpi_insn[0] net2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_39_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_36_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3005_ _0159_ clknet_4_10_0_clk picorv32_pcpi_div_inst_0.dividend\[25\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_61_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_34_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2979__CLK clknet_4_1_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_25_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1884_ _1345_ _0059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_28_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1953_ _1398_ _1401_ _1404_ _1405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_22_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2505_ _1391_ _0645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_11_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2367_ _0418_ _0520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2436_ _0581_ _0582_ _0583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2298_ net19 net30 net41 net44 _0457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XPHY_EDGE_ROW_22_Left_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_66_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2213__I _1315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3007__CLK clknet_4_3_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_22_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1695__A1 _1037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_45_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1998__A2 _1095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2152_ picorv32_pcpi_div_inst_0.quotient_msk\[1\] _1360_ _0346_ picorv32_pcpi_div_inst_0.quotient_msk\[2\]
+ _0347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2221_ _0389_ _0128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_17_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2083_ _0298_ _0304_ _0075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1989__A2 _1074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1610__A1 _1100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1936_ _1341_ _1172_ _1383_ _1388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_33_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1867_ _1316_ _1334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_8_425 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2985_ _0139_ clknet_4_2_0_clk picorv32_pcpi_div_inst_0.dividend\[5\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_16_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1798_ picorv32_pcpi_div_inst_0.quotient_msk\[26\] picorv32_pcpi_div_inst_0.quotient_msk\[25\]
+ picorv32_pcpi_div_inst_0.quotient_msk\[24\] picorv32_pcpi_div_inst_0.quotient_msk\[23\]
+ _1282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XANTENNA__1913__A2 _1364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput82 pcpi_rs2[9] net82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput71 pcpi_rs2[28] net71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput60 pcpi_rs2[18] net60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_12_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_4_13_0_clk_I clknet_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1677__A1 _1037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input21_I pcpi_rs1[11] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2419_ _0562_ _0563_ _0567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_output108_I net108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2208__I _0362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_50_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_7_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2118__I _0313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_58_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1721_ _1201_ picorv32_pcpi_div_inst_0.dividend\[24\] _1193_ _1214_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_38_361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2770_ _0861_ _0727_ _0840_ _0879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1583_ picorv32_pcpi_div_inst_0.quotient\[12\] _1089_ _1090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1652_ _1150_ _1151_ _1152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_0_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2204_ picorv32_pcpi_div_inst_0.quotient_msk\[21\] _0375_ _0378_ picorv32_pcpi_div_inst_0.quotient_msk\[22\]
+ _0379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2135_ picorv32_pcpi_div_inst_0.quotient_msk\[26\] _0336_ _1209_ _0337_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_28_73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2066_ _1367_ _0293_ _0069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1867__I _1316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2968_ _0122_ clknet_4_15_0_clk picorv32_pcpi_div_inst_0.quotient_msk\[21\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_63_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1919_ _1369_ _1370_ _1371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input69_I pcpi_rs2[26] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2899_ _0053_ clknet_4_9_0_clk picorv32_pcpi_div_inst_0.divisor\[15\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_12_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_55_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_4_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_39_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1726__B _1202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1461__B _0977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2862__CLK clknet_4_13_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1704_ _0977_ _1198_ _1199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_41_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2684_ _0803_ _0804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2822_ picorv32_pcpi_div_inst_0.divisor\[57\] _0923_ _0924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2753_ picorv32_pcpi_div_inst_0.divisor\[48\] _0855_ _0864_ _0865_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1497_ _0999_ _0998_ _1011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_1635_ _1134_ _1136_ _1137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_39_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1566_ picorv32_pcpi_div_inst_0.dividend\[11\] _1074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_2
X_2118_ _0313_ _0326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_55_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2049_ picorv32_pcpi_div_inst_0.divisor\[55\] picorv32_pcpi_div_inst_0.divisor\[54\]
+ picorv32_pcpi_div_inst_0.divisor\[53\] picorv32_pcpi_div_inst_0.divisor\[52\] _0277_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XTAP_TAPCELL_ROW_52_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2885__CLK clknet_4_3_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_15_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2220__A1 picorv32_pcpi_div_inst_0.quotient_msk\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_4_1_0_clk_I clknet_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_66_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3021_ _0173_ clknet_4_4_0_clk picorv32_pcpi_div_inst_0.divisor\[35\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2287__A1 net44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2805_ net67 _0908_ _0909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_41_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2667_ _0720_ _0721_ _0789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_1618_ picorv32_pcpi_div_inst_0.dividend\[16\] _1121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__3040__CLK clknet_4_0_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2736_ net56 _0849_ _0850_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_5_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1549_ picorv32_pcpi_div_inst_0.dividend\[9\] _1059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2598_ net64 net63 _0729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_49_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2450__A1 _0469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_12_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_20_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_28_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2521_ _0658_ _0659_ _0660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_23_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_11_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2900__CLK clknet_4_9_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2452_ _0597_ _0151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2383_ _1322_ _1079_ _0529_ _0535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_EDGE_ROW_18_Right_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xinput3 pcpi_insn[12] net3 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3004_ _0158_ clknet_4_12_0_clk picorv32_pcpi_div_inst_0.dividend\[24\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_27_Right_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_34_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_42_495 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_36_Right_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_input51_I pcpi_rs2[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2719_ net54 _0834_ _0835_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XPHY_EDGE_ROW_45_Right_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_37_245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_25_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2423__A1 net24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2923__CLK clknet_4_13_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_54_Right_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_52_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_63_Right_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_48_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1883_ _1341_ _1343_ _1340_ _1344_ _1345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1952_ _1402_ _1403_ _1404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2504_ _1177_ _0402_ _0644_ _0156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_24_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2435_ _0579_ _0460_ _0578_ _0582_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_11_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2297_ _0455_ _0456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2366_ _0518_ _0519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__1456__A2 _0973_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2946__CLK clknet_4_4_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_22_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2405__A1 _0439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2151_ _1349_ _0346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2082_ picorv32_pcpi_div_inst_0.quotient_msk\[6\] _0302_ picorv32_pcpi_div_inst_0.quotient\[6\]
+ _0304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2220_ picorv32_pcpi_div_inst_0.quotient_msk\[27\] _0388_ _0384_ picorv32_pcpi_div_inst_0.quotient_msk\[28\]
+ _0389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__2969__CLK clknet_4_15_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2635__A1 _0747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2984_ _0138_ clknet_4_2_0_clk picorv32_pcpi_div_inst_0.dividend\[4\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1797_ picorv32_pcpi_div_inst_0.quotient_msk\[22\] picorv32_pcpi_div_inst_0.quotient_msk\[21\]
+ picorv32_pcpi_div_inst_0.quotient_msk\[20\] picorv32_pcpi_div_inst_0.quotient_msk\[19\]
+ _1281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_56_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1610__A2 _1102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1935_ _1341_ _1172_ _1387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_3_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput50 pcpi_rs1[9] net50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput61 pcpi_rs2[19] net61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_12_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_16_215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1866_ _1333_ _0053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xinput72 pcpi_rs2[29] net72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput83 resetn net83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2418_ _0454_ _0565_ _0566_ _0148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_12_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input14_I pcpi_insn[31] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2349_ _0502_ _0503_ _0406_ _0504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_66_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_0_Right_0 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_62_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1601__A2 _1031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_50_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_54_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_7_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_58_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2134__I _0329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_41_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1651_ _1142_ _1144_ _1135_ _1151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1720_ picorv32_pcpi_div_inst_0.dividend\[26\] _1213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_13_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1582_ _1086_ _1088_ _1089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_28_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2203_ _0358_ _0378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2134_ _0329_ _0336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_input6_I pcpi_insn[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2065_ picorv32_pcpi_div_inst_0.quotient_msk\[0\] _0292_ _0953_ _0293_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2967_ _0121_ clknet_4_15_0_clk picorv32_pcpi_div_inst_0.quotient_msk\[20\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_63_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1918_ picorv32_pcpi_div_inst_0.divisor\[18\] picorv32_pcpi_div_inst_0.dividend\[18\]
+ _1370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_4_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1849_ _1318_ _1321_ _1317_ _1322_ _1323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_8_289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2898_ _0052_ clknet_4_9_0_clk picorv32_pcpi_div_inst_0.divisor\[14\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_67_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_55_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2219__I _0387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_4_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2129__I _0313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1813__A2 _1291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2821_ _0394_ _0923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1703_ picorv32_pcpi_div_inst_0.quotient\[22\] picorv32_pcpi_div_inst_0.quotient\[23\]
+ _1183_ _1198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_1634_ _1122_ _1124_ _1135_ _1136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2683_ _0737_ _0416_ _0803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2752_ _0846_ _0863_ _0864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_14_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1565_ picorv32_pcpi_div_inst_0.quotient\[11\] _1072_ _1073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1496_ _1000_ _1003_ _1009_ _1010_ _0026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_39_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2117_ _0320_ _0325_ _0088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_55_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1501__A1 _0947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2048_ picorv32_pcpi_div_inst_0.divisor\[51\] picorv32_pcpi_div_inst_0.divisor\[50\]
+ picorv32_pcpi_div_inst_0.divisor\[49\] picorv32_pcpi_div_inst_0.divisor\[48\] _0276_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_64_427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1568__A1 _1074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input81_I pcpi_rs2[8] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_15_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_41_Left_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_23_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_50_Left_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1731__A1 _1116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_66_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3020_ _0172_ clknet_4_4_0_clk picorv32_pcpi_div_inst_0.divisor\[34\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_61_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1647__B _0973_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2804_ _0731_ _0812_ _0908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1617_ _1112_ _1115_ _1120_ _0006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_41_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2666_ _0769_ _0787_ _0788_ _0174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_1_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2597_ net61 _0726_ _0727_ _0728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_2735_ _0847_ _0848_ _0849_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1548_ _1056_ _1057_ _1058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1479_ _0992_ _0994_ _0985_ _0995_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_37_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2232__I _0395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_20_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1713__A1 _1153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_390 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2852__CLK clknet_4_12_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_28_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1795__A4 picorv32_pcpi_div_inst_0.quotient_msk\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1467__B _0983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2520_ _0655_ _0656_ _0659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2451_ _1134_ _0596_ _0574_ _0597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__1704__A1 _0977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput4 pcpi_insn[13] net4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3003_ _0157_ clknet_4_10_0_clk picorv32_pcpi_div_inst_0.dividend\[23\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2382_ net21 _0533_ _0534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_36_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2718_ _0833_ _0756_ _0834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_6_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2875__CLK clknet_4_14_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2649_ picorv32_pcpi_div_inst_0.divisor\[34\] _0751_ _0774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1891__I _1349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input44_I pcpi_rs1[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_25_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3030__CLK clknet_4_1_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1882_ picorv32_pcpi_div_inst_0.divisor\[22\] _1344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_24_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1951_ picorv32_pcpi_div_inst_0.divisor\[3\] picorv32_pcpi_div_inst_0.dividend\[3\]
+ _1403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_2503_ _0305_ _0638_ _0643_ _0644_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_3_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2434_ _0406_ _0581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__2898__CLK clknet_4_9_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2365_ _1364_ _0518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2296_ _0418_ _0455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_63_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_47_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_22_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2081_ _0298_ _0303_ _0074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2150_ _0345_ _0101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2332__A1 _0454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1934_ _1376_ _1381_ _1382_ _1385_ _1386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_2983_ _0137_ clknet_4_3_0_clk picorv32_pcpi_div_inst_0.dividend\[3\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_8_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1796_ picorv32_pcpi_div_inst_0.running _1278_ _1279_ _1280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
Xinput62 pcpi_rs2[1] net62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput51 pcpi_rs2[0] net51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput73 pcpi_rs2[2] net73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput40 pcpi_rs1[29] net40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_3_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1865_ picorv32_pcpi_div_inst_0.divisor\[15\] _1330_ _1327_ picorv32_pcpi_div_inst_0.divisor\[16\]
+ _1333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__2571__A1 net40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2417_ _1100_ _0292_ _0566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2348_ _0208_ _0503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2913__CLK clknet_4_4_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2279_ _0437_ _1402_ _0440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_50_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1437__I0 _0952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2240__I net19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_58_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_7_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_41_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2617__A2 _0297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1581_ _1051_ _1031_ _1087_ _1088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_1650_ picorv32_pcpi_div_inst_0.dividend\[19\] _1150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2202_ _0377_ _0121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2936__CLK clknet_4_14_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2553__A1 net38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2133_ _0333_ _0335_ _0094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2064_ _0291_ _0292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_2966_ _0120_ clknet_4_15_0_clk picorv32_pcpi_div_inst_0.quotient_msk\[19\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_48_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1917_ picorv32_pcpi_div_inst_0.divisor\[19\] picorv32_pcpi_div_inst_0.dividend\[19\]
+ _1369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_2897_ _0051_ clknet_4_9_0_clk picorv32_pcpi_div_inst_0.divisor\[13\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1779_ net15 _1256_ _1258_ _1265_ _1266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_44_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1848_ picorv32_pcpi_div_inst_0.divisor\[10\] _1322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_12_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_67_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_55_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2235__I _0398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2959__CLK clknet_4_13_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2535__A1 net37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2820_ picorv32_pcpi_div_inst_0.divisor\[58\] _0890_ _0921_ _0922_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2751_ net58 _0862_ _0863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_18_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1564_ _0993_ _1071_ _1072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1633_ _1020_ _1135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1702_ _1196_ _1197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_30_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2682_ _0722_ _0802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1495_ _0955_ _1010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_39_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2116_ picorv32_pcpi_div_inst_0.quotient_msk\[19\] _0323_ picorv32_pcpi_div_inst_0.quotient\[19\]
+ _0325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2047_ _1362_ _1249_ _0274_ _0275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2949_ _0103_ clknet_4_5_0_clk picorv32_pcpi_div_inst_0.quotient_msk\[2\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2214__B1 _0384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1894__I _1297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input74_I pcpi_rs2[30] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2508__A1 net33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_66_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1753__B _0955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2734_ _0755_ _0848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2803_ picorv32_pcpi_div_inst_0.divisor\[55\] _0907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1547_ _1050_ _1052_ _1021_ _1057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1616_ _1116_ _1119_ _1120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2665_ picorv32_pcpi_div_inst_0.divisor\[36\] _0780_ _0788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_22_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2596_ net59 net58 net60 _0727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_1478_ picorv32_pcpi_div_inst_0.dividend\[2\] _0961_ _0951_ _0993_ _0994_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_49_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_32_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_20_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_28_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_11_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2450_ _0469_ _0590_ _0595_ _0596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_23_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2381_ net20 _0521_ _0520_ _0533_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xinput5 pcpi_insn[14] net5 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3002_ _0156_ clknet_4_10_0_clk picorv32_pcpi_div_inst_0.dividend\[22\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_52_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2333__I _0432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2717_ _0802_ _0723_ _0833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_65_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2648_ picorv32_pcpi_div_inst_0.divisor\[35\] _0753_ _0772_ _0773_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2579_ _0274_ _0711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA_input37_I pcpi_rs1[26] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2489__B _0449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_25_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1478__B _0993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1950_ picorv32_pcpi_div_inst_0.divisor\[2\] picorv32_pcpi_div_inst_0.dividend\[2\]
+ _1402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_22_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2502_ net33 _0640_ _0642_ _0643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1881_ _1320_ _1343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_24_431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1689__B2 _1169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2433_ _0456_ _0578_ _0579_ _0580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2364_ _1060_ _0508_ _0517_ _0143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_66_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2295_ _0401_ _0454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__2063__I _0290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1916__A2 _1249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2992__CLK clknet_4_8_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2238__I _0329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1907__A2 _1360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_4_9_0_clk clknet_0_clk clknet_4_9_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_2080_ picorv32_pcpi_div_inst_0.quotient_msk\[5\] _0302_ _1012_ _0303_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_56_353 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2865__CLK clknet_4_14_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_44_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1933_ _1383_ _1384_ _1385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XPHY_EDGE_ROW_26_Left_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2982_ _0136_ clknet_4_8_0_clk picorv32_pcpi_div_inst_0.dividend\[2\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_16_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1795_ picorv32_pcpi_div_inst_0.quotient_msk\[30\] picorv32_pcpi_div_inst_0.quotient_msk\[29\]
+ picorv32_pcpi_div_inst_0.quotient_msk\[28\] picorv32_pcpi_div_inst_0.quotient_msk\[27\]
+ _1279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
Xinput52 pcpi_rs2[10] net52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput74 pcpi_rs2[30] net74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput30 pcpi_rs1[1] net30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput41 pcpi_rs1[2] net41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_12_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xinput63 pcpi_rs2[20] net63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1864_ _1332_ _0052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_58_73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2278_ _0423_ _0439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2416_ _0559_ _0561_ _0564_ _0469_ _0565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XPHY_EDGE_ROW_10_Left_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2347_ _0501_ _0502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_50_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3020__CLK clknet_4_4_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2314__A2 _1005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_58_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_7_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_41_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2888__CLK clknet_4_2_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1580_ picorv32_pcpi_div_inst_0.quotient\[8\] picorv32_pcpi_div_inst_0.quotient\[9\]
+ picorv32_pcpi_div_inst_0.quotient\[10\] picorv32_pcpi_div_inst_0.quotient\[11\]
+ _1087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_53_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2201_ picorv32_pcpi_div_inst_0.quotient_msk\[20\] _0375_ _0372_ picorv32_pcpi_div_inst_0.quotient_msk\[21\]
+ _0377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2132_ picorv32_pcpi_div_inst_0.quotient_msk\[25\] _0330_ picorv32_pcpi_div_inst_0.quotient\[25\]
+ _0335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_28_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2063_ _0290_ _0291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2965_ _0119_ clknet_4_15_0_clk picorv32_pcpi_div_inst_0.quotient_msk\[18\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_56_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1916_ _1362_ _1249_ _1368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3043__CLK clknet_4_2_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2896_ _0050_ clknet_4_9_0_clk picorv32_pcpi_div_inst_0.divisor\[12\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1847_ _1320_ _1321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1778_ _1259_ _1261_ _1264_ _1265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XTAP_TAPCELL_ROW_63_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2471__A1 _0581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2426__I _0430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1701_ _1192_ _1194_ _0965_ _1196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2681_ picorv32_pcpi_div_inst_0.divisor\[39\] _0801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_5_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2750_ _0861_ _0848_ _0862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2161__I _1349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1563_ picorv32_pcpi_div_inst_0.quotient\[8\] _1056_ _1067_ _1052_ _1071_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_0_41_326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1494_ _1005_ _1008_ _1009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__2903__CLK clknet_4_10_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1632_ picorv32_pcpi_div_inst_0.dividend\[17\] _1134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2115_ _0320_ _0324_ _0087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2046_ _0270_ picorv32_pcpi_div_inst_0.dividend\[30\] _0274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2462__A1 _0407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2948_ _0102_ clknet_4_5_0_clk picorv32_pcpi_div_inst_0.quotient_msk\[1\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_57_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2879_ _0020_ clknet_4_12_0_clk net104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_32_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2765__A2 _0581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input67_I pcpi_rs2[24] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_13_Left_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2926__CLK clknet_4_13_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_66_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2156__I _1352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2444__A1 net27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2664_ picorv32_pcpi_div_inst_0.divisor\[37\] _0783_ _0786_ _0787_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_26_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2802_ _0867_ _0905_ _0906_ _0192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2733_ _0722_ _0723_ _0724_ _0847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_1546_ picorv32_pcpi_div_inst_0.quotient\[9\] _1056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1615_ picorv32_pcpi_div_inst_0.quotient\[15\] _1118_ _1119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1477_ _0958_ _0993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_1_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2595_ _0722_ _0723_ _0724_ _0725_ _0726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_0_49_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_45_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2029_ _0253_ picorv32_pcpi_div_inst_0.dividend\[25\] _0257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_9_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_20_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_28_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_11_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2380_ _1079_ _0508_ _0532_ _0144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xinput6 pcpi_insn[1] net6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3001_ _0155_ clknet_4_11_0_clk picorv32_pcpi_div_inst_0.dividend\[21\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_36_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2417__A1 _1100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2647_ _0519_ _0771_ _0772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2716_ _0795_ _0831_ _0832_ _0180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2578_ _0710_ _0164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1529_ picorv32_pcpi_div_inst_0.dividend\[8\] _1040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_10_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_25_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2408__A1 _1095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_14_Right_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_23_Right_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_20_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2647__A1 _0519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1759__B _1202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_38_Left_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_32_Right_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1880_ _1342_ _0058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_22_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2434__I _0406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_47_Left_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2501_ net33 _0640_ _0641_ _0642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_24_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_41_Right_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_39_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2432_ net26 _0579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2294_ _0992_ _0429_ _0453_ _0137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2363_ _0509_ _0516_ _0517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_56_Left_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_50_Right_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_65_Left_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_62_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_2_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_44_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1932_ picorv32_pcpi_div_inst_0.divisor\[20\] _1158_ _1384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xinput31 pcpi_rs1[20] net31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2981_ _0135_ clknet_4_3_0_clk picorv32_pcpi_div_inst_0.dividend\[1\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xinput20 pcpi_rs1[10] net20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1863_ picorv32_pcpi_div_inst_0.divisor\[14\] _1330_ _1327_ picorv32_pcpi_div_inst_0.divisor\[15\]
+ _1332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1794_ picorv32_pcpi_div_inst_0.quotient_msk\[31\] _1278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xinput42 pcpi_rs1[30] net42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput75 pcpi_rs2[31] net75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput53 pcpi_rs2[11] net53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_12_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xinput64 pcpi_rs2[21] net64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2415_ _0562_ _0563_ _0564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2277_ _0437_ _1402_ _0438_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2346_ _1413_ _1421_ _0501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_66_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_47_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_50_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1598__A1 _0977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_58_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_41_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2200_ _0376_ _0120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2131_ _0333_ _0334_ _0093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2062_ _0289_ _0290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__1513__A1 _1016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2964_ _0118_ clknet_4_15_0_clk picorv32_pcpi_div_inst_0.quotient_msk\[17\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_44_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2982__CLK clknet_4_8_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1915_ _1366_ _1367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1777_ net18 _1263_ _1264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_29_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1846_ _1290_ _1320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2895_ _0049_ clknet_4_8_0_clk picorv32_pcpi_div_inst_0.divisor\[11\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_40_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_4_Right_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_input12_I pcpi_insn[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2329_ _0484_ _0485_ _0407_ _0486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xclkbuf_4_8_0_clk clknet_0_clk clknet_4_8_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_62_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_390 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2855__CLK clknet_4_6_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1631_ _1126_ _1128_ _1133_ _1055_ _0007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1700_ _1192_ _1194_ _1195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_41_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2680_ _0795_ _0799_ _0800_ _0176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_26_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1562_ _0976_ _1066_ _1070_ _0001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1493_ _1006_ _1007_ _1008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_39_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2114_ picorv32_pcpi_div_inst_0.quotient_msk\[18\] _0323_ picorv32_pcpi_div_inst_0.quotient\[18\]
+ _0324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_55_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input4_I pcpi_insn[13] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2045_ _0264_ _0268_ _0272_ _0273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__3010__CLK clknet_4_1_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_460 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2947_ _0101_ clknet_4_5_0_clk picorv32_pcpi_div_inst_0.quotient_msk\[0\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_29_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2878__CLK clknet_4_12_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2878_ _0019_ clknet_4_12_0_clk net103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_4_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_9_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1829_ _1307_ _0042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_17_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_66_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3033__CLK clknet_4_0_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1798__A4 picorv32_pcpi_div_inst_0.quotient_msk\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2801_ picorv32_pcpi_div_inst_0.divisor\[54\] _0883_ _0906_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_14_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1614_ _1117_ _1107_ _1030_ _1118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2663_ _0775_ _0785_ _0786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2732_ _0518_ _0846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2594_ net57 net56 _0725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1545_ _1045_ _1049_ _1054_ _1055_ _0030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1476_ _0991_ _0992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_5_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2028_ _0255_ picorv32_pcpi_div_inst_0.dividend\[24\] _0256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_64_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_20_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_28_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_11_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput7 pcpi_insn[25] net7 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_52_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3000_ _0154_ clknet_4_10_0_clk picorv32_pcpi_div_inst_0.dividend\[20\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2417__A2 _0292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2646_ net76 _0770_ _0771_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2577_ _1239_ _0709_ _0401_ _0710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2715_ picorv32_pcpi_div_inst_0.divisor\[42\] _0819_ _0832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_6_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2353__A1 _1041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1690__B _1135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1459_ _0963_ _0970_ _0975_ _0976_ _0011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_1528_ _1029_ _1033_ _1036_ _1039_ _0029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_45_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_33_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2939__CLK clknet_4_12_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2583__A1 net40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2431_ _0577_ _0578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_24_433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2500_ _0412_ _0641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_11_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_39_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2293_ _0431_ _0452_ _0453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_2_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2362_ _0489_ _0511_ _0515_ _0516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_59_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_47_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_42_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2629_ _0755_ _0756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_input42_I pcpi_rs1[30] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2565__A1 net38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2270__I _0430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_44_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2980_ _0134_ clknet_4_3_0_clk picorv32_pcpi_div_inst_0.dividend\[0\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1793_ _1274_ _1275_ _1276_ _1277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
Xinput10 pcpi_insn[28] net10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_56_355 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1931_ picorv32_pcpi_div_inst_0.divisor\[20\] _1158_ _1383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
Xinput32 pcpi_rs1[21] net32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput43 pcpi_rs1[31] net43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput21 pcpi_rs1[11] net21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_12_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1862_ _1331_ _0051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xinput54 pcpi_rs2[12] net54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_58_75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput76 pcpi_rs2[3] net76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput65 pcpi_rs2[22] net65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2414_ _0203_ _0544_ _0227_ _0563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2276_ _1398_ _1401_ _0437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2345_ net49 _0499_ _0500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_59_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1598__A2 _1102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2355__I _0430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2265__I _0329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_41_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2130_ picorv32_pcpi_div_inst_0.quotient_msk\[24\] _0330_ picorv32_pcpi_div_inst_0.quotient\[24\]
+ _0334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2061_ _0287_ _0288_ _1288_ _0289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2963_ _0117_ clknet_4_15_0_clk picorv32_pcpi_div_inst_0.quotient_msk\[16\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_60_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1914_ _1365_ _1366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2226__B1 _1294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_388 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1776_ _1262_ net16 net17 _1263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__2529__A1 net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2894_ _0048_ clknet_4_8_0_clk picorv32_pcpi_div_inst_0.divisor\[10\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1845_ _1319_ _0046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_8_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1963__B _1025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2328_ _0481_ _0482_ _0485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_12_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2259_ net30 _0420_ _0421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_62_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_3_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1630_ _1129_ _1132_ _1133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_34_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1561_ _1067_ _1068_ _1069_ _1070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_39_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_39_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1492_ picorv32_pcpi_div_inst_0.dividend\[3\] picorv32_pcpi_div_inst_0.dividend\[2\]
+ picorv32_pcpi_div_inst_0.dividend\[1\] picorv32_pcpi_div_inst_0.dividend\[0\] _1007_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or4_1
X_2113_ _0301_ _0323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_55_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_52_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2044_ _0269_ _0271_ _0272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2877_ _0018_ clknet_4_12_0_clk net102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2946_ _0100_ clknet_4_4_0_clk picorv32_pcpi_div_inst_0.quotient\[31\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_29_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1759_ picorv32_pcpi_div_inst_0.quotient\[30\] _1244_ _1202_ _1247_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_40_350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_9_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1828_ _1304_ _1299_ _1306_ picorv32_pcpi_div_inst_0.divisor\[5\] _1307_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__1661__A1 _1113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2972__CLK clknet_4_13_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2453__I _0404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2800_ picorv32_pcpi_div_inst_0.divisor\[55\] _0890_ _0904_ _0905_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_14_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2731_ _0839_ _0844_ _0845_ _0182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1613_ _1108_ _1117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1544_ _1048_ _1055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_41_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2662_ net78 _0784_ _0785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2593_ net55 net54 _0724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_1_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_4_7_0_clk clknet_0_clk clknet_4_7_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_1475_ picorv32_pcpi_div_inst_0.dividend\[3\] _0991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_5_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1643__A1 _1134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2027_ picorv32_pcpi_div_inst_0.divisor\[24\] _0255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_9_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2929_ _0083_ clknet_4_14_0_clk picorv32_pcpi_div_inst_0.quotient\[14\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_45_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input72_I pcpi_rs2[29] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_20_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_394 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2995__CLK clknet_4_9_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_28_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3000__CLK clknet_4_10_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_11_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_11_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput8 pcpi_insn[26] net8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2868__CLK clknet_4_11_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2714_ picorv32_pcpi_div_inst_0.divisor\[43\] _0826_ _0830_ _0831_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_6_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1527_ _1037_ _1038_ _1039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2645_ net62 _0748_ net73 _0755_ _0770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_2576_ _0444_ _0705_ _0707_ _0708_ _0709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_22_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1458_ _0966_ _0976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__1616__A1 _1116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3023__CLK clknet_4_1_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_423 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2280__A1 _0439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2583__A2 net42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2430_ net22 net23 _0540_ _0576_ _0577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or4_1
X_2361_ _0439_ _0514_ _0515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2178__I _0362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_39_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2292_ _0444_ _0447_ _0451_ _0452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_59_320 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_47_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3046__CLK clknet_4_3_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_6_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_6_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2559_ _0444_ _0689_ _0691_ _0693_ _0694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA_input35_I pcpi_rs1[24] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2628_ _0754_ _0755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_33_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2565__A2 net39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_17_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_44_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1930_ picorv32_pcpi_div_inst_0.divisor\[21\] _1172_ _1382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1792_ picorv32_pcpi_div_inst_0.quotient_msk\[10\] picorv32_pcpi_div_inst_0.quotient_msk\[9\]
+ picorv32_pcpi_div_inst_0.quotient_msk\[8\] picorv32_pcpi_div_inst_0.quotient_msk\[7\]
+ _1276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
Xinput11 pcpi_insn[29] net11 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput33 pcpi_rs1[22] net33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2906__CLK clknet_4_10_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput77 pcpi_rs2[4] net77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_24_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput44 pcpi_rs1[3] net44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput22 pcpi_rs1[12] net22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput66 pcpi_rs2[23] net66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1861_ _1328_ _1330_ _1327_ picorv32_pcpi_div_inst_0.divisor\[14\] _1331_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_16_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput55 pcpi_rs2[13] net55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_58_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2344_ _0419_ _0498_ _0499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2413_ _1423_ _0562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2275_ net41 _0435_ _0436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_59_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_57_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2929__CLK clknet_4_14_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2483__A1 _0407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_41_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2060_ _1292_ _1286_ _0288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_44_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_6_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2962_ _0116_ clknet_4_15_0_clk picorv32_pcpi_div_inst_0.quotient_msk\[15\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_56_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1913_ _1271_ _1364_ _1365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_29_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2893_ _0047_ clknet_4_8_0_clk picorv32_pcpi_div_inst_0.divisor\[9\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_52_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1775_ net12 _1262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_4_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1844_ _1313_ _1308_ _1317_ _1318_ _1319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_8_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2258_ _0403_ _0419_ _0420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2327_ _1309_ _1024_ _0484_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2189_ picorv32_pcpi_div_inst_0.quotient_msk\[15\] _0369_ _0366_ picorv32_pcpi_div_inst_0.quotient_msk\[16\]
+ _0370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_62_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_47_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1560_ _1067_ _1068_ _0946_ _1069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2112_ _0320_ _0322_ _0086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1491_ _0972_ _1006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_39_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_52_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2043_ _0270_ picorv32_pcpi_div_inst_0.dividend\[30\] _0271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_17_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_60_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2876_ _0017_ clknet_4_12_0_clk net101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2945_ _0099_ clknet_4_4_0_clk picorv32_pcpi_div_inst_0.quotient\[30\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_32_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1827_ _1294_ _1306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1689_ _1179_ _1181_ _1185_ _1169_ _0014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1758_ _1241_ _1242_ _1246_ _1169_ _0023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_40_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_9_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1903__I _1349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2429__A1 net24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2661_ net77 _0720_ _0762_ _0784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_26_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_14_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2730_ picorv32_pcpi_div_inst_0.divisor\[44\] _0819_ _0845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1474_ picorv32_pcpi_div_inst_0.quotient\[3\] _0989_ _0990_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1543_ _1050_ _1053_ _1054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1612_ _0946_ _1116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2592_ net82 net81 net53 net52 _0723_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_1_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_65_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2026_ _0253_ _1201_ _0254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2644__I _0768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2928_ _0082_ clknet_4_13_0_clk picorv32_pcpi_div_inst_0.quotient\[13\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2859_ _0030_ clknet_4_12_0_clk net114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_32_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_input65_I pcpi_rs2[22] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_17_Left_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_36_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_11_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput9 pcpi_insn[27] net9 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_52_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2644_ _0768_ _0769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2713_ _0811_ _0829_ _0830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_14_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1457_ _0971_ _0974_ _0975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1526_ _1035_ _0968_ _1034_ _1038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_2575_ _0706_ _0271_ _0641_ _0708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_22_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2962__CLK clknet_4_15_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2009_ _0236_ _1391_ _0237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_9_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2041__A2 _1249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1552__A1 _1060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_4_6_0_clk clknet_0_clk clknet_4_6_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_22_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2291_ _0448_ _1403_ _0450_ _0451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2360_ _0207_ _0513_ _0514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_63_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_39_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_10_Right_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_59_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_47_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2985__CLK clknet_4_2_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput110 net110 pcpi_div_rd[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_2627_ net75 _0415_ _0754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_12_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1509_ _1012_ _1011_ _1021_ _1022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1534__A1 _1041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2558_ _0658_ _0692_ _0693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_34_Left_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2489_ _1382_ _0630_ _0449_ _0631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_input28_I pcpi_rs1[18] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_43_Left_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_53_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_52_Left_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2858__CLK clknet_4_12_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2228__B _0297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_44_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2742__I _0782_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1860_ _1320_ _1330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1791_ picorv32_pcpi_div_inst_0.quotient_msk\[6\] picorv32_pcpi_div_inst_0.quotient_msk\[5\]
+ picorv32_pcpi_div_inst_0.quotient_msk\[4\] picorv32_pcpi_div_inst_0.quotient_msk\[3\]
+ _1275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
Xinput12 pcpi_insn[2] net12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1764__A1 _1249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput34 pcpi_rs1[23] net34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput78 pcpi_rs2[5] net78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_24_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput23 pcpi_rs1[13] net23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput45 pcpi_rs1[4] net45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_12_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput67 pcpi_rs2[24] net67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput56 pcpi_rs2[14] net56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2274_ _0403_ net30 _0434_ _0435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2412_ _0459_ _0560_ _0561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2343_ net47 net48 _0478_ _0498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XANTENNA__3013__CLK clknet_4_4_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1989_ _1324_ _1074_ _1079_ _1322_ _0217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__1522__A4 _1007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_41_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_316 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1906__I _1352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3036__CLK clknet_4_0_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_5_Left_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_6_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2961_ _0115_ clknet_4_15_0_clk picorv32_pcpi_div_inst_0.quotient_msk\[14\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_60_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1912_ _1273_ _1364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_44_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1843_ picorv32_pcpi_div_inst_0.divisor\[9\] _1318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2892_ _0046_ clknet_4_8_0_clk picorv32_pcpi_div_inst_0.divisor\[8\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_17_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1774_ net8 _1260_ net10 net9 _1261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XANTENNA__1816__I _1297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_12_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2257_ _0418_ _0419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2326_ _0481_ _0482_ _1407_ _0483_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_18_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2188_ _0362_ _0369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_55_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_31_Left_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_14_27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1719__A1 _0947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1490_ _1004_ _1005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2111_ picorv32_pcpi_div_inst_0.quotient_msk\[17\] _0317_ _1138_ _0322_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_55_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2042_ picorv32_pcpi_div_inst_0.divisor\[30\] _0270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_52_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_8_Right_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_17_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_60_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2944_ _0098_ clknet_4_5_0_clk picorv32_pcpi_div_inst_0.quotient\[29\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2875_ _0016_ clknet_4_14_0_clk net100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_44_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1826_ _1305_ _0041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_17_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1688_ picorv32_pcpi_div_inst_0.quotient\[22\] _1184_ _1185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1757_ picorv32_pcpi_div_inst_0.quotient\[30\] _1245_ _1246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_40_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_39_Right_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_9_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input10_I pcpi_insn[28] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_0_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2309_ _1005_ _0305_ _0468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_EDGE_ROW_48_Right_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1661__A3 _1102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_57_Right_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_31_385 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_66_Right_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_39_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2429__A2 net25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1611_ _1113_ _1114_ _1115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_41_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2660_ _0782_ _0783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_14_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1473_ picorv32_pcpi_div_inst_0.quotient\[0\] _0971_ picorv32_pcpi_div_inst_0.quotient\[2\]
+ _0973_ _0989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_1542_ _0993_ _1052_ _1053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2591_ net80 net79 _0720_ _0721_ _0722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_5_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_65_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input2_I pcpi_insn[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2025_ picorv32_pcpi_div_inst_0.divisor\[25\] _0253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2927_ _0081_ clknet_4_15_0_clk picorv32_pcpi_div_inst_0.quotient\[12\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_57_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1809_ net117 _1272_ _1292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2858_ _0029_ clknet_4_12_0_clk net113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_31_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2660__I _0782_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2789_ picorv32_pcpi_div_inst_0.divisor\[52\] _0883_ _0896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input58_I pcpi_rs2[16] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2891__CLK clknet_4_2_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_11_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2574_ _0706_ _0271_ _0707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2643_ _1290_ _0768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2712_ net53 _0828_ _0829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_6_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1456_ _0953_ _0973_ _0974_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1525_ _0965_ _1037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2008_ _1344_ _1177_ _0236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_9_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2501__A1 net33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2290_ _0448_ _1403_ _0449_ _0450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_59_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_47_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_42_211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2559__A1 _0444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_30_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput111 net111 pcpi_div_rd[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput100 net100 pcpi_div_rd[24] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_42_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1534__A2 _1042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2557_ _0690_ _0262_ _0692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2626_ _0641_ _0753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1508_ _1020_ _1021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1439_ picorv32_pcpi_div_inst_0.outsign _0957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2488_ _0618_ _0620_ _1383_ _0630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1470__A1 _0981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1790_ picorv32_pcpi_div_inst_0.quotient_msk\[2\] picorv32_pcpi_div_inst_0.quotient_msk\[1\]
+ picorv32_pcpi_div_inst_0.quotient_msk\[0\] _1274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XTAP_TAPCELL_ROW_44_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput13 pcpi_insn[30] net13 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_4_8_0_clk_I clknet_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xinput35 pcpi_rs1[24] net35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput79 pcpi_rs2[6] net79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_24_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2411_ _0460_ _0558_ net24 _0560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_20_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput24 pcpi_rs1[14] net24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput46 pcpi_rs1[5] net46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput68 pcpi_rs2[25] net68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput57 pcpi_rs2[15] net57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2273_ _0417_ _0434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2342_ _1414_ _0429_ _0497_ _0141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_59_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1988_ _1324_ _1074_ _0216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1549__I picorv32_pcpi_div_inst_0.dividend\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2609_ picorv32_pcpi_div_inst_0.instr_div _0739_ _0740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_30_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input40_I pcpi_rs1[29] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_4_5_0_clk clknet_0_clk clknet_4_5_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__2329__B _0407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2960_ _0114_ clknet_4_13_0_clk picorv32_pcpi_div_inst_0.quotient_msk\[13\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_29_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1773_ net7 _1260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_44_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1911_ _1363_ _0068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2891_ _0045_ clknet_4_2_0_clk picorv32_pcpi_div_inst_0.divisor\[7\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1985__A2 _1060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1842_ _1316_ _1317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2187_ _0368_ _0115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_55_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2256_ _0417_ _0418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2325_ _1417_ _1419_ _0482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_18_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_63_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2848__CLK clknet_4_4_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2998__CLK clknet_4_10_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3003__CLK clknet_4_10_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2110_ _0320_ _0321_ _0085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_55_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2041_ picorv32_pcpi_div_inst_0.divisor\[31\] _1249_ _0269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_60_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_464 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2943_ _0097_ clknet_4_5_0_clk picorv32_pcpi_div_inst_0.quotient\[28\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_49_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_17_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1756_ _0977_ _1244_ _1245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2874_ _0015_ clknet_4_11_0_clk net99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_17_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1827__I _1294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1825_ _1302_ _1299_ _1295_ _1304_ _1305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1687_ _1086_ _1183_ _1184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_40_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2308_ _0458_ _0462_ _0465_ _0466_ _0467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2239_ _0401_ _0402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_0_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3026__CLK clknet_4_1_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_50_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_16_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_14_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1610_ _1100_ _1102_ _1021_ _1114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2590_ net78 net77 _0721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_66_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1541_ _1051_ _1031_ _1052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1472_ _0966_ _0988_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_1_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_65_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2024_ _0241_ _1217_ picorv32_pcpi_div_inst_0.dividend\[26\] _0251_ _0252_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_2926_ _0080_ clknet_4_13_0_clk picorv32_pcpi_div_inst_0.quotient\[11\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2857_ _0028_ clknet_4_13_0_clk net112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_45_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1739_ _1217_ picorv32_pcpi_div_inst_0.dividend\[26\] _1214_ _1230_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_40_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_32_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1808_ _1290_ _1291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2788_ picorv32_pcpi_div_inst_0.divisor\[53\] _0890_ _0894_ _0895_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2292__A1 _0444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_11_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_39_250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2909__CLK clknet_4_11_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2283__A1 _0981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2711_ _0802_ _0827_ _0804_ _0828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_6_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1524_ _0997_ _1034_ _1035_ _1036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2642_ _0747_ _0766_ _0767_ _0171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2573_ _0264_ _0268_ _0706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_10_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1455_ _0972_ _0973_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_37_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2007_ _1369_ _1370_ _0234_ _0235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XTAP_TAPCELL_ROW_25_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2909_ _0063_ clknet_4_11_0_clk picorv32_pcpi_div_inst_0.divisor\[25\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_5_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_input70_I pcpi_rs2[27] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_28_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_4_4_0_clk_I clknet_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2756__I _0768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_47_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2881__CLK clknet_4_6_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_30_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput112 net112 pcpi_div_rd[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput101 net101 pcpi_div_rd[25] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_1507_ picorv32_pcpi_div_inst_0.outsign _1020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_42_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2625_ _0747_ _0750_ _0752_ _0169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2556_ _0690_ _0262_ _0691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2487_ net32 _0628_ _0629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_23_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1438_ _0956_ _0000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_38_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3039_ _0191_ clknet_4_2_0_clk picorv32_pcpi_div_inst_0.divisor\[53\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_33_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2486__A1 net31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_44_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput14 pcpi_insn[31] net14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput36 pcpi_rs1[25] net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_24_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2410__A1 net24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput25 pcpi_rs1[15] net25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2410_ net24 _0456_ _0558_ _0559_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_20_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_3_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput69 pcpi_rs2[26] net69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput47 pcpi_rs1[6] net47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput58 pcpi_rs2[16] net58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2341_ _0431_ _0496_ _0497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2272_ _0432_ _0433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_59_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_59_175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2401__A1 net22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1987_ _0212_ _0213_ _0214_ _0215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_15_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_61_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1514__B _0985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2539_ _0658_ _0675_ _0676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input33_I pcpi_rs1[22] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2608_ _0714_ _0737_ _0739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_58_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1682__A2 _0997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1910_ picorv32_pcpi_div_inst_0.divisor\[30\] _1360_ _1358_ _1362_ _1363_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2890_ _0044_ clknet_4_2_0_clk picorv32_pcpi_div_inst_0.divisor\[6\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_52_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1772_ net13 net11 net14 _1259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_1841_ _1315_ _1316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_37_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2324_ _0463_ _1411_ _0481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2186_ picorv32_pcpi_div_inst_0.quotient_msk\[14\] _0363_ _0366_ picorv32_pcpi_div_inst_0.quotient_msk\[15\]
+ _0368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2255_ net43 _0416_ _0417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_63_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_4_12_0_clk_I clknet_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1509__B _1021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_7_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2040_ _0265_ picorv32_pcpi_div_inst_0.dividend\[29\] _0267_ _0268_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_60_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2942_ _0096_ clknet_4_7_0_clk picorv32_pcpi_div_inst_0.quotient\[27\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2873_ _0014_ clknet_4_11_0_clk net98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_44_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_17_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1686_ _1165_ _1182_ _1183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1755_ _1243_ _1244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xclkbuf_4_4_0_clk clknet_0_clk clknet_4_4_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__1591__A1 picorv32_pcpi_div_inst_0.dividend\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1824_ picorv32_pcpi_div_inst_0.divisor\[4\] _1304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2238_ _0329_ _0401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2307_ _0413_ _0466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2965__CLK clknet_4_15_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2169_ picorv32_pcpi_div_inst_0.quotient_msk\[8\] _0355_ _0352_ picorv32_pcpi_div_inst_0.quotient_msk\[9\]
+ _0357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_51_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2674__I _0768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_8_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_14_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1540_ picorv32_pcpi_div_inst_0.quotient\[7\] _1051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_41_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1573__A1 _1074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1471_ _0976_ _0979_ _0987_ _0022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_65_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2023_ picorv32_pcpi_div_inst_0.divisor\[26\] _0251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2988__CLK clknet_4_8_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2925_ _0079_ clknet_4_13_0_clk picorv32_pcpi_div_inst_0.quotient\[10\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2856_ _0027_ clknet_4_6_0_clk net111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1807_ _1289_ _1290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_17_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1564__A1 _0993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1669_ picorv32_pcpi_div_inst_0.quotient\[20\] _1167_ _1168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1738_ _1228_ _1229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_25_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2787_ _0878_ _0893_ _0894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_13_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output102_I net102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1555__A1 picorv32_pcpi_div_inst_0.dividend\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2528__B _0612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2710_ net82 net81 net52 _0827_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_14_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_4_0_0_clk_I clknet_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1454_ picorv32_pcpi_div_inst_0.outsign _0972_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2641_ picorv32_pcpi_div_inst_0.divisor\[33\] _0751_ _0767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2572_ net42 _0704_ _0705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_22_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1523_ picorv32_pcpi_div_inst_0.dividend\[7\] _1035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__3016__CLK clknet_4_3_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_25_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2006_ _0232_ _0233_ _0234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2274__A2 net30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2908_ _0062_ clknet_4_11_0_clk picorv32_pcpi_div_inst_0.divisor\[24\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_33_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_33_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input63_I pcpi_rs2[20] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_468 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2839_ picorv32_pcpi_div_inst_0.divisor\[61\] _0466_ _0937_ _0938_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_51_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_493 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3039__CLK clknet_4_2_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_47_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2624_ _1362_ _0751_ _0752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_30_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_6_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput102 net102 pcpi_div_rd[26] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_1437_ _0952_ _0953_ _0955_ _0956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xoutput113 net113 pcpi_div_rd[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_1506_ _1013_ _1015_ _1019_ _1010_ _0027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_2555_ _0250_ _0260_ _0690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2486_ net31 _0623_ _0520_ _0628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_2_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_10_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2319__I0 _1016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_38_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2247__A2 _0405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3038_ _0190_ clknet_4_0_0_clk picorv32_pcpi_div_inst_0.divisor\[52\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1758__B2 _1169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput15 pcpi_insn[3] net15 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1749__A1 _1116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput37 pcpi_rs1[26] net37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput26 pcpi_rs1[16] net26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput48 pcpi_rs1[7] net48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput59 pcpi_rs2[17] net59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_58_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2271_ _0412_ _0432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_20_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2340_ _0489_ _0492_ _0495_ _0496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_62_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1986_ _1318_ _1060_ _1041_ _1313_ _0214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_2607_ _0714_ _0736_ _0737_ _0738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_23_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2538_ _0244_ _0673_ _0675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2469_ net28 _0604_ _0612_ _0613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_input26_I pcpi_rs1[16] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2871__CLK clknet_4_11_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_44_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1840_ _1293_ _1315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_29_316 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1771_ _1257_ net2 net6 _1258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_12_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2254_ _0415_ _0416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2323_ net47 _0479_ _0480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_2185_ _0367_ _0114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_63_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2622__A2 _0598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1969_ _1415_ _1420_ _1421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__2894__CLK clknet_4_8_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_3_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2310__A1 _0454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_9_Left_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2356__B _0490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1486__I _0973_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2377__A1 _0439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_9_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_60_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2941_ _0095_ clknet_4_6_0_clk picorv32_pcpi_div_inst_0.quotient\[26\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2872_ _0013_ clknet_4_11_0_clk net97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_25_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1823_ _1303_ _0040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_17_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1685_ picorv32_pcpi_div_inst_0.quotient\[20\] picorv32_pcpi_div_inst_0.quotient\[21\]
+ _1182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_52_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1754_ picorv32_pcpi_div_inst_0.quotient\[28\] picorv32_pcpi_div_inst_0.quotient\[29\]
+ _1223_ _1243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_25_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2540__A1 _0444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2237_ _0396_ _0400_ _0133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2306_ _0463_ _0464_ _0465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2168_ _0356_ _0108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2099_ picorv32_pcpi_div_inst_0.quotient_msk\[12\] _0310_ picorv32_pcpi_div_inst_0.quotient\[12\]
+ _0315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_51_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_0_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_17_Right_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_26_Right_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_8_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_425 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_35_Right_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_14_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1470_ _0981_ _0984_ _0986_ _0987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_34_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_65_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_44_Right_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2522__A1 _0414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_59_Left_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_53_Right_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2022_ _1394_ _0240_ _0249_ _0250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_9_316 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2924_ _0078_ clknet_4_13_0_clk picorv32_pcpi_div_inst_0.quotient\[9\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2855_ _0026_ clknet_4_6_0_clk net110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_45_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1806_ _1288_ _1289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_31_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2786_ net64 _0892_ _0893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XPHY_EDGE_ROW_62_Right_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1668_ _1086_ _1166_ _1167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1599_ _1100_ _1103_ _1104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1737_ picorv32_pcpi_div_inst_0.dividend\[28\] _1228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_40_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2513__A1 net33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2932__CLK clknet_4_14_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_28_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1555__A2 _1046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_36_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_4_3_0_clk clknet_0_clk clknet_4_3_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_6_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_42_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2640_ picorv32_pcpi_div_inst_0.divisor\[34\] _0753_ _0765_ _0766_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1453_ picorv32_pcpi_div_inst_0.quotient\[1\] _0971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2571_ net40 _0699_ _0490_ _0704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_10_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1522_ _1024_ picorv32_pcpi_div_inst_0.dividend\[5\] _1004_ _1007_ _1034_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__or4_2
X_2005_ picorv32_pcpi_div_inst_0.divisor\[16\] picorv32_pcpi_div_inst_0.dividend\[16\]
+ _0233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2907_ _0061_ clknet_4_10_0_clk picorv32_pcpi_div_inst_0.divisor\[23\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_33_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2769_ _0518_ _0878_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2838_ _0918_ _0936_ _0937_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_input56_I pcpi_rs2[14] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_51_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2978__CLK clknet_4_4_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_47_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput103 net103 pcpi_div_rd[27] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_42_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput114 net114 pcpi_div_rd[8] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_2623_ _0387_ _0751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2554_ net39 _0688_ _0689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_30_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1436_ _0954_ _0955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1505_ _1016_ _1018_ _1019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2485_ _1158_ _0402_ _0627_ _0154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_10_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_38_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3037_ _0189_ clknet_4_0_0_clk picorv32_pcpi_div_inst_0.divisor\[51\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__1997__A2 _1078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput16 pcpi_insn[4] net16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3006__CLK clknet_4_6_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput27 pcpi_rs1[17] net27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput38 pcpi_rs1[27] net38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput49 pcpi_rs1[8] net49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_58_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_32_280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1921__A2 _1134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2270_ _0430_ _0431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2783__I _0782_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1985_ _1318_ _1060_ _0213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1988__A2 _1074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2537_ _0244_ _0673_ _0674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2606_ net75 _0737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_15_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2468_ _0417_ _0612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_3_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_11_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2399_ _0509_ _0549_ _0550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_38_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3029__CLK clknet_4_1_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input19_I pcpi_rs1[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1979__A2 picorv32_pcpi_div_inst_0.dividend\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_44_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2108__I _0313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1770_ net116 _1257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2147__A2 _0342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2184_ picorv32_pcpi_div_inst_0.quotient_msk\[13\] _0363_ _0366_ picorv32_pcpi_div_inst_0.quotient_msk\[14\]
+ _0367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2253_ picorv32_pcpi_div_inst_0.instr_div picorv32_pcpi_div_inst_0.instr_rem _0415_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_20_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2322_ _0445_ _0478_ _0479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_63_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_40_Left_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_25_Left_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_1899_ _1355_ _0064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_7_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1968_ _1408_ _1417_ _1419_ _1414_ _1311_ _1420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XANTENNA__2386__A2 _0292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2688__I _0641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_54_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_3_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_26_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2547__B net38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2940_ _0094_ clknet_4_13_0_clk picorv32_pcpi_div_inst_0.quotient\[25\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_29_114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_17_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_60_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1753_ _1239_ _1240_ _0955_ _1242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2612__I0 _1042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2871_ _0012_ clknet_4_11_0_clk net96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_40_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_386 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1822_ _1300_ _1299_ _1295_ _1302_ _1303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_4_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1684_ picorv32_pcpi_div_inst_0.dividend\[22\] _1180_ _1084_ _1181_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_40_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2167_ picorv32_pcpi_div_inst_0.quotient_msk\[7\] _0355_ _0352_ picorv32_pcpi_div_inst_0.quotient_msk\[8\]
+ _0356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2236_ picorv32_pcpi_div_inst_0.running _0399_ _0400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2305_ _1304_ _1004_ _0464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2098_ _0313_ _0314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_51_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2861__CLK clknet_4_12_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_8_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_456 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2021_ _0245_ _0248_ _0249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2923_ _0077_ clknet_4_13_0_clk picorv32_pcpi_div_inst_0.quotient\[8\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_57_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2884__CLK clknet_4_3_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2854_ _0025_ clknet_4_12_0_clk net109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_53_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_53_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1805_ net83 _1287_ _1288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1736_ _1048_ _1226_ _1227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_31_40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2785_ net63 _0891_ _0886_ _0892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1667_ _1165_ _1166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1598_ _0977_ _1102_ _1103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1870__I _1320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2219_ _0387_ _0388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_63_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_36_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_12_Left_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2504__A2 _0402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2570_ _0703_ _0163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2440__B2 _0586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1521_ picorv32_pcpi_div_inst_0.quotient\[7\] _1032_ _1033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1452_ _0966_ _0969_ _0970_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2259__A1 net30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2004_ picorv32_pcpi_div_inst_0.divisor\[17\] picorv32_pcpi_div_inst_0.dividend\[17\]
+ _0232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2906_ _0060_ clknet_4_10_0_clk picorv32_pcpi_div_inst_0.divisor\[22\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_33_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1719_ _0947_ _1211_ _1212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_41_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2699_ picorv32_pcpi_div_inst_0.divisor\[41\] _0783_ _0817_ _0818_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_6_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2768_ _0877_ _0187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2837_ net72 _0935_ _0936_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__2498__A1 net31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input49_I pcpi_rs1[8] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_24_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_17_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2422__A1 _0459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput104 net104 pcpi_div_rd[28] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput115 net115 pcpi_div_rd[9] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__2922__CLK clknet_4_13_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1504_ _1006_ _1017_ _1018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2622_ _0748_ _0598_ _0749_ _0750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2510__S _0398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_30_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2553_ net38 _0682_ _0490_ _0688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2290__B _0449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1435_ _0945_ _0954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1634__B _1135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2484_ _0598_ _0621_ _0626_ _0342_ _0627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_53_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_38_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3036_ _0188_ clknet_4_0_0_clk picorv32_pcpi_div_inst_0.divisor\[50\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_4_2_0_clk clknet_0_clk clknet_4_2_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__2945__CLK clknet_4_4_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput17 pcpi_insn[5] net17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput39 pcpi_rs1[28] net39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_32_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput28 pcpi_rs1[18] net28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_20_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1984_ _0205_ _0206_ _0212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_15_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2536_ _0655_ _0248_ _0258_ _0673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2467_ _1369_ _0610_ _0611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2605_ _0719_ _0735_ _0736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2398_ _0489_ _0542_ _0548_ _0549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2968__CLK clknet_4_15_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3019_ _0171_ clknet_4_4_0_clk picorv32_pcpi_div_inst_0.divisor\[33\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2625__A1 _0747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_6_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2124__I _0329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2321_ net45 net46 _0457_ _0478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_2183_ _0358_ _0366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2252_ _0413_ _0414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_18_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_63_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1594__A1 _1091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1898_ picorv32_pcpi_div_inst_0.divisor\[26\] _1353_ _1350_ picorv32_pcpi_div_inst_0.divisor\[27\]
+ _1355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_28_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1967_ _1416_ picorv32_pcpi_div_inst_0.dividend\[5\] _1004_ _1418_ _1419_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2519_ _0423_ _0658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA_input31_I pcpi_rs1[20] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_54_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_3_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_19_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_22_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1888__A2 _1343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2065__A2 _0292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2870_ _0010_ clknet_4_11_0_clk net94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_17_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_60_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1752_ _1239_ _1240_ _1241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_44_118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1683_ _1123_ _1178_ _1180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_25_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1821_ picorv32_pcpi_div_inst_0.divisor\[3\] _1302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__3019__CLK clknet_4_4_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2304_ _1395_ _1396_ _1405_ _0463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_0_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_20_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2166_ _1352_ _0355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2097_ _1365_ _0313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_45_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2235_ _0398_ _0399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_0_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_51_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2999_ _0153_ clknet_4_9_0_clk picorv32_pcpi_div_inst_0.dividend\[19\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_28_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_3_Right_3 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1567__A1 picorv32_pcpi_div_inst_0.dividend\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input79_I pcpi_rs2[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_8_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2047__A2 _1249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1730__A1 _1153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2020_ _0246_ _0247_ _0248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2286__A2 net30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2922_ _0076_ clknet_4_13_0_clk picorv32_pcpi_div_inst_0.quotient\[7\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2853_ _0022_ clknet_4_12_0_clk net106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_31_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1666_ _1106_ _1130_ _1164_ _1165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_1735_ _1001_ _1224_ _1223_ _1226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_1804_ _1271_ _1287_ _0037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2784_ _0754_ _0891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_56_71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1597_ _1035_ _1034_ _1080_ _1101_ _1102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or4_2
XFILLER_0_0_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2149_ picorv32_pcpi_div_inst_0.quotient_msk\[0\] _1271_ _1358_ picorv32_pcpi_div_inst_0.quotient_msk\[1\]
+ _0345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2218_ _1297_ _0387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_36_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1547__B _1021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_59_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1520_ _1030_ _1031_ _1032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_2_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1451_ _0962_ _0952_ _0968_ _0969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__2851__CLK clknet_4_4_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2003_ _1382_ _1385_ _0231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_42_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_33_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2905_ _0059_ clknet_4_10_0_clk picorv32_pcpi_div_inst_0.divisor\[21\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_18_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2836_ _0734_ _0762_ _0935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1718_ _1001_ _1209_ _1208_ _1211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_1649_ _1145_ _1147_ _1149_ _1055_ _0009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_41_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1881__I _1320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2698_ _0811_ _0816_ _0817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2767_ _0876_ picorv32_pcpi_div_inst_0.divisor\[49\] _0395_ _0877_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_67_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2498__A2 net32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_24_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2874__CLK clknet_4_11_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_30_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2571__B _0490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_15_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput105 net105 pcpi_div_rd[29] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput116 net116 pcpi_div_ready vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_56_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1503_ _1005_ _1007_ _1017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_2621_ picorv32_pcpi_div_inst_0.divisor\[32\] _0658_ _0749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2552_ _0687_ _0161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2483_ _0407_ _0625_ _0626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_23_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1434_ picorv32_pcpi_div_inst_0.quotient\[0\] _0953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_38_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3035_ _0187_ clknet_4_0_0_clk picorv32_pcpi_div_inst_0.divisor\[49\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_58_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_58_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2819_ _0918_ _0920_ _0921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_14_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input61_I pcpi_rs2[19] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2897__CLK clknet_4_9_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput18 pcpi_insn[6] net18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_58_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput29 pcpi_rs1[19] net29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_17_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_59_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_43_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1983_ _1413_ _1421_ _0210_ _0211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_2604_ net72 _0734_ _0735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2535_ net37 _0671_ _0672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2466_ _1379_ _1142_ _0609_ _0610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_23_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1428__A3 _0947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3018_ _0170_ clknet_4_4_0_clk picorv32_pcpi_div_inst_0.divisor\[32\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2397_ _0545_ _0547_ _0548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_61_388 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2230__I _1289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_6_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_57_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2912__CLK clknet_4_4_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2251_ _0412_ _0413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2320_ _0477_ _0139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2182_ _0365_ _0113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_18_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_4_1_0_clk clknet_0_clk clknet_4_1_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_TAPCELL_ROW_63_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1966_ _1304_ _1418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_59_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1897_ _1354_ _0063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_28_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2935__CLK clknet_4_15_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2518_ _0655_ _0656_ _0657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2449_ _0424_ _0594_ _0595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input24_I pcpi_rs1[14] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_54_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_3_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_38_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_385 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1820_ _1301_ _0039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2222__B1 _0384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1751_ _1233_ _1229_ _1230_ _0983_ _1240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_1682_ _1177_ _0997_ _1178_ _1179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_40_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2958__CLK clknet_4_13_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2234_ _0397_ _0398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_0_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2303_ _0459_ _0461_ _0462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2096_ _0307_ _0312_ _0080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2165_ _0354_ _0107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_51_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_48_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2998_ _0152_ clknet_4_10_0_clk picorv32_pcpi_div_inst_0.dividend\[18\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1949_ _1399_ picorv32_pcpi_div_inst_0.dividend\[0\] _1400_ _1401_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_28_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2516__A1 _1394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_8_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2204__B1 _0378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1494__A1 _1005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2286__A3 net41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_13_Right_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_15_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2921_ _0075_ clknet_4_7_0_clk picorv32_pcpi_div_inst_0.quotient\[6\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2852_ _0011_ clknet_4_12_0_clk net95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1803_ _1273_ _1286_ _1287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_45_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_22_Right_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2783_ _0782_ _0890_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_15_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1665_ picorv32_pcpi_div_inst_0.quotient\[16\] picorv32_pcpi_div_inst_0.quotient\[17\]
+ picorv32_pcpi_div_inst_0.quotient\[18\] picorv32_pcpi_div_inst_0.quotient\[19\]
+ _1164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_1734_ _0960_ _1223_ _1224_ _1225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_40_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_40_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1596_ _1094_ _1078_ _1101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_0_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_13_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2217_ _0386_ _0127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_EDGE_ROW_37_Left_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_31_Right_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2079_ _0301_ _0302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__1485__A1 _0997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2148_ _0339_ _0344_ _0100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_EDGE_ROW_46_Left_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_36_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_40_Right_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_36_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_55_Left_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_64_Left_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_54_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3009__CLK clknet_4_3_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1450_ _0967_ _0968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_22_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1473__B _0973_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2002_ _0219_ _0229_ _0230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_41_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_33_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2904_ _0058_ clknet_4_10_0_clk picorv32_pcpi_div_inst_0.divisor\[20\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_5_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2766_ _0405_ _0874_ _0875_ _0876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2835_ _0912_ _0933_ _0934_ _0197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_13_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1648_ picorv32_pcpi_div_inst_0.quotient\[18\] _1148_ _1149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1579_ _1020_ _1086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1717_ _0960_ _1208_ _1209_ _1210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2697_ net82 _0815_ _0816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_36_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_24_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_59_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1621__A1 _1113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2620_ net51 _0748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_30_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput106 net106 pcpi_div_rd[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput117 net117 pcpi_div_wait vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_1433_ _0951_ _0952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2551_ _1217_ _0686_ _0678_ _0687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2482_ net31 _0624_ _0625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_10_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1502_ picorv32_pcpi_div_inst_0.dividend\[5\] _1016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_49_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_38_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3034_ _0186_ clknet_4_0_0_clk picorv32_pcpi_div_inst_0.divisor\[48\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_58_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_46_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2818_ net69 _0919_ _0920_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2749_ _0726_ _0861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_input54_I pcpi_rs2[12] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_394 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput19 pcpi_rs1[0] net19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2991__CLK clknet_4_8_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1751__B _0983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2331__A2 _0292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1982_ _0204_ _0209_ _0210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2534_ _0455_ _0670_ _0671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2603_ net70 net71 _0733_ _0734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_2465_ _0599_ _0601_ _0609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_2_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2396_ _0404_ _0546_ _0547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3017_ _0169_ clknet_4_4_0_clk picorv32_pcpi_div_inst_0.divisor\[31\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2864__CLK clknet_4_14_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_353 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_57_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1481__B _0996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2250_ _1364_ _0412_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_20_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2181_ picorv32_pcpi_div_inst_0.quotient_msk\[12\] _0363_ _0359_ picorv32_pcpi_div_inst_0.quotient_msk\[13\]
+ _0365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_34_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2887__CLK clknet_4_3_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_43_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1965_ _1416_ _1016_ _1417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_59_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1896_ picorv32_pcpi_div_inst_0.divisor\[25\] _1353_ _1350_ picorv32_pcpi_div_inst_0.divisor\[26\]
+ _1354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2517_ _0247_ _0656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_3_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2448_ _0232_ _0593_ _0594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_3_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2379_ _0509_ _0531_ _0532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input17_I pcpi_insn[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_54_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2707__S _0395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_46_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3042__CLK clknet_4_2_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output85_I net85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2298__A1 net19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_44_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1750_ picorv32_pcpi_div_inst_0.dividend\[30\] _1239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_29_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2470__A1 net29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2151__I _1349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1681_ picorv32_pcpi_div_inst_0.dividend\[21\] picorv32_pcpi_div_inst_0.dividend\[20\]
+ _1160_ _1178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XPHY_EDGE_ROW_29_Left_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_25_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2164_ picorv32_pcpi_div_inst_0.quotient_msk\[6\] _0349_ _0352_ picorv32_pcpi_div_inst_0.quotient_msk\[7\]
+ _0354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_input9_I pcpi_insn[27] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2233_ _1292_ _0397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2302_ _0460_ _0457_ net45 _0461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_0_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2095_ picorv32_pcpi_div_inst_0.quotient_msk\[11\] _0310_ picorv32_pcpi_div_inst_0.quotient\[11\]
+ _0312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_TAPCELL_ROW_51_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_0_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1879_ picorv32_pcpi_div_inst_0.divisor\[20\] _1336_ _1340_ _1341_ _1342_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1948_ picorv32_pcpi_div_inst_0.divisor\[1\] _0961_ _1400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_28_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2997_ _0151_ clknet_4_9_0_clk picorv32_pcpi_div_inst_0.dividend\[17\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_16_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2902__CLK clknet_4_9_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_8_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_429 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_4_0_0_clk clknet_0_clk clknet_4_0_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_2920_ _0074_ clknet_4_7_0_clk picorv32_pcpi_div_inst_0.quotient\[5\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2925__CLK clknet_4_13_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1802_ _1277_ _1280_ _1285_ _1286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_57_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1733_ picorv32_pcpi_div_inst_0.quotient\[28\] _1224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2851_ _0000_ clknet_4_4_0_clk net84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_45_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2782_ _0885_ _0396_ _0888_ _0889_ _0189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_TAPCELL_ROW_13_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1664_ picorv32_pcpi_div_inst_0.dividend\[20\] _1162_ _1084_ _1163_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1595_ picorv32_pcpi_div_inst_0.dividend\[14\] _1100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_25_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2216_ picorv32_pcpi_div_inst_0.quotient_msk\[26\] _0381_ _0384_ picorv32_pcpi_div_inst_0.quotient_msk\[27\]
+ _0386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2147_ picorv32_pcpi_div_inst_0.quotient_msk\[31\] _0342_ picorv32_pcpi_div_inst_0.quotient\[31\]
+ _0344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2484__C _0342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2078_ _0290_ _0301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_48_289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1895__I _1352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_36_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_27_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2425__B2 _0433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2001_ _0221_ _0223_ _0200_ _0227_ _0228_ _0229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_0_42_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2903_ _0057_ clknet_4_10_0_clk picorv32_pcpi_div_inst_0.divisor\[19\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2416__B2 _0469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1716_ picorv32_pcpi_div_inst_0.quotient\[26\] _1209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_33_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2696_ _0812_ _0814_ _0815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2765_ picorv32_pcpi_div_inst_0.divisor\[50\] _0581_ _0875_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2834_ picorv32_pcpi_div_inst_0.divisor\[59\] _0923_ _0934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_13_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1647_ _1129_ _1138_ _1131_ _0973_ _1148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_1578_ picorv32_pcpi_div_inst_0.dividend\[12\] _1083_ _1084_ _1085_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_6_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_49_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_16_Left_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_51_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_24_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1621__A2 _1100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput107 net107 pcpi_div_rd[30] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_2550_ _0586_ _0681_ _0683_ _0685_ _0686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_23_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput118 net118 pcpi_div_wr vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_1501_ _0947_ _1014_ _1015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_37_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1432_ picorv32_pcpi_div_inst_0.dividend\[0\] _0951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2481_ _0434_ _0623_ _0624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3033_ _0185_ clknet_4_0_0_clk picorv32_pcpi_div_inst_0.divisor\[47\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_46_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2679_ picorv32_pcpi_div_inst_0.divisor\[38\] _0780_ _0800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_5_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2748_ _0839_ _0859_ _0860_ _0184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_14_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2817_ _0732_ _0848_ _0919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_input47_I pcpi_rs1[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_1_Left_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_64_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2244__I _0406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1479__B _0985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1981_ _0205_ _0206_ _0207_ _0208_ _0209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_2533_ net35 net36 _0652_ _0670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_2_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2602_ net69 _0732_ _0733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_2464_ _1143_ _0402_ _0608_ _0152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2395_ _0202_ _0544_ _0546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3016_ _0168_ clknet_4_3_0_clk picorv32_pcpi_div_inst_0.divisor\[62\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_46_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1597__A1 _1035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_57_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_37_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2180_ _0364_ _0112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_20_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1895_ _1352_ _1353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_28_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1964_ picorv32_pcpi_div_inst_0.divisor\[5\] _1416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__1672__B _1135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2516_ _1394_ _0240_ _0655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2447_ _1374_ _1121_ _0592_ _0593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_11_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1503__A1 _1005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_3_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2378_ _0519_ _0523_ _0528_ _0530_ _0531_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XTAP_TAPCELL_ROW_62_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_54_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2981__CLK clknet_4_3_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2298__A2 net30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2432__I net26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_4_Left_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_13_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1680_ _1176_ _1177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2301_ _0445_ _0460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_20_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2163_ _0353_ _0106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2854__CLK clknet_4_12_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2232_ _0395_ _0396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2094_ _0307_ _0311_ _0079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_51_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_16_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1878_ picorv32_pcpi_div_inst_0.divisor\[21\] _1341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1947_ picorv32_pcpi_div_inst_0.divisor\[0\] _1399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_2996_ _0150_ clknet_4_9_0_clk picorv32_pcpi_div_inst_0.dividend\[16\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_9_20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2877__CLK clknet_4_12_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_30_Left_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2850_ _0036_ clknet_4_4_0_clk picorv32_pcpi_div_inst_0.instr_div vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_15_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1801_ _1281_ _1282_ _1283_ _1284_ _1285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_0_53_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1732_ picorv32_pcpi_div_inst_0.quotient\[26\] picorv32_pcpi_div_inst_0.quotient\[27\]
+ _1208_ _1223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_1663_ _1123_ _1160_ _1162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_31_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2781_ picorv32_pcpi_div_inst_0.divisor\[52\] _0808_ _0809_ _0889_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_13_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1594_ _1091_ _1093_ _1099_ _0004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1706__B2 _1169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_7_Right_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2215_ _0385_ _0126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2077_ _0298_ _0300_ _0073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2146_ _0339_ _0343_ _0099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3032__CLK clknet_4_0_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_36_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2979_ _0133_ clknet_4_1_0_clk picorv32_pcpi_div_inst_0.running vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_8_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input77_I pcpi_rs2[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_27_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2361__A1 _0439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2000_ _0220_ picorv32_pcpi_div_inst_0.dividend\[15\] _0228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2902_ _0056_ clknet_4_9_0_clk picorv32_pcpi_div_inst_0.divisor\[18\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2833_ picorv32_pcpi_div_inst_0.divisor\[60\] _0466_ _0932_ _0933_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1715_ picorv32_pcpi_div_inst_0.quotient\[24\] picorv32_pcpi_div_inst_0.quotient\[25\]
+ _1198_ _1208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XANTENNA__1437__S _0955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1646_ _1142_ _1146_ _1084_ _1147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_41_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2695_ _0813_ _0802_ _0814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2764_ net60 _0873_ _0874_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_13_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1577_ _0954_ _1084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2129_ _0313_ _0333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_TAPCELL_ROW_49_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_24_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_32_499 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2915__CLK clknet_4_6_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput108 net108 pcpi_div_rd[31] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_1500_ _1001_ _1012_ _1011_ _1014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_50_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1621__A3 _1102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2480_ _0578_ _0622_ _0623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_23_499 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput90 net90 pcpi_div_rd[15] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_1431_ _0950_ _0033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3032_ _0184_ clknet_4_0_0_clk picorv32_pcpi_div_inst_0.divisor\[46\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_46_503 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2816_ _0518_ _0918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2938__CLK clknet_4_14_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1629_ _1086_ _1131_ _1132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2678_ picorv32_pcpi_div_inst_0.divisor\[39\] _0783_ _0798_ _0799_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2747_ picorv32_pcpi_div_inst_0.divisor\[46\] _0853_ _0860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_49_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1980_ picorv32_pcpi_div_inst_0.divisor\[8\] _1046_ _0208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_0_7_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2532_ _0669_ _0159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2463_ _0598_ _0602_ _0607_ _0342_ _0608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_23_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2601_ net68 net67 _0731_ _0732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_3015_ _0167_ clknet_4_4_0_clk picorv32_pcpi_div_inst_0.instr_remu vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_3_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2394_ _0202_ _0544_ _0545_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_46_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_46_355 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2546__A1 net37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1597__A2 _1034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_57_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_40_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_388 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1894_ _1297_ _1352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_43_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2528__A1 net35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_355 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_1963_ _1311_ _1414_ _1025_ picorv32_pcpi_div_inst_0.divisor\[6\] _1415_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_2515_ net35 _0653_ _0654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2446_ _0591_ _0233_ _0592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_11_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_54_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1503__A2 _1007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2377_ _0439_ _0529_ _0530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_TAPCELL_ROW_62_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2216__B1 _0384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_19_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2298__A3 net41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2300_ _0412_ _0459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2231_ _0394_ _0395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_2162_ picorv32_pcpi_div_inst_0.quotient_msk\[5\] _0349_ _0352_ picorv32_pcpi_div_inst_0.quotient_msk\[6\]
+ _0353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2093_ picorv32_pcpi_div_inst_0.quotient_msk\[10\] _0310_ _1067_ _0311_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_45_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2623__I _0387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_16_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2995_ _0149_ clknet_4_9_0_clk picorv32_pcpi_div_inst_0.dividend\[15\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_43_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1877_ _1316_ _1340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_28_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1946_ _1397_ _0961_ _1398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_24_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1488__A1 _0947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2429_ net24 net25 _0576_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA_input22_I pcpi_rs1[12] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_66_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_62_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_22_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_497 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1800_ picorv32_pcpi_div_inst_0.quotient_msk\[14\] picorv32_pcpi_div_inst_0.quotient_msk\[13\]
+ picorv32_pcpi_div_inst_0.quotient_msk\[12\] picorv32_pcpi_div_inst_0.quotient_msk\[11\]
+ _1284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_0_38_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1731_ _1116_ _1219_ _1222_ _0019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1662_ _1158_ _0997_ _1160_ _1161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_25_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2451__I0 _1134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2780_ _0399_ _0887_ _0888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2971__CLK clknet_4_13_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2214_ picorv32_pcpi_div_inst_0.quotient_msk\[25\] _0381_ _0384_ picorv32_pcpi_div_inst_0.quotient_msk\[26\]
+ _0385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1593_ _1029_ _1098_ _1099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_0_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2076_ picorv32_pcpi_div_inst_0.quotient_msk\[4\] _0294_ _0999_ _0300_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2145_ picorv32_pcpi_div_inst_0.quotient_msk\[30\] _0342_ picorv32_pcpi_div_inst_0.quotient\[30\]
+ _0343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_48_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2978_ _0132_ clknet_4_4_0_clk picorv32_pcpi_div_inst_0.quotient_msk\[31\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_36_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1929_ _1378_ _1380_ _1381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_31_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_27_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_33_Left_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_22_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_42_Left_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2994__CLK clknet_4_8_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2901_ _0055_ clknet_4_9_0_clk picorv32_pcpi_div_inst_0.divisor\[17\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2763_ net59 net58 _0861_ _0812_ _0873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_2832_ _0918_ _0931_ _0932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1714_ _1112_ _1204_ _1207_ _0017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1517__I _0964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1576_ _0968_ _1081_ _1083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1645_ _1123_ _1144_ _1146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2694_ net81 _0813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2128_ _0326_ _0332_ _0092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_49_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2867__CLK clknet_4_11_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2059_ _1368_ _0273_ _0275_ _0286_ _0287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XTAP_TAPCELL_ROW_24_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_423 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_32_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput109 net109 pcpi_div_rd[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_50_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1430_ net117 _0948_ _0950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__3022__CLK clknet_4_1_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput91 net91 pcpi_div_rd[16] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_37_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3031_ _0183_ clknet_4_0_0_clk picorv32_pcpi_div_inst_0.divisor\[45\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_58_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2022__A1 _1394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2815_ _0912_ _0916_ _0917_ _0194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2746_ picorv32_pcpi_div_inst_0.divisor\[47\] _0855_ _0858_ _0859_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_14_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1628_ _1107_ _1130_ _1131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1559_ _1050_ _1056_ _1052_ _0959_ _1068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_2677_ _0775_ _0797_ _0798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_14_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2078__I _0290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3045__CLK clknet_4_2_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_67_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2600_ _0728_ _0729_ _0730_ _0731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_2531_ _1201_ _0668_ _0634_ _0669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2462_ _0407_ _0606_ _0607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_23_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2393_ _0501_ _0209_ _0543_ _0544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_47_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3014_ _0166_ clknet_4_4_0_clk picorv32_pcpi_div_inst_0.outsign vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_58_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_58_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2626__I _0641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2491__A1 _0414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2905__CLK clknet_4_10_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1597__A3 _1080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2729_ picorv32_pcpi_div_inst_0.divisor\[45\] _0826_ _0843_ _0844_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_input52_I pcpi_rs2[10] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_57_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1440__I _0957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_29_Right_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2482__A1 net31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_40_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_38_Right_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_37_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_4_7_0_clk_I clknet_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_47_Right_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2928__CLK clknet_4_13_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_56_Right_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_50_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_28_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1962_ picorv32_pcpi_div_inst_0.dividend\[7\] _1414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_16_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1893_ _1351_ _0062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_28_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_65_Right_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2445_ _0211_ _0230_ _0591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2514_ _0455_ _0652_ _0653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2376_ _0524_ _0527_ _0529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_11_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_54_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_19_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_62_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2216__B2 picorv32_pcpi_div_inst_0.quotient_msk\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1435__I _0945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2298__A4 net44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_2_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_315 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2230_ _1289_ _0394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2161_ _1349_ _0352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2092_ _0301_ _0310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_48_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1945_ picorv32_pcpi_div_inst_0.divisor\[1\] _1397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2994_ _0148_ clknet_4_8_0_clk picorv32_pcpi_div_inst_0.dividend\[14\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_43_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1876_ _1339_ _0057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2428_ _0575_ _0149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2359_ _0502_ _0503_ _0512_ _0513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_66_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input15_I pcpi_insn[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2437__A1 _0211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_34_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_22_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2724__I _0768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1730_ _1153_ _1221_ _1222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_40_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1592_ _1095_ _1097_ _1098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1661_ _1113_ picorv32_pcpi_div_inst_0.dividend\[14\] _1102_ _1159_ _1160_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__or4_2
XFILLER_0_21_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2213_ _1315_ _0384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_56_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input7_I pcpi_insn[25] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2144_ _0290_ _0342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2075_ _0298_ _0299_ _0072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_48_215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2977_ _0131_ clknet_4_5_0_clk picorv32_pcpi_div_inst_0.quotient_msk\[30\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1928_ _1377_ _1150_ picorv32_pcpi_div_inst_0.dividend\[18\] _1379_ _1380_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_1859_ _1329_ _0050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_16_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_4_15_0_clk_I clknet_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2809__I _1298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_35_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_27_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_10_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2900_ _0054_ clknet_4_9_0_clk picorv32_pcpi_div_inst_0.divisor\[16\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1713_ _1153_ _1206_ _1207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_5_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2762_ _0867_ _0871_ _0872_ _0186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2831_ net71 _0930_ _0931_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1575_ _1078_ _1042_ _1081_ _1082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_1644_ _1143_ _1042_ _1144_ _1145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_6_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2693_ _0755_ _0812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2127_ picorv32_pcpi_div_inst_0.quotient_msk\[23\] _0330_ picorv32_pcpi_div_inst_0.quotient\[23\]
+ _0332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_64_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2058_ _0280_ _0285_ _0286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_24_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_32_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input82_I pcpi_rs2[9] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1551__A1 _1046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2961__CLK clknet_4_15_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1542__A1 _0993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput92 net92 pcpi_div_rd[17] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__2385__S _0459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3030_ _0182_ clknet_4_1_0_clk picorv32_pcpi_div_inst_0.divisor\[44\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_58_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_61_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2676_ net80 _0796_ _0797_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_26_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2814_ picorv32_pcpi_div_inst_0.divisor\[56\] _0883_ _0917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2745_ _0846_ _0857_ _0858_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_14_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_1558_ picorv32_pcpi_div_inst_0.quotient\[10\] _1067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1627_ picorv32_pcpi_div_inst_0.quotient\[14\] picorv32_pcpi_div_inst_0.quotient\[15\]
+ _1130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1489_ picorv32_pcpi_div_inst_0.dividend\[4\] _1004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_61_Left_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_49_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2984__CLK clknet_4_2_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2269__I _0290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1524__A1 _0997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_43_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2530_ _0663_ _0665_ _0667_ _0433_ _0668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_0_23_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_4_3_0_clk_I clknet_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2857__CLK clknet_4_13_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1515__A1 _1025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2461_ net28 _0605_ _0606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2392_ _0215_ _0218_ _0543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3013_ _0033_ clknet_4_4_0_clk picorv32_pcpi_div_inst_0.pcpi_wait_q vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_58_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2659_ _0423_ _0782_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2728_ _0811_ _0842_ _0843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3012__CLK clknet_4_4_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input45_I pcpi_rs1[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_57_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_40_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2501__B _0641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_5_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1892_ picorv32_pcpi_div_inst_0.divisor\[24\] _1343_ _1350_ picorv32_pcpi_div_inst_0.divisor\[25\]
+ _1351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_34_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1961_ _1395_ _1396_ _1405_ _1412_ _1413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_0_51_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2513_ net33 net34 _0639_ _0652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XANTENNA__2411__B net24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2444_ net27 _0589_ _0590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__3035__CLK clknet_4_0_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2375_ _0524_ _0527_ _0528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2464__A2 _0402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_19_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_62_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_2_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2160_ _0351_ _0105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_45_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_29_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2391__A1 net22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2091_ _0307_ _0309_ _0078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_45_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_45_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_61_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1875_ picorv32_pcpi_div_inst_0.divisor\[19\] _1336_ _1334_ picorv32_pcpi_div_inst_0.divisor\[20\]
+ _1339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_28_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1944_ _1302_ _0991_ _0980_ _1300_ _1396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_8_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2993_ _0147_ clknet_4_8_0_clk picorv32_pcpi_div_inst_0.dividend\[13\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2568__S _0404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2427_ _1113_ _0573_ _0574_ _0575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_3_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_67_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_4_15_0_clk clknet_0_clk clknet_4_15_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_2289_ _0397_ _0449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2358_ _1313_ _1041_ _0512_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_clkbuf_4_11_0_clk_I clknet_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2316__B _0449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_22_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_8_Left_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_53_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_31_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1591_ picorv32_pcpi_div_inst_0.dividend\[12\] _1081_ _1096_ _1097_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1660_ picorv32_pcpi_div_inst_0.dividend\[19\] picorv32_pcpi_div_inst_0.dividend\[18\]
+ picorv32_pcpi_div_inst_0.dividend\[17\] _1121_ _1159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_0_21_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2364__A1 _1060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2212_ _0383_ _0125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2143_ _0339_ _0341_ _0098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2074_ picorv32_pcpi_div_inst_0.quotient_msk\[3\] _0294_ picorv32_pcpi_div_inst_0.quotient\[3\]
+ _0299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_48_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2976_ _0130_ clknet_4_5_0_clk picorv32_pcpi_div_inst_0.quotient_msk\[29\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_29_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1927_ picorv32_pcpi_div_inst_0.divisor\[18\] _1379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_24_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_12_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1858_ picorv32_pcpi_div_inst_0.divisor\[12\] _1321_ _1327_ _1328_ _1329_ vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1789_ net117 _1272_ _1273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_12_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output114_I net114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_27_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_35_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_10_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2890__CLK clknet_4_2_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2830_ net70 _0733_ _0891_ _0930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_53_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1712_ picorv32_pcpi_div_inst_0.quotient\[25\] _1205_ _1206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_1643_ _1134_ _1121_ _1124_ _1144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XANTENNA__2585__A1 _0586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2692_ _0432_ _0811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2761_ picorv32_pcpi_div_inst_0.divisor\[48\] _0853_ _0872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1574_ _1044_ _1080_ _1081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_0_6_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2126_ _0326_ _0331_ _0091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2057_ _0281_ _0282_ _0283_ _0284_ _0285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__2846__S _0395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2959_ _0113_ clknet_4_13_0_clk picorv32_pcpi_div_inst_0.quotient_msk\[12\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_44_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_32_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_24_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2576__A1 _0444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input75_I pcpi_rs2[31] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2567__A1 net40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_458 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput93 net93 pcpi_div_rd[18] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_53_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_38_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2813_ picorv32_pcpi_div_inst_0.divisor\[57\] _0890_ _0915_ _0916_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1626_ picorv32_pcpi_div_inst_0.quotient\[16\] _1129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_41_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2558__A1 _0658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2675_ net79 _0789_ _0762_ _0796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_26_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2744_ net57 _0856_ _0857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1488_ _0947_ _1002_ _1003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1557_ picorv32_pcpi_div_inst_0.dividend\[10\] _1065_ _1066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2109_ picorv32_pcpi_div_inst_0.quotient_msk\[16\] _0317_ _1129_ _0321_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_49_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2549__A1 _0398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1454__I picorv32_pcpi_div_inst_0.outsign vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1524__A2 _1034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_43_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2460_ _0434_ _0604_ _0605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_EDGE_ROW_21_Left_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_48_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2391_ net22 _0541_ _0542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_58_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3012_ _0032_ clknet_4_4_0_clk net117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_58_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2658_ _0769_ _0779_ _0781_ _0173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2589_ net62 net51 net76 net73 _0720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or4_2
X_1609_ picorv32_pcpi_div_inst_0.dividend\[15\] _1113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_14_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2727_ net55 _0841_ _0842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_TAPCELL_ROW_57_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input38_I pcpi_rs1[27] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_40_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_45_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1449__I _0957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_5_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1891_ _1349_ _1350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_36_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1960_ _1408_ _1411_ _1412_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_59_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2512_ _0651_ _0157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2443_ _0579_ _0578_ _0520_ _0589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2374_ _0525_ _0207_ _0208_ _0526_ _0527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_0_46_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2152__A2 _1360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_2_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_464 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2997__CLK clknet_4_9_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2090_ picorv32_pcpi_div_inst_0.quotient_msk\[9\] _0302_ _1056_ _0309_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_48_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2992_ _0146_ clknet_4_8_0_clk picorv32_pcpi_div_inst_0.dividend\[12\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3002__CLK clknet_4_10_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1874_ _1338_ _0056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1943_ _1302_ _0992_ _1395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_9_24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1817__I _1298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_24_Left_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2426_ _0430_ _0574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_TAPCELL_ROW_67_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2288_ _1300_ _0981_ _0440_ _0448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2357_ net50 _0510_ _0511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_66_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3025__CLK clknet_4_1_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_13_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1590_ _0957_ _1096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_0_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2211_ picorv32_pcpi_div_inst_0.quotient_msk\[24\] _0381_ _0378_ picorv32_pcpi_div_inst_0.quotient_msk\[25\]
+ _0383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2073_ _0297_ _0298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_56_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2142_ picorv32_pcpi_div_inst_0.quotient_msk\[29\] _0336_ picorv32_pcpi_div_inst_0.quotient\[29\]
+ _0341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2975_ _0129_ clknet_4_5_0_clk picorv32_pcpi_div_inst_0.quotient_msk\[28\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_29_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2427__I0 _1113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1788_ picorv32_pcpi_div_inst_0.pcpi_wait_q _1272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_44_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1926_ _1377_ _1150_ _1378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1857_ picorv32_pcpi_div_inst_0.divisor\[13\] _1328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2409_ net22 net23 _0540_ _0558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XANTENNA_input20_I pcpi_rs1[10] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_27_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_35_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_10_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_4_14_0_clk clknet_0_clk clknet_4_14_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_53_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1711_ picorv32_pcpi_div_inst_0.quotient\[24\] _1198_ _0982_ _1205_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1642_ _1142_ _1143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2691_ _0801_ _0396_ _0807_ _0810_ _0177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2760_ picorv32_pcpi_div_inst_0.divisor\[49\] _0855_ _0870_ _0871_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2337__A2 _1025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2198__I _0362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1573_ _1074_ _1079_ _1059_ _1040_ _1080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_2125_ picorv32_pcpi_div_inst_0.quotient_msk\[22\] _0330_ picorv32_pcpi_div_inst_0.quotient\[22\]
+ _0331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2056_ picorv32_pcpi_div_inst_0.divisor\[35\] picorv32_pcpi_div_inst_0.divisor\[34\]
+ picorv32_pcpi_div_inst_0.divisor\[33\] picorv32_pcpi_div_inst_0.divisor\[32\] _0284_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XANTENNA__1830__I _1298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2958_ _0112_ clknet_4_13_0_clk picorv32_pcpi_div_inst_0.quotient_msk\[11\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_1909_ picorv32_pcpi_div_inst_0.divisor\[31\] _1362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2908__CLK clknet_4_11_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_32_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2889_ _0043_ clknet_4_2_0_clk picorv32_pcpi_div_inst_0.divisor\[5\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_input68_I pcpi_rs2[25] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2264__A1 _0414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput94 net94 pcpi_div_rd[19] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_31_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_46_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2255__A1 net43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2812_ _0878_ _0914_ _0915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2743_ net56 _0847_ _0840_ _0856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1625_ _1127_ _1128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1556_ _0993_ _1064_ _1065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2674_ _0768_ _0795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_1_320 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1487_ _1001_ _0999_ _0998_ _1002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__2656__I _0387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2108_ _0313_ _0320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2039_ _1356_ _0266_ _0267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2246__A1 _0407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2880__CLK clknet_4_12_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2767__S _0395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_67_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_43_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3011_ _0165_ clknet_4_3_0_clk picorv32_pcpi_div_inst_0.dividend\[31\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_2390_ _0419_ _0540_ _0541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_46_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1451__A2 _0952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_6_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2400__A1 _1078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2726_ net54 _0833_ _0840_ _0841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1539_ picorv32_pcpi_div_inst_0.quotient\[8\] _1050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1608_ _0955_ _1112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2657_ picorv32_pcpi_div_inst_0.divisor\[35\] _0780_ _0781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2588_ net74 _0719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_1_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_64_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_40_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2335__B _0490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1465__I _0957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_5_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_16_Right_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_50_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1890_ _1315_ _1349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_36_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_25_Right_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_59_12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2511_ picorv32_pcpi_div_inst_0.dividend\[23\] _0650_ _0634_ _0651_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2442_ _0588_ _0150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2373_ _0213_ _0214_ _0526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_45_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_34_Right_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2449__A1 _0424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_49_Left_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_46_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_43_Right_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_42_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2709_ _0782_ _0826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_58_Left_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_52_Right_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_input50_I pcpi_rs1[9] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_2_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_67_Left_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_61_Right_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_52_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1942_ _1390_ _1392_ _1393_ _1394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_28_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2991_ _0145_ clknet_4_8_0_clk picorv32_pcpi_div_inst_0.dividend\[11\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__2941__CLK clknet_4_6_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1873_ picorv32_pcpi_div_inst_0.divisor\[18\] _1336_ _1334_ picorv32_pcpi_div_inst_0.divisor\[19\]
+ _1338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_3_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_10_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2425_ _0568_ _0570_ _0572_ _0433_ _0573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_2356_ net49 _0498_ _0490_ _0510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_67_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2287_ net44 _0446_ _0447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_62_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2964__CLK clknet_4_15_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_21_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_13_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2210_ _0382_ _0124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2141_ _0339_ _0340_ _0097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2072_ _1366_ _0297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2974_ _0128_ clknet_4_5_0_clk picorv32_pcpi_div_inst_0.quotient_msk\[27\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_44_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1925_ picorv32_pcpi_div_inst_0.divisor\[19\] _1377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_8_326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1787_ _0948_ _1271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_12_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1856_ _1316_ _1327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_EDGE_ROW_2_Right_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2339_ _1406_ _0493_ _0494_ _0495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2408_ _1095_ _0508_ _0557_ _0147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_input13_I pcpi_insn[30] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_27_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2987__CLK clknet_4_8_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_35_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_10_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2806__A1 _0598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_38_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1710_ _1201_ _1203_ _1204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1641_ picorv32_pcpi_div_inst_0.dividend\[18\] _1142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2690_ picorv32_pcpi_div_inst_0.divisor\[40\] _0808_ _0809_ _0810_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_6_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1572_ picorv32_pcpi_div_inst_0.dividend\[10\] _1079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_2124_ _0329_ _0330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_input5_I pcpi_insn[14] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2055_ picorv32_pcpi_div_inst_0.divisor\[39\] picorv32_pcpi_div_inst_0.divisor\[38\]
+ picorv32_pcpi_div_inst_0.divisor\[37\] picorv32_pcpi_div_inst_0.divisor\[36\] _0283_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_0_16_71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2957_ _0111_ clknet_4_13_0_clk picorv32_pcpi_div_inst_0.quotient_msk\[10\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_44_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1908_ _1361_ _0067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1839_ _1314_ _0045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_8_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2888_ _0042_ clknet_4_2_0_clk picorv32_pcpi_div_inst_0.divisor\[4\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_17_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3015__CLK clknet_4_4_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2338__B _0406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1527__A1 _1037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput84 net84 pcpi_div_rd[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput95 net95 pcpi_div_rd[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_46_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1766__A1 _1091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2742_ _0782_ _0855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2811_ net68 _0913_ _0914_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1624_ _1122_ _1125_ _0965_ _1127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_41_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1555_ picorv32_pcpi_div_inst_0.dividend\[9\] _1046_ _1043_ _1064_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__or3_1
X_2673_ _0769_ _0793_ _0794_ _0175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3038__CLK clknet_4_0_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2107_ _0314_ _0319_ _0084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1486_ _0973_ _1001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1841__I _1315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_390 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2038_ _0265_ picorv32_pcpi_div_inst_0.dividend\[29\] _1228_ _0266_ vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_input80_I pcpi_rs2[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_4_13_0_clk clknet_0_clk clknet_4_13_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_40_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2485__A2 _0402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2582__I net43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1748__A1 _1153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_43_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3010_ _0164_ clknet_4_1_0_clk picorv32_pcpi_div_inst_0.dividend\[30\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_58_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1610__B _1021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2228__A2 _1291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2492__I _0430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2656_ _0387_ _0780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_6_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2725_ _0754_ _0840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1607_ _0976_ _1104_ _1109_ _1111_ _0005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1538_ _1046_ _1047_ _1048_ _1049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1469_ _0981_ _0984_ _0985_ _0986_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2587_ _0718_ _0165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1571__I picorv32_pcpi_div_inst_0.dividend\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_64_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_40_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2458__A2 net27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_5_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2510_ _0647_ _0649_ _0398_ _0650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_3_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1605__B _0985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2441_ _1122_ _0587_ _0574_ _0588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_2372_ _0502_ _0525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_59_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2870__CLK clknet_4_11_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2621__A2 _0658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2137__A1 picorv32_pcpi_div_inst_0.quotient_msk\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2639_ _0519_ _0764_ _0765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2708_ _0825_ _0179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1896__B1 _1350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input43_I pcpi_rs1[31] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_53_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_37_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_33_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2893__CLK clknet_4_8_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1941_ _1346_ _1188_ _1393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_28_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1872_ _1337_ _0055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2990_ _0144_ clknet_4_8_0_clk picorv32_pcpi_div_inst_0.dividend\[10\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_TAPCELL_ROW_16_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_67_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_67_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2286_ _0403_ net30 net41 _0445_ _0446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_2424_ net25 _0571_ _0572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_19_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2355_ _0430_ _0509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_47_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1581__A2 _1031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2530__B2 _0433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_13_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2140_ picorv32_pcpi_div_inst_0.quotient_msk\[28\] _0336_ _1224_ _0340_ vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2521__A1 _0658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2071_ _1367_ _0296_ _0071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2973_ _0127_ clknet_4_7_0_clk picorv32_pcpi_div_inst_0.quotient_msk\[26\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_56_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1924_ _1371_ _1373_ _1375_ _1376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_21_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1855_ _1326_ _0049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1786_ _1270_ _0036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2269_ _0290_ _0430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2338_ _1406_ _0493_ _0406_ _0494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2407_ _0509_ _0556_ _0557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_67_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_35_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_10_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2503__A1 _0305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2931__CLK clknet_4_14_0_clk vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1640_ _1112_ _1137_ _1141_ _0008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1571_ picorv32_pcpi_div_inst_0.dividend\[12\] _1078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_13_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2123_ _0289_ _0329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_TAPCELL_ROW_49_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2054_ picorv32_pcpi_div_inst_0.divisor\[47\] picorv32_pcpi_div_inst_0.divisor\[46\]
+ picorv32_pcpi_div_inst_0.divisor\[45\] picorv32_pcpi_div_inst_0.divisor\[44\] _0282_
+ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
X_2956_ _0110_ clknet_4_13_0_clk picorv32_pcpi_div_inst_0.quotient_msk\[9\] vdd vdd
+ vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_44_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1907_ picorv32_pcpi_div_inst_0.divisor\[29\] _1360_ _1358_ picorv32_pcpi_div_inst_0.divisor\[30\]
+ _1361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1838_ _1311_ _1308_ _1306_ _1313_ _1314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2887_ _0041_ clknet_4_3_0_clk picorv32_pcpi_div_inst_0.divisor\[3\] vdd vdd vss
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_1769_ _0948_ net1 _1256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_12_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput85 net85 pcpi_div_rd[10] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
Xoutput96 net96 pcpi_div_rd[20] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_58_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_46_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2672_ picorv32_pcpi_div_inst_0.divisor\[37\] _0780_ _0794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_26_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2741_ _0839_ _0852_ _0854_ _0183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2810_ net67 _0731_ _0891_ _0913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1554_ _0988_ _1058_ _1063_ _0031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1485_ _0997_ _0998_ _0999_ _1000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1623_ _1122_ _1125_ _1126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
.ends


magic
tech gf180mcuD
magscale 1 10
timestamp 1702206049
<< metal1 >>
rect 1344 76858 58576 76892
rect 1344 76806 19838 76858
rect 19890 76806 19942 76858
rect 19994 76806 20046 76858
rect 20098 76806 50558 76858
rect 50610 76806 50662 76858
rect 50714 76806 50766 76858
rect 50818 76806 58576 76858
rect 1344 76772 58576 76806
rect 1344 76074 58576 76108
rect 1344 76022 4478 76074
rect 4530 76022 4582 76074
rect 4634 76022 4686 76074
rect 4738 76022 35198 76074
rect 35250 76022 35302 76074
rect 35354 76022 35406 76074
rect 35458 76022 58576 76074
rect 1344 75988 58576 76022
rect 1344 75290 58576 75324
rect 1344 75238 19838 75290
rect 19890 75238 19942 75290
rect 19994 75238 20046 75290
rect 20098 75238 50558 75290
rect 50610 75238 50662 75290
rect 50714 75238 50766 75290
rect 50818 75238 58576 75290
rect 1344 75204 58576 75238
rect 1344 74506 58576 74540
rect 1344 74454 4478 74506
rect 4530 74454 4582 74506
rect 4634 74454 4686 74506
rect 4738 74454 35198 74506
rect 35250 74454 35302 74506
rect 35354 74454 35406 74506
rect 35458 74454 58576 74506
rect 1344 74420 58576 74454
rect 1344 73722 58576 73756
rect 1344 73670 19838 73722
rect 19890 73670 19942 73722
rect 19994 73670 20046 73722
rect 20098 73670 50558 73722
rect 50610 73670 50662 73722
rect 50714 73670 50766 73722
rect 50818 73670 58576 73722
rect 1344 73636 58576 73670
rect 1344 72938 58576 72972
rect 1344 72886 4478 72938
rect 4530 72886 4582 72938
rect 4634 72886 4686 72938
rect 4738 72886 35198 72938
rect 35250 72886 35302 72938
rect 35354 72886 35406 72938
rect 35458 72886 58576 72938
rect 1344 72852 58576 72886
rect 1344 72154 58576 72188
rect 1344 72102 19838 72154
rect 19890 72102 19942 72154
rect 19994 72102 20046 72154
rect 20098 72102 50558 72154
rect 50610 72102 50662 72154
rect 50714 72102 50766 72154
rect 50818 72102 58576 72154
rect 1344 72068 58576 72102
rect 40238 71986 40290 71998
rect 40238 71922 40290 71934
rect 39106 71822 39118 71874
rect 39170 71822 39182 71874
rect 39890 71710 39902 71762
rect 39954 71710 39966 71762
rect 40350 71650 40402 71662
rect 36978 71598 36990 71650
rect 37042 71598 37054 71650
rect 40350 71586 40402 71598
rect 40910 71650 40962 71662
rect 40910 71586 40962 71598
rect 41022 71538 41074 71550
rect 41022 71474 41074 71486
rect 1344 71370 58576 71404
rect 1344 71318 4478 71370
rect 4530 71318 4582 71370
rect 4634 71318 4686 71370
rect 4738 71318 35198 71370
rect 35250 71318 35302 71370
rect 35354 71318 35406 71370
rect 35458 71318 58576 71370
rect 1344 71284 58576 71318
rect 34402 71038 34414 71090
rect 34466 71038 34478 71090
rect 31602 70926 31614 70978
rect 31666 70926 31678 70978
rect 41906 70926 41918 70978
rect 41970 70926 41982 70978
rect 34862 70866 34914 70878
rect 32274 70814 32286 70866
rect 32338 70814 32350 70866
rect 37202 70814 37214 70866
rect 37266 70814 37278 70866
rect 34862 70802 34914 70814
rect 34750 70754 34802 70766
rect 34750 70690 34802 70702
rect 42702 70754 42754 70766
rect 42702 70690 42754 70702
rect 1344 70586 58576 70620
rect 1344 70534 19838 70586
rect 19890 70534 19942 70586
rect 19994 70534 20046 70586
rect 20098 70534 50558 70586
rect 50610 70534 50662 70586
rect 50714 70534 50766 70586
rect 50818 70534 58576 70586
rect 1344 70500 58576 70534
rect 31054 70418 31106 70430
rect 31054 70354 31106 70366
rect 32398 70418 32450 70430
rect 32398 70354 32450 70366
rect 40238 70418 40290 70430
rect 40238 70354 40290 70366
rect 33954 70254 33966 70306
rect 34018 70254 34030 70306
rect 41682 70254 41694 70306
rect 41746 70254 41758 70306
rect 31166 70194 31218 70206
rect 40126 70194 40178 70206
rect 27794 70142 27806 70194
rect 27858 70142 27870 70194
rect 33170 70142 33182 70194
rect 33234 70142 33246 70194
rect 36418 70142 36430 70194
rect 36482 70142 36494 70194
rect 39778 70142 39790 70194
rect 39842 70142 39854 70194
rect 31166 70130 31218 70142
rect 40126 70130 40178 70142
rect 40350 70194 40402 70206
rect 40898 70142 40910 70194
rect 40962 70142 40974 70194
rect 40350 70130 40402 70142
rect 23998 70082 24050 70094
rect 23998 70018 24050 70030
rect 25454 70082 25506 70094
rect 25454 70018 25506 70030
rect 25790 70082 25842 70094
rect 32510 70082 32562 70094
rect 28578 70030 28590 70082
rect 28642 70030 28654 70082
rect 30706 70030 30718 70082
rect 30770 70030 30782 70082
rect 36082 70030 36094 70082
rect 36146 70030 36158 70082
rect 37202 70030 37214 70082
rect 37266 70030 37278 70082
rect 39330 70030 39342 70082
rect 39394 70030 39406 70082
rect 43810 70030 43822 70082
rect 43874 70030 43886 70082
rect 25790 70018 25842 70030
rect 32510 70018 32562 70030
rect 23886 69970 23938 69982
rect 23886 69906 23938 69918
rect 25902 69970 25954 69982
rect 25902 69906 25954 69918
rect 1344 69802 58576 69836
rect 1344 69750 4478 69802
rect 4530 69750 4582 69802
rect 4634 69750 4686 69802
rect 4738 69750 35198 69802
rect 35250 69750 35302 69802
rect 35354 69750 35406 69802
rect 35458 69750 58576 69802
rect 1344 69716 58576 69750
rect 31278 69634 31330 69646
rect 31278 69570 31330 69582
rect 35646 69634 35698 69646
rect 35646 69570 35698 69582
rect 36430 69634 36482 69646
rect 36430 69570 36482 69582
rect 32958 69522 33010 69534
rect 22866 69470 22878 69522
rect 22930 69470 22942 69522
rect 24994 69470 25006 69522
rect 25058 69470 25070 69522
rect 26114 69470 26126 69522
rect 26178 69470 26190 69522
rect 28242 69470 28254 69522
rect 28306 69470 28318 69522
rect 30930 69470 30942 69522
rect 30994 69470 31006 69522
rect 32958 69458 33010 69470
rect 34302 69522 34354 69534
rect 34302 69458 34354 69470
rect 38446 69522 38498 69534
rect 42578 69470 42590 69522
rect 42642 69470 42654 69522
rect 38446 69458 38498 69470
rect 30382 69410 30434 69422
rect 34414 69410 34466 69422
rect 22194 69358 22206 69410
rect 22258 69358 22270 69410
rect 25330 69358 25342 69410
rect 25394 69358 25406 69410
rect 33394 69358 33406 69410
rect 33458 69358 33470 69410
rect 30382 69346 30434 69358
rect 34414 69346 34466 69358
rect 35310 69410 35362 69422
rect 39666 69358 39678 69410
rect 39730 69358 39742 69410
rect 35310 69346 35362 69358
rect 29038 69298 29090 69310
rect 29038 69234 29090 69246
rect 29374 69298 29426 69310
rect 29374 69234 29426 69246
rect 30606 69298 30658 69310
rect 30606 69234 30658 69246
rect 31390 69298 31442 69310
rect 31390 69234 31442 69246
rect 31838 69298 31890 69310
rect 31838 69234 31890 69246
rect 34974 69298 35026 69310
rect 34974 69234 35026 69246
rect 35534 69298 35586 69310
rect 35534 69234 35586 69246
rect 36318 69298 36370 69310
rect 36318 69234 36370 69246
rect 37550 69298 37602 69310
rect 37550 69234 37602 69246
rect 39230 69298 39282 69310
rect 39230 69234 39282 69246
rect 39342 69298 39394 69310
rect 43710 69298 43762 69310
rect 40450 69246 40462 69298
rect 40514 69246 40526 69298
rect 39342 69234 39394 69246
rect 43710 69234 43762 69246
rect 45278 69298 45330 69310
rect 45278 69234 45330 69246
rect 29262 69186 29314 69198
rect 29262 69122 29314 69134
rect 29710 69186 29762 69198
rect 29710 69122 29762 69134
rect 29822 69186 29874 69198
rect 29822 69122 29874 69134
rect 29934 69186 29986 69198
rect 29934 69122 29986 69134
rect 30830 69186 30882 69198
rect 30830 69122 30882 69134
rect 31054 69186 31106 69198
rect 31054 69122 31106 69134
rect 31614 69186 31666 69198
rect 31614 69122 31666 69134
rect 32846 69186 32898 69198
rect 32846 69122 32898 69134
rect 33070 69186 33122 69198
rect 33070 69122 33122 69134
rect 33966 69186 34018 69198
rect 33966 69122 34018 69134
rect 34190 69186 34242 69198
rect 34190 69122 34242 69134
rect 34638 69186 34690 69198
rect 34638 69122 34690 69134
rect 34750 69186 34802 69198
rect 34750 69122 34802 69134
rect 35646 69186 35698 69198
rect 35646 69122 35698 69134
rect 37214 69186 37266 69198
rect 37214 69122 37266 69134
rect 37438 69186 37490 69198
rect 37438 69122 37490 69134
rect 37662 69186 37714 69198
rect 37662 69122 37714 69134
rect 38110 69186 38162 69198
rect 38110 69122 38162 69134
rect 38334 69186 38386 69198
rect 38334 69122 38386 69134
rect 38558 69186 38610 69198
rect 38558 69122 38610 69134
rect 42926 69186 42978 69198
rect 43598 69186 43650 69198
rect 43250 69134 43262 69186
rect 43314 69134 43326 69186
rect 42926 69122 42978 69134
rect 43598 69122 43650 69134
rect 44158 69186 44210 69198
rect 44158 69122 44210 69134
rect 45390 69186 45442 69198
rect 45390 69122 45442 69134
rect 1344 69018 58576 69052
rect 1344 68966 19838 69018
rect 19890 68966 19942 69018
rect 19994 68966 20046 69018
rect 20098 68966 50558 69018
rect 50610 68966 50662 69018
rect 50714 68966 50766 69018
rect 50818 68966 58576 69018
rect 1344 68932 58576 68966
rect 24558 68850 24610 68862
rect 24558 68786 24610 68798
rect 24670 68850 24722 68862
rect 24670 68786 24722 68798
rect 33294 68850 33346 68862
rect 33294 68786 33346 68798
rect 33518 68850 33570 68862
rect 33518 68786 33570 68798
rect 37326 68850 37378 68862
rect 37326 68786 37378 68798
rect 38110 68850 38162 68862
rect 38110 68786 38162 68798
rect 38222 68850 38274 68862
rect 38222 68786 38274 68798
rect 41358 68850 41410 68862
rect 41358 68786 41410 68798
rect 41470 68850 41522 68862
rect 41470 68786 41522 68798
rect 23774 68738 23826 68750
rect 35982 68738 36034 68750
rect 27794 68686 27806 68738
rect 27858 68686 27870 68738
rect 34402 68686 34414 68738
rect 34466 68686 34478 68738
rect 23774 68674 23826 68686
rect 35982 68674 36034 68686
rect 36430 68738 36482 68750
rect 36430 68674 36482 68686
rect 36654 68738 36706 68750
rect 39230 68738 39282 68750
rect 38770 68686 38782 68738
rect 38834 68686 38846 68738
rect 36654 68674 36706 68686
rect 39230 68674 39282 68686
rect 40350 68738 40402 68750
rect 40350 68674 40402 68686
rect 41246 68738 41298 68750
rect 42354 68686 42366 68738
rect 42418 68686 42430 68738
rect 41246 68674 41298 68686
rect 23998 68626 24050 68638
rect 22754 68574 22766 68626
rect 22818 68574 22830 68626
rect 23314 68574 23326 68626
rect 23378 68574 23390 68626
rect 23538 68574 23550 68626
rect 23602 68574 23614 68626
rect 23998 68562 24050 68574
rect 24446 68626 24498 68638
rect 32958 68626 33010 68638
rect 25442 68574 25454 68626
rect 25506 68574 25518 68626
rect 24446 68562 24498 68574
rect 32958 68562 33010 68574
rect 34750 68626 34802 68638
rect 34750 68562 34802 68574
rect 35646 68626 35698 68638
rect 35646 68562 35698 68574
rect 36318 68626 36370 68638
rect 36318 68562 36370 68574
rect 36766 68626 36818 68638
rect 37550 68626 37602 68638
rect 39118 68626 39170 68638
rect 37090 68574 37102 68626
rect 37154 68574 37166 68626
rect 37874 68574 37886 68626
rect 37938 68574 37950 68626
rect 38546 68574 38558 68626
rect 38610 68574 38622 68626
rect 36766 68562 36818 68574
rect 37550 68562 37602 68574
rect 39118 68562 39170 68574
rect 39454 68626 39506 68638
rect 39454 68562 39506 68574
rect 39790 68626 39842 68638
rect 40114 68574 40126 68626
rect 40178 68574 40190 68626
rect 40898 68574 40910 68626
rect 40962 68574 40974 68626
rect 45826 68574 45838 68626
rect 45890 68574 45902 68626
rect 39790 68562 39842 68574
rect 23886 68514 23938 68526
rect 35310 68514 35362 68526
rect 40014 68514 40066 68526
rect 19842 68462 19854 68514
rect 19906 68462 19918 68514
rect 21970 68462 21982 68514
rect 22034 68462 22046 68514
rect 33394 68462 33406 68514
rect 33458 68462 33470 68514
rect 37202 68462 37214 68514
rect 37266 68462 37278 68514
rect 23886 68450 23938 68462
rect 35310 68450 35362 68462
rect 40014 68450 40066 68462
rect 1344 68234 58576 68268
rect 1344 68182 4478 68234
rect 4530 68182 4582 68234
rect 4634 68182 4686 68234
rect 4738 68182 35198 68234
rect 35250 68182 35302 68234
rect 35354 68182 35406 68234
rect 35458 68182 58576 68234
rect 1344 68148 58576 68182
rect 21422 68066 21474 68078
rect 21422 68002 21474 68014
rect 37438 68066 37490 68078
rect 37438 68002 37490 68014
rect 40910 68066 40962 68078
rect 40910 68002 40962 68014
rect 20750 67954 20802 67966
rect 20750 67890 20802 67902
rect 24782 67954 24834 67966
rect 24782 67890 24834 67902
rect 25678 67954 25730 67966
rect 25678 67890 25730 67902
rect 29150 67954 29202 67966
rect 29150 67890 29202 67902
rect 29262 67954 29314 67966
rect 30370 67902 30382 67954
rect 30434 67902 30446 67954
rect 32498 67902 32510 67954
rect 32562 67902 32574 67954
rect 41346 67902 41358 67954
rect 41410 67902 41422 67954
rect 43474 67902 43486 67954
rect 43538 67902 43550 67954
rect 44818 67902 44830 67954
rect 44882 67902 44894 67954
rect 46946 67902 46958 67954
rect 47010 67902 47022 67954
rect 29262 67890 29314 67902
rect 21870 67842 21922 67854
rect 21870 67778 21922 67790
rect 22542 67842 22594 67854
rect 23438 67842 23490 67854
rect 22866 67790 22878 67842
rect 22930 67790 22942 67842
rect 22542 67778 22594 67790
rect 23438 67778 23490 67790
rect 25118 67842 25170 67854
rect 25118 67778 25170 67790
rect 26126 67842 26178 67854
rect 26126 67778 26178 67790
rect 28030 67842 28082 67854
rect 28030 67778 28082 67790
rect 28254 67842 28306 67854
rect 37550 67842 37602 67854
rect 29698 67790 29710 67842
rect 29762 67790 29774 67842
rect 40786 67790 40798 67842
rect 40850 67790 40862 67842
rect 44146 67790 44158 67842
rect 44210 67790 44222 67842
rect 47618 67790 47630 67842
rect 47682 67790 47694 67842
rect 28254 67778 28306 67790
rect 37550 67778 37602 67790
rect 21310 67730 21362 67742
rect 21310 67666 21362 67678
rect 21982 67730 22034 67742
rect 21982 67666 22034 67678
rect 24894 67730 24946 67742
rect 37438 67730 37490 67742
rect 41022 67730 41074 67742
rect 36194 67678 36206 67730
rect 36258 67678 36270 67730
rect 38434 67678 38446 67730
rect 38498 67678 38510 67730
rect 24894 67666 24946 67678
rect 37438 67666 37490 67678
rect 41022 67666 41074 67678
rect 22094 67618 22146 67630
rect 22094 67554 22146 67566
rect 23102 67618 23154 67630
rect 24446 67618 24498 67630
rect 23762 67566 23774 67618
rect 23826 67566 23838 67618
rect 23102 67554 23154 67566
rect 24446 67554 24498 67566
rect 24670 67618 24722 67630
rect 24670 67554 24722 67566
rect 25566 67618 25618 67630
rect 25566 67554 25618 67566
rect 25790 67618 25842 67630
rect 25790 67554 25842 67566
rect 26238 67618 26290 67630
rect 26238 67554 26290 67566
rect 26462 67618 26514 67630
rect 33406 67618 33458 67630
rect 28578 67566 28590 67618
rect 28642 67566 28654 67618
rect 33058 67566 33070 67618
rect 33122 67566 33134 67618
rect 26462 67554 26514 67566
rect 33406 67554 33458 67566
rect 35646 67618 35698 67630
rect 35646 67554 35698 67566
rect 35870 67618 35922 67630
rect 35870 67554 35922 67566
rect 38110 67618 38162 67630
rect 38110 67554 38162 67566
rect 38782 67618 38834 67630
rect 38782 67554 38834 67566
rect 40238 67618 40290 67630
rect 40238 67554 40290 67566
rect 40574 67618 40626 67630
rect 40574 67554 40626 67566
rect 1344 67450 58576 67484
rect 1344 67398 19838 67450
rect 19890 67398 19942 67450
rect 19994 67398 20046 67450
rect 20098 67398 50558 67450
rect 50610 67398 50662 67450
rect 50714 67398 50766 67450
rect 50818 67398 58576 67450
rect 1344 67364 58576 67398
rect 21982 67282 22034 67294
rect 20514 67230 20526 67282
rect 20578 67230 20590 67282
rect 21982 67218 22034 67230
rect 22542 67282 22594 67294
rect 22542 67218 22594 67230
rect 22878 67282 22930 67294
rect 22878 67218 22930 67230
rect 29262 67282 29314 67294
rect 29262 67218 29314 67230
rect 39678 67282 39730 67294
rect 39678 67218 39730 67230
rect 21310 67170 21362 67182
rect 21310 67106 21362 67118
rect 22654 67170 22706 67182
rect 22654 67106 22706 67118
rect 23550 67170 23602 67182
rect 23550 67106 23602 67118
rect 23998 67170 24050 67182
rect 23998 67106 24050 67118
rect 24222 67170 24274 67182
rect 24222 67106 24274 67118
rect 29150 67170 29202 67182
rect 29150 67106 29202 67118
rect 29486 67170 29538 67182
rect 30382 67170 30434 67182
rect 29698 67118 29710 67170
rect 29762 67118 29774 67170
rect 29486 67106 29538 67118
rect 30382 67106 30434 67118
rect 30494 67170 30546 67182
rect 32062 67170 32114 67182
rect 31266 67118 31278 67170
rect 31330 67118 31342 67170
rect 30494 67106 30546 67118
rect 32062 67106 32114 67118
rect 41470 67170 41522 67182
rect 42478 67170 42530 67182
rect 41794 67118 41806 67170
rect 41858 67118 41870 67170
rect 41470 67106 41522 67118
rect 42478 67106 42530 67118
rect 43262 67170 43314 67182
rect 43262 67106 43314 67118
rect 43486 67170 43538 67182
rect 43486 67106 43538 67118
rect 44494 67170 44546 67182
rect 44494 67106 44546 67118
rect 45502 67170 45554 67182
rect 45502 67106 45554 67118
rect 21086 67058 21138 67070
rect 20290 67006 20302 67058
rect 20354 67006 20366 67058
rect 21086 66994 21138 67006
rect 21422 67058 21474 67070
rect 21422 66994 21474 67006
rect 21758 67058 21810 67070
rect 24334 67058 24386 67070
rect 22306 67006 22318 67058
rect 22370 67006 22382 67058
rect 23090 67006 23102 67058
rect 23154 67006 23166 67058
rect 21758 66994 21810 67006
rect 24334 66994 24386 67006
rect 30046 67058 30098 67070
rect 30046 66994 30098 67006
rect 30606 67058 30658 67070
rect 41134 67058 41186 67070
rect 43038 67058 43090 67070
rect 30930 67006 30942 67058
rect 30994 67006 31006 67058
rect 31490 67006 31502 67058
rect 31554 67006 31566 67058
rect 42018 67006 42030 67058
rect 42082 67006 42094 67058
rect 42690 67006 42702 67058
rect 42754 67006 42766 67058
rect 30606 66994 30658 67006
rect 41134 66994 41186 67006
rect 43038 66994 43090 67006
rect 43934 67058 43986 67070
rect 43934 66994 43986 67006
rect 44046 67058 44098 67070
rect 44046 66994 44098 67006
rect 44718 67058 44770 67070
rect 44718 66994 44770 67006
rect 44942 67058 44994 67070
rect 44942 66994 44994 67006
rect 45390 67058 45442 67070
rect 45390 66994 45442 67006
rect 45614 67058 45666 67070
rect 45614 66994 45666 67006
rect 15374 66946 15426 66958
rect 15374 66882 15426 66894
rect 19854 66946 19906 66958
rect 19854 66882 19906 66894
rect 21870 66946 21922 66958
rect 21870 66882 21922 66894
rect 25678 66946 25730 66958
rect 25678 66882 25730 66894
rect 26126 66946 26178 66958
rect 26126 66882 26178 66894
rect 26462 66946 26514 66958
rect 26462 66882 26514 66894
rect 27022 66946 27074 66958
rect 27022 66882 27074 66894
rect 28702 66946 28754 66958
rect 28702 66882 28754 66894
rect 34414 66946 34466 66958
rect 34414 66882 34466 66894
rect 36766 66946 36818 66958
rect 36766 66882 36818 66894
rect 40238 66946 40290 66958
rect 40238 66882 40290 66894
rect 42814 66946 42866 66958
rect 42814 66882 42866 66894
rect 43374 66946 43426 66958
rect 43374 66882 43426 66894
rect 44606 66946 44658 66958
rect 44606 66882 44658 66894
rect 15262 66834 15314 66846
rect 25666 66782 25678 66834
rect 25730 66831 25742 66834
rect 26450 66831 26462 66834
rect 25730 66785 26462 66831
rect 25730 66782 25742 66785
rect 26450 66782 26462 66785
rect 26514 66782 26526 66834
rect 15262 66770 15314 66782
rect 1344 66666 58576 66700
rect 1344 66614 4478 66666
rect 4530 66614 4582 66666
rect 4634 66614 4686 66666
rect 4738 66614 35198 66666
rect 35250 66614 35302 66666
rect 35354 66614 35406 66666
rect 35458 66614 58576 66666
rect 1344 66580 58576 66614
rect 14030 66498 14082 66510
rect 14030 66434 14082 66446
rect 22318 66498 22370 66510
rect 22318 66434 22370 66446
rect 26126 66498 26178 66510
rect 26126 66434 26178 66446
rect 31054 66498 31106 66510
rect 31054 66434 31106 66446
rect 41134 66498 41186 66510
rect 41134 66434 41186 66446
rect 43374 66498 43426 66510
rect 43374 66434 43426 66446
rect 43934 66498 43986 66510
rect 43934 66434 43986 66446
rect 21422 66386 21474 66398
rect 17378 66334 17390 66386
rect 17442 66334 17454 66386
rect 21422 66322 21474 66334
rect 25566 66386 25618 66398
rect 25566 66322 25618 66334
rect 34526 66386 34578 66398
rect 48066 66334 48078 66386
rect 48130 66334 48142 66386
rect 34526 66322 34578 66334
rect 21646 66274 21698 66286
rect 25790 66274 25842 66286
rect 14466 66222 14478 66274
rect 14530 66222 14542 66274
rect 19954 66222 19966 66274
rect 20018 66222 20030 66274
rect 21970 66222 21982 66274
rect 22034 66222 22046 66274
rect 21646 66210 21698 66222
rect 25790 66210 25842 66222
rect 26238 66274 26290 66286
rect 26238 66210 26290 66222
rect 27806 66274 27858 66286
rect 27806 66210 27858 66222
rect 28142 66274 28194 66286
rect 28142 66210 28194 66222
rect 35198 66274 35250 66286
rect 35198 66210 35250 66222
rect 35422 66274 35474 66286
rect 35422 66210 35474 66222
rect 37326 66274 37378 66286
rect 37326 66210 37378 66222
rect 37662 66274 37714 66286
rect 37662 66210 37714 66222
rect 38670 66274 38722 66286
rect 38670 66210 38722 66222
rect 41246 66274 41298 66286
rect 41246 66210 41298 66222
rect 41582 66274 41634 66286
rect 42702 66274 42754 66286
rect 42242 66222 42254 66274
rect 42306 66222 42318 66274
rect 41582 66210 41634 66222
rect 42702 66210 42754 66222
rect 44158 66274 44210 66286
rect 45154 66222 45166 66274
rect 45218 66222 45230 66274
rect 44158 66210 44210 66222
rect 13918 66162 13970 66174
rect 24670 66162 24722 66174
rect 15250 66110 15262 66162
rect 15314 66110 15326 66162
rect 13918 66098 13970 66110
rect 24670 66098 24722 66110
rect 25454 66162 25506 66174
rect 25454 66098 25506 66110
rect 26126 66162 26178 66174
rect 26126 66098 26178 66110
rect 28366 66162 28418 66174
rect 28366 66098 28418 66110
rect 30270 66162 30322 66174
rect 30270 66098 30322 66110
rect 30606 66162 30658 66174
rect 30606 66098 30658 66110
rect 30942 66162 30994 66174
rect 30942 66098 30994 66110
rect 31054 66162 31106 66174
rect 31054 66098 31106 66110
rect 33630 66162 33682 66174
rect 33630 66098 33682 66110
rect 34078 66162 34130 66174
rect 34078 66098 34130 66110
rect 36206 66162 36258 66174
rect 36206 66098 36258 66110
rect 36430 66162 36482 66174
rect 36430 66098 36482 66110
rect 36990 66162 37042 66174
rect 36990 66098 37042 66110
rect 39902 66162 39954 66174
rect 39902 66098 39954 66110
rect 41918 66162 41970 66174
rect 43262 66162 43314 66174
rect 42466 66110 42478 66162
rect 42530 66110 42542 66162
rect 41918 66098 41970 66110
rect 43262 66098 43314 66110
rect 43598 66162 43650 66174
rect 45938 66110 45950 66162
rect 46002 66110 46014 66162
rect 43598 66098 43650 66110
rect 14030 66050 14082 66062
rect 20638 66050 20690 66062
rect 20178 65998 20190 66050
rect 20242 65998 20254 66050
rect 14030 65986 14082 65998
rect 20638 65986 20690 65998
rect 21310 66050 21362 66062
rect 21310 65986 21362 65998
rect 22206 66050 22258 66062
rect 22206 65986 22258 65998
rect 24446 66050 24498 66062
rect 24446 65986 24498 65998
rect 24782 66050 24834 66062
rect 24782 65986 24834 65998
rect 25006 66050 25058 66062
rect 25006 65986 25058 65998
rect 25230 66050 25282 66062
rect 25230 65986 25282 65998
rect 27022 66050 27074 66062
rect 27022 65986 27074 65998
rect 27246 66050 27298 66062
rect 27246 65986 27298 65998
rect 27358 66050 27410 66062
rect 27358 65986 27410 65998
rect 27470 66050 27522 66062
rect 27470 65986 27522 65998
rect 27918 66050 27970 66062
rect 27918 65986 27970 65998
rect 29374 66050 29426 66062
rect 29374 65986 29426 65998
rect 30046 66050 30098 66062
rect 30046 65986 30098 65998
rect 32734 66050 32786 66062
rect 32734 65986 32786 65998
rect 33294 66050 33346 66062
rect 33294 65986 33346 65998
rect 33518 66050 33570 66062
rect 33518 65986 33570 65998
rect 33966 66050 34018 66062
rect 36318 66050 36370 66062
rect 35746 65998 35758 66050
rect 35810 65998 35822 66050
rect 33966 65986 34018 65998
rect 36318 65986 36370 65998
rect 37326 66050 37378 66062
rect 37326 65986 37378 65998
rect 39118 66050 39170 66062
rect 39118 65986 39170 65998
rect 39230 66050 39282 66062
rect 39230 65986 39282 65998
rect 39342 66050 39394 66062
rect 39342 65986 39394 65998
rect 39566 66050 39618 66062
rect 39566 65986 39618 65998
rect 39790 66050 39842 66062
rect 39790 65986 39842 65998
rect 40350 66050 40402 66062
rect 40350 65986 40402 65998
rect 41134 66050 41186 66062
rect 41134 65986 41186 65998
rect 41694 66050 41746 66062
rect 41694 65986 41746 65998
rect 43038 66050 43090 66062
rect 43038 65986 43090 65998
rect 43822 66050 43874 66062
rect 43822 65986 43874 65998
rect 1344 65882 58576 65916
rect 1344 65830 19838 65882
rect 19890 65830 19942 65882
rect 19994 65830 20046 65882
rect 20098 65830 50558 65882
rect 50610 65830 50662 65882
rect 50714 65830 50766 65882
rect 50818 65830 58576 65882
rect 1344 65796 58576 65830
rect 16382 65714 16434 65726
rect 16382 65650 16434 65662
rect 25790 65714 25842 65726
rect 25790 65650 25842 65662
rect 43598 65714 43650 65726
rect 43598 65650 43650 65662
rect 43822 65714 43874 65726
rect 43822 65650 43874 65662
rect 44158 65714 44210 65726
rect 44158 65650 44210 65662
rect 44382 65714 44434 65726
rect 44382 65650 44434 65662
rect 45390 65714 45442 65726
rect 45390 65650 45442 65662
rect 16494 65602 16546 65614
rect 16494 65538 16546 65550
rect 18510 65602 18562 65614
rect 24222 65602 24274 65614
rect 30270 65602 30322 65614
rect 20738 65550 20750 65602
rect 20802 65550 20814 65602
rect 23202 65550 23214 65602
rect 23266 65550 23278 65602
rect 27346 65550 27358 65602
rect 27410 65550 27422 65602
rect 18510 65538 18562 65550
rect 24222 65538 24274 65550
rect 30270 65538 30322 65550
rect 32174 65602 32226 65614
rect 32174 65538 32226 65550
rect 34190 65602 34242 65614
rect 34190 65538 34242 65550
rect 43934 65602 43986 65614
rect 43934 65538 43986 65550
rect 44494 65602 44546 65614
rect 44494 65538 44546 65550
rect 45278 65602 45330 65614
rect 47506 65550 47518 65602
rect 47570 65550 47582 65602
rect 45278 65538 45330 65550
rect 16158 65490 16210 65502
rect 17614 65490 17666 65502
rect 9874 65438 9886 65490
rect 9938 65438 9950 65490
rect 13122 65438 13134 65490
rect 13186 65438 13198 65490
rect 17378 65438 17390 65490
rect 17442 65438 17454 65490
rect 16158 65426 16210 65438
rect 17614 65426 17666 65438
rect 17726 65490 17778 65502
rect 17726 65426 17778 65438
rect 17838 65490 17890 65502
rect 18398 65490 18450 65502
rect 25566 65490 25618 65502
rect 30046 65490 30098 65502
rect 18050 65438 18062 65490
rect 18114 65438 18126 65490
rect 19954 65438 19966 65490
rect 20018 65438 20030 65490
rect 23426 65438 23438 65490
rect 23490 65438 23502 65490
rect 24434 65438 24446 65490
rect 24498 65438 24510 65490
rect 25218 65438 25230 65490
rect 25282 65438 25294 65490
rect 26562 65438 26574 65490
rect 26626 65438 26638 65490
rect 17838 65426 17890 65438
rect 18398 65426 18450 65438
rect 25566 65426 25618 65438
rect 30046 65426 30098 65438
rect 30158 65490 30210 65502
rect 30158 65426 30210 65438
rect 30718 65490 30770 65502
rect 30718 65426 30770 65438
rect 31950 65490 32002 65502
rect 31950 65426 32002 65438
rect 32510 65490 32562 65502
rect 32510 65426 32562 65438
rect 32958 65490 33010 65502
rect 32958 65426 33010 65438
rect 33406 65490 33458 65502
rect 33406 65426 33458 65438
rect 33630 65490 33682 65502
rect 33630 65426 33682 65438
rect 33966 65490 34018 65502
rect 47854 65490 47906 65502
rect 34514 65438 34526 65490
rect 34578 65438 34590 65490
rect 40226 65438 40238 65490
rect 40290 65438 40302 65490
rect 41234 65438 41246 65490
rect 41298 65438 41310 65490
rect 33966 65426 34018 65438
rect 47854 65426 47906 65438
rect 25678 65378 25730 65390
rect 10546 65326 10558 65378
rect 10610 65326 10622 65378
rect 12674 65326 12686 65378
rect 12738 65326 12750 65378
rect 13794 65326 13806 65378
rect 13858 65326 13870 65378
rect 15922 65326 15934 65378
rect 15986 65326 15998 65378
rect 22866 65326 22878 65378
rect 22930 65326 22942 65378
rect 25678 65314 25730 65326
rect 26126 65378 26178 65390
rect 26126 65314 26178 65326
rect 26238 65378 26290 65390
rect 26238 65314 26290 65326
rect 29486 65378 29538 65390
rect 29486 65314 29538 65326
rect 33518 65378 33570 65390
rect 33518 65314 33570 65326
rect 34078 65378 34130 65390
rect 41022 65378 41074 65390
rect 37426 65326 37438 65378
rect 37490 65326 37502 65378
rect 34078 65314 34130 65326
rect 41022 65314 41074 65326
rect 41806 65378 41858 65390
rect 41806 65314 41858 65326
rect 42142 65378 42194 65390
rect 42142 65314 42194 65326
rect 42590 65378 42642 65390
rect 42590 65314 42642 65326
rect 43038 65378 43090 65390
rect 43038 65314 43090 65326
rect 40910 65266 40962 65278
rect 41458 65214 41470 65266
rect 41522 65263 41534 65266
rect 41794 65263 41806 65266
rect 41522 65217 41806 65263
rect 41522 65214 41534 65217
rect 41794 65214 41806 65217
rect 41858 65214 41870 65266
rect 42354 65214 42366 65266
rect 42418 65263 42430 65266
rect 42578 65263 42590 65266
rect 42418 65217 42590 65263
rect 42418 65214 42430 65217
rect 42578 65214 42590 65217
rect 42642 65214 42654 65266
rect 40910 65202 40962 65214
rect 1344 65098 58576 65132
rect 1344 65046 4478 65098
rect 4530 65046 4582 65098
rect 4634 65046 4686 65098
rect 4738 65046 35198 65098
rect 35250 65046 35302 65098
rect 35354 65046 35406 65098
rect 35458 65046 58576 65098
rect 1344 65012 58576 65046
rect 26574 64930 26626 64942
rect 34974 64930 35026 64942
rect 26898 64878 26910 64930
rect 26962 64878 26974 64930
rect 29922 64878 29934 64930
rect 29986 64927 29998 64930
rect 30930 64927 30942 64930
rect 29986 64881 30942 64927
rect 29986 64878 29998 64881
rect 30930 64878 30942 64881
rect 30994 64878 31006 64930
rect 36418 64878 36430 64930
rect 36482 64878 36494 64930
rect 41682 64878 41694 64930
rect 41746 64878 41758 64930
rect 43026 64878 43038 64930
rect 43090 64927 43102 64930
rect 43586 64927 43598 64930
rect 43090 64881 43598 64927
rect 43090 64878 43102 64881
rect 43586 64878 43598 64881
rect 43650 64878 43662 64930
rect 26574 64866 26626 64878
rect 34974 64866 35026 64878
rect 13918 64818 13970 64830
rect 12898 64766 12910 64818
rect 12962 64766 12974 64818
rect 17490 64766 17502 64818
rect 17554 64766 17566 64818
rect 20738 64766 20750 64818
rect 20802 64766 20814 64818
rect 23762 64766 23774 64818
rect 23826 64766 23838 64818
rect 25890 64766 25902 64818
rect 25954 64766 25966 64818
rect 31938 64766 31950 64818
rect 32002 64766 32014 64818
rect 34066 64766 34078 64818
rect 34130 64766 34142 64818
rect 13918 64754 13970 64766
rect 13694 64706 13746 64718
rect 21646 64706 21698 64718
rect 27246 64706 27298 64718
rect 10098 64654 10110 64706
rect 10162 64654 10174 64706
rect 14242 64654 14254 64706
rect 14306 64654 14318 64706
rect 14578 64654 14590 64706
rect 14642 64654 14654 64706
rect 17938 64654 17950 64706
rect 18002 64654 18014 64706
rect 22978 64654 22990 64706
rect 23042 64654 23054 64706
rect 13694 64642 13746 64654
rect 21646 64642 21698 64654
rect 27246 64642 27298 64654
rect 27470 64706 27522 64718
rect 28030 64706 28082 64718
rect 27794 64654 27806 64706
rect 27858 64654 27870 64706
rect 27470 64642 27522 64654
rect 28030 64642 28082 64654
rect 29374 64706 29426 64718
rect 29374 64642 29426 64654
rect 29822 64706 29874 64718
rect 34638 64706 34690 64718
rect 31154 64654 31166 64706
rect 31218 64654 31230 64706
rect 29822 64642 29874 64654
rect 34638 64642 34690 64654
rect 35758 64706 35810 64718
rect 35758 64642 35810 64654
rect 35870 64706 35922 64718
rect 41134 64706 41186 64718
rect 37426 64654 37438 64706
rect 37490 64654 37502 64706
rect 35870 64642 35922 64654
rect 41134 64642 41186 64654
rect 42030 64706 42082 64718
rect 42030 64642 42082 64654
rect 42702 64706 42754 64718
rect 42702 64642 42754 64654
rect 44718 64706 44770 64718
rect 44718 64642 44770 64654
rect 45166 64706 45218 64718
rect 45166 64642 45218 64654
rect 21310 64594 21362 64606
rect 10770 64542 10782 64594
rect 10834 64542 10846 64594
rect 15362 64542 15374 64594
rect 15426 64542 15438 64594
rect 18610 64542 18622 64594
rect 18674 64542 18686 64594
rect 21310 64530 21362 64542
rect 21422 64594 21474 64606
rect 21422 64530 21474 64542
rect 28142 64594 28194 64606
rect 29150 64594 29202 64606
rect 28578 64542 28590 64594
rect 28642 64542 28654 64594
rect 28142 64530 28194 64542
rect 29150 64530 29202 64542
rect 34414 64594 34466 64606
rect 34414 64530 34466 64542
rect 35982 64594 36034 64606
rect 35982 64530 36034 64542
rect 37214 64594 37266 64606
rect 41022 64594 41074 64606
rect 38210 64542 38222 64594
rect 38274 64542 38286 64594
rect 37214 64530 37266 64542
rect 41022 64530 41074 64542
rect 41246 64594 41298 64606
rect 41246 64530 41298 64542
rect 42254 64594 42306 64606
rect 42254 64530 42306 64542
rect 43038 64594 43090 64606
rect 43038 64530 43090 64542
rect 44046 64594 44098 64606
rect 44046 64530 44098 64542
rect 13806 64482 13858 64494
rect 13806 64418 13858 64430
rect 14030 64482 14082 64494
rect 14030 64418 14082 64430
rect 22766 64482 22818 64494
rect 22766 64418 22818 64430
rect 26350 64482 26402 64494
rect 26350 64418 26402 64430
rect 26462 64482 26514 64494
rect 26462 64418 26514 64430
rect 29598 64482 29650 64494
rect 29598 64418 29650 64430
rect 30158 64482 30210 64494
rect 30158 64418 30210 64430
rect 30606 64482 30658 64494
rect 42478 64482 42530 64494
rect 40450 64430 40462 64482
rect 40514 64430 40526 64482
rect 30606 64418 30658 64430
rect 42478 64418 42530 64430
rect 43598 64482 43650 64494
rect 43598 64418 43650 64430
rect 43934 64482 43986 64494
rect 43934 64418 43986 64430
rect 45278 64482 45330 64494
rect 45278 64418 45330 64430
rect 45390 64482 45442 64494
rect 45390 64418 45442 64430
rect 45950 64482 46002 64494
rect 45950 64418 46002 64430
rect 46846 64482 46898 64494
rect 46846 64418 46898 64430
rect 1344 64314 58576 64348
rect 1344 64262 19838 64314
rect 19890 64262 19942 64314
rect 19994 64262 20046 64314
rect 20098 64262 50558 64314
rect 50610 64262 50662 64314
rect 50714 64262 50766 64314
rect 50818 64262 58576 64314
rect 1344 64228 58576 64262
rect 11678 64146 11730 64158
rect 11678 64082 11730 64094
rect 11790 64146 11842 64158
rect 11790 64082 11842 64094
rect 12798 64146 12850 64158
rect 12798 64082 12850 64094
rect 14814 64146 14866 64158
rect 14814 64082 14866 64094
rect 15598 64146 15650 64158
rect 15598 64082 15650 64094
rect 16158 64146 16210 64158
rect 16158 64082 16210 64094
rect 16270 64146 16322 64158
rect 16270 64082 16322 64094
rect 16382 64146 16434 64158
rect 16382 64082 16434 64094
rect 17950 64146 18002 64158
rect 17950 64082 18002 64094
rect 19294 64146 19346 64158
rect 19294 64082 19346 64094
rect 20302 64146 20354 64158
rect 20302 64082 20354 64094
rect 22542 64146 22594 64158
rect 26126 64146 26178 64158
rect 22978 64094 22990 64146
rect 23042 64094 23054 64146
rect 22542 64082 22594 64094
rect 26126 64082 26178 64094
rect 26574 64146 26626 64158
rect 26574 64082 26626 64094
rect 28590 64146 28642 64158
rect 28590 64082 28642 64094
rect 30382 64146 30434 64158
rect 30382 64082 30434 64094
rect 31726 64146 31778 64158
rect 31726 64082 31778 64094
rect 33518 64146 33570 64158
rect 33518 64082 33570 64094
rect 33854 64146 33906 64158
rect 33854 64082 33906 64094
rect 37774 64146 37826 64158
rect 37774 64082 37826 64094
rect 37998 64146 38050 64158
rect 37998 64082 38050 64094
rect 38670 64146 38722 64158
rect 38670 64082 38722 64094
rect 38894 64146 38946 64158
rect 41022 64146 41074 64158
rect 39554 64094 39566 64146
rect 39618 64094 39630 64146
rect 38894 64082 38946 64094
rect 41022 64082 41074 64094
rect 42478 64146 42530 64158
rect 42478 64082 42530 64094
rect 47182 64146 47234 64158
rect 47182 64082 47234 64094
rect 12462 64034 12514 64046
rect 12462 63970 12514 63982
rect 13470 64034 13522 64046
rect 13470 63970 13522 63982
rect 13918 64034 13970 64046
rect 13918 63970 13970 63982
rect 14030 64034 14082 64046
rect 14030 63970 14082 63982
rect 14926 64034 14978 64046
rect 23550 64034 23602 64046
rect 15250 63982 15262 64034
rect 15314 63982 15326 64034
rect 14926 63970 14978 63982
rect 23550 63970 23602 63982
rect 26686 64034 26738 64046
rect 26686 63970 26738 63982
rect 28814 64034 28866 64046
rect 28814 63970 28866 63982
rect 28926 64034 28978 64046
rect 28926 63970 28978 63982
rect 29374 64034 29426 64046
rect 29374 63970 29426 63982
rect 31614 64034 31666 64046
rect 31614 63970 31666 63982
rect 31950 64034 32002 64046
rect 31950 63970 32002 63982
rect 32510 64034 32562 64046
rect 32510 63970 32562 63982
rect 33630 64034 33682 64046
rect 33630 63970 33682 63982
rect 34078 64034 34130 64046
rect 34078 63970 34130 63982
rect 34190 64034 34242 64046
rect 34190 63970 34242 63982
rect 41918 64034 41970 64046
rect 41918 63970 41970 63982
rect 42590 64034 42642 64046
rect 47630 64034 47682 64046
rect 43810 63982 43822 64034
rect 43874 63982 43886 64034
rect 42590 63970 42642 63982
rect 47630 63970 47682 63982
rect 48974 64034 49026 64046
rect 48974 63970 49026 63982
rect 11454 63922 11506 63934
rect 11454 63858 11506 63870
rect 11566 63922 11618 63934
rect 12574 63922 12626 63934
rect 13358 63922 13410 63934
rect 12002 63870 12014 63922
rect 12066 63870 12078 63922
rect 13010 63870 13022 63922
rect 13074 63870 13086 63922
rect 11566 63858 11618 63870
rect 12574 63858 12626 63870
rect 13358 63858 13410 63870
rect 13694 63922 13746 63934
rect 13694 63858 13746 63870
rect 16046 63922 16098 63934
rect 17390 63922 17442 63934
rect 16594 63870 16606 63922
rect 16658 63870 16670 63922
rect 16046 63858 16098 63870
rect 17390 63858 17442 63870
rect 20190 63922 20242 63934
rect 20190 63858 20242 63870
rect 20526 63922 20578 63934
rect 20526 63858 20578 63870
rect 22318 63922 22370 63934
rect 22318 63858 22370 63870
rect 22654 63922 22706 63934
rect 22654 63858 22706 63870
rect 23774 63922 23826 63934
rect 23774 63858 23826 63870
rect 24222 63922 24274 63934
rect 24222 63858 24274 63870
rect 24446 63922 24498 63934
rect 24446 63858 24498 63870
rect 25454 63922 25506 63934
rect 25454 63858 25506 63870
rect 25902 63922 25954 63934
rect 25902 63858 25954 63870
rect 26014 63922 26066 63934
rect 26014 63858 26066 63870
rect 27694 63922 27746 63934
rect 29598 63922 29650 63934
rect 28354 63870 28366 63922
rect 28418 63870 28430 63922
rect 27694 63858 27746 63870
rect 29598 63858 29650 63870
rect 30046 63922 30098 63934
rect 33182 63922 33234 63934
rect 30482 63870 30494 63922
rect 30546 63870 30558 63922
rect 32162 63870 32174 63922
rect 32226 63870 32238 63922
rect 30046 63858 30098 63870
rect 33182 63858 33234 63870
rect 33294 63922 33346 63934
rect 39342 63922 39394 63934
rect 37426 63870 37438 63922
rect 37490 63870 37502 63922
rect 38322 63870 38334 63922
rect 38386 63870 38398 63922
rect 33294 63858 33346 63870
rect 39342 63858 39394 63870
rect 40126 63922 40178 63934
rect 40126 63858 40178 63870
rect 40798 63922 40850 63934
rect 40798 63858 40850 63870
rect 41134 63922 41186 63934
rect 41134 63858 41186 63870
rect 41358 63922 41410 63934
rect 41358 63858 41410 63870
rect 42030 63922 42082 63934
rect 42030 63858 42082 63870
rect 42254 63922 42306 63934
rect 47070 63922 47122 63934
rect 43138 63870 43150 63922
rect 43202 63870 43214 63922
rect 42254 63858 42306 63870
rect 47070 63858 47122 63870
rect 47854 63922 47906 63934
rect 47854 63858 47906 63870
rect 48302 63922 48354 63934
rect 48302 63858 48354 63870
rect 49422 63922 49474 63934
rect 49422 63858 49474 63870
rect 17502 63810 17554 63822
rect 12450 63758 12462 63810
rect 12514 63758 12526 63810
rect 17502 63746 17554 63758
rect 19406 63810 19458 63822
rect 19406 63746 19458 63758
rect 22206 63810 22258 63822
rect 22206 63746 22258 63758
rect 24334 63810 24386 63822
rect 29486 63810 29538 63822
rect 32398 63810 32450 63822
rect 37886 63810 37938 63822
rect 27570 63758 27582 63810
rect 27634 63758 27646 63810
rect 30370 63758 30382 63810
rect 30434 63758 30446 63810
rect 34514 63758 34526 63810
rect 34578 63758 34590 63810
rect 36642 63758 36654 63810
rect 36706 63758 36718 63810
rect 24334 63746 24386 63758
rect 14814 63698 14866 63710
rect 23326 63698 23378 63710
rect 21970 63646 21982 63698
rect 22034 63695 22046 63698
rect 22194 63695 22206 63698
rect 22034 63649 22206 63695
rect 22034 63646 22046 63649
rect 22194 63646 22206 63649
rect 22258 63646 22270 63698
rect 14814 63634 14866 63646
rect 23326 63634 23378 63646
rect 26574 63698 26626 63710
rect 27585 63695 27631 63758
rect 29486 63746 29538 63758
rect 32398 63746 32450 63758
rect 37886 63746 37938 63758
rect 38782 63810 38834 63822
rect 38782 63746 38834 63758
rect 39902 63810 39954 63822
rect 46398 63810 46450 63822
rect 45938 63758 45950 63810
rect 46002 63758 46014 63810
rect 39902 63746 39954 63758
rect 46398 63746 46450 63758
rect 47742 63810 47794 63822
rect 47742 63746 47794 63758
rect 28030 63698 28082 63710
rect 27794 63695 27806 63698
rect 27585 63649 27806 63695
rect 27794 63646 27806 63649
rect 27858 63646 27870 63698
rect 26574 63634 26626 63646
rect 28030 63634 28082 63646
rect 28366 63698 28418 63710
rect 28366 63634 28418 63646
rect 41918 63698 41970 63710
rect 41918 63634 41970 63646
rect 47182 63698 47234 63710
rect 47182 63634 47234 63646
rect 48862 63698 48914 63710
rect 48862 63634 48914 63646
rect 1344 63530 58576 63564
rect 1344 63478 4478 63530
rect 4530 63478 4582 63530
rect 4634 63478 4686 63530
rect 4738 63478 35198 63530
rect 35250 63478 35302 63530
rect 35354 63478 35406 63530
rect 35458 63478 58576 63530
rect 1344 63444 58576 63478
rect 12574 63362 12626 63374
rect 44382 63362 44434 63374
rect 24546 63310 24558 63362
rect 24610 63310 24622 63362
rect 12574 63298 12626 63310
rect 44382 63298 44434 63310
rect 12686 63250 12738 63262
rect 12686 63186 12738 63198
rect 19854 63250 19906 63262
rect 25118 63250 25170 63262
rect 35982 63250 36034 63262
rect 24210 63198 24222 63250
rect 24274 63198 24286 63250
rect 31154 63198 31166 63250
rect 31218 63198 31230 63250
rect 19854 63186 19906 63198
rect 25118 63186 25170 63198
rect 35982 63186 36034 63198
rect 38334 63250 38386 63262
rect 38334 63186 38386 63198
rect 38894 63250 38946 63262
rect 38894 63186 38946 63198
rect 39454 63250 39506 63262
rect 40226 63198 40238 63250
rect 40290 63198 40302 63250
rect 39454 63186 39506 63198
rect 19182 63138 19234 63150
rect 18722 63086 18734 63138
rect 18786 63086 18798 63138
rect 19182 63074 19234 63086
rect 19742 63138 19794 63150
rect 19742 63074 19794 63086
rect 21982 63138 22034 63150
rect 21982 63074 22034 63086
rect 22094 63138 22146 63150
rect 22990 63138 23042 63150
rect 24334 63138 24386 63150
rect 22754 63086 22766 63138
rect 22818 63086 22830 63138
rect 23538 63086 23550 63138
rect 23602 63086 23614 63138
rect 22094 63074 22146 63086
rect 22990 63074 23042 63086
rect 24334 63074 24386 63086
rect 25006 63138 25058 63150
rect 25006 63074 25058 63086
rect 25230 63138 25282 63150
rect 25230 63074 25282 63086
rect 25566 63138 25618 63150
rect 35870 63138 35922 63150
rect 34738 63086 34750 63138
rect 34802 63086 34814 63138
rect 25566 63074 25618 63086
rect 35870 63074 35922 63086
rect 36094 63138 36146 63150
rect 36094 63074 36146 63086
rect 37214 63138 37266 63150
rect 37214 63074 37266 63086
rect 37886 63138 37938 63150
rect 37886 63074 37938 63086
rect 38110 63138 38162 63150
rect 38110 63074 38162 63086
rect 40014 63138 40066 63150
rect 43138 63086 43150 63138
rect 43202 63086 43214 63138
rect 48738 63086 48750 63138
rect 48802 63086 48814 63138
rect 40014 63074 40066 63086
rect 11790 63026 11842 63038
rect 21646 63026 21698 63038
rect 14242 62974 14254 63026
rect 14306 62974 14318 63026
rect 11790 62962 11842 62974
rect 21646 62962 21698 62974
rect 22430 63026 22482 63038
rect 22430 62962 22482 62974
rect 23102 63026 23154 63038
rect 23102 62962 23154 62974
rect 37102 63026 37154 63038
rect 37102 62962 37154 62974
rect 38446 63026 38498 63038
rect 43822 63026 43874 63038
rect 42354 62974 42366 63026
rect 42418 62974 42430 63026
rect 45378 62974 45390 63026
rect 45442 62974 45454 63026
rect 38446 62962 38498 62974
rect 43822 62962 43874 62974
rect 11454 62914 11506 62926
rect 11454 62850 11506 62862
rect 11678 62914 11730 62926
rect 11678 62850 11730 62862
rect 19966 62914 20018 62926
rect 19966 62850 20018 62862
rect 20190 62914 20242 62926
rect 20190 62850 20242 62862
rect 22318 62914 22370 62926
rect 22318 62850 22370 62862
rect 26014 62914 26066 62926
rect 26014 62850 26066 62862
rect 28478 62914 28530 62926
rect 28478 62850 28530 62862
rect 35198 62914 35250 62926
rect 35198 62850 35250 62862
rect 35646 62914 35698 62926
rect 35646 62850 35698 62862
rect 36878 62914 36930 62926
rect 36878 62850 36930 62862
rect 39342 62914 39394 62926
rect 39342 62850 39394 62862
rect 39566 62914 39618 62926
rect 39566 62850 39618 62862
rect 44046 62914 44098 62926
rect 44046 62850 44098 62862
rect 44270 62914 44322 62926
rect 44270 62850 44322 62862
rect 1344 62746 58576 62780
rect 1344 62694 19838 62746
rect 19890 62694 19942 62746
rect 19994 62694 20046 62746
rect 20098 62694 50558 62746
rect 50610 62694 50662 62746
rect 50714 62694 50766 62746
rect 50818 62694 58576 62746
rect 1344 62660 58576 62694
rect 12686 62578 12738 62590
rect 12686 62514 12738 62526
rect 12910 62578 12962 62590
rect 12910 62514 12962 62526
rect 15822 62578 15874 62590
rect 15822 62514 15874 62526
rect 16046 62578 16098 62590
rect 16046 62514 16098 62526
rect 17950 62578 18002 62590
rect 24670 62578 24722 62590
rect 24210 62526 24222 62578
rect 24274 62575 24286 62578
rect 24546 62575 24558 62578
rect 24274 62529 24558 62575
rect 24274 62526 24286 62529
rect 24546 62526 24558 62529
rect 24610 62526 24622 62578
rect 17950 62514 18002 62526
rect 24670 62514 24722 62526
rect 33070 62578 33122 62590
rect 33070 62514 33122 62526
rect 33294 62578 33346 62590
rect 33294 62514 33346 62526
rect 34078 62578 34130 62590
rect 34078 62514 34130 62526
rect 36542 62578 36594 62590
rect 36542 62514 36594 62526
rect 37662 62578 37714 62590
rect 37662 62514 37714 62526
rect 38110 62578 38162 62590
rect 38110 62514 38162 62526
rect 39118 62578 39170 62590
rect 39118 62514 39170 62526
rect 41022 62578 41074 62590
rect 41022 62514 41074 62526
rect 41134 62578 41186 62590
rect 41134 62514 41186 62526
rect 41694 62578 41746 62590
rect 41694 62514 41746 62526
rect 42030 62578 42082 62590
rect 42030 62514 42082 62526
rect 42590 62578 42642 62590
rect 42590 62514 42642 62526
rect 43262 62578 43314 62590
rect 43262 62514 43314 62526
rect 43822 62578 43874 62590
rect 43822 62514 43874 62526
rect 44606 62578 44658 62590
rect 44606 62514 44658 62526
rect 16718 62466 16770 62478
rect 16718 62402 16770 62414
rect 16830 62466 16882 62478
rect 28142 62466 28194 62478
rect 18610 62414 18622 62466
rect 18674 62414 18686 62466
rect 16830 62402 16882 62414
rect 28142 62402 28194 62414
rect 28254 62466 28306 62478
rect 28254 62402 28306 62414
rect 33518 62466 33570 62478
rect 33518 62402 33570 62414
rect 34302 62466 34354 62478
rect 34302 62402 34354 62414
rect 39454 62466 39506 62478
rect 39454 62402 39506 62414
rect 40350 62466 40402 62478
rect 40350 62402 40402 62414
rect 41358 62466 41410 62478
rect 41358 62402 41410 62414
rect 41806 62466 41858 62478
rect 44046 62466 44098 62478
rect 43586 62414 43598 62466
rect 43650 62414 43662 62466
rect 41806 62402 41858 62414
rect 44046 62402 44098 62414
rect 44158 62466 44210 62478
rect 44158 62402 44210 62414
rect 13022 62354 13074 62366
rect 9650 62302 9662 62354
rect 9714 62302 9726 62354
rect 13022 62290 13074 62302
rect 15710 62354 15762 62366
rect 16494 62354 16546 62366
rect 28478 62354 28530 62366
rect 35198 62354 35250 62366
rect 16258 62302 16270 62354
rect 16322 62302 16334 62354
rect 18386 62302 18398 62354
rect 18450 62302 18462 62354
rect 24210 62302 24222 62354
rect 24274 62302 24286 62354
rect 28802 62302 28814 62354
rect 28866 62302 28878 62354
rect 29474 62302 29486 62354
rect 29538 62302 29550 62354
rect 33842 62302 33854 62354
rect 33906 62302 33918 62354
rect 15710 62290 15762 62302
rect 16494 62290 16546 62302
rect 28478 62290 28530 62302
rect 35198 62290 35250 62302
rect 39678 62354 39730 62366
rect 39678 62290 39730 62302
rect 40014 62354 40066 62366
rect 40014 62290 40066 62302
rect 40910 62354 40962 62366
rect 40910 62290 40962 62302
rect 42366 62354 42418 62366
rect 42802 62302 42814 62354
rect 42866 62302 42878 62354
rect 45378 62302 45390 62354
rect 45442 62302 45454 62354
rect 48738 62302 48750 62354
rect 48802 62302 48814 62354
rect 42366 62290 42418 62302
rect 15934 62242 15986 62254
rect 25342 62242 25394 62254
rect 10322 62190 10334 62242
rect 10386 62190 10398 62242
rect 12450 62190 12462 62242
rect 12514 62190 12526 62242
rect 21298 62190 21310 62242
rect 21362 62190 21374 62242
rect 15934 62178 15986 62190
rect 25342 62178 25394 62190
rect 26014 62242 26066 62254
rect 26014 62178 26066 62190
rect 27470 62242 27522 62254
rect 27470 62178 27522 62190
rect 27918 62242 27970 62254
rect 27918 62178 27970 62190
rect 31614 62242 31666 62254
rect 31614 62178 31666 62190
rect 32286 62242 32338 62254
rect 32286 62178 32338 62190
rect 34750 62242 34802 62254
rect 34750 62178 34802 62190
rect 35646 62242 35698 62254
rect 35646 62178 35698 62190
rect 36094 62242 36146 62254
rect 36094 62178 36146 62190
rect 37326 62242 37378 62254
rect 37326 62178 37378 62190
rect 39902 62242 39954 62254
rect 46050 62190 46062 62242
rect 46114 62190 46126 62242
rect 48178 62190 48190 62242
rect 48242 62190 48254 62242
rect 50754 62190 50766 62242
rect 50818 62190 50830 62242
rect 39902 62178 39954 62190
rect 32958 62130 33010 62142
rect 27122 62078 27134 62130
rect 27186 62127 27198 62130
rect 27794 62127 27806 62130
rect 27186 62081 27806 62127
rect 27186 62078 27198 62081
rect 27794 62078 27806 62081
rect 27858 62078 27870 62130
rect 32958 62066 33010 62078
rect 33966 62130 34018 62142
rect 33966 62066 34018 62078
rect 1344 61962 58576 61996
rect 1344 61910 4478 61962
rect 4530 61910 4582 61962
rect 4634 61910 4686 61962
rect 4738 61910 35198 61962
rect 35250 61910 35302 61962
rect 35354 61910 35406 61962
rect 35458 61910 58576 61962
rect 1344 61876 58576 61910
rect 40798 61794 40850 61806
rect 30482 61742 30494 61794
rect 30546 61742 30558 61794
rect 40798 61730 40850 61742
rect 41134 61794 41186 61806
rect 41134 61730 41186 61742
rect 41470 61794 41522 61806
rect 41470 61730 41522 61742
rect 41806 61794 41858 61806
rect 41806 61730 41858 61742
rect 42142 61794 42194 61806
rect 42142 61730 42194 61742
rect 45726 61794 45778 61806
rect 45726 61730 45778 61742
rect 9998 61682 10050 61694
rect 32398 61682 32450 61694
rect 40574 61682 40626 61694
rect 10546 61630 10558 61682
rect 10610 61630 10622 61682
rect 15026 61630 15038 61682
rect 15090 61630 15102 61682
rect 17154 61630 17166 61682
rect 17218 61630 17230 61682
rect 20402 61630 20414 61682
rect 20466 61630 20478 61682
rect 22082 61630 22094 61682
rect 22146 61630 22158 61682
rect 24210 61630 24222 61682
rect 24274 61630 24286 61682
rect 25106 61630 25118 61682
rect 25170 61630 25182 61682
rect 31826 61630 31838 61682
rect 31890 61630 31902 61682
rect 33618 61630 33630 61682
rect 33682 61630 33694 61682
rect 38098 61630 38110 61682
rect 38162 61630 38174 61682
rect 9998 61618 10050 61630
rect 32398 61618 32450 61630
rect 40574 61618 40626 61630
rect 43598 61682 43650 61694
rect 43598 61618 43650 61630
rect 45278 61682 45330 61694
rect 45278 61618 45330 61630
rect 46286 61682 46338 61694
rect 48066 61630 48078 61682
rect 48130 61630 48142 61682
rect 50194 61630 50206 61682
rect 50258 61630 50270 61682
rect 46286 61618 46338 61630
rect 10110 61570 10162 61582
rect 10670 61570 10722 61582
rect 11902 61570 11954 61582
rect 27470 61570 27522 61582
rect 10434 61518 10446 61570
rect 10498 61518 10510 61570
rect 11106 61518 11118 61570
rect 11170 61518 11182 61570
rect 12114 61518 12126 61570
rect 12178 61518 12190 61570
rect 14242 61518 14254 61570
rect 14306 61518 14318 61570
rect 17602 61518 17614 61570
rect 17666 61518 17678 61570
rect 21298 61518 21310 61570
rect 21362 61518 21374 61570
rect 24546 61518 24558 61570
rect 24610 61518 24622 61570
rect 25330 61518 25342 61570
rect 25394 61518 25406 61570
rect 10110 61506 10162 61518
rect 10670 61506 10722 61518
rect 11902 61506 11954 61518
rect 27470 61506 27522 61518
rect 27694 61570 27746 61582
rect 27694 61506 27746 61518
rect 27918 61570 27970 61582
rect 27918 61506 27970 61518
rect 28366 61570 28418 61582
rect 28366 61506 28418 61518
rect 29038 61570 29090 61582
rect 29038 61506 29090 61518
rect 29934 61570 29986 61582
rect 32174 61570 32226 61582
rect 30818 61518 30830 61570
rect 30882 61518 30894 61570
rect 31378 61518 31390 61570
rect 31442 61518 31454 61570
rect 29934 61506 29986 61518
rect 32174 61506 32226 61518
rect 32510 61570 32562 61582
rect 32510 61506 32562 61518
rect 32734 61570 32786 61582
rect 39902 61570 39954 61582
rect 33954 61518 33966 61570
rect 34018 61518 34030 61570
rect 34626 61518 34638 61570
rect 34690 61518 34702 61570
rect 35074 61518 35086 61570
rect 35138 61518 35150 61570
rect 37538 61518 37550 61570
rect 37602 61518 37614 61570
rect 38658 61518 38670 61570
rect 38722 61518 38734 61570
rect 32734 61506 32786 61518
rect 39902 61506 39954 61518
rect 40238 61570 40290 61582
rect 40238 61506 40290 61518
rect 45950 61570 46002 61582
rect 45950 61506 46002 61518
rect 46398 61570 46450 61582
rect 50878 61570 50930 61582
rect 47282 61518 47294 61570
rect 47346 61518 47358 61570
rect 46398 61506 46450 61518
rect 50878 61506 50930 61518
rect 11454 61458 11506 61470
rect 26238 61458 26290 61470
rect 12562 61406 12574 61458
rect 12626 61406 12638 61458
rect 13906 61406 13918 61458
rect 13970 61406 13982 61458
rect 18274 61406 18286 61458
rect 18338 61406 18350 61458
rect 25666 61406 25678 61458
rect 25730 61406 25742 61458
rect 11454 61394 11506 61406
rect 26238 61394 26290 61406
rect 26350 61458 26402 61470
rect 26350 61394 26402 61406
rect 29262 61458 29314 61470
rect 29262 61394 29314 61406
rect 29374 61458 29426 61470
rect 29374 61394 29426 61406
rect 29822 61458 29874 61470
rect 29822 61394 29874 61406
rect 30046 61458 30098 61470
rect 40126 61458 40178 61470
rect 31490 61406 31502 61458
rect 31554 61406 31566 61458
rect 33730 61406 33742 61458
rect 33794 61406 33806 61458
rect 37986 61406 37998 61458
rect 38050 61406 38062 61458
rect 30046 61394 30098 61406
rect 40126 61394 40178 61406
rect 42254 61458 42306 61470
rect 42254 61394 42306 61406
rect 42702 61458 42754 61470
rect 42702 61394 42754 61406
rect 44942 61458 44994 61470
rect 44942 61394 44994 61406
rect 46174 61458 46226 61470
rect 46174 61394 46226 61406
rect 10894 61346 10946 61358
rect 10894 61282 10946 61294
rect 11678 61346 11730 61358
rect 11678 61282 11730 61294
rect 11790 61346 11842 61358
rect 11790 61282 11842 61294
rect 12910 61346 12962 61358
rect 12910 61282 12962 61294
rect 13582 61346 13634 61358
rect 13582 61282 13634 61294
rect 26574 61346 26626 61358
rect 26574 61282 26626 61294
rect 26798 61346 26850 61358
rect 26798 61282 26850 61294
rect 26910 61346 26962 61358
rect 26910 61282 26962 61294
rect 27022 61346 27074 61358
rect 27022 61282 27074 61294
rect 28142 61346 28194 61358
rect 35758 61346 35810 61358
rect 35298 61294 35310 61346
rect 35362 61294 35374 61346
rect 28142 61282 28194 61294
rect 35758 61282 35810 61294
rect 36206 61346 36258 61358
rect 36206 61282 36258 61294
rect 37326 61346 37378 61358
rect 37326 61282 37378 61294
rect 39006 61346 39058 61358
rect 41582 61346 41634 61358
rect 39330 61294 39342 61346
rect 39394 61294 39406 61346
rect 39006 61282 39058 61294
rect 41582 61282 41634 61294
rect 43150 61346 43202 61358
rect 43150 61282 43202 61294
rect 44382 61346 44434 61358
rect 44382 61282 44434 61294
rect 45166 61346 45218 61358
rect 45166 61282 45218 61294
rect 45390 61346 45442 61358
rect 45390 61282 45442 61294
rect 46958 61346 47010 61358
rect 50530 61294 50542 61346
rect 50594 61294 50606 61346
rect 46958 61282 47010 61294
rect 1344 61178 58576 61212
rect 1344 61126 19838 61178
rect 19890 61126 19942 61178
rect 19994 61126 20046 61178
rect 20098 61126 50558 61178
rect 50610 61126 50662 61178
rect 50714 61126 50766 61178
rect 50818 61126 58576 61178
rect 1344 61092 58576 61126
rect 14478 61010 14530 61022
rect 18846 61010 18898 61022
rect 12786 60958 12798 61010
rect 12850 60958 12862 61010
rect 14802 60958 14814 61010
rect 14866 60958 14878 61010
rect 14478 60946 14530 60958
rect 18846 60946 18898 60958
rect 19630 61010 19682 61022
rect 19630 60946 19682 60958
rect 20862 61010 20914 61022
rect 20862 60946 20914 60958
rect 21758 61010 21810 61022
rect 21758 60946 21810 60958
rect 22430 61010 22482 61022
rect 22430 60946 22482 60958
rect 23102 61010 23154 61022
rect 28926 61010 28978 61022
rect 24658 60958 24670 61010
rect 24722 60958 24734 61010
rect 23102 60946 23154 60958
rect 28926 60946 28978 60958
rect 30382 61010 30434 61022
rect 30382 60946 30434 60958
rect 31502 61010 31554 61022
rect 31502 60946 31554 60958
rect 41694 61010 41746 61022
rect 41694 60946 41746 60958
rect 50318 61010 50370 61022
rect 50318 60946 50370 60958
rect 16046 60898 16098 60910
rect 10322 60846 10334 60898
rect 10386 60846 10398 60898
rect 16046 60834 16098 60846
rect 16158 60898 16210 60910
rect 18958 60898 19010 60910
rect 16818 60846 16830 60898
rect 16882 60846 16894 60898
rect 16158 60834 16210 60846
rect 18958 60834 19010 60846
rect 22206 60898 22258 60910
rect 22206 60834 22258 60846
rect 22654 60898 22706 60910
rect 22654 60834 22706 60846
rect 23214 60898 23266 60910
rect 23214 60834 23266 60846
rect 28478 60898 28530 60910
rect 28478 60834 28530 60846
rect 30270 60898 30322 60910
rect 30270 60834 30322 60846
rect 30606 60898 30658 60910
rect 30606 60834 30658 60846
rect 32062 60898 32114 60910
rect 48850 60846 48862 60898
rect 48914 60846 48926 60898
rect 32062 60834 32114 60846
rect 13134 60786 13186 60798
rect 17950 60786 18002 60798
rect 9538 60734 9550 60786
rect 9602 60734 9614 60786
rect 16594 60734 16606 60786
rect 16658 60734 16670 60786
rect 13134 60722 13186 60734
rect 17950 60722 18002 60734
rect 19518 60786 19570 60798
rect 19518 60722 19570 60734
rect 19742 60786 19794 60798
rect 19742 60722 19794 60734
rect 20190 60786 20242 60798
rect 20190 60722 20242 60734
rect 20302 60786 20354 60798
rect 21198 60786 21250 60798
rect 22094 60786 22146 60798
rect 20626 60734 20638 60786
rect 20690 60734 20702 60786
rect 21522 60734 21534 60786
rect 21586 60734 21598 60786
rect 20302 60722 20354 60734
rect 21198 60722 21250 60734
rect 22094 60722 22146 60734
rect 22990 60786 23042 60798
rect 22990 60722 23042 60734
rect 24334 60786 24386 60798
rect 28702 60786 28754 60798
rect 28130 60734 28142 60786
rect 28194 60734 28206 60786
rect 24334 60722 24386 60734
rect 28702 60722 28754 60734
rect 30158 60786 30210 60798
rect 30158 60722 30210 60734
rect 32286 60786 32338 60798
rect 32286 60722 32338 60734
rect 32510 60786 32562 60798
rect 34750 60786 34802 60798
rect 32946 60734 32958 60786
rect 33010 60734 33022 60786
rect 33730 60734 33742 60786
rect 33794 60734 33806 60786
rect 32510 60722 32562 60734
rect 34750 60722 34802 60734
rect 34974 60786 35026 60798
rect 34974 60722 35026 60734
rect 35422 60786 35474 60798
rect 38894 60786 38946 60798
rect 35746 60734 35758 60786
rect 35810 60734 35822 60786
rect 35422 60722 35474 60734
rect 38894 60722 38946 60734
rect 39118 60786 39170 60798
rect 39118 60722 39170 60734
rect 39566 60786 39618 60798
rect 46162 60734 46174 60786
rect 46226 60734 46238 60786
rect 46946 60734 46958 60786
rect 47010 60734 47022 60786
rect 47506 60734 47518 60786
rect 47570 60734 47582 60786
rect 49074 60734 49086 60786
rect 49138 60734 49150 60786
rect 49858 60734 49870 60786
rect 49922 60734 49934 60786
rect 39566 60722 39618 60734
rect 17502 60674 17554 60686
rect 12450 60622 12462 60674
rect 12514 60622 12526 60674
rect 17502 60610 17554 60622
rect 21422 60674 21474 60686
rect 21422 60610 21474 60622
rect 23998 60674 24050 60686
rect 28590 60674 28642 60686
rect 25218 60622 25230 60674
rect 25282 60622 25294 60674
rect 27346 60622 27358 60674
rect 27410 60622 27422 60674
rect 23998 60610 24050 60622
rect 28590 60610 28642 60622
rect 29710 60674 29762 60686
rect 29710 60610 29762 60622
rect 31054 60674 31106 60686
rect 31054 60610 31106 60622
rect 32398 60674 32450 60686
rect 34862 60674 34914 60686
rect 39006 60674 39058 60686
rect 33170 60622 33182 60674
rect 33234 60622 33246 60674
rect 33618 60622 33630 60674
rect 33682 60622 33694 60674
rect 36418 60622 36430 60674
rect 36482 60622 36494 60674
rect 38546 60622 38558 60674
rect 38610 60622 38622 60674
rect 32398 60610 32450 60622
rect 34862 60610 34914 60622
rect 39006 60610 39058 60622
rect 40014 60674 40066 60686
rect 40014 60610 40066 60622
rect 40350 60674 40402 60686
rect 40350 60610 40402 60622
rect 41022 60674 41074 60686
rect 41022 60610 41074 60622
rect 42366 60674 42418 60686
rect 42366 60610 42418 60622
rect 43038 60674 43090 60686
rect 43250 60622 43262 60674
rect 43314 60622 43326 60674
rect 45378 60622 45390 60674
rect 45442 60622 45454 60674
rect 47394 60622 47406 60674
rect 47458 60622 47470 60674
rect 48850 60622 48862 60674
rect 48914 60622 48926 60674
rect 43038 60610 43090 60622
rect 16046 60562 16098 60574
rect 16046 60498 16098 60510
rect 17390 60562 17442 60574
rect 17390 60498 17442 60510
rect 20526 60562 20578 60574
rect 20526 60498 20578 60510
rect 47294 60562 47346 60574
rect 47294 60498 47346 60510
rect 1344 60394 58576 60428
rect 1344 60342 4478 60394
rect 4530 60342 4582 60394
rect 4634 60342 4686 60394
rect 4738 60342 35198 60394
rect 35250 60342 35302 60394
rect 35354 60342 35406 60394
rect 35458 60342 58576 60394
rect 1344 60308 58576 60342
rect 12126 60226 12178 60238
rect 12126 60162 12178 60174
rect 26238 60226 26290 60238
rect 28030 60226 28082 60238
rect 26562 60174 26574 60226
rect 26626 60174 26638 60226
rect 26238 60162 26290 60174
rect 28030 60162 28082 60174
rect 28366 60226 28418 60238
rect 28366 60162 28418 60174
rect 36206 60226 36258 60238
rect 48750 60226 48802 60238
rect 48066 60174 48078 60226
rect 48130 60174 48142 60226
rect 36206 60162 36258 60174
rect 48750 60162 48802 60174
rect 49086 60226 49138 60238
rect 49086 60162 49138 60174
rect 49198 60226 49250 60238
rect 49198 60162 49250 60174
rect 12238 60114 12290 60126
rect 12238 60050 12290 60062
rect 23102 60114 23154 60126
rect 29598 60114 29650 60126
rect 35982 60114 36034 60126
rect 24322 60062 24334 60114
rect 24386 60062 24398 60114
rect 32834 60062 32846 60114
rect 32898 60062 32910 60114
rect 34962 60062 34974 60114
rect 35026 60062 35038 60114
rect 23102 60050 23154 60062
rect 29598 60050 29650 60062
rect 35982 60050 36034 60062
rect 38110 60114 38162 60126
rect 39554 60062 39566 60114
rect 39618 60062 39630 60114
rect 46946 60062 46958 60114
rect 47010 60062 47022 60114
rect 38110 60050 38162 60062
rect 11454 60002 11506 60014
rect 11454 59938 11506 59950
rect 15486 60002 15538 60014
rect 19630 60002 19682 60014
rect 23662 60002 23714 60014
rect 16034 59950 16046 60002
rect 16098 59950 16110 60002
rect 20514 59950 20526 60002
rect 20578 59950 20590 60002
rect 22082 59950 22094 60002
rect 22146 59950 22158 60002
rect 15486 59938 15538 59950
rect 19630 59938 19682 59950
rect 23662 59938 23714 59950
rect 23886 60002 23938 60014
rect 23886 59938 23938 59950
rect 26014 60002 26066 60014
rect 27134 60002 27186 60014
rect 37102 60002 37154 60014
rect 26898 59950 26910 60002
rect 26962 59950 26974 60002
rect 28018 59950 28030 60002
rect 28082 59950 28094 60002
rect 32162 59950 32174 60002
rect 32226 59950 32238 60002
rect 26014 59938 26066 59950
rect 27134 59938 27186 59950
rect 37102 59938 37154 59950
rect 37326 60002 37378 60014
rect 42366 60002 42418 60014
rect 37538 59950 37550 60002
rect 37602 59950 37614 60002
rect 38210 59950 38222 60002
rect 38274 59950 38286 60002
rect 39330 59950 39342 60002
rect 39394 59950 39406 60002
rect 39778 59950 39790 60002
rect 39842 59950 39854 60002
rect 40002 59950 40014 60002
rect 40066 59950 40078 60002
rect 42018 59950 42030 60002
rect 42082 59950 42094 60002
rect 37326 59938 37378 59950
rect 42366 59938 42418 59950
rect 42590 60002 42642 60014
rect 43710 60002 43762 60014
rect 42914 59950 42926 60002
rect 42978 59950 42990 60002
rect 42590 59938 42642 59950
rect 43710 59938 43762 59950
rect 46398 60002 46450 60014
rect 47518 60002 47570 60014
rect 46722 59950 46734 60002
rect 46786 59950 46798 60002
rect 46398 59938 46450 59950
rect 47518 59938 47570 59950
rect 48862 60002 48914 60014
rect 48862 59938 48914 59950
rect 11678 59890 11730 59902
rect 11678 59826 11730 59838
rect 11790 59890 11842 59902
rect 11790 59826 11842 59838
rect 16494 59890 16546 59902
rect 27246 59890 27298 59902
rect 40574 59890 40626 59902
rect 20738 59838 20750 59890
rect 20802 59838 20814 59890
rect 21858 59838 21870 59890
rect 21922 59838 21934 59890
rect 30930 59838 30942 59890
rect 30994 59838 31006 59890
rect 38546 59838 38558 59890
rect 38610 59838 38622 59890
rect 16494 59826 16546 59838
rect 27246 59826 27298 59838
rect 40574 59826 40626 59838
rect 42254 59890 42306 59902
rect 42254 59826 42306 59838
rect 43486 59890 43538 59902
rect 43486 59826 43538 59838
rect 44830 59890 44882 59902
rect 44830 59826 44882 59838
rect 45166 59890 45218 59902
rect 45166 59826 45218 59838
rect 45502 59890 45554 59902
rect 45502 59826 45554 59838
rect 45614 59890 45666 59902
rect 45614 59826 45666 59838
rect 46958 59890 47010 59902
rect 46958 59826 47010 59838
rect 47406 59890 47458 59902
rect 47406 59826 47458 59838
rect 47630 59890 47682 59902
rect 47630 59826 47682 59838
rect 15598 59778 15650 59790
rect 15598 59714 15650 59726
rect 15710 59778 15762 59790
rect 15710 59714 15762 59726
rect 15822 59778 15874 59790
rect 15822 59714 15874 59726
rect 16382 59778 16434 59790
rect 16382 59714 16434 59726
rect 20078 59778 20130 59790
rect 20078 59714 20130 59726
rect 21534 59778 21586 59790
rect 21534 59714 21586 59726
rect 22654 59778 22706 59790
rect 22654 59714 22706 59726
rect 25230 59778 25282 59790
rect 25230 59714 25282 59726
rect 25790 59778 25842 59790
rect 31278 59778 31330 59790
rect 27682 59726 27694 59778
rect 27746 59726 27758 59778
rect 25790 59714 25842 59726
rect 31278 59714 31330 59726
rect 31838 59778 31890 59790
rect 31838 59714 31890 59726
rect 35534 59778 35586 59790
rect 35534 59714 35586 59726
rect 35646 59778 35698 59790
rect 35646 59714 35698 59726
rect 35758 59778 35810 59790
rect 35758 59714 35810 59726
rect 37438 59778 37490 59790
rect 37438 59714 37490 59726
rect 39566 59778 39618 59790
rect 39566 59714 39618 59726
rect 40238 59778 40290 59790
rect 40238 59714 40290 59726
rect 40462 59778 40514 59790
rect 40462 59714 40514 59726
rect 41022 59778 41074 59790
rect 41022 59714 41074 59726
rect 41470 59778 41522 59790
rect 41470 59714 41522 59726
rect 43150 59778 43202 59790
rect 43150 59714 43202 59726
rect 43262 59778 43314 59790
rect 46062 59778 46114 59790
rect 44034 59726 44046 59778
rect 44098 59726 44110 59778
rect 43262 59714 43314 59726
rect 46062 59714 46114 59726
rect 49758 59778 49810 59790
rect 49758 59714 49810 59726
rect 50206 59778 50258 59790
rect 50206 59714 50258 59726
rect 1344 59610 58576 59644
rect 1344 59558 19838 59610
rect 19890 59558 19942 59610
rect 19994 59558 20046 59610
rect 20098 59558 50558 59610
rect 50610 59558 50662 59610
rect 50714 59558 50766 59610
rect 50818 59558 58576 59610
rect 1344 59524 58576 59558
rect 17502 59442 17554 59454
rect 17502 59378 17554 59390
rect 18846 59442 18898 59454
rect 18846 59378 18898 59390
rect 19070 59442 19122 59454
rect 19966 59442 20018 59454
rect 19394 59390 19406 59442
rect 19458 59390 19470 59442
rect 19070 59378 19122 59390
rect 19966 59378 20018 59390
rect 24110 59442 24162 59454
rect 24110 59378 24162 59390
rect 24558 59442 24610 59454
rect 24558 59378 24610 59390
rect 27134 59442 27186 59454
rect 34526 59442 34578 59454
rect 39342 59442 39394 59454
rect 33058 59390 33070 59442
rect 33122 59390 33134 59442
rect 27134 59378 27186 59390
rect 34190 59386 34242 59398
rect 19742 59330 19794 59342
rect 26238 59330 26290 59342
rect 14690 59278 14702 59330
rect 14754 59278 14766 59330
rect 19742 59266 19794 59278
rect 20190 59274 20242 59286
rect 21410 59278 21422 59330
rect 21474 59278 21486 59330
rect 26238 59266 26290 59278
rect 27470 59330 27522 59342
rect 27470 59266 27522 59278
rect 33518 59330 33570 59342
rect 33518 59266 33570 59278
rect 33630 59330 33682 59342
rect 37986 59390 37998 59442
rect 38050 59390 38062 59442
rect 34526 59378 34578 59390
rect 39342 59378 39394 59390
rect 39566 59442 39618 59454
rect 39566 59378 39618 59390
rect 39678 59442 39730 59454
rect 39678 59378 39730 59390
rect 39902 59442 39954 59454
rect 42590 59442 42642 59454
rect 41122 59390 41134 59442
rect 41186 59390 41198 59442
rect 39902 59378 39954 59390
rect 42590 59378 42642 59390
rect 43710 59442 43762 59454
rect 43710 59378 43762 59390
rect 47518 59442 47570 59454
rect 47518 59378 47570 59390
rect 48638 59442 48690 59454
rect 48638 59378 48690 59390
rect 48862 59442 48914 59454
rect 48862 59378 48914 59390
rect 49422 59442 49474 59454
rect 49422 59378 49474 59390
rect 49870 59442 49922 59454
rect 49870 59378 49922 59390
rect 34190 59322 34242 59334
rect 34302 59330 34354 59342
rect 38446 59330 38498 59342
rect 33630 59266 33682 59278
rect 35522 59278 35534 59330
rect 35586 59278 35598 59330
rect 34302 59266 34354 59278
rect 38446 59266 38498 59278
rect 38558 59330 38610 59342
rect 47742 59330 47794 59342
rect 41570 59278 41582 59330
rect 41634 59278 41646 59330
rect 38558 59266 38610 59278
rect 47742 59266 47794 59278
rect 9538 59166 9550 59218
rect 9602 59166 9614 59218
rect 14018 59166 14030 59218
rect 14082 59166 14094 59218
rect 20190 59210 20242 59222
rect 22766 59218 22818 59230
rect 20738 59166 20750 59218
rect 20802 59166 20814 59218
rect 21522 59166 21534 59218
rect 21586 59166 21598 59218
rect 22766 59154 22818 59166
rect 24670 59218 24722 59230
rect 24670 59154 24722 59166
rect 26126 59218 26178 59230
rect 26126 59154 26178 59166
rect 26798 59218 26850 59230
rect 26798 59154 26850 59166
rect 27134 59218 27186 59230
rect 32286 59218 32338 59230
rect 29026 59166 29038 59218
rect 29090 59166 29102 59218
rect 27134 59154 27186 59166
rect 32286 59154 32338 59166
rect 33742 59218 33794 59230
rect 38670 59218 38722 59230
rect 34850 59166 34862 59218
rect 34914 59166 34926 59218
rect 33742 59154 33794 59166
rect 38670 59154 38722 59166
rect 39230 59218 39282 59230
rect 39230 59154 39282 59166
rect 40014 59218 40066 59230
rect 42478 59218 42530 59230
rect 41122 59166 41134 59218
rect 41186 59166 41198 59218
rect 41794 59166 41806 59218
rect 41858 59166 41870 59218
rect 40014 59154 40066 59166
rect 42478 59154 42530 59166
rect 42814 59218 42866 59230
rect 42814 59154 42866 59166
rect 43486 59218 43538 59230
rect 43486 59154 43538 59166
rect 43822 59218 43874 59230
rect 43822 59154 43874 59166
rect 44046 59218 44098 59230
rect 46174 59218 46226 59230
rect 46958 59218 47010 59230
rect 44258 59166 44270 59218
rect 44322 59166 44334 59218
rect 45154 59166 45166 59218
rect 45218 59166 45230 59218
rect 46498 59166 46510 59218
rect 46562 59166 46574 59218
rect 44046 59154 44098 59166
rect 46174 59154 46226 59166
rect 46958 59154 47010 59166
rect 47294 59218 47346 59230
rect 47294 59154 47346 59166
rect 48974 59218 49026 59230
rect 48974 59154 49026 59166
rect 8990 59106 9042 59118
rect 22430 59106 22482 59118
rect 10322 59054 10334 59106
rect 10386 59054 10398 59106
rect 12450 59054 12462 59106
rect 12514 59054 12526 59106
rect 16818 59054 16830 59106
rect 16882 59054 16894 59106
rect 20066 59054 20078 59106
rect 20130 59054 20142 59106
rect 21410 59054 21422 59106
rect 21474 59054 21486 59106
rect 8990 59042 9042 59054
rect 22430 59042 22482 59054
rect 23662 59106 23714 59118
rect 23662 59042 23714 59054
rect 27918 59106 27970 59118
rect 27918 59042 27970 59054
rect 28814 59106 28866 59118
rect 43150 59106 43202 59118
rect 29810 59054 29822 59106
rect 29874 59054 29886 59106
rect 31938 59054 31950 59106
rect 32002 59054 32014 59106
rect 37650 59054 37662 59106
rect 37714 59054 37726 59106
rect 28814 59042 28866 59054
rect 43150 59042 43202 59054
rect 45502 59106 45554 59118
rect 45502 59042 45554 59054
rect 47406 59106 47458 59118
rect 47406 59042 47458 59054
rect 50318 59106 50370 59118
rect 50318 59042 50370 59054
rect 8878 58994 8930 59006
rect 8878 58930 8930 58942
rect 24558 58994 24610 59006
rect 24558 58930 24610 58942
rect 25230 58994 25282 59006
rect 25230 58930 25282 58942
rect 25342 58994 25394 59006
rect 25342 58930 25394 58942
rect 25566 58994 25618 59006
rect 25566 58930 25618 58942
rect 25678 58994 25730 59006
rect 25678 58930 25730 58942
rect 26238 58994 26290 59006
rect 26238 58930 26290 58942
rect 32398 58994 32450 59006
rect 45266 58942 45278 58994
rect 45330 58942 45342 58994
rect 32398 58930 32450 58942
rect 1344 58826 58576 58860
rect 1344 58774 4478 58826
rect 4530 58774 4582 58826
rect 4634 58774 4686 58826
rect 4738 58774 35198 58826
rect 35250 58774 35302 58826
rect 35354 58774 35406 58826
rect 35458 58774 58576 58826
rect 1344 58740 58576 58774
rect 27694 58658 27746 58670
rect 27694 58594 27746 58606
rect 29486 58658 29538 58670
rect 29486 58594 29538 58606
rect 33182 58658 33234 58670
rect 33182 58594 33234 58606
rect 33518 58658 33570 58670
rect 33518 58594 33570 58606
rect 34302 58658 34354 58670
rect 40786 58606 40798 58658
rect 40850 58606 40862 58658
rect 41794 58606 41806 58658
rect 41858 58606 41870 58658
rect 34302 58594 34354 58606
rect 21534 58546 21586 58558
rect 30046 58546 30098 58558
rect 9650 58494 9662 58546
rect 9714 58494 9726 58546
rect 14914 58494 14926 58546
rect 14978 58494 14990 58546
rect 15922 58494 15934 58546
rect 15986 58494 15998 58546
rect 24658 58494 24670 58546
rect 24722 58494 24734 58546
rect 25778 58494 25790 58546
rect 25842 58494 25854 58546
rect 21534 58482 21586 58494
rect 30046 58482 30098 58494
rect 30942 58546 30994 58558
rect 30942 58482 30994 58494
rect 32734 58546 32786 58558
rect 32734 58482 32786 58494
rect 33406 58546 33458 58558
rect 33406 58482 33458 58494
rect 39566 58546 39618 58558
rect 45278 58546 45330 58558
rect 41458 58494 41470 58546
rect 41522 58494 41534 58546
rect 50082 58494 50094 58546
rect 50146 58494 50158 58546
rect 39566 58482 39618 58494
rect 45278 58482 45330 58494
rect 15038 58434 15090 58446
rect 16046 58434 16098 58446
rect 12226 58382 12238 58434
rect 12290 58382 12302 58434
rect 14802 58382 14814 58434
rect 14866 58382 14878 58434
rect 15474 58382 15486 58434
rect 15538 58382 15550 58434
rect 15038 58370 15090 58382
rect 16046 58370 16098 58382
rect 17166 58434 17218 58446
rect 17166 58370 17218 58382
rect 17614 58434 17666 58446
rect 19854 58434 19906 58446
rect 30158 58434 30210 58446
rect 34190 58434 34242 58446
rect 18834 58382 18846 58434
rect 18898 58382 18910 58434
rect 21858 58382 21870 58434
rect 21922 58382 21934 58434
rect 24882 58382 24894 58434
rect 24946 58382 24958 58434
rect 25666 58382 25678 58434
rect 25730 58382 25742 58434
rect 26898 58382 26910 58434
rect 26962 58382 26974 58434
rect 28018 58382 28030 58434
rect 28082 58382 28094 58434
rect 29810 58382 29822 58434
rect 29874 58382 29886 58434
rect 32946 58382 32958 58434
rect 33010 58382 33022 58434
rect 17614 58370 17666 58382
rect 19854 58370 19906 58382
rect 30158 58370 30210 58382
rect 34190 58370 34242 58382
rect 37102 58434 37154 58446
rect 37102 58370 37154 58382
rect 37550 58434 37602 58446
rect 37550 58370 37602 58382
rect 38446 58434 38498 58446
rect 38446 58370 38498 58382
rect 39230 58434 39282 58446
rect 39230 58370 39282 58382
rect 39454 58434 39506 58446
rect 39454 58370 39506 58382
rect 39790 58434 39842 58446
rect 39790 58370 39842 58382
rect 40238 58434 40290 58446
rect 41346 58382 41358 58434
rect 41410 58382 41422 58434
rect 45938 58382 45950 58434
rect 46002 58382 46014 58434
rect 46834 58382 46846 58434
rect 46898 58382 46910 58434
rect 47170 58382 47182 58434
rect 47234 58382 47246 58434
rect 40238 58370 40290 58382
rect 16494 58322 16546 58334
rect 16494 58258 16546 58270
rect 17502 58322 17554 58334
rect 17502 58258 17554 58270
rect 17950 58322 18002 58334
rect 17950 58258 18002 58270
rect 20190 58322 20242 58334
rect 20190 58258 20242 58270
rect 20526 58322 20578 58334
rect 20526 58258 20578 58270
rect 20750 58322 20802 58334
rect 28142 58322 28194 58334
rect 36094 58322 36146 58334
rect 22530 58270 22542 58322
rect 22594 58270 22606 58322
rect 26338 58270 26350 58322
rect 26402 58270 26414 58322
rect 26674 58270 26686 58322
rect 26738 58270 26750 58322
rect 35186 58270 35198 58322
rect 35250 58270 35262 58322
rect 20750 58258 20802 58270
rect 28142 58258 28194 58270
rect 36094 58258 36146 58270
rect 38110 58322 38162 58334
rect 38110 58258 38162 58270
rect 38222 58322 38274 58334
rect 38222 58258 38274 58270
rect 40126 58322 40178 58334
rect 40126 58258 40178 58270
rect 40350 58322 40402 58334
rect 44382 58322 44434 58334
rect 42914 58270 42926 58322
rect 42978 58270 42990 58322
rect 40350 58258 40402 58270
rect 43598 58266 43650 58278
rect 12686 58210 12738 58222
rect 12686 58146 12738 58158
rect 14030 58210 14082 58222
rect 15262 58210 15314 58222
rect 14354 58158 14366 58210
rect 14418 58158 14430 58210
rect 14030 58146 14082 58158
rect 15262 58146 15314 58158
rect 15934 58210 15986 58222
rect 15934 58146 15986 58158
rect 16270 58210 16322 58222
rect 16270 58146 16322 58158
rect 17278 58210 17330 58222
rect 17278 58146 17330 58158
rect 17838 58210 17890 58222
rect 17838 58146 17890 58158
rect 18622 58210 18674 58222
rect 18622 58146 18674 58158
rect 19518 58210 19570 58222
rect 19518 58146 19570 58158
rect 19742 58210 19794 58222
rect 19742 58146 19794 58158
rect 20302 58210 20354 58222
rect 20302 58146 20354 58158
rect 28254 58210 28306 58222
rect 28254 58146 28306 58158
rect 28366 58210 28418 58222
rect 28366 58146 28418 58158
rect 29934 58210 29986 58222
rect 29934 58146 29986 58158
rect 31502 58210 31554 58222
rect 31502 58146 31554 58158
rect 31950 58210 32002 58222
rect 31950 58146 32002 58158
rect 34302 58210 34354 58222
rect 34302 58146 34354 58158
rect 34862 58210 34914 58222
rect 34862 58146 34914 58158
rect 35646 58210 35698 58222
rect 35646 58146 35698 58158
rect 37662 58210 37714 58222
rect 37662 58146 37714 58158
rect 37774 58210 37826 58222
rect 37774 58146 37826 58158
rect 38782 58210 38834 58222
rect 38782 58146 38834 58158
rect 42590 58210 42642 58222
rect 43598 58202 43650 58214
rect 43710 58266 43762 58278
rect 46722 58270 46734 58322
rect 46786 58270 46798 58322
rect 47954 58270 47966 58322
rect 48018 58270 48030 58322
rect 44382 58258 44434 58270
rect 43710 58202 43762 58214
rect 43934 58210 43986 58222
rect 42590 58146 42642 58158
rect 43934 58146 43986 58158
rect 44942 58210 44994 58222
rect 44942 58146 44994 58158
rect 45166 58210 45218 58222
rect 45166 58146 45218 58158
rect 45390 58210 45442 58222
rect 45826 58158 45838 58210
rect 45890 58158 45902 58210
rect 45390 58146 45442 58158
rect 1344 58042 58576 58076
rect 1344 57990 19838 58042
rect 19890 57990 19942 58042
rect 19994 57990 20046 58042
rect 20098 57990 50558 58042
rect 50610 57990 50662 58042
rect 50714 57990 50766 58042
rect 50818 57990 58576 58042
rect 1344 57956 58576 57990
rect 10670 57874 10722 57886
rect 10670 57810 10722 57822
rect 20750 57874 20802 57886
rect 20750 57810 20802 57822
rect 20974 57874 21026 57886
rect 20974 57810 21026 57822
rect 21422 57874 21474 57886
rect 21422 57810 21474 57822
rect 21534 57874 21586 57886
rect 21534 57810 21586 57822
rect 22766 57874 22818 57886
rect 22766 57810 22818 57822
rect 22878 57874 22930 57886
rect 30830 57874 30882 57886
rect 24546 57822 24558 57874
rect 24610 57822 24622 57874
rect 22878 57810 22930 57822
rect 30830 57810 30882 57822
rect 32622 57874 32674 57886
rect 32622 57810 32674 57822
rect 41806 57874 41858 57886
rect 41806 57810 41858 57822
rect 41918 57874 41970 57886
rect 41918 57810 41970 57822
rect 42030 57874 42082 57886
rect 42030 57810 42082 57822
rect 43486 57874 43538 57886
rect 43486 57810 43538 57822
rect 43710 57874 43762 57886
rect 43710 57810 43762 57822
rect 45166 57874 45218 57886
rect 47182 57874 47234 57886
rect 46722 57822 46734 57874
rect 46786 57822 46798 57874
rect 45166 57810 45218 57822
rect 47182 57810 47234 57822
rect 9662 57762 9714 57774
rect 21086 57762 21138 57774
rect 41134 57762 41186 57774
rect 13458 57710 13470 57762
rect 13522 57710 13534 57762
rect 18386 57710 18398 57762
rect 18450 57710 18462 57762
rect 23538 57710 23550 57762
rect 23602 57710 23614 57762
rect 9662 57698 9714 57710
rect 21086 57698 21138 57710
rect 41134 57698 41186 57710
rect 42254 57762 42306 57774
rect 42254 57698 42306 57710
rect 43822 57762 43874 57774
rect 43822 57698 43874 57710
rect 48078 57762 48130 57774
rect 48078 57698 48130 57710
rect 9550 57650 9602 57662
rect 6178 57598 6190 57650
rect 6242 57598 6254 57650
rect 9550 57586 9602 57598
rect 9886 57650 9938 57662
rect 9886 57586 9938 57598
rect 10446 57650 10498 57662
rect 10446 57586 10498 57598
rect 10558 57650 10610 57662
rect 10558 57586 10610 57598
rect 10782 57650 10834 57662
rect 21646 57650 21698 57662
rect 22654 57650 22706 57662
rect 10994 57598 11006 57650
rect 11058 57598 11070 57650
rect 12786 57598 12798 57650
rect 12850 57598 12862 57650
rect 17602 57598 17614 57650
rect 17666 57598 17678 57650
rect 21970 57598 21982 57650
rect 22034 57598 22046 57650
rect 10782 57586 10834 57598
rect 21646 57586 21698 57598
rect 22654 57586 22706 57598
rect 23326 57650 23378 57662
rect 30942 57650 30994 57662
rect 41022 57650 41074 57662
rect 23986 57598 23998 57650
rect 24050 57598 24062 57650
rect 24658 57598 24670 57650
rect 24722 57598 24734 57650
rect 25218 57598 25230 57650
rect 25282 57598 25294 57650
rect 33506 57598 33518 57650
rect 33570 57598 33582 57650
rect 38546 57598 38558 57650
rect 38610 57598 38622 57650
rect 23326 57586 23378 57598
rect 30942 57586 30994 57598
rect 41022 57586 41074 57598
rect 41358 57650 41410 57662
rect 41358 57586 41410 57598
rect 41582 57650 41634 57662
rect 41582 57586 41634 57598
rect 44942 57650 44994 57662
rect 44942 57586 44994 57598
rect 45278 57650 45330 57662
rect 45278 57586 45330 57598
rect 45614 57650 45666 57662
rect 45614 57586 45666 57598
rect 46062 57650 46114 57662
rect 46062 57586 46114 57598
rect 46174 57650 46226 57662
rect 46174 57586 46226 57598
rect 46286 57650 46338 57662
rect 46286 57586 46338 57598
rect 46958 57650 47010 57662
rect 46958 57586 47010 57598
rect 47406 57650 47458 57662
rect 47406 57586 47458 57598
rect 47630 57650 47682 57662
rect 47630 57586 47682 57598
rect 47854 57650 47906 57662
rect 47854 57586 47906 57598
rect 48190 57650 48242 57662
rect 48190 57586 48242 57598
rect 31390 57538 31442 57550
rect 34078 57538 34130 57550
rect 40350 57538 40402 57550
rect 6850 57486 6862 57538
rect 6914 57486 6926 57538
rect 8978 57486 8990 57538
rect 9042 57486 9054 57538
rect 20514 57486 20526 57538
rect 20578 57486 20590 57538
rect 27234 57486 27246 57538
rect 27298 57486 27310 57538
rect 33170 57486 33182 57538
rect 33234 57486 33246 57538
rect 36866 57486 36878 57538
rect 36930 57486 36942 57538
rect 31390 57474 31442 57486
rect 34078 57474 34130 57486
rect 40350 57474 40402 57486
rect 48862 57538 48914 57550
rect 48862 57474 48914 57486
rect 49310 57538 49362 57550
rect 49310 57474 49362 57486
rect 49758 57538 49810 57550
rect 49758 57474 49810 57486
rect 1344 57258 58576 57292
rect 1344 57206 4478 57258
rect 4530 57206 4582 57258
rect 4634 57206 4686 57258
rect 4738 57206 35198 57258
rect 35250 57206 35302 57258
rect 35354 57206 35406 57258
rect 35458 57206 58576 57258
rect 1344 57172 58576 57206
rect 11678 57090 11730 57102
rect 11678 57026 11730 57038
rect 13806 57090 13858 57102
rect 13806 57026 13858 57038
rect 18510 57090 18562 57102
rect 18510 57026 18562 57038
rect 18846 57090 18898 57102
rect 18846 57026 18898 57038
rect 19182 57090 19234 57102
rect 19182 57026 19234 57038
rect 20302 57090 20354 57102
rect 20302 57026 20354 57038
rect 21422 57090 21474 57102
rect 21422 57026 21474 57038
rect 22990 57090 23042 57102
rect 36318 57090 36370 57102
rect 24882 57038 24894 57090
rect 24946 57038 24958 57090
rect 22990 57026 23042 57038
rect 36318 57026 36370 57038
rect 11790 56978 11842 56990
rect 20414 56978 20466 56990
rect 8530 56926 8542 56978
rect 8594 56926 8606 56978
rect 8978 56926 8990 56978
rect 9042 56926 9054 56978
rect 15698 56926 15710 56978
rect 15762 56926 15774 56978
rect 17826 56926 17838 56978
rect 17890 56926 17902 56978
rect 11790 56914 11842 56926
rect 20414 56914 20466 56926
rect 23662 56978 23714 56990
rect 33966 56978 34018 56990
rect 45838 56978 45890 56990
rect 26450 56926 26462 56978
rect 26514 56926 26526 56978
rect 28578 56926 28590 56978
rect 28642 56926 28654 56978
rect 39330 56926 39342 56978
rect 39394 56926 39406 56978
rect 41458 56926 41470 56978
rect 41522 56926 41534 56978
rect 23662 56914 23714 56926
rect 33966 56914 34018 56926
rect 45838 56914 45890 56926
rect 48750 56978 48802 56990
rect 48750 56914 48802 56926
rect 9438 56866 9490 56878
rect 5730 56814 5742 56866
rect 5794 56814 5806 56866
rect 8866 56814 8878 56866
rect 8930 56814 8942 56866
rect 9438 56802 9490 56814
rect 11006 56866 11058 56878
rect 21310 56866 21362 56878
rect 14242 56814 14254 56866
rect 14306 56814 14318 56866
rect 14914 56814 14926 56866
rect 14978 56814 14990 56866
rect 18162 56814 18174 56866
rect 18226 56814 18238 56866
rect 11006 56802 11058 56814
rect 21310 56802 21362 56814
rect 22094 56866 22146 56878
rect 22094 56802 22146 56814
rect 22318 56866 22370 56878
rect 23550 56866 23602 56878
rect 23202 56814 23214 56866
rect 23266 56814 23278 56866
rect 22318 56802 22370 56814
rect 23550 56802 23602 56814
rect 23774 56866 23826 56878
rect 23774 56802 23826 56814
rect 24222 56866 24274 56878
rect 29150 56866 29202 56878
rect 32846 56866 32898 56878
rect 36430 56866 36482 56878
rect 47294 56866 47346 56878
rect 25666 56814 25678 56866
rect 25730 56814 25742 56866
rect 31826 56814 31838 56866
rect 31890 56814 31902 56866
rect 34402 56814 34414 56866
rect 34466 56814 34478 56866
rect 42242 56814 42254 56866
rect 42306 56814 42318 56866
rect 24222 56802 24274 56814
rect 29150 56802 29202 56814
rect 32846 56802 32898 56814
rect 36430 56802 36482 56814
rect 47294 56802 47346 56814
rect 9102 56754 9154 56766
rect 6402 56702 6414 56754
rect 6466 56702 6478 56754
rect 9102 56690 9154 56702
rect 10334 56754 10386 56766
rect 10334 56690 10386 56702
rect 10782 56754 10834 56766
rect 10782 56690 10834 56702
rect 11230 56754 11282 56766
rect 11230 56690 11282 56702
rect 11342 56754 11394 56766
rect 11342 56690 11394 56702
rect 13694 56754 13746 56766
rect 13694 56690 13746 56702
rect 18398 56754 18450 56766
rect 18398 56690 18450 56702
rect 19406 56754 19458 56766
rect 19406 56690 19458 56702
rect 21422 56754 21474 56766
rect 21422 56690 21474 56702
rect 22654 56754 22706 56766
rect 22654 56690 22706 56702
rect 22878 56754 22930 56766
rect 22878 56690 22930 56702
rect 24334 56754 24386 56766
rect 24334 56690 24386 56702
rect 24446 56754 24498 56766
rect 36990 56754 37042 56766
rect 30146 56702 30158 56754
rect 30210 56702 30222 56754
rect 33506 56702 33518 56754
rect 33570 56702 33582 56754
rect 35186 56702 35198 56754
rect 35250 56702 35262 56754
rect 24446 56690 24498 56702
rect 36990 56690 37042 56702
rect 37438 56754 37490 56766
rect 37438 56690 37490 56702
rect 38670 56754 38722 56766
rect 38670 56690 38722 56702
rect 44046 56754 44098 56766
rect 44046 56690 44098 56702
rect 47406 56754 47458 56766
rect 47406 56690 47458 56702
rect 47630 56754 47682 56766
rect 48302 56754 48354 56766
rect 47630 56690 47682 56702
rect 47966 56698 48018 56710
rect 9326 56642 9378 56654
rect 9326 56578 9378 56590
rect 9998 56642 10050 56654
rect 9998 56578 10050 56590
rect 10222 56642 10274 56654
rect 10222 56578 10274 56590
rect 10670 56642 10722 56654
rect 25342 56642 25394 56654
rect 30494 56642 30546 56654
rect 14466 56590 14478 56642
rect 14530 56590 14542 56642
rect 29474 56590 29486 56642
rect 29538 56590 29550 56642
rect 10670 56578 10722 56590
rect 25342 56578 25394 56590
rect 30494 56578 30546 56590
rect 30942 56642 30994 56654
rect 32286 56642 32338 56654
rect 31602 56590 31614 56642
rect 31666 56590 31678 56642
rect 30942 56578 30994 56590
rect 32286 56578 32338 56590
rect 33182 56642 33234 56654
rect 33182 56578 33234 56590
rect 34862 56642 34914 56654
rect 34862 56578 34914 56590
rect 37102 56642 37154 56654
rect 37102 56578 37154 56590
rect 37550 56642 37602 56654
rect 37550 56578 37602 56590
rect 37998 56642 38050 56654
rect 39006 56642 39058 56654
rect 38322 56590 38334 56642
rect 38386 56590 38398 56642
rect 37998 56578 38050 56590
rect 39006 56578 39058 56590
rect 43710 56642 43762 56654
rect 43710 56578 43762 56590
rect 43934 56642 43986 56654
rect 43934 56578 43986 56590
rect 46734 56642 46786 56654
rect 48302 56690 48354 56702
rect 47966 56634 48018 56646
rect 46734 56578 46786 56590
rect 1344 56474 58576 56508
rect 1344 56422 19838 56474
rect 19890 56422 19942 56474
rect 19994 56422 20046 56474
rect 20098 56422 50558 56474
rect 50610 56422 50662 56474
rect 50714 56422 50766 56474
rect 50818 56422 58576 56474
rect 1344 56388 58576 56422
rect 9102 56306 9154 56318
rect 15710 56306 15762 56318
rect 11554 56254 11566 56306
rect 11618 56254 11630 56306
rect 9102 56242 9154 56254
rect 15710 56242 15762 56254
rect 17390 56306 17442 56318
rect 17390 56242 17442 56254
rect 17950 56306 18002 56318
rect 17950 56242 18002 56254
rect 21646 56306 21698 56318
rect 21646 56242 21698 56254
rect 22094 56306 22146 56318
rect 25230 56306 25282 56318
rect 24434 56254 24446 56306
rect 24498 56254 24510 56306
rect 22094 56242 22146 56254
rect 25230 56242 25282 56254
rect 30382 56306 30434 56318
rect 30382 56242 30434 56254
rect 32510 56306 32562 56318
rect 32510 56242 32562 56254
rect 42366 56306 42418 56318
rect 42366 56242 42418 56254
rect 44158 56306 44210 56318
rect 44158 56242 44210 56254
rect 44494 56306 44546 56318
rect 44494 56242 44546 56254
rect 45390 56306 45442 56318
rect 45390 56242 45442 56254
rect 46398 56306 46450 56318
rect 46398 56242 46450 56254
rect 46958 56306 47010 56318
rect 46958 56242 47010 56254
rect 47294 56306 47346 56318
rect 47294 56242 47346 56254
rect 7198 56194 7250 56206
rect 7198 56130 7250 56142
rect 8430 56194 8482 56206
rect 8430 56130 8482 56142
rect 8766 56194 8818 56206
rect 8766 56130 8818 56142
rect 8878 56194 8930 56206
rect 8878 56130 8930 56142
rect 9886 56194 9938 56206
rect 16606 56194 16658 56206
rect 13010 56142 13022 56194
rect 13074 56142 13086 56194
rect 9886 56130 9938 56142
rect 16606 56130 16658 56142
rect 16718 56194 16770 56206
rect 16718 56130 16770 56142
rect 17502 56194 17554 56206
rect 42702 56194 42754 56206
rect 22306 56142 22318 56194
rect 22370 56142 22382 56194
rect 23538 56142 23550 56194
rect 23602 56142 23614 56194
rect 34290 56142 34302 56194
rect 34354 56142 34366 56194
rect 38546 56142 38558 56194
rect 38610 56142 38622 56194
rect 17502 56130 17554 56142
rect 42702 56130 42754 56142
rect 43710 56194 43762 56206
rect 43710 56130 43762 56142
rect 45166 56194 45218 56206
rect 45166 56130 45218 56142
rect 45502 56194 45554 56206
rect 45502 56130 45554 56142
rect 47854 56194 47906 56206
rect 47854 56130 47906 56142
rect 48078 56194 48130 56206
rect 48078 56130 48130 56142
rect 48974 56194 49026 56206
rect 48974 56130 49026 56142
rect 49086 56194 49138 56206
rect 49086 56130 49138 56142
rect 6974 56082 7026 56094
rect 6974 56018 7026 56030
rect 7086 56082 7138 56094
rect 7086 56018 7138 56030
rect 7310 56082 7362 56094
rect 7310 56018 7362 56030
rect 7422 56082 7474 56094
rect 7422 56018 7474 56030
rect 8318 56082 8370 56094
rect 8318 56018 8370 56030
rect 10110 56082 10162 56094
rect 10110 56018 10162 56030
rect 10334 56082 10386 56094
rect 15934 56082 15986 56094
rect 16382 56082 16434 56094
rect 25454 56082 25506 56094
rect 10546 56030 10558 56082
rect 10610 56030 10622 56082
rect 11330 56030 11342 56082
rect 11394 56030 11406 56082
rect 12226 56030 12238 56082
rect 12290 56030 12302 56082
rect 15474 56030 15486 56082
rect 15538 56030 15550 56082
rect 16146 56030 16158 56082
rect 16210 56030 16222 56082
rect 22530 56030 22542 56082
rect 22594 56030 22606 56082
rect 23986 56030 23998 56082
rect 24050 56030 24062 56082
rect 24322 56030 24334 56082
rect 24386 56030 24398 56082
rect 10334 56018 10386 56030
rect 15934 56018 15986 56030
rect 16382 56018 16434 56030
rect 25454 56018 25506 56030
rect 25902 56082 25954 56094
rect 33070 56082 33122 56094
rect 33966 56082 34018 56094
rect 43262 56082 43314 56094
rect 45054 56082 45106 56094
rect 48862 56082 48914 56094
rect 26562 56030 26574 56082
rect 26626 56030 26638 56082
rect 33506 56030 33518 56082
rect 33570 56030 33582 56082
rect 34962 56030 34974 56082
rect 35026 56030 35038 56082
rect 42914 56030 42926 56082
rect 42978 56030 42990 56082
rect 43922 56030 43934 56082
rect 43986 56030 43998 56082
rect 44706 56030 44718 56082
rect 44770 56030 44782 56082
rect 47618 56030 47630 56082
rect 47682 56030 47694 56082
rect 25902 56018 25954 56030
rect 33070 56018 33122 56030
rect 33966 56018 34018 56030
rect 43262 56018 43314 56030
rect 45054 56018 45106 56030
rect 48862 56018 48914 56030
rect 7982 55970 8034 55982
rect 15822 55970 15874 55982
rect 10434 55918 10446 55970
rect 10498 55918 10510 55970
rect 15138 55918 15150 55970
rect 15202 55918 15214 55970
rect 7982 55906 8034 55918
rect 15822 55906 15874 55918
rect 20414 55970 20466 55982
rect 20414 55906 20466 55918
rect 23102 55970 23154 55982
rect 23102 55906 23154 55918
rect 25342 55970 25394 55982
rect 25342 55906 25394 55918
rect 26350 55970 26402 55982
rect 29934 55970 29986 55982
rect 27346 55918 27358 55970
rect 27410 55918 27422 55970
rect 29474 55918 29486 55970
rect 29538 55918 29550 55970
rect 26350 55906 26402 55918
rect 29934 55906 29986 55918
rect 31838 55970 31890 55982
rect 31838 55906 31890 55918
rect 40350 55970 40402 55982
rect 40350 55906 40402 55918
rect 41022 55970 41074 55982
rect 45838 55970 45890 55982
rect 42690 55918 42702 55970
rect 42754 55918 42766 55970
rect 41022 55906 41074 55918
rect 45838 55906 45890 55918
rect 7870 55858 7922 55870
rect 7870 55794 7922 55806
rect 20302 55858 20354 55870
rect 20302 55794 20354 55806
rect 44270 55858 44322 55870
rect 44270 55794 44322 55806
rect 44382 55858 44434 55870
rect 44382 55794 44434 55806
rect 45950 55858 46002 55870
rect 45950 55794 46002 55806
rect 47742 55858 47794 55870
rect 49522 55806 49534 55858
rect 49586 55806 49598 55858
rect 47742 55794 47794 55806
rect 1344 55690 58576 55724
rect 1344 55638 4478 55690
rect 4530 55638 4582 55690
rect 4634 55638 4686 55690
rect 4738 55638 35198 55690
rect 35250 55638 35302 55690
rect 35354 55638 35406 55690
rect 35458 55638 58576 55690
rect 1344 55604 58576 55638
rect 28030 55410 28082 55422
rect 8530 55358 8542 55410
rect 8594 55358 8606 55410
rect 9314 55358 9326 55410
rect 9378 55358 9390 55410
rect 13458 55358 13470 55410
rect 13522 55358 13534 55410
rect 15586 55358 15598 55410
rect 15650 55358 15662 55410
rect 17826 55358 17838 55410
rect 17890 55358 17902 55410
rect 28030 55346 28082 55358
rect 31726 55410 31778 55422
rect 34974 55410 35026 55422
rect 43822 55410 43874 55422
rect 34402 55358 34414 55410
rect 34466 55358 34478 55410
rect 37762 55358 37774 55410
rect 37826 55358 37838 55410
rect 39890 55358 39902 55410
rect 39954 55358 39966 55410
rect 45938 55358 45950 55410
rect 46002 55358 46014 55410
rect 48066 55358 48078 55410
rect 48130 55358 48142 55410
rect 48626 55358 48638 55410
rect 48690 55358 48702 55410
rect 31726 55346 31778 55358
rect 34974 55346 35026 55358
rect 43822 55346 43874 55358
rect 19630 55298 19682 55310
rect 28142 55298 28194 55310
rect 5730 55246 5742 55298
rect 5794 55246 5806 55298
rect 12226 55246 12238 55298
rect 12290 55246 12302 55298
rect 16370 55246 16382 55298
rect 16434 55246 16446 55298
rect 26338 55246 26350 55298
rect 26402 55246 26414 55298
rect 27010 55246 27022 55298
rect 27074 55246 27086 55298
rect 19630 55234 19682 55246
rect 28142 55234 28194 55246
rect 28366 55298 28418 55310
rect 28366 55234 28418 55246
rect 28590 55298 28642 55310
rect 28590 55234 28642 55246
rect 29262 55298 29314 55310
rect 29262 55234 29314 55246
rect 32062 55298 32114 55310
rect 32062 55234 32114 55246
rect 33966 55298 34018 55310
rect 36542 55298 36594 55310
rect 43374 55298 43426 55310
rect 36194 55246 36206 55298
rect 36258 55246 36270 55298
rect 36978 55246 36990 55298
rect 37042 55246 37054 55298
rect 41570 55246 41582 55298
rect 41634 55246 41646 55298
rect 42690 55246 42702 55298
rect 42754 55246 42766 55298
rect 33966 55234 34018 55246
rect 36542 55234 36594 55246
rect 43374 55234 43426 55246
rect 43710 55298 43762 55310
rect 43710 55234 43762 55246
rect 44382 55298 44434 55310
rect 45154 55246 45166 55298
rect 45218 55246 45230 55298
rect 48738 55246 48750 55298
rect 48802 55246 48814 55298
rect 49298 55246 49310 55298
rect 49362 55246 49374 55298
rect 50418 55246 50430 55298
rect 50482 55246 50494 55298
rect 44382 55234 44434 55246
rect 19966 55186 20018 55198
rect 6402 55134 6414 55186
rect 6466 55134 6478 55186
rect 11442 55134 11454 55186
rect 11506 55134 11518 55186
rect 19966 55122 20018 55134
rect 20526 55186 20578 55198
rect 20526 55122 20578 55134
rect 20638 55186 20690 55198
rect 32398 55186 32450 55198
rect 23426 55134 23438 55186
rect 23490 55134 23502 55186
rect 27234 55134 27246 55186
rect 27298 55134 27310 55186
rect 30258 55134 30270 55186
rect 30322 55134 30334 55186
rect 20638 55122 20690 55134
rect 32398 55122 32450 55134
rect 35646 55186 35698 55198
rect 35646 55122 35698 55134
rect 41022 55186 41074 55198
rect 41022 55122 41074 55134
rect 42254 55186 42306 55198
rect 48514 55134 48526 55186
rect 48578 55134 48590 55186
rect 42254 55122 42306 55134
rect 17390 55074 17442 55086
rect 17390 55010 17442 55022
rect 18398 55074 18450 55086
rect 18398 55010 18450 55022
rect 19854 55074 19906 55086
rect 19854 55010 19906 55022
rect 20302 55074 20354 55086
rect 20302 55010 20354 55022
rect 27918 55074 27970 55086
rect 27918 55010 27970 55022
rect 29150 55074 29202 55086
rect 29150 55010 29202 55022
rect 29934 55074 29986 55086
rect 29934 55010 29986 55022
rect 30718 55074 30770 55086
rect 30718 55010 30770 55022
rect 31166 55074 31218 55086
rect 31166 55010 31218 55022
rect 35310 55074 35362 55086
rect 35310 55010 35362 55022
rect 35870 55074 35922 55086
rect 35870 55010 35922 55022
rect 35982 55074 36034 55086
rect 35982 55010 36034 55022
rect 41134 55074 41186 55086
rect 41134 55010 41186 55022
rect 41806 55074 41858 55086
rect 41806 55010 41858 55022
rect 42142 55074 42194 55086
rect 42142 55010 42194 55022
rect 42366 55074 42418 55086
rect 43934 55074 43986 55086
rect 43026 55022 43038 55074
rect 43090 55022 43102 55074
rect 42366 55010 42418 55022
rect 43934 55010 43986 55022
rect 49870 55074 49922 55086
rect 49870 55010 49922 55022
rect 49982 55074 50034 55086
rect 49982 55010 50034 55022
rect 50094 55074 50146 55086
rect 50094 55010 50146 55022
rect 1344 54906 58576 54940
rect 1344 54854 19838 54906
rect 19890 54854 19942 54906
rect 19994 54854 20046 54906
rect 20098 54854 50558 54906
rect 50610 54854 50662 54906
rect 50714 54854 50766 54906
rect 50818 54854 58576 54906
rect 1344 54820 58576 54854
rect 6638 54738 6690 54750
rect 6638 54674 6690 54686
rect 6750 54738 6802 54750
rect 6750 54674 6802 54686
rect 6974 54738 7026 54750
rect 6974 54674 7026 54686
rect 7422 54738 7474 54750
rect 7422 54674 7474 54686
rect 7646 54738 7698 54750
rect 15598 54738 15650 54750
rect 8642 54686 8654 54738
rect 8706 54686 8718 54738
rect 7646 54674 7698 54686
rect 15598 54674 15650 54686
rect 24558 54738 24610 54750
rect 24558 54674 24610 54686
rect 26462 54738 26514 54750
rect 26462 54674 26514 54686
rect 31166 54738 31218 54750
rect 34078 54738 34130 54750
rect 31826 54686 31838 54738
rect 31890 54686 31902 54738
rect 31166 54674 31218 54686
rect 34078 54674 34130 54686
rect 34414 54738 34466 54750
rect 34414 54674 34466 54686
rect 36318 54738 36370 54750
rect 36318 54674 36370 54686
rect 47966 54738 48018 54750
rect 47966 54674 48018 54686
rect 2046 54626 2098 54638
rect 2046 54562 2098 54574
rect 7758 54626 7810 54638
rect 7758 54562 7810 54574
rect 15150 54626 15202 54638
rect 15150 54562 15202 54574
rect 15262 54626 15314 54638
rect 26798 54626 26850 54638
rect 16482 54574 16494 54626
rect 16546 54574 16558 54626
rect 26114 54574 26126 54626
rect 26178 54574 26190 54626
rect 15262 54562 15314 54574
rect 26798 54562 26850 54574
rect 26910 54626 26962 54638
rect 26910 54562 26962 54574
rect 29150 54626 29202 54638
rect 29150 54562 29202 54574
rect 29486 54626 29538 54638
rect 29486 54562 29538 54574
rect 29822 54626 29874 54638
rect 29822 54562 29874 54574
rect 30158 54626 30210 54638
rect 30158 54562 30210 54574
rect 30494 54626 30546 54638
rect 35086 54626 35138 54638
rect 48190 54626 48242 54638
rect 34738 54574 34750 54626
rect 34802 54574 34814 54626
rect 37538 54574 37550 54626
rect 37602 54574 37614 54626
rect 41682 54574 41694 54626
rect 41746 54574 41758 54626
rect 50866 54574 50878 54626
rect 50930 54574 50942 54626
rect 30494 54562 30546 54574
rect 35086 54562 35138 54574
rect 48190 54562 48242 54574
rect 1710 54514 1762 54526
rect 14926 54514 14978 54526
rect 7186 54462 7198 54514
rect 7250 54462 7262 54514
rect 8866 54462 8878 54514
rect 8930 54462 8942 54514
rect 9650 54462 9662 54514
rect 9714 54462 9726 54514
rect 1710 54450 1762 54462
rect 14926 54450 14978 54462
rect 15710 54514 15762 54526
rect 24446 54514 24498 54526
rect 16258 54462 16270 54514
rect 16322 54462 16334 54514
rect 23426 54462 23438 54514
rect 23490 54462 23502 54514
rect 15710 54450 15762 54462
rect 24446 54450 24498 54462
rect 24782 54514 24834 54526
rect 24782 54450 24834 54462
rect 25678 54514 25730 54526
rect 32174 54514 32226 54526
rect 35646 54514 35698 54526
rect 30930 54462 30942 54514
rect 30994 54462 31006 54514
rect 35298 54462 35310 54514
rect 35362 54462 35374 54514
rect 25678 54450 25730 54462
rect 32174 54450 32226 54462
rect 35646 54450 35698 54462
rect 35758 54514 35810 54526
rect 35758 54450 35810 54462
rect 36206 54514 36258 54526
rect 36206 54450 36258 54462
rect 36430 54514 36482 54526
rect 36754 54462 36766 54514
rect 36818 54462 36830 54514
rect 41010 54462 41022 54514
rect 41074 54462 41086 54514
rect 44146 54462 44158 54514
rect 44210 54462 44222 54514
rect 47618 54462 47630 54514
rect 47682 54462 47694 54514
rect 51650 54462 51662 54514
rect 51714 54462 51726 54514
rect 36430 54450 36482 54462
rect 2494 54402 2546 54414
rect 17502 54402 17554 54414
rect 6626 54350 6638 54402
rect 6690 54350 6702 54402
rect 10322 54350 10334 54402
rect 10386 54350 10398 54402
rect 12450 54350 12462 54402
rect 12514 54350 12526 54402
rect 2494 54338 2546 54350
rect 17502 54338 17554 54350
rect 18062 54402 18114 54414
rect 27470 54402 27522 54414
rect 21298 54350 21310 54402
rect 21362 54350 21374 54402
rect 18062 54338 18114 54350
rect 27470 54338 27522 54350
rect 27918 54402 27970 54414
rect 27918 54338 27970 54350
rect 28366 54402 28418 54414
rect 28366 54338 28418 54350
rect 33294 54402 33346 54414
rect 48078 54402 48130 54414
rect 39666 54350 39678 54402
rect 39730 54350 39742 54402
rect 43810 54350 43822 54402
rect 43874 54350 43886 54402
rect 44930 54350 44942 54402
rect 44994 54350 45006 54402
rect 47058 54350 47070 54402
rect 47122 54350 47134 54402
rect 48738 54350 48750 54402
rect 48802 54350 48814 54402
rect 33294 54338 33346 54350
rect 48078 54338 48130 54350
rect 25342 54290 25394 54302
rect 25342 54226 25394 54238
rect 25454 54290 25506 54302
rect 25454 54226 25506 54238
rect 25790 54290 25842 54302
rect 25790 54226 25842 54238
rect 26910 54290 26962 54302
rect 26910 54226 26962 54238
rect 33406 54290 33458 54302
rect 33406 54226 33458 54238
rect 35422 54290 35474 54302
rect 35422 54226 35474 54238
rect 1344 54122 58576 54156
rect 1344 54070 4478 54122
rect 4530 54070 4582 54122
rect 4634 54070 4686 54122
rect 4738 54070 35198 54122
rect 35250 54070 35302 54122
rect 35354 54070 35406 54122
rect 35458 54070 58576 54122
rect 1344 54036 58576 54070
rect 44942 53954 44994 53966
rect 44942 53890 44994 53902
rect 49534 53954 49586 53966
rect 49534 53890 49586 53902
rect 49758 53954 49810 53966
rect 49758 53890 49810 53902
rect 49870 53954 49922 53966
rect 49870 53890 49922 53902
rect 10446 53842 10498 53854
rect 26686 53842 26738 53854
rect 6626 53790 6638 53842
rect 6690 53790 6702 53842
rect 20738 53790 20750 53842
rect 20802 53790 20814 53842
rect 22082 53790 22094 53842
rect 22146 53790 22158 53842
rect 24210 53790 24222 53842
rect 24274 53790 24286 53842
rect 25330 53790 25342 53842
rect 25394 53790 25406 53842
rect 10446 53778 10498 53790
rect 26686 53778 26738 53790
rect 27918 53842 27970 53854
rect 34974 53842 35026 53854
rect 31602 53790 31614 53842
rect 31666 53790 31678 53842
rect 27918 53778 27970 53790
rect 34974 53778 35026 53790
rect 37438 53842 37490 53854
rect 49422 53842 49474 53854
rect 47842 53790 47854 53842
rect 47906 53790 47918 53842
rect 48626 53790 48638 53842
rect 48690 53790 48702 53842
rect 37438 53778 37490 53790
rect 49422 53778 49474 53790
rect 6750 53730 6802 53742
rect 6750 53666 6802 53678
rect 6974 53730 7026 53742
rect 6974 53666 7026 53678
rect 7422 53730 7474 53742
rect 7422 53666 7474 53678
rect 7758 53730 7810 53742
rect 7758 53666 7810 53678
rect 8206 53730 8258 53742
rect 10222 53730 10274 53742
rect 9650 53678 9662 53730
rect 9714 53678 9726 53730
rect 8206 53666 8258 53678
rect 10222 53666 10274 53678
rect 10558 53730 10610 53742
rect 11118 53730 11170 53742
rect 10770 53678 10782 53730
rect 10834 53678 10846 53730
rect 10558 53666 10610 53678
rect 11118 53666 11170 53678
rect 11230 53730 11282 53742
rect 26126 53730 26178 53742
rect 17938 53678 17950 53730
rect 18002 53678 18014 53730
rect 18610 53678 18622 53730
rect 18674 53678 18686 53730
rect 21298 53678 21310 53730
rect 21362 53678 21374 53730
rect 24434 53678 24446 53730
rect 24498 53678 24510 53730
rect 25554 53678 25566 53730
rect 25618 53678 25630 53730
rect 11230 53666 11282 53678
rect 26126 53666 26178 53678
rect 26798 53730 26850 53742
rect 26798 53666 26850 53678
rect 27470 53730 27522 53742
rect 27470 53666 27522 53678
rect 27694 53730 27746 53742
rect 35086 53730 35138 53742
rect 28018 53678 28030 53730
rect 28082 53678 28094 53730
rect 33730 53678 33742 53730
rect 33794 53678 33806 53730
rect 34402 53678 34414 53730
rect 34466 53678 34478 53730
rect 27694 53666 27746 53678
rect 35086 53666 35138 53678
rect 35534 53730 35586 53742
rect 35534 53666 35586 53678
rect 35758 53730 35810 53742
rect 35758 53666 35810 53678
rect 35982 53730 36034 53742
rect 35982 53666 36034 53678
rect 36430 53730 36482 53742
rect 36430 53666 36482 53678
rect 37886 53730 37938 53742
rect 37886 53666 37938 53678
rect 38222 53730 38274 53742
rect 38222 53666 38274 53678
rect 40126 53730 40178 53742
rect 40126 53666 40178 53678
rect 40798 53730 40850 53742
rect 40798 53666 40850 53678
rect 42478 53730 42530 53742
rect 42478 53666 42530 53678
rect 43038 53730 43090 53742
rect 43038 53666 43090 53678
rect 43934 53730 43986 53742
rect 46734 53730 46786 53742
rect 50542 53730 50594 53742
rect 44258 53678 44270 53730
rect 44322 53678 44334 53730
rect 47058 53678 47070 53730
rect 47122 53678 47134 53730
rect 47730 53678 47742 53730
rect 47794 53678 47806 53730
rect 48514 53678 48526 53730
rect 48578 53678 48590 53730
rect 43934 53666 43986 53678
rect 46734 53666 46786 53678
rect 50542 53666 50594 53678
rect 1710 53618 1762 53630
rect 1710 53554 1762 53566
rect 7198 53618 7250 53630
rect 16270 53618 16322 53630
rect 27134 53618 27186 53630
rect 9426 53566 9438 53618
rect 9490 53566 9502 53618
rect 25218 53566 25230 53618
rect 25282 53566 25294 53618
rect 7198 53554 7250 53566
rect 16270 53554 16322 53566
rect 27134 53554 27186 53566
rect 27246 53618 27298 53630
rect 27246 53554 27298 53566
rect 30046 53618 30098 53630
rect 37102 53618 37154 53630
rect 30370 53566 30382 53618
rect 30434 53566 30446 53618
rect 30046 53554 30098 53566
rect 37102 53554 37154 53566
rect 41358 53618 41410 53630
rect 41358 53554 41410 53566
rect 41694 53618 41746 53630
rect 41694 53554 41746 53566
rect 42702 53618 42754 53630
rect 42702 53554 42754 53566
rect 43262 53618 43314 53630
rect 43262 53554 43314 53566
rect 43374 53618 43426 53630
rect 43374 53554 43426 53566
rect 43822 53618 43874 53630
rect 43822 53554 43874 53566
rect 44830 53618 44882 53630
rect 44830 53554 44882 53566
rect 50206 53618 50258 53630
rect 50206 53554 50258 53566
rect 50318 53618 50370 53630
rect 50318 53554 50370 53566
rect 50878 53618 50930 53630
rect 50878 53554 50930 53566
rect 2046 53506 2098 53518
rect 2046 53442 2098 53454
rect 2494 53506 2546 53518
rect 2494 53442 2546 53454
rect 6638 53506 6690 53518
rect 6638 53442 6690 53454
rect 7646 53506 7698 53518
rect 7646 53442 7698 53454
rect 8094 53506 8146 53518
rect 8094 53442 8146 53454
rect 10334 53506 10386 53518
rect 10334 53442 10386 53454
rect 16382 53506 16434 53518
rect 16382 53442 16434 53454
rect 16606 53506 16658 53518
rect 16606 53442 16658 53454
rect 16942 53506 16994 53518
rect 16942 53442 16994 53454
rect 17614 53506 17666 53518
rect 17614 53442 17666 53454
rect 26574 53506 26626 53518
rect 26574 53442 26626 53454
rect 28254 53506 28306 53518
rect 28254 53442 28306 53454
rect 29710 53506 29762 53518
rect 29710 53442 29762 53454
rect 34862 53506 34914 53518
rect 34862 53442 34914 53454
rect 35870 53506 35922 53518
rect 35870 53442 35922 53454
rect 37326 53506 37378 53518
rect 37326 53442 37378 53454
rect 37550 53506 37602 53518
rect 37550 53442 37602 53454
rect 37998 53506 38050 53518
rect 41022 53506 41074 53518
rect 40450 53454 40462 53506
rect 40514 53454 40526 53506
rect 37998 53442 38050 53454
rect 41022 53442 41074 53454
rect 41246 53506 41298 53518
rect 41246 53442 41298 53454
rect 41806 53506 41858 53518
rect 41806 53442 41858 53454
rect 42030 53506 42082 53518
rect 42030 53442 42082 53454
rect 42254 53506 42306 53518
rect 42254 53442 42306 53454
rect 42366 53506 42418 53518
rect 42366 53442 42418 53454
rect 43710 53506 43762 53518
rect 43710 53442 43762 53454
rect 46510 53506 46562 53518
rect 46510 53442 46562 53454
rect 46622 53506 46674 53518
rect 46622 53442 46674 53454
rect 1344 53338 58576 53372
rect 1344 53286 19838 53338
rect 19890 53286 19942 53338
rect 19994 53286 20046 53338
rect 20098 53286 50558 53338
rect 50610 53286 50662 53338
rect 50714 53286 50766 53338
rect 50818 53286 58576 53338
rect 1344 53252 58576 53286
rect 11678 53170 11730 53182
rect 8418 53118 8430 53170
rect 8482 53118 8494 53170
rect 9986 53118 9998 53170
rect 10050 53118 10062 53170
rect 11678 53106 11730 53118
rect 14478 53170 14530 53182
rect 14478 53106 14530 53118
rect 15598 53170 15650 53182
rect 15598 53106 15650 53118
rect 22990 53170 23042 53182
rect 22990 53106 23042 53118
rect 23326 53170 23378 53182
rect 27246 53170 27298 53182
rect 24658 53118 24670 53170
rect 24722 53118 24734 53170
rect 26674 53118 26686 53170
rect 26738 53118 26750 53170
rect 23326 53106 23378 53118
rect 27246 53106 27298 53118
rect 28366 53170 28418 53182
rect 28366 53106 28418 53118
rect 30046 53170 30098 53182
rect 30046 53106 30098 53118
rect 30270 53170 30322 53182
rect 30270 53106 30322 53118
rect 30830 53170 30882 53182
rect 30830 53106 30882 53118
rect 31054 53170 31106 53182
rect 31054 53106 31106 53118
rect 32286 53170 32338 53182
rect 32286 53106 32338 53118
rect 33070 53170 33122 53182
rect 33070 53106 33122 53118
rect 35198 53170 35250 53182
rect 35198 53106 35250 53118
rect 35422 53170 35474 53182
rect 35422 53106 35474 53118
rect 35534 53170 35586 53182
rect 35534 53106 35586 53118
rect 36430 53170 36482 53182
rect 36430 53106 36482 53118
rect 36766 53170 36818 53182
rect 36766 53106 36818 53118
rect 37438 53170 37490 53182
rect 37438 53106 37490 53118
rect 46958 53170 47010 53182
rect 46958 53106 47010 53118
rect 48302 53170 48354 53182
rect 49074 53118 49086 53170
rect 49138 53118 49150 53170
rect 48302 53106 48354 53118
rect 2046 53058 2098 53070
rect 13582 53058 13634 53070
rect 14926 53058 14978 53070
rect 5282 53006 5294 53058
rect 5346 53006 5358 53058
rect 7746 53006 7758 53058
rect 7810 53006 7822 53058
rect 13906 53006 13918 53058
rect 13970 53006 13982 53058
rect 2046 52994 2098 53006
rect 13582 52994 13634 53006
rect 14926 52994 14978 53006
rect 15934 53058 15986 53070
rect 20974 53058 21026 53070
rect 16482 53006 16494 53058
rect 16546 53006 16558 53058
rect 15934 52994 15986 53006
rect 20974 52994 21026 53006
rect 23214 53058 23266 53070
rect 23214 52994 23266 53006
rect 24110 53058 24162 53070
rect 29038 53058 29090 53070
rect 34526 53058 34578 53070
rect 26002 53006 26014 53058
rect 26066 53006 26078 53058
rect 33394 53006 33406 53058
rect 33458 53006 33470 53058
rect 24110 52994 24162 53006
rect 29038 52994 29090 53006
rect 34526 52994 34578 53006
rect 34638 53058 34690 53070
rect 34638 52994 34690 53006
rect 36542 53058 36594 53070
rect 36542 52994 36594 53006
rect 39454 53058 39506 53070
rect 39454 52994 39506 53006
rect 42590 53058 42642 53070
rect 43150 53058 43202 53070
rect 42590 52994 42642 53006
rect 42814 53002 42866 53014
rect 1710 52946 1762 52958
rect 8094 52946 8146 52958
rect 4610 52894 4622 52946
rect 4674 52894 4686 52946
rect 1710 52882 1762 52894
rect 8094 52882 8146 52894
rect 8766 52946 8818 52958
rect 12014 52946 12066 52958
rect 9762 52894 9774 52946
rect 9826 52894 9838 52946
rect 8766 52882 8818 52894
rect 12014 52882 12066 52894
rect 14366 52946 14418 52958
rect 14366 52882 14418 52894
rect 14702 52946 14754 52958
rect 14702 52882 14754 52894
rect 15374 52946 15426 52958
rect 15374 52882 15426 52894
rect 15486 52946 15538 52958
rect 15486 52882 15538 52894
rect 15710 52946 15762 52958
rect 21198 52946 21250 52958
rect 16706 52894 16718 52946
rect 16770 52894 16782 52946
rect 17490 52894 17502 52946
rect 17554 52894 17566 52946
rect 20738 52894 20750 52946
rect 20802 52894 20814 52946
rect 15710 52882 15762 52894
rect 21198 52882 21250 52894
rect 21646 52946 21698 52958
rect 21646 52882 21698 52894
rect 21870 52946 21922 52958
rect 23998 52946 24050 52958
rect 22754 52894 22766 52946
rect 22818 52894 22830 52946
rect 21870 52882 21922 52894
rect 23998 52882 24050 52894
rect 24222 52946 24274 52958
rect 24222 52882 24274 52894
rect 25678 52946 25730 52958
rect 25678 52882 25730 52894
rect 26350 52946 26402 52958
rect 26350 52882 26402 52894
rect 27470 52946 27522 52958
rect 27470 52882 27522 52894
rect 27918 52946 27970 52958
rect 27918 52882 27970 52894
rect 28478 52946 28530 52958
rect 28478 52882 28530 52894
rect 28814 52946 28866 52958
rect 28814 52882 28866 52894
rect 29486 52946 29538 52958
rect 29486 52882 29538 52894
rect 30606 52946 30658 52958
rect 30606 52882 30658 52894
rect 31390 52946 31442 52958
rect 31390 52882 31442 52894
rect 34862 52946 34914 52958
rect 34862 52882 34914 52894
rect 37102 52946 37154 52958
rect 37102 52882 37154 52894
rect 37214 52946 37266 52958
rect 37214 52882 37266 52894
rect 37550 52946 37602 52958
rect 37550 52882 37602 52894
rect 39006 52946 39058 52958
rect 39006 52882 39058 52894
rect 39678 52946 39730 52958
rect 39678 52882 39730 52894
rect 42254 52946 42306 52958
rect 43150 52994 43202 53006
rect 45390 53058 45442 53070
rect 45390 52994 45442 53006
rect 45950 53058 46002 53070
rect 45950 52994 46002 53006
rect 46062 53058 46114 53070
rect 46062 52994 46114 53006
rect 47966 53058 48018 53070
rect 47966 52994 48018 53006
rect 48078 53058 48130 53070
rect 48078 52994 48130 53006
rect 42814 52938 42866 52950
rect 45714 52894 45726 52946
rect 45778 52894 45790 52946
rect 47170 52894 47182 52946
rect 47234 52894 47246 52946
rect 49298 52894 49310 52946
rect 49362 52894 49374 52946
rect 42254 52882 42306 52894
rect 2494 52834 2546 52846
rect 14590 52834 14642 52846
rect 21758 52834 21810 52846
rect 7410 52782 7422 52834
rect 7474 52782 7486 52834
rect 18162 52782 18174 52834
rect 18226 52782 18238 52834
rect 20290 52782 20302 52834
rect 20354 52782 20366 52834
rect 2494 52770 2546 52782
rect 14590 52770 14642 52782
rect 21758 52770 21810 52782
rect 25342 52834 25394 52846
rect 25342 52770 25394 52782
rect 27358 52834 27410 52846
rect 27358 52770 27410 52782
rect 28926 52834 28978 52846
rect 39230 52834 39282 52846
rect 29474 52782 29486 52834
rect 29538 52831 29550 52834
rect 29810 52831 29822 52834
rect 29538 52785 29822 52831
rect 29538 52782 29550 52785
rect 29810 52782 29822 52785
rect 29874 52782 29886 52834
rect 31826 52782 31838 52834
rect 31890 52782 31902 52834
rect 28926 52770 28978 52782
rect 39230 52770 39282 52782
rect 42478 52834 42530 52846
rect 47282 52782 47294 52834
rect 47346 52782 47358 52834
rect 42478 52770 42530 52782
rect 28366 52722 28418 52734
rect 28366 52658 28418 52670
rect 29934 52722 29986 52734
rect 29934 52658 29986 52670
rect 30718 52722 30770 52734
rect 30718 52658 30770 52670
rect 34526 52722 34578 52734
rect 34526 52658 34578 52670
rect 43262 52722 43314 52734
rect 46498 52670 46510 52722
rect 46562 52670 46574 52722
rect 43262 52658 43314 52670
rect 1344 52554 58576 52588
rect 1344 52502 4478 52554
rect 4530 52502 4582 52554
rect 4634 52502 4686 52554
rect 4738 52502 35198 52554
rect 35250 52502 35302 52554
rect 35354 52502 35406 52554
rect 35458 52502 58576 52554
rect 1344 52468 58576 52502
rect 8094 52386 8146 52398
rect 8094 52322 8146 52334
rect 11902 52386 11954 52398
rect 11902 52322 11954 52334
rect 19182 52386 19234 52398
rect 19182 52322 19234 52334
rect 20526 52386 20578 52398
rect 25342 52386 25394 52398
rect 21186 52334 21198 52386
rect 21250 52383 21262 52386
rect 21746 52383 21758 52386
rect 21250 52337 21758 52383
rect 21250 52334 21262 52337
rect 21746 52334 21758 52337
rect 21810 52334 21822 52386
rect 20526 52322 20578 52334
rect 25342 52322 25394 52334
rect 29262 52386 29314 52398
rect 29262 52322 29314 52334
rect 20078 52274 20130 52286
rect 6626 52222 6638 52274
rect 6690 52222 6702 52274
rect 15250 52222 15262 52274
rect 15314 52222 15326 52274
rect 17378 52222 17390 52274
rect 17442 52222 17454 52274
rect 20078 52210 20130 52222
rect 20638 52274 20690 52286
rect 20638 52210 20690 52222
rect 21422 52274 21474 52286
rect 23550 52274 23602 52286
rect 22418 52222 22430 52274
rect 22482 52222 22494 52274
rect 21422 52210 21474 52222
rect 23550 52210 23602 52222
rect 25230 52274 25282 52286
rect 33294 52274 33346 52286
rect 28578 52222 28590 52274
rect 28642 52222 28654 52274
rect 25230 52210 25282 52222
rect 33294 52210 33346 52222
rect 34862 52274 34914 52286
rect 34862 52210 34914 52222
rect 38894 52274 38946 52286
rect 45490 52222 45502 52274
rect 45554 52222 45566 52274
rect 38894 52210 38946 52222
rect 1710 52162 1762 52174
rect 1710 52098 1762 52110
rect 2494 52162 2546 52174
rect 6750 52162 6802 52174
rect 6514 52110 6526 52162
rect 6578 52110 6590 52162
rect 2494 52098 2546 52110
rect 6750 52098 6802 52110
rect 6974 52162 7026 52174
rect 6974 52098 7026 52110
rect 7086 52162 7138 52174
rect 7086 52098 7138 52110
rect 7422 52162 7474 52174
rect 7422 52098 7474 52110
rect 8206 52162 8258 52174
rect 8206 52098 8258 52110
rect 11454 52162 11506 52174
rect 11454 52098 11506 52110
rect 12574 52162 12626 52174
rect 12574 52098 12626 52110
rect 13022 52162 13074 52174
rect 18286 52162 18338 52174
rect 13906 52110 13918 52162
rect 13970 52110 13982 52162
rect 14578 52110 14590 52162
rect 14642 52110 14654 52162
rect 13022 52098 13074 52110
rect 18286 52098 18338 52110
rect 19406 52162 19458 52174
rect 20190 52162 20242 52174
rect 29038 52162 29090 52174
rect 19618 52110 19630 52162
rect 19682 52110 19694 52162
rect 22194 52110 22206 52162
rect 22258 52110 22270 52162
rect 22866 52110 22878 52162
rect 22930 52110 22942 52162
rect 24210 52110 24222 52162
rect 24274 52110 24286 52162
rect 25666 52110 25678 52162
rect 25730 52110 25742 52162
rect 19406 52098 19458 52110
rect 20190 52098 20242 52110
rect 29038 52098 29090 52110
rect 30158 52162 30210 52174
rect 30158 52098 30210 52110
rect 30718 52162 30770 52174
rect 30718 52098 30770 52110
rect 32398 52162 32450 52174
rect 32398 52098 32450 52110
rect 33518 52162 33570 52174
rect 33518 52098 33570 52110
rect 38222 52162 38274 52174
rect 38222 52098 38274 52110
rect 38446 52162 38498 52174
rect 38446 52098 38498 52110
rect 39790 52162 39842 52174
rect 39790 52098 39842 52110
rect 39902 52162 39954 52174
rect 39902 52098 39954 52110
rect 40014 52162 40066 52174
rect 40014 52098 40066 52110
rect 44270 52162 44322 52174
rect 49410 52110 49422 52162
rect 49474 52110 49486 52162
rect 44270 52098 44322 52110
rect 7646 52050 7698 52062
rect 7646 51986 7698 51998
rect 7758 52050 7810 52062
rect 7758 51986 7810 51998
rect 11118 52050 11170 52062
rect 11118 51986 11170 51998
rect 12014 52050 12066 52062
rect 19070 52050 19122 52062
rect 14130 51998 14142 52050
rect 14194 51998 14206 52050
rect 12014 51986 12066 51998
rect 19070 51986 19122 51998
rect 19966 52050 20018 52062
rect 23998 52050 24050 52062
rect 29374 52050 29426 52062
rect 23090 51998 23102 52050
rect 23154 51998 23166 52050
rect 26450 51998 26462 52050
rect 26514 51998 26526 52050
rect 19966 51986 20018 51998
rect 23998 51986 24050 51998
rect 29374 51986 29426 51998
rect 29598 52050 29650 52062
rect 29598 51986 29650 51998
rect 30382 52050 30434 52062
rect 30382 51986 30434 51998
rect 30942 52050 30994 52062
rect 30942 51986 30994 51998
rect 31054 52050 31106 52062
rect 31054 51986 31106 51998
rect 32734 52050 32786 52062
rect 38670 52050 38722 52062
rect 33842 51998 33854 52050
rect 33906 51998 33918 52050
rect 32734 51986 32786 51998
rect 38670 51986 38722 51998
rect 39006 52050 39058 52062
rect 39006 51986 39058 51998
rect 2046 51938 2098 51950
rect 2046 51874 2098 51886
rect 11902 51938 11954 51950
rect 11902 51874 11954 51886
rect 17950 51938 18002 51950
rect 17950 51874 18002 51886
rect 18398 51938 18450 51950
rect 18398 51874 18450 51886
rect 18622 51938 18674 51950
rect 18622 51874 18674 51886
rect 18846 51938 18898 51950
rect 18846 51874 18898 51886
rect 29934 51938 29986 51950
rect 29934 51874 29986 51886
rect 30046 51938 30098 51950
rect 30046 51874 30098 51886
rect 32622 51938 32674 51950
rect 32622 51874 32674 51886
rect 34750 51938 34802 51950
rect 39330 51886 39342 51938
rect 39394 51886 39406 51938
rect 34750 51874 34802 51886
rect 1344 51770 58576 51804
rect 1344 51718 19838 51770
rect 19890 51718 19942 51770
rect 19994 51718 20046 51770
rect 20098 51718 50558 51770
rect 50610 51718 50662 51770
rect 50714 51718 50766 51770
rect 50818 51718 58576 51770
rect 1344 51684 58576 51718
rect 16270 51602 16322 51614
rect 16270 51538 16322 51550
rect 16718 51602 16770 51614
rect 16718 51538 16770 51550
rect 17838 51602 17890 51614
rect 17838 51538 17890 51550
rect 19742 51602 19794 51614
rect 19742 51538 19794 51550
rect 20526 51602 20578 51614
rect 20526 51538 20578 51550
rect 28478 51602 28530 51614
rect 28478 51538 28530 51550
rect 36430 51602 36482 51614
rect 36430 51538 36482 51550
rect 38558 51602 38610 51614
rect 38558 51538 38610 51550
rect 39006 51602 39058 51614
rect 39006 51538 39058 51550
rect 45054 51602 45106 51614
rect 45054 51538 45106 51550
rect 47742 51602 47794 51614
rect 47742 51538 47794 51550
rect 48078 51602 48130 51614
rect 48078 51538 48130 51550
rect 48862 51602 48914 51614
rect 48862 51538 48914 51550
rect 49758 51602 49810 51614
rect 49758 51538 49810 51550
rect 2046 51490 2098 51502
rect 9886 51490 9938 51502
rect 5282 51438 5294 51490
rect 5346 51438 5358 51490
rect 2046 51426 2098 51438
rect 9886 51426 9938 51438
rect 16830 51490 16882 51502
rect 19966 51490 20018 51502
rect 18050 51438 18062 51490
rect 18114 51438 18126 51490
rect 16830 51426 16882 51438
rect 19966 51426 20018 51438
rect 21198 51490 21250 51502
rect 21198 51426 21250 51438
rect 22878 51490 22930 51502
rect 22878 51426 22930 51438
rect 23214 51490 23266 51502
rect 28590 51490 28642 51502
rect 37998 51490 38050 51502
rect 44830 51490 44882 51502
rect 26002 51438 26014 51490
rect 26066 51438 26078 51490
rect 33954 51438 33966 51490
rect 34018 51438 34030 51490
rect 43362 51438 43374 51490
rect 43426 51438 43438 51490
rect 23214 51426 23266 51438
rect 28590 51426 28642 51438
rect 37998 51426 38050 51438
rect 44830 51426 44882 51438
rect 45166 51490 45218 51502
rect 45166 51426 45218 51438
rect 45390 51490 45442 51502
rect 47518 51490 47570 51502
rect 46722 51438 46734 51490
rect 46786 51438 46798 51490
rect 45390 51426 45442 51438
rect 47518 51426 47570 51438
rect 48750 51490 48802 51502
rect 48750 51426 48802 51438
rect 49310 51490 49362 51502
rect 49310 51426 49362 51438
rect 1710 51378 1762 51390
rect 16046 51378 16098 51390
rect 4610 51326 4622 51378
rect 4674 51326 4686 51378
rect 10098 51326 10110 51378
rect 10162 51326 10174 51378
rect 15810 51326 15822 51378
rect 15874 51326 15886 51378
rect 1710 51314 1762 51326
rect 16046 51314 16098 51326
rect 16382 51378 16434 51390
rect 19406 51378 19458 51390
rect 18274 51326 18286 51378
rect 18338 51326 18350 51378
rect 16382 51314 16434 51326
rect 19406 51314 19458 51326
rect 20302 51378 20354 51390
rect 20302 51314 20354 51326
rect 20638 51378 20690 51390
rect 20638 51314 20690 51326
rect 20750 51378 20802 51390
rect 20750 51314 20802 51326
rect 21422 51378 21474 51390
rect 21422 51314 21474 51326
rect 21870 51378 21922 51390
rect 21870 51314 21922 51326
rect 22094 51378 22146 51390
rect 22094 51314 22146 51326
rect 22542 51378 22594 51390
rect 22542 51314 22594 51326
rect 23326 51378 23378 51390
rect 23326 51314 23378 51326
rect 23438 51378 23490 51390
rect 23438 51314 23490 51326
rect 23774 51378 23826 51390
rect 23774 51314 23826 51326
rect 24222 51378 24274 51390
rect 36766 51378 36818 51390
rect 25218 51326 25230 51378
rect 25282 51326 25294 51378
rect 29026 51326 29038 51378
rect 29090 51326 29102 51378
rect 33170 51326 33182 51378
rect 33234 51326 33246 51378
rect 24222 51314 24274 51326
rect 36766 51314 36818 51326
rect 37886 51378 37938 51390
rect 37886 51314 37938 51326
rect 38782 51378 38834 51390
rect 38782 51314 38834 51326
rect 38894 51378 38946 51390
rect 47406 51378 47458 51390
rect 39442 51326 39454 51378
rect 39506 51326 39518 51378
rect 39890 51326 39902 51378
rect 39954 51326 39966 51378
rect 44146 51326 44158 51378
rect 44210 51326 44222 51378
rect 46162 51326 46174 51378
rect 46226 51326 46238 51378
rect 46946 51326 46958 51378
rect 47010 51326 47022 51378
rect 38894 51314 38946 51326
rect 47406 51314 47458 51326
rect 47966 51378 48018 51390
rect 47966 51314 48018 51326
rect 48974 51378 49026 51390
rect 48974 51314 49026 51326
rect 2494 51266 2546 51278
rect 2494 51202 2546 51214
rect 2942 51266 2994 51278
rect 19294 51266 19346 51278
rect 7410 51214 7422 51266
rect 7474 51214 7486 51266
rect 11778 51214 11790 51266
rect 11842 51214 11854 51266
rect 2942 51202 2994 51214
rect 19294 51202 19346 51214
rect 19630 51266 19682 51278
rect 19630 51202 19682 51214
rect 21310 51266 21362 51278
rect 37214 51266 37266 51278
rect 28130 51214 28142 51266
rect 28194 51214 28206 51266
rect 29698 51214 29710 51266
rect 29762 51214 29774 51266
rect 31826 51214 31838 51266
rect 31890 51214 31902 51266
rect 36082 51214 36094 51266
rect 36146 51214 36158 51266
rect 41234 51214 41246 51266
rect 41298 51214 41310 51266
rect 46386 51214 46398 51266
rect 46450 51214 46462 51266
rect 21310 51202 21362 51214
rect 37214 51202 37266 51214
rect 37998 51154 38050 51166
rect 48078 51154 48130 51166
rect 39442 51102 39454 51154
rect 39506 51102 39518 51154
rect 37998 51090 38050 51102
rect 48078 51090 48130 51102
rect 1344 50986 58576 51020
rect 1344 50934 4478 50986
rect 4530 50934 4582 50986
rect 4634 50934 4686 50986
rect 4738 50934 35198 50986
rect 35250 50934 35302 50986
rect 35354 50934 35406 50986
rect 35458 50934 58576 50986
rect 1344 50900 58576 50934
rect 7086 50818 7138 50830
rect 7086 50754 7138 50766
rect 14478 50818 14530 50830
rect 29934 50818 29986 50830
rect 22754 50766 22766 50818
rect 22818 50766 22830 50818
rect 14478 50754 14530 50766
rect 29934 50754 29986 50766
rect 36542 50818 36594 50830
rect 36542 50754 36594 50766
rect 41806 50818 41858 50830
rect 41806 50754 41858 50766
rect 14590 50706 14642 50718
rect 23326 50706 23378 50718
rect 10882 50654 10894 50706
rect 10946 50654 10958 50706
rect 16594 50654 16606 50706
rect 16658 50654 16670 50706
rect 14590 50642 14642 50654
rect 23326 50642 23378 50654
rect 30046 50706 30098 50718
rect 30046 50642 30098 50654
rect 33854 50706 33906 50718
rect 33854 50642 33906 50654
rect 35646 50706 35698 50718
rect 42366 50706 42418 50718
rect 39218 50654 39230 50706
rect 39282 50654 39294 50706
rect 41346 50654 41358 50706
rect 41410 50654 41422 50706
rect 35646 50642 35698 50654
rect 42366 50642 42418 50654
rect 46734 50706 46786 50718
rect 47058 50654 47070 50706
rect 47122 50654 47134 50706
rect 49186 50654 49198 50706
rect 49250 50654 49262 50706
rect 46734 50642 46786 50654
rect 7198 50594 7250 50606
rect 12910 50594 12962 50606
rect 20750 50594 20802 50606
rect 1810 50542 1822 50594
rect 1874 50542 1886 50594
rect 12226 50542 12238 50594
rect 12290 50542 12302 50594
rect 13682 50542 13694 50594
rect 13746 50542 13758 50594
rect 20066 50542 20078 50594
rect 20130 50542 20142 50594
rect 7198 50530 7250 50542
rect 12910 50530 12962 50542
rect 20750 50530 20802 50542
rect 22206 50594 22258 50606
rect 22206 50530 22258 50542
rect 22318 50594 22370 50606
rect 22318 50530 22370 50542
rect 26350 50594 26402 50606
rect 26350 50530 26402 50542
rect 27022 50594 27074 50606
rect 27022 50530 27074 50542
rect 31278 50594 31330 50606
rect 35870 50594 35922 50606
rect 41694 50594 41746 50606
rect 33394 50542 33406 50594
rect 33458 50542 33470 50594
rect 36978 50542 36990 50594
rect 37042 50542 37054 50594
rect 37986 50542 37998 50594
rect 38050 50542 38062 50594
rect 38546 50542 38558 50594
rect 38610 50542 38622 50594
rect 31278 50530 31330 50542
rect 35870 50530 35922 50542
rect 41694 50530 41746 50542
rect 43150 50594 43202 50606
rect 43822 50594 43874 50606
rect 43474 50542 43486 50594
rect 43538 50542 43550 50594
rect 49970 50542 49982 50594
rect 50034 50542 50046 50594
rect 43150 50530 43202 50542
rect 43822 50530 43874 50542
rect 2046 50482 2098 50494
rect 2046 50418 2098 50430
rect 2382 50482 2434 50494
rect 2382 50418 2434 50430
rect 2718 50482 2770 50494
rect 2718 50418 2770 50430
rect 3166 50482 3218 50494
rect 3166 50418 3218 50430
rect 7086 50482 7138 50494
rect 7086 50418 7138 50430
rect 9438 50482 9490 50494
rect 10110 50482 10162 50494
rect 10894 50482 10946 50494
rect 9762 50430 9774 50482
rect 9826 50430 9838 50482
rect 10434 50430 10446 50482
rect 10498 50430 10510 50482
rect 9438 50418 9490 50430
rect 10110 50418 10162 50430
rect 10894 50418 10946 50430
rect 11006 50482 11058 50494
rect 11006 50418 11058 50430
rect 11230 50482 11282 50494
rect 11230 50418 11282 50430
rect 11454 50482 11506 50494
rect 11454 50418 11506 50430
rect 12462 50482 12514 50494
rect 12462 50418 12514 50430
rect 12798 50482 12850 50494
rect 12798 50418 12850 50430
rect 13470 50482 13522 50494
rect 13470 50418 13522 50430
rect 20638 50482 20690 50494
rect 20638 50418 20690 50430
rect 22094 50482 22146 50494
rect 22094 50418 22146 50430
rect 23662 50482 23714 50494
rect 41806 50482 41858 50494
rect 37090 50430 37102 50482
rect 37154 50430 37166 50482
rect 23662 50418 23714 50430
rect 41806 50418 41858 50430
rect 43934 50482 43986 50494
rect 43934 50418 43986 50430
rect 20414 50370 20466 50382
rect 21646 50370 21698 50382
rect 21298 50318 21310 50370
rect 21362 50318 21374 50370
rect 20414 50306 20466 50318
rect 21646 50306 21698 50318
rect 26462 50370 26514 50382
rect 26462 50306 26514 50318
rect 26574 50370 26626 50382
rect 26574 50306 26626 50318
rect 30942 50370 30994 50382
rect 30942 50306 30994 50318
rect 36206 50370 36258 50382
rect 36206 50306 36258 50318
rect 36430 50370 36482 50382
rect 44046 50370 44098 50382
rect 37874 50318 37886 50370
rect 37938 50318 37950 50370
rect 36430 50306 36482 50318
rect 44046 50306 44098 50318
rect 1344 50202 58576 50236
rect 1344 50150 19838 50202
rect 19890 50150 19942 50202
rect 19994 50150 20046 50202
rect 20098 50150 50558 50202
rect 50610 50150 50662 50202
rect 50714 50150 50766 50202
rect 50818 50150 58576 50202
rect 1344 50116 58576 50150
rect 7086 50034 7138 50046
rect 7086 49970 7138 49982
rect 7870 50034 7922 50046
rect 16270 50034 16322 50046
rect 27470 50034 27522 50046
rect 8194 49982 8206 50034
rect 8258 49982 8270 50034
rect 17490 49982 17502 50034
rect 17554 49982 17566 50034
rect 7870 49970 7922 49982
rect 16270 49970 16322 49982
rect 27470 49970 27522 49982
rect 28142 50034 28194 50046
rect 28142 49970 28194 49982
rect 36542 50034 36594 50046
rect 40114 49982 40126 50034
rect 40178 49982 40190 50034
rect 36542 49970 36594 49982
rect 2046 49922 2098 49934
rect 16046 49922 16098 49934
rect 7522 49870 7534 49922
rect 7586 49870 7598 49922
rect 13570 49870 13582 49922
rect 13634 49870 13646 49922
rect 2046 49858 2098 49870
rect 16046 49858 16098 49870
rect 25342 49922 25394 49934
rect 25342 49858 25394 49870
rect 27694 49922 27746 49934
rect 27694 49858 27746 49870
rect 28254 49922 28306 49934
rect 28254 49858 28306 49870
rect 30382 49922 30434 49934
rect 30382 49858 30434 49870
rect 30606 49922 30658 49934
rect 30606 49858 30658 49870
rect 31726 49922 31778 49934
rect 31726 49858 31778 49870
rect 35198 49922 35250 49934
rect 42254 49922 42306 49934
rect 36194 49870 36206 49922
rect 36258 49870 36270 49922
rect 38210 49870 38222 49922
rect 38274 49870 38286 49922
rect 39218 49870 39230 49922
rect 39282 49870 39294 49922
rect 35198 49858 35250 49870
rect 42254 49858 42306 49870
rect 45838 49922 45890 49934
rect 51650 49870 51662 49922
rect 51714 49870 51726 49922
rect 45838 49858 45890 49870
rect 1710 49810 1762 49822
rect 1710 49746 1762 49758
rect 6862 49810 6914 49822
rect 6862 49746 6914 49758
rect 7198 49810 7250 49822
rect 7198 49746 7250 49758
rect 8542 49810 8594 49822
rect 16494 49810 16546 49822
rect 26350 49810 26402 49822
rect 9650 49758 9662 49810
rect 9714 49758 9726 49810
rect 12786 49758 12798 49810
rect 12850 49758 12862 49810
rect 16706 49758 16718 49810
rect 16770 49758 16782 49810
rect 18498 49758 18510 49810
rect 18562 49758 18574 49810
rect 19282 49758 19294 49810
rect 19346 49758 19358 49810
rect 8542 49746 8594 49758
rect 16494 49746 16546 49758
rect 26350 49746 26402 49758
rect 26574 49810 26626 49822
rect 26574 49746 26626 49758
rect 27022 49810 27074 49822
rect 31390 49810 31442 49822
rect 27234 49758 27246 49810
rect 27298 49758 27310 49810
rect 30146 49758 30158 49810
rect 30210 49758 30222 49810
rect 27022 49746 27074 49758
rect 31390 49746 31442 49758
rect 35310 49810 35362 49822
rect 42142 49810 42194 49822
rect 36754 49758 36766 49810
rect 36818 49758 36830 49810
rect 37538 49758 37550 49810
rect 37602 49758 37614 49810
rect 39442 49758 39454 49810
rect 39506 49758 39518 49810
rect 40002 49758 40014 49810
rect 40066 49758 40078 49810
rect 35310 49746 35362 49758
rect 42142 49746 42194 49758
rect 42478 49810 42530 49822
rect 43486 49810 43538 49822
rect 43138 49758 43150 49810
rect 43202 49758 43214 49810
rect 42478 49746 42530 49758
rect 43486 49746 43538 49758
rect 43710 49810 43762 49822
rect 43710 49746 43762 49758
rect 43934 49810 43986 49822
rect 43934 49746 43986 49758
rect 44270 49810 44322 49822
rect 44270 49746 44322 49758
rect 44494 49810 44546 49822
rect 44494 49746 44546 49758
rect 49310 49810 49362 49822
rect 49634 49758 49646 49810
rect 49698 49758 49710 49810
rect 49310 49746 49362 49758
rect 2494 49698 2546 49710
rect 16382 49698 16434 49710
rect 10322 49646 10334 49698
rect 10386 49646 10398 49698
rect 12450 49646 12462 49698
rect 12514 49646 12526 49698
rect 15698 49646 15710 49698
rect 15762 49646 15774 49698
rect 2494 49634 2546 49646
rect 16382 49634 16434 49646
rect 18062 49698 18114 49710
rect 26462 49698 26514 49710
rect 18834 49646 18846 49698
rect 18898 49646 18910 49698
rect 20066 49646 20078 49698
rect 20130 49646 20142 49698
rect 22194 49646 22206 49698
rect 22258 49646 22270 49698
rect 18062 49634 18114 49646
rect 26462 49634 26514 49646
rect 28702 49698 28754 49710
rect 28702 49634 28754 49646
rect 29598 49698 29650 49710
rect 29598 49634 29650 49646
rect 34750 49698 34802 49710
rect 34750 49634 34802 49646
rect 35870 49698 35922 49710
rect 43598 49698 43650 49710
rect 37426 49646 37438 49698
rect 37490 49646 37502 49698
rect 35870 49634 35922 49646
rect 43598 49634 43650 49646
rect 44158 49698 44210 49710
rect 44158 49634 44210 49646
rect 45390 49698 45442 49710
rect 45390 49634 45442 49646
rect 17838 49586 17890 49598
rect 17838 49522 17890 49534
rect 25230 49586 25282 49598
rect 25230 49522 25282 49534
rect 27358 49586 27410 49598
rect 27358 49522 27410 49534
rect 28142 49586 28194 49598
rect 30270 49586 30322 49598
rect 29362 49534 29374 49586
rect 29426 49583 29438 49586
rect 29586 49583 29598 49586
rect 29426 49537 29598 49583
rect 29426 49534 29438 49537
rect 29586 49534 29598 49537
rect 29650 49534 29662 49586
rect 28142 49522 28194 49534
rect 30270 49522 30322 49534
rect 35198 49586 35250 49598
rect 35198 49522 35250 49534
rect 1344 49418 58576 49452
rect 1344 49366 4478 49418
rect 4530 49366 4582 49418
rect 4634 49366 4686 49418
rect 4738 49366 35198 49418
rect 35250 49366 35302 49418
rect 35354 49366 35406 49418
rect 35458 49366 58576 49418
rect 1344 49332 58576 49366
rect 43822 49250 43874 49262
rect 43822 49186 43874 49198
rect 45950 49250 46002 49262
rect 45950 49186 46002 49198
rect 1934 49138 1986 49150
rect 8990 49138 9042 49150
rect 21422 49138 21474 49150
rect 27246 49138 27298 49150
rect 37102 49138 37154 49150
rect 8530 49086 8542 49138
rect 8594 49086 8606 49138
rect 10210 49086 10222 49138
rect 10274 49086 10286 49138
rect 12338 49086 12350 49138
rect 12402 49086 12414 49138
rect 13570 49086 13582 49138
rect 13634 49086 13646 49138
rect 15362 49086 15374 49138
rect 15426 49086 15438 49138
rect 17490 49086 17502 49138
rect 17554 49086 17566 49138
rect 24322 49086 24334 49138
rect 24386 49086 24398 49138
rect 26450 49086 26462 49138
rect 26514 49086 26526 49138
rect 28130 49086 28142 49138
rect 28194 49086 28206 49138
rect 32610 49086 32622 49138
rect 32674 49086 32686 49138
rect 1934 49074 1986 49086
rect 8990 49074 9042 49086
rect 21422 49074 21474 49086
rect 27246 49074 27298 49086
rect 37102 49074 37154 49086
rect 38670 49138 38722 49150
rect 38670 49074 38722 49086
rect 40238 49138 40290 49150
rect 40238 49074 40290 49086
rect 41134 49138 41186 49150
rect 44942 49138 44994 49150
rect 43138 49086 43150 49138
rect 43202 49086 43214 49138
rect 49970 49086 49982 49138
rect 50034 49086 50046 49138
rect 41134 49074 41186 49086
rect 44942 49074 44994 49086
rect 12574 49026 12626 49038
rect 13918 49026 13970 49038
rect 4274 48974 4286 49026
rect 4338 48974 4350 49026
rect 5618 48974 5630 49026
rect 5682 48974 5694 49026
rect 9538 48974 9550 49026
rect 9602 48974 9614 49026
rect 13458 48974 13470 49026
rect 13522 48974 13534 49026
rect 12574 48962 12626 48974
rect 13918 48962 13970 48974
rect 14030 49026 14082 49038
rect 18286 49026 18338 49038
rect 14690 48974 14702 49026
rect 14754 48974 14766 49026
rect 14030 48962 14082 48974
rect 18286 48962 18338 48974
rect 20414 49026 20466 49038
rect 20414 48962 20466 48974
rect 20750 49026 20802 49038
rect 33406 49026 33458 49038
rect 23650 48974 23662 49026
rect 23714 48974 23726 49026
rect 27682 48974 27694 49026
rect 27746 48974 27758 49026
rect 29810 48974 29822 49026
rect 29874 48974 29886 49026
rect 20750 48962 20802 48974
rect 33406 48962 33458 48974
rect 34638 49026 34690 49038
rect 34638 48962 34690 48974
rect 35758 49026 35810 49038
rect 35758 48962 35810 48974
rect 35870 49026 35922 49038
rect 38110 49026 38162 49038
rect 37538 48974 37550 49026
rect 37602 48974 37614 49026
rect 35870 48962 35922 48974
rect 38110 48962 38162 48974
rect 39006 49026 39058 49038
rect 39006 48962 39058 48974
rect 39454 49026 39506 49038
rect 39454 48962 39506 48974
rect 41806 49026 41858 49038
rect 46174 49026 46226 49038
rect 50430 49026 50482 49038
rect 42018 48974 42030 49026
rect 42082 48974 42094 49026
rect 42690 48974 42702 49026
rect 42754 48974 42766 49026
rect 47170 48974 47182 49026
rect 47234 48974 47246 49026
rect 41806 48962 41858 48974
rect 46174 48962 46226 48974
rect 50430 48962 50482 48974
rect 4734 48914 4786 48926
rect 12910 48914 12962 48926
rect 6402 48862 6414 48914
rect 6466 48862 6478 48914
rect 4734 48850 4786 48862
rect 12910 48850 12962 48862
rect 13694 48914 13746 48926
rect 13694 48850 13746 48862
rect 17838 48914 17890 48926
rect 17838 48850 17890 48862
rect 18062 48914 18114 48926
rect 20638 48914 20690 48926
rect 20178 48862 20190 48914
rect 20242 48862 20254 48914
rect 18062 48850 18114 48862
rect 20638 48850 20690 48862
rect 29374 48914 29426 48926
rect 35982 48914 36034 48926
rect 30482 48862 30494 48914
rect 30546 48862 30558 48914
rect 33730 48862 33742 48914
rect 33794 48862 33806 48914
rect 29374 48850 29426 48862
rect 35982 48850 36034 48862
rect 39678 48914 39730 48926
rect 39678 48850 39730 48862
rect 39790 48914 39842 48926
rect 39790 48850 39842 48862
rect 41470 48914 41522 48926
rect 41470 48850 41522 48862
rect 42254 48914 42306 48926
rect 42254 48850 42306 48862
rect 42366 48914 42418 48926
rect 42366 48850 42418 48862
rect 43598 48914 43650 48926
rect 43598 48850 43650 48862
rect 45278 48914 45330 48926
rect 45278 48850 45330 48862
rect 46510 48914 46562 48926
rect 47842 48862 47854 48914
rect 47906 48862 47918 48914
rect 46510 48850 46562 48862
rect 8878 48802 8930 48814
rect 8878 48738 8930 48750
rect 12798 48802 12850 48814
rect 12798 48738 12850 48750
rect 18174 48802 18226 48814
rect 18174 48738 18226 48750
rect 18398 48802 18450 48814
rect 18398 48738 18450 48750
rect 19070 48802 19122 48814
rect 19070 48738 19122 48750
rect 19630 48802 19682 48814
rect 19630 48738 19682 48750
rect 19854 48802 19906 48814
rect 19854 48738 19906 48750
rect 29038 48802 29090 48814
rect 29038 48738 29090 48750
rect 29262 48802 29314 48814
rect 29262 48738 29314 48750
rect 34414 48802 34466 48814
rect 36990 48802 37042 48814
rect 34962 48750 34974 48802
rect 35026 48750 35038 48802
rect 36418 48750 36430 48802
rect 36482 48750 36494 48802
rect 34414 48738 34466 48750
rect 36990 48738 37042 48750
rect 37214 48802 37266 48814
rect 37214 48738 37266 48750
rect 37774 48802 37826 48814
rect 37774 48738 37826 48750
rect 37998 48802 38050 48814
rect 37998 48738 38050 48750
rect 39118 48802 39170 48814
rect 39118 48738 39170 48750
rect 39342 48802 39394 48814
rect 39342 48738 39394 48750
rect 41582 48802 41634 48814
rect 41582 48738 41634 48750
rect 42926 48802 42978 48814
rect 42926 48738 42978 48750
rect 43150 48802 43202 48814
rect 45614 48802 45666 48814
rect 44146 48750 44158 48802
rect 44210 48750 44222 48802
rect 43150 48738 43202 48750
rect 45614 48738 45666 48750
rect 46398 48802 46450 48814
rect 46398 48738 46450 48750
rect 46622 48802 46674 48814
rect 46622 48738 46674 48750
rect 50318 48802 50370 48814
rect 50318 48738 50370 48750
rect 1344 48634 58576 48668
rect 1344 48582 19838 48634
rect 19890 48582 19942 48634
rect 19994 48582 20046 48634
rect 20098 48582 50558 48634
rect 50610 48582 50662 48634
rect 50714 48582 50766 48634
rect 50818 48582 58576 48634
rect 1344 48548 58576 48582
rect 6974 48466 7026 48478
rect 6974 48402 7026 48414
rect 7086 48466 7138 48478
rect 7086 48402 7138 48414
rect 8094 48466 8146 48478
rect 8094 48402 8146 48414
rect 11678 48466 11730 48478
rect 11678 48402 11730 48414
rect 16718 48466 16770 48478
rect 16718 48402 16770 48414
rect 17502 48466 17554 48478
rect 17502 48402 17554 48414
rect 17726 48466 17778 48478
rect 17726 48402 17778 48414
rect 21198 48466 21250 48478
rect 21198 48402 21250 48414
rect 22094 48466 22146 48478
rect 22094 48402 22146 48414
rect 23774 48466 23826 48478
rect 23774 48402 23826 48414
rect 33742 48466 33794 48478
rect 33742 48402 33794 48414
rect 38222 48466 38274 48478
rect 38222 48402 38274 48414
rect 39118 48466 39170 48478
rect 39118 48402 39170 48414
rect 40014 48466 40066 48478
rect 40014 48402 40066 48414
rect 41022 48466 41074 48478
rect 41022 48402 41074 48414
rect 43374 48466 43426 48478
rect 43374 48402 43426 48414
rect 43598 48466 43650 48478
rect 43598 48402 43650 48414
rect 43822 48466 43874 48478
rect 43822 48402 43874 48414
rect 44830 48466 44882 48478
rect 44830 48402 44882 48414
rect 7198 48354 7250 48366
rect 10110 48354 10162 48366
rect 7746 48302 7758 48354
rect 7810 48302 7822 48354
rect 8642 48302 8654 48354
rect 8706 48302 8718 48354
rect 7198 48290 7250 48302
rect 10110 48290 10162 48302
rect 16830 48354 16882 48366
rect 16830 48290 16882 48302
rect 17390 48354 17442 48366
rect 17390 48290 17442 48302
rect 22206 48354 22258 48366
rect 37998 48354 38050 48366
rect 31266 48302 31278 48354
rect 31330 48302 31342 48354
rect 33058 48302 33070 48354
rect 33122 48302 33134 48354
rect 22206 48290 22258 48302
rect 37998 48290 38050 48302
rect 38446 48354 38498 48366
rect 38446 48290 38498 48302
rect 43262 48354 43314 48366
rect 46050 48302 46062 48354
rect 46114 48302 46126 48354
rect 43262 48290 43314 48302
rect 6862 48242 6914 48254
rect 9886 48242 9938 48254
rect 4274 48190 4286 48242
rect 4338 48190 4350 48242
rect 7410 48190 7422 48242
rect 7474 48190 7486 48242
rect 8866 48190 8878 48242
rect 8930 48190 8942 48242
rect 6862 48178 6914 48190
rect 9886 48178 9938 48190
rect 10222 48242 10274 48254
rect 10222 48178 10274 48190
rect 11454 48242 11506 48254
rect 11454 48178 11506 48190
rect 11790 48242 11842 48254
rect 18062 48242 18114 48254
rect 15250 48190 15262 48242
rect 15314 48190 15326 48242
rect 16034 48190 16046 48242
rect 16098 48190 16110 48242
rect 11790 48178 11842 48190
rect 18062 48178 18114 48190
rect 20974 48242 21026 48254
rect 20974 48178 21026 48190
rect 21310 48242 21362 48254
rect 21310 48178 21362 48190
rect 21534 48242 21586 48254
rect 21534 48178 21586 48190
rect 21758 48242 21810 48254
rect 21758 48178 21810 48190
rect 22430 48242 22482 48254
rect 38670 48242 38722 48254
rect 24210 48190 24222 48242
rect 24274 48190 24286 48242
rect 25218 48190 25230 48242
rect 25282 48190 25294 48242
rect 30930 48190 30942 48242
rect 30994 48190 31006 48242
rect 32050 48190 32062 48242
rect 32114 48190 32126 48242
rect 33282 48190 33294 48242
rect 33346 48190 33358 48242
rect 22430 48178 22482 48190
rect 34626 48178 34638 48230
rect 34690 48178 34702 48230
rect 38670 48178 38722 48190
rect 39342 48242 39394 48254
rect 40238 48242 40290 48254
rect 39666 48190 39678 48242
rect 39730 48190 39742 48242
rect 39342 48178 39394 48190
rect 40238 48178 40290 48190
rect 41470 48242 41522 48254
rect 45378 48190 45390 48242
rect 45442 48190 45454 48242
rect 41470 48178 41522 48190
rect 4846 48130 4898 48142
rect 4846 48066 4898 48078
rect 6302 48130 6354 48142
rect 6302 48066 6354 48078
rect 11118 48130 11170 48142
rect 15710 48130 15762 48142
rect 12450 48078 12462 48130
rect 12514 48078 12526 48130
rect 14578 48078 14590 48130
rect 14642 48078 14654 48130
rect 11118 48066 11170 48078
rect 15710 48066 15762 48078
rect 15822 48130 15874 48142
rect 15822 48066 15874 48078
rect 17950 48130 18002 48142
rect 17950 48066 18002 48078
rect 18510 48130 18562 48142
rect 18510 48066 18562 48078
rect 22878 48130 22930 48142
rect 22878 48066 22930 48078
rect 24670 48130 24722 48142
rect 32510 48130 32562 48142
rect 27234 48078 27246 48130
rect 27298 48078 27310 48130
rect 31602 48078 31614 48130
rect 31666 48078 31678 48130
rect 24670 48066 24722 48078
rect 32510 48066 32562 48078
rect 34302 48130 34354 48142
rect 39230 48130 39282 48142
rect 35410 48078 35422 48130
rect 35474 48078 35486 48130
rect 37538 48078 37550 48130
rect 37602 48078 37614 48130
rect 38434 48078 38446 48130
rect 38498 48078 38510 48130
rect 34302 48066 34354 48078
rect 39230 48066 39282 48078
rect 40126 48130 40178 48142
rect 40126 48066 40178 48078
rect 40910 48130 40962 48142
rect 40910 48066 40962 48078
rect 42478 48130 42530 48142
rect 42478 48066 42530 48078
rect 42926 48130 42978 48142
rect 42926 48066 42978 48078
rect 43934 48130 43986 48142
rect 43934 48066 43986 48078
rect 44382 48130 44434 48142
rect 48178 48078 48190 48130
rect 48242 48078 48254 48130
rect 44382 48066 44434 48078
rect 1934 48018 1986 48030
rect 1934 47954 1986 47966
rect 6414 48018 6466 48030
rect 42466 47966 42478 48018
rect 42530 48015 42542 48018
rect 42690 48015 42702 48018
rect 42530 47969 42702 48015
rect 42530 47966 42542 47969
rect 42690 47966 42702 47969
rect 42754 47966 42766 48018
rect 6414 47954 6466 47966
rect 1344 47850 58576 47884
rect 1344 47798 4478 47850
rect 4530 47798 4582 47850
rect 4634 47798 4686 47850
rect 4738 47798 35198 47850
rect 35250 47798 35302 47850
rect 35354 47798 35406 47850
rect 35458 47798 58576 47850
rect 1344 47764 58576 47798
rect 12798 47682 12850 47694
rect 12798 47618 12850 47630
rect 14478 47682 14530 47694
rect 14478 47618 14530 47630
rect 38110 47682 38162 47694
rect 38110 47618 38162 47630
rect 41022 47682 41074 47694
rect 42018 47630 42030 47682
rect 42082 47679 42094 47682
rect 42242 47679 42254 47682
rect 42082 47633 42254 47679
rect 42082 47630 42094 47633
rect 42242 47630 42254 47633
rect 42306 47630 42318 47682
rect 41022 47618 41074 47630
rect 1934 47570 1986 47582
rect 12686 47570 12738 47582
rect 5842 47518 5854 47570
rect 5906 47518 5918 47570
rect 1934 47506 1986 47518
rect 12686 47506 12738 47518
rect 14366 47570 14418 47582
rect 32622 47570 32674 47582
rect 38894 47570 38946 47582
rect 16258 47518 16270 47570
rect 16322 47518 16334 47570
rect 18386 47518 18398 47570
rect 18450 47518 18462 47570
rect 27682 47518 27694 47570
rect 27746 47518 27758 47570
rect 37426 47518 37438 47570
rect 37490 47518 37502 47570
rect 14366 47506 14418 47518
rect 32622 47506 32674 47518
rect 38894 47506 38946 47518
rect 39566 47570 39618 47582
rect 39566 47506 39618 47518
rect 40574 47570 40626 47582
rect 40574 47506 40626 47518
rect 42254 47570 42306 47582
rect 42254 47506 42306 47518
rect 48302 47570 48354 47582
rect 48302 47506 48354 47518
rect 48750 47570 48802 47582
rect 48750 47506 48802 47518
rect 57934 47570 57986 47582
rect 57934 47506 57986 47518
rect 11342 47458 11394 47470
rect 21982 47458 22034 47470
rect 4274 47406 4286 47458
rect 4338 47406 4350 47458
rect 10098 47406 10110 47458
rect 10162 47406 10174 47458
rect 19170 47406 19182 47458
rect 19234 47406 19246 47458
rect 21522 47406 21534 47458
rect 21586 47406 21598 47458
rect 11342 47394 11394 47406
rect 21982 47394 22034 47406
rect 22654 47458 22706 47470
rect 22654 47394 22706 47406
rect 23326 47458 23378 47470
rect 28030 47458 28082 47470
rect 24770 47406 24782 47458
rect 24834 47406 24846 47458
rect 23326 47394 23378 47406
rect 28030 47394 28082 47406
rect 28702 47458 28754 47470
rect 28702 47394 28754 47406
rect 29822 47458 29874 47470
rect 31054 47458 31106 47470
rect 31838 47458 31890 47470
rect 30146 47406 30158 47458
rect 30210 47406 30222 47458
rect 30482 47406 30494 47458
rect 30546 47406 30558 47458
rect 31266 47406 31278 47458
rect 31330 47406 31342 47458
rect 31602 47406 31614 47458
rect 31666 47406 31678 47458
rect 29822 47394 29874 47406
rect 31054 47394 31106 47406
rect 31838 47394 31890 47406
rect 32062 47458 32114 47470
rect 32062 47394 32114 47406
rect 32174 47458 32226 47470
rect 32174 47394 32226 47406
rect 32734 47458 32786 47470
rect 32734 47394 32786 47406
rect 33742 47458 33794 47470
rect 33742 47394 33794 47406
rect 34302 47458 34354 47470
rect 34302 47394 34354 47406
rect 35198 47458 35250 47470
rect 35198 47394 35250 47406
rect 35758 47458 35810 47470
rect 35758 47394 35810 47406
rect 36206 47458 36258 47470
rect 36206 47394 36258 47406
rect 36990 47458 37042 47470
rect 38334 47458 38386 47470
rect 37874 47406 37886 47458
rect 37938 47406 37950 47458
rect 36990 47394 37042 47406
rect 38334 47394 38386 47406
rect 40126 47458 40178 47470
rect 40126 47394 40178 47406
rect 40350 47458 40402 47470
rect 40350 47394 40402 47406
rect 40798 47458 40850 47470
rect 40798 47394 40850 47406
rect 43598 47458 43650 47470
rect 43598 47394 43650 47406
rect 44046 47458 44098 47470
rect 44046 47394 44098 47406
rect 45166 47458 45218 47470
rect 45166 47394 45218 47406
rect 45278 47458 45330 47470
rect 46398 47458 46450 47470
rect 45714 47406 45726 47458
rect 45778 47406 45790 47458
rect 45278 47394 45330 47406
rect 46398 47394 46450 47406
rect 46622 47458 46674 47470
rect 55570 47406 55582 47458
rect 55634 47406 55646 47458
rect 46622 47394 46674 47406
rect 14254 47346 14306 47358
rect 14254 47282 14306 47294
rect 16046 47346 16098 47358
rect 16046 47282 16098 47294
rect 21758 47346 21810 47358
rect 21758 47282 21810 47294
rect 23102 47346 23154 47358
rect 23102 47282 23154 47294
rect 23662 47346 23714 47358
rect 29598 47346 29650 47358
rect 25554 47294 25566 47346
rect 25618 47294 25630 47346
rect 23662 47282 23714 47294
rect 29598 47282 29650 47294
rect 30942 47346 30994 47358
rect 30942 47282 30994 47294
rect 32958 47346 33010 47358
rect 32958 47282 33010 47294
rect 34750 47346 34802 47358
rect 34750 47282 34802 47294
rect 39790 47346 39842 47358
rect 39790 47282 39842 47294
rect 41134 47346 41186 47358
rect 41134 47282 41186 47294
rect 41246 47346 41298 47358
rect 41246 47282 41298 47294
rect 42926 47346 42978 47358
rect 42926 47282 42978 47294
rect 43374 47346 43426 47358
rect 43374 47282 43426 47294
rect 44270 47346 44322 47358
rect 44270 47282 44322 47294
rect 45054 47346 45106 47358
rect 45054 47282 45106 47294
rect 46062 47346 46114 47358
rect 46062 47282 46114 47294
rect 46958 47346 47010 47358
rect 46958 47282 47010 47294
rect 47182 47346 47234 47358
rect 47182 47282 47234 47294
rect 47630 47346 47682 47358
rect 47630 47282 47682 47294
rect 47742 47346 47794 47358
rect 47742 47282 47794 47294
rect 4734 47234 4786 47246
rect 4734 47170 4786 47182
rect 11454 47234 11506 47246
rect 11454 47170 11506 47182
rect 11566 47234 11618 47246
rect 11566 47170 11618 47182
rect 11678 47234 11730 47246
rect 11678 47170 11730 47182
rect 11790 47234 11842 47246
rect 11790 47170 11842 47182
rect 20078 47234 20130 47246
rect 20078 47170 20130 47182
rect 20526 47234 20578 47246
rect 20526 47170 20578 47182
rect 21870 47234 21922 47246
rect 21870 47170 21922 47182
rect 22094 47234 22146 47246
rect 22094 47170 22146 47182
rect 22542 47234 22594 47246
rect 22542 47170 22594 47182
rect 23214 47234 23266 47246
rect 23214 47170 23266 47182
rect 24446 47234 24498 47246
rect 24446 47170 24498 47182
rect 28142 47234 28194 47246
rect 28142 47170 28194 47182
rect 28254 47234 28306 47246
rect 28254 47170 28306 47182
rect 29262 47234 29314 47246
rect 29262 47170 29314 47182
rect 29710 47234 29762 47246
rect 29710 47170 29762 47182
rect 32510 47234 32562 47246
rect 32510 47170 32562 47182
rect 34974 47234 35026 47246
rect 34974 47170 35026 47182
rect 35086 47234 35138 47246
rect 35086 47170 35138 47182
rect 35534 47234 35586 47246
rect 35534 47170 35586 47182
rect 35646 47234 35698 47246
rect 35646 47170 35698 47182
rect 37998 47234 38050 47246
rect 41806 47234 41858 47246
rect 39218 47182 39230 47234
rect 39282 47182 39294 47234
rect 37998 47170 38050 47182
rect 41806 47170 41858 47182
rect 42702 47234 42754 47246
rect 42702 47170 42754 47182
rect 42814 47234 42866 47246
rect 42814 47170 42866 47182
rect 43262 47234 43314 47246
rect 43262 47170 43314 47182
rect 43934 47234 43986 47246
rect 43934 47170 43986 47182
rect 46286 47234 46338 47246
rect 46286 47170 46338 47182
rect 47070 47234 47122 47246
rect 47070 47170 47122 47182
rect 47966 47234 48018 47246
rect 47966 47170 48018 47182
rect 1344 47066 58576 47100
rect 1344 47014 19838 47066
rect 19890 47014 19942 47066
rect 19994 47014 20046 47066
rect 20098 47014 50558 47066
rect 50610 47014 50662 47066
rect 50714 47014 50766 47066
rect 50818 47014 58576 47066
rect 1344 46980 58576 47014
rect 8206 46898 8258 46910
rect 8206 46834 8258 46846
rect 17838 46898 17890 46910
rect 27470 46898 27522 46910
rect 27122 46846 27134 46898
rect 27186 46846 27198 46898
rect 17838 46834 17890 46846
rect 27470 46834 27522 46846
rect 27694 46898 27746 46910
rect 35758 46898 35810 46910
rect 32274 46846 32286 46898
rect 32338 46846 32350 46898
rect 27694 46834 27746 46846
rect 35758 46834 35810 46846
rect 40798 46898 40850 46910
rect 40798 46834 40850 46846
rect 41022 46898 41074 46910
rect 41022 46834 41074 46846
rect 41582 46898 41634 46910
rect 41582 46834 41634 46846
rect 44494 46898 44546 46910
rect 44494 46834 44546 46846
rect 45950 46898 46002 46910
rect 45950 46834 46002 46846
rect 2046 46786 2098 46798
rect 28590 46786 28642 46798
rect 33966 46786 34018 46798
rect 11666 46734 11678 46786
rect 11730 46734 11742 46786
rect 29922 46734 29934 46786
rect 29986 46734 29998 46786
rect 2046 46722 2098 46734
rect 28590 46722 28642 46734
rect 33966 46722 34018 46734
rect 34078 46786 34130 46798
rect 34078 46722 34130 46734
rect 34974 46786 35026 46798
rect 34974 46722 35026 46734
rect 41134 46786 41186 46798
rect 41134 46722 41186 46734
rect 44382 46786 44434 46798
rect 44382 46722 44434 46734
rect 46174 46786 46226 46798
rect 47630 46786 47682 46798
rect 47058 46734 47070 46786
rect 47122 46734 47134 46786
rect 46174 46722 46226 46734
rect 47630 46722 47682 46734
rect 1710 46674 1762 46686
rect 7982 46674 8034 46686
rect 17614 46674 17666 46686
rect 4610 46622 4622 46674
rect 4674 46622 4686 46674
rect 7746 46622 7758 46674
rect 7810 46622 7822 46674
rect 8418 46622 8430 46674
rect 8482 46622 8494 46674
rect 12338 46622 12350 46674
rect 12402 46622 12414 46674
rect 1710 46610 1762 46622
rect 7982 46610 8034 46622
rect 17614 46610 17666 46622
rect 17838 46674 17890 46686
rect 17838 46610 17890 46622
rect 18174 46674 18226 46686
rect 25342 46674 25394 46686
rect 21298 46622 21310 46674
rect 21362 46622 21374 46674
rect 24658 46622 24670 46674
rect 24722 46622 24734 46674
rect 18174 46610 18226 46622
rect 25342 46610 25394 46622
rect 25790 46674 25842 46686
rect 25790 46610 25842 46622
rect 26574 46674 26626 46686
rect 26574 46610 26626 46622
rect 26798 46674 26850 46686
rect 26798 46610 26850 46622
rect 28142 46674 28194 46686
rect 28142 46610 28194 46622
rect 28366 46674 28418 46686
rect 28366 46610 28418 46622
rect 28702 46674 28754 46686
rect 28702 46610 28754 46622
rect 29262 46674 29314 46686
rect 34190 46674 34242 46686
rect 29698 46622 29710 46674
rect 29762 46622 29774 46674
rect 30370 46622 30382 46674
rect 30434 46622 30446 46674
rect 31266 46622 31278 46674
rect 31330 46622 31342 46674
rect 31490 46622 31502 46674
rect 31554 46622 31566 46674
rect 32050 46622 32062 46674
rect 32114 46622 32126 46674
rect 29262 46610 29314 46622
rect 34190 46610 34242 46622
rect 34638 46674 34690 46686
rect 34638 46610 34690 46622
rect 35198 46674 35250 46686
rect 35198 46610 35250 46622
rect 35982 46674 36034 46686
rect 35982 46610 36034 46622
rect 36430 46674 36482 46686
rect 41806 46674 41858 46686
rect 37426 46622 37438 46674
rect 37490 46622 37502 46674
rect 36430 46610 36482 46622
rect 41806 46610 41858 46622
rect 42030 46674 42082 46686
rect 42030 46610 42082 46622
rect 42478 46674 42530 46686
rect 42478 46610 42530 46622
rect 42926 46674 42978 46686
rect 42926 46610 42978 46622
rect 43038 46674 43090 46686
rect 43038 46610 43090 46622
rect 43486 46674 43538 46686
rect 43486 46610 43538 46622
rect 44606 46674 44658 46686
rect 44606 46610 44658 46622
rect 44942 46674 44994 46686
rect 44942 46610 44994 46622
rect 45502 46674 45554 46686
rect 45502 46610 45554 46622
rect 46062 46674 46114 46686
rect 46062 46610 46114 46622
rect 46510 46674 46562 46686
rect 46510 46610 46562 46622
rect 46734 46674 46786 46686
rect 46734 46610 46786 46622
rect 47406 46674 47458 46686
rect 47954 46622 47966 46674
rect 48018 46622 48030 46674
rect 53442 46622 53454 46674
rect 53506 46622 53518 46674
rect 47406 46610 47458 46622
rect 2494 46562 2546 46574
rect 2494 46498 2546 46510
rect 2942 46562 2994 46574
rect 8094 46562 8146 46574
rect 16942 46562 16994 46574
rect 27582 46562 27634 46574
rect 5282 46510 5294 46562
rect 5346 46510 5358 46562
rect 7410 46510 7422 46562
rect 7474 46510 7486 46562
rect 9538 46510 9550 46562
rect 9602 46510 9614 46562
rect 18498 46510 18510 46562
rect 18562 46510 18574 46562
rect 20626 46510 20638 46562
rect 20690 46510 20702 46562
rect 21746 46510 21758 46562
rect 21810 46510 21822 46562
rect 23874 46510 23886 46562
rect 23938 46510 23950 46562
rect 2942 46498 2994 46510
rect 8094 46498 8146 46510
rect 16942 46498 16994 46510
rect 27582 46498 27634 46510
rect 33182 46562 33234 46574
rect 33182 46498 33234 46510
rect 34750 46562 34802 46574
rect 34750 46498 34802 46510
rect 35870 46562 35922 46574
rect 35870 46498 35922 46510
rect 36766 46562 36818 46574
rect 41694 46562 41746 46574
rect 38210 46510 38222 46562
rect 38274 46510 38286 46562
rect 40338 46510 40350 46562
rect 40402 46510 40414 46562
rect 36766 46498 36818 46510
rect 41694 46498 41746 46510
rect 42254 46562 42306 46574
rect 42254 46498 42306 46510
rect 42702 46562 42754 46574
rect 42702 46498 42754 46510
rect 47518 46562 47570 46574
rect 47518 46498 47570 46510
rect 53230 46562 53282 46574
rect 53230 46498 53282 46510
rect 25230 46450 25282 46462
rect 25230 46386 25282 46398
rect 30382 46450 30434 46462
rect 43710 46450 43762 46462
rect 33506 46398 33518 46450
rect 33570 46398 33582 46450
rect 36530 46398 36542 46450
rect 36594 46447 36606 46450
rect 36866 46447 36878 46450
rect 36594 46401 36878 46447
rect 36594 46398 36606 46401
rect 36866 46398 36878 46401
rect 36930 46398 36942 46450
rect 44034 46398 44046 46450
rect 44098 46398 44110 46450
rect 55346 46398 55358 46450
rect 55410 46398 55422 46450
rect 30382 46386 30434 46398
rect 43710 46386 43762 46398
rect 1344 46282 58576 46316
rect 1344 46230 4478 46282
rect 4530 46230 4582 46282
rect 4634 46230 4686 46282
rect 4738 46230 35198 46282
rect 35250 46230 35302 46282
rect 35354 46230 35406 46282
rect 35458 46230 58576 46282
rect 1344 46196 58576 46230
rect 8990 46114 9042 46126
rect 8990 46050 9042 46062
rect 11678 46114 11730 46126
rect 11678 46050 11730 46062
rect 21534 46114 21586 46126
rect 35858 46062 35870 46114
rect 35922 46062 35934 46114
rect 43250 46062 43262 46114
rect 43314 46062 43326 46114
rect 21534 46050 21586 46062
rect 11566 46002 11618 46014
rect 36430 46002 36482 46014
rect 55022 46002 55074 46014
rect 6402 45950 6414 46002
rect 6466 45950 6478 46002
rect 10658 45950 10670 46002
rect 10722 45950 10734 46002
rect 16594 45950 16606 46002
rect 16658 45950 16670 46002
rect 17154 45950 17166 46002
rect 17218 45950 17230 46002
rect 22418 45950 22430 46002
rect 22482 45950 22494 46002
rect 23650 45950 23662 46002
rect 23714 45950 23726 46002
rect 28466 45950 28478 46002
rect 28530 45950 28542 46002
rect 46386 45950 46398 46002
rect 46450 45950 46462 46002
rect 48514 45950 48526 46002
rect 48578 45950 48590 46002
rect 57810 45950 57822 46002
rect 57874 45950 57886 46002
rect 11566 45938 11618 45950
rect 36430 45938 36482 45950
rect 55022 45938 55074 45950
rect 6750 45890 6802 45902
rect 8206 45890 8258 45902
rect 10334 45890 10386 45902
rect 1810 45838 1822 45890
rect 1874 45838 1886 45890
rect 6962 45838 6974 45890
rect 7026 45838 7038 45890
rect 10098 45838 10110 45890
rect 10162 45838 10174 45890
rect 6750 45826 6802 45838
rect 8206 45826 8258 45838
rect 10334 45826 10386 45838
rect 10558 45890 10610 45902
rect 11118 45890 11170 45902
rect 21982 45890 22034 45902
rect 10770 45838 10782 45890
rect 10834 45838 10846 45890
rect 12898 45838 12910 45890
rect 12962 45838 12974 45890
rect 13794 45838 13806 45890
rect 13858 45838 13870 45890
rect 20066 45838 20078 45890
rect 20130 45838 20142 45890
rect 10558 45826 10610 45838
rect 11118 45826 11170 45838
rect 21982 45826 22034 45838
rect 22318 45890 22370 45902
rect 23214 45890 23266 45902
rect 22530 45838 22542 45890
rect 22594 45838 22606 45890
rect 22318 45826 22370 45838
rect 23214 45826 23266 45838
rect 23550 45890 23602 45902
rect 35310 45890 35362 45902
rect 23762 45838 23774 45890
rect 23826 45838 23838 45890
rect 27682 45838 27694 45890
rect 27746 45838 27758 45890
rect 28018 45838 28030 45890
rect 28082 45838 28094 45890
rect 34626 45838 34638 45890
rect 34690 45838 34702 45890
rect 23550 45826 23602 45838
rect 35310 45826 35362 45838
rect 36206 45890 36258 45902
rect 36206 45826 36258 45838
rect 36878 45890 36930 45902
rect 43822 45890 43874 45902
rect 44830 45890 44882 45902
rect 42802 45838 42814 45890
rect 42866 45838 42878 45890
rect 44034 45838 44046 45890
rect 44098 45838 44110 45890
rect 36878 45826 36930 45838
rect 43822 45826 43874 45838
rect 44830 45826 44882 45838
rect 45054 45890 45106 45902
rect 45838 45890 45890 45902
rect 45378 45838 45390 45890
rect 45442 45838 45454 45890
rect 49186 45838 49198 45890
rect 49250 45838 49262 45890
rect 52658 45838 52670 45890
rect 52722 45838 52734 45890
rect 55570 45838 55582 45890
rect 55634 45838 55646 45890
rect 45054 45826 45106 45838
rect 45838 45826 45890 45838
rect 2382 45778 2434 45790
rect 2382 45714 2434 45726
rect 3166 45778 3218 45790
rect 3166 45714 3218 45726
rect 6526 45778 6578 45790
rect 6526 45714 6578 45726
rect 7534 45778 7586 45790
rect 7534 45714 7586 45726
rect 7982 45778 8034 45790
rect 7982 45714 8034 45726
rect 8430 45778 8482 45790
rect 8430 45714 8482 45726
rect 8542 45778 8594 45790
rect 8542 45714 8594 45726
rect 8878 45778 8930 45790
rect 8878 45714 8930 45726
rect 8990 45778 9042 45790
rect 8990 45714 9042 45726
rect 11230 45778 11282 45790
rect 11230 45714 11282 45726
rect 12574 45778 12626 45790
rect 20750 45778 20802 45790
rect 14466 45726 14478 45778
rect 14530 45726 14542 45778
rect 19282 45726 19294 45778
rect 19346 45726 19358 45778
rect 12574 45714 12626 45726
rect 20750 45714 20802 45726
rect 21422 45778 21474 45790
rect 34974 45778 35026 45790
rect 28466 45726 28478 45778
rect 28530 45726 28542 45778
rect 30258 45726 30270 45778
rect 30322 45726 30334 45778
rect 21422 45714 21474 45726
rect 34974 45714 35026 45726
rect 35534 45778 35586 45790
rect 35534 45714 35586 45726
rect 37214 45778 37266 45790
rect 43710 45778 43762 45790
rect 37762 45726 37774 45778
rect 37826 45726 37838 45778
rect 37214 45714 37266 45726
rect 43710 45714 43762 45726
rect 2046 45666 2098 45678
rect 2046 45602 2098 45614
rect 2718 45666 2770 45678
rect 2718 45602 2770 45614
rect 6414 45666 6466 45678
rect 6414 45602 6466 45614
rect 7422 45666 7474 45678
rect 7422 45602 7474 45614
rect 7646 45666 7698 45678
rect 7646 45602 7698 45614
rect 7758 45666 7810 45678
rect 7758 45602 7810 45614
rect 12686 45666 12738 45678
rect 12686 45602 12738 45614
rect 20526 45666 20578 45678
rect 20526 45602 20578 45614
rect 20638 45666 20690 45678
rect 20638 45602 20690 45614
rect 22094 45666 22146 45678
rect 22094 45602 22146 45614
rect 23326 45666 23378 45678
rect 23326 45602 23378 45614
rect 35310 45666 35362 45678
rect 35310 45602 35362 45614
rect 37102 45666 37154 45678
rect 37102 45602 37154 45614
rect 44942 45666 44994 45678
rect 44942 45602 44994 45614
rect 1344 45498 58576 45532
rect 1344 45446 19838 45498
rect 19890 45446 19942 45498
rect 19994 45446 20046 45498
rect 20098 45446 50558 45498
rect 50610 45446 50662 45498
rect 50714 45446 50766 45498
rect 50818 45446 58576 45498
rect 1344 45412 58576 45446
rect 8654 45330 8706 45342
rect 8654 45266 8706 45278
rect 8878 45330 8930 45342
rect 8878 45266 8930 45278
rect 18286 45330 18338 45342
rect 18286 45266 18338 45278
rect 18734 45330 18786 45342
rect 18734 45266 18786 45278
rect 18958 45330 19010 45342
rect 18958 45266 19010 45278
rect 27358 45330 27410 45342
rect 27358 45266 27410 45278
rect 27582 45330 27634 45342
rect 31502 45330 31554 45342
rect 28018 45278 28030 45330
rect 28082 45278 28094 45330
rect 27582 45266 27634 45278
rect 31502 45266 31554 45278
rect 32622 45330 32674 45342
rect 32622 45266 32674 45278
rect 33406 45330 33458 45342
rect 33406 45266 33458 45278
rect 33518 45330 33570 45342
rect 33518 45266 33570 45278
rect 34638 45330 34690 45342
rect 34638 45266 34690 45278
rect 38558 45330 38610 45342
rect 38558 45266 38610 45278
rect 44158 45330 44210 45342
rect 44158 45266 44210 45278
rect 44382 45330 44434 45342
rect 45838 45330 45890 45342
rect 45378 45278 45390 45330
rect 45442 45278 45454 45330
rect 44382 45266 44434 45278
rect 45838 45266 45890 45278
rect 46398 45330 46450 45342
rect 46398 45266 46450 45278
rect 2046 45218 2098 45230
rect 8990 45218 9042 45230
rect 13470 45218 13522 45230
rect 5954 45166 5966 45218
rect 6018 45166 6030 45218
rect 11666 45166 11678 45218
rect 11730 45166 11742 45218
rect 2046 45154 2098 45166
rect 8990 45154 9042 45166
rect 13470 45154 13522 45166
rect 18174 45218 18226 45230
rect 18174 45154 18226 45166
rect 27134 45218 27186 45230
rect 27134 45154 27186 45166
rect 28590 45218 28642 45230
rect 28590 45154 28642 45166
rect 29374 45218 29426 45230
rect 29374 45154 29426 45166
rect 31278 45218 31330 45230
rect 31278 45154 31330 45166
rect 32398 45218 32450 45230
rect 32398 45154 32450 45166
rect 33630 45218 33682 45230
rect 33630 45154 33682 45166
rect 33966 45218 34018 45230
rect 38894 45218 38946 45230
rect 35634 45166 35646 45218
rect 35698 45166 35710 45218
rect 41682 45166 41694 45218
rect 41746 45166 41758 45218
rect 33966 45154 34018 45166
rect 38894 45154 38946 45166
rect 1710 45106 1762 45118
rect 18510 45106 18562 45118
rect 5170 45054 5182 45106
rect 5234 45054 5246 45106
rect 12338 45054 12350 45106
rect 12402 45054 12414 45106
rect 14018 45054 14030 45106
rect 14082 45054 14094 45106
rect 17714 45054 17726 45106
rect 17778 45054 17790 45106
rect 1710 45042 1762 45054
rect 18510 45042 18562 45054
rect 19070 45106 19122 45118
rect 25342 45106 25394 45118
rect 23202 45054 23214 45106
rect 23266 45054 23278 45106
rect 19070 45042 19122 45054
rect 25342 45042 25394 45054
rect 28478 45106 28530 45118
rect 28478 45042 28530 45054
rect 28702 45106 28754 45118
rect 28702 45042 28754 45054
rect 29150 45106 29202 45118
rect 29150 45042 29202 45054
rect 29822 45106 29874 45118
rect 31950 45106 32002 45118
rect 31602 45054 31614 45106
rect 31666 45054 31678 45106
rect 29822 45042 29874 45054
rect 31950 45042 32002 45054
rect 32286 45106 32338 45118
rect 32286 45042 32338 45054
rect 34078 45106 34130 45118
rect 44830 45106 44882 45118
rect 34850 45054 34862 45106
rect 34914 45054 34926 45106
rect 40898 45054 40910 45106
rect 40962 45054 40974 45106
rect 34078 45042 34130 45054
rect 44830 45042 44882 45054
rect 45054 45106 45106 45118
rect 45054 45042 45106 45054
rect 45614 45106 45666 45118
rect 45614 45042 45666 45054
rect 45950 45106 46002 45118
rect 45950 45042 46002 45054
rect 2494 44994 2546 45006
rect 27470 44994 27522 45006
rect 8082 44942 8094 44994
rect 8146 44942 8158 44994
rect 9538 44942 9550 44994
rect 9602 44942 9614 44994
rect 13570 44942 13582 44994
rect 13634 44942 13646 44994
rect 14690 44942 14702 44994
rect 14754 44942 14766 44994
rect 16818 44942 16830 44994
rect 16882 44942 16894 44994
rect 18274 44942 18286 44994
rect 18338 44942 18350 44994
rect 21746 44942 21758 44994
rect 21810 44942 21822 44994
rect 2494 44930 2546 44942
rect 27470 44930 27522 44942
rect 29598 44994 29650 45006
rect 29598 44930 29650 44942
rect 30942 44994 30994 45006
rect 30942 44930 30994 44942
rect 31390 44994 31442 45006
rect 44270 44994 44322 45006
rect 37762 44942 37774 44994
rect 37826 44942 37838 44994
rect 43810 44942 43822 44994
rect 43874 44942 43886 44994
rect 31390 44930 31442 44942
rect 44270 44930 44322 44942
rect 13246 44882 13298 44894
rect 13246 44818 13298 44830
rect 1344 44714 58576 44748
rect 1344 44662 4478 44714
rect 4530 44662 4582 44714
rect 4634 44662 4686 44714
rect 4738 44662 35198 44714
rect 35250 44662 35302 44714
rect 35354 44662 35406 44714
rect 35458 44662 58576 44714
rect 1344 44628 58576 44662
rect 12462 44546 12514 44558
rect 12462 44482 12514 44494
rect 12910 44546 12962 44558
rect 21310 44546 21362 44558
rect 19618 44494 19630 44546
rect 19682 44494 19694 44546
rect 42802 44494 42814 44546
rect 42866 44543 42878 44546
rect 43362 44543 43374 44546
rect 42866 44497 43374 44543
rect 42866 44494 42878 44497
rect 43362 44494 43374 44497
rect 43426 44494 43438 44546
rect 12910 44482 12962 44494
rect 21310 44482 21362 44494
rect 9102 44434 9154 44446
rect 6514 44382 6526 44434
rect 6578 44382 6590 44434
rect 8642 44382 8654 44434
rect 8706 44382 8718 44434
rect 9102 44370 9154 44382
rect 11118 44434 11170 44446
rect 11118 44370 11170 44382
rect 11454 44434 11506 44446
rect 11454 44370 11506 44382
rect 11902 44434 11954 44446
rect 11902 44370 11954 44382
rect 21422 44434 21474 44446
rect 21422 44370 21474 44382
rect 22094 44434 22146 44446
rect 22094 44370 22146 44382
rect 27134 44434 27186 44446
rect 27134 44370 27186 44382
rect 27582 44434 27634 44446
rect 34526 44434 34578 44446
rect 31266 44382 31278 44434
rect 31330 44382 31342 44434
rect 33394 44382 33406 44434
rect 33458 44382 33470 44434
rect 27582 44370 27634 44382
rect 34526 44370 34578 44382
rect 35870 44434 35922 44446
rect 35870 44370 35922 44382
rect 42926 44434 42978 44446
rect 42926 44370 42978 44382
rect 45502 44434 45554 44446
rect 45502 44370 45554 44382
rect 57934 44434 57986 44446
rect 57934 44370 57986 44382
rect 12574 44322 12626 44334
rect 5730 44270 5742 44322
rect 5794 44270 5806 44322
rect 12574 44258 12626 44270
rect 12798 44322 12850 44334
rect 19854 44322 19906 44334
rect 17602 44270 17614 44322
rect 17666 44270 17678 44322
rect 19394 44270 19406 44322
rect 19458 44270 19470 44322
rect 12798 44258 12850 44270
rect 19854 44258 19906 44270
rect 22654 44322 22706 44334
rect 27022 44322 27074 44334
rect 25106 44270 25118 44322
rect 25170 44270 25182 44322
rect 22654 44258 22706 44270
rect 27022 44258 27074 44270
rect 27358 44322 27410 44334
rect 27358 44258 27410 44270
rect 27918 44322 27970 44334
rect 27918 44258 27970 44270
rect 28366 44322 28418 44334
rect 44942 44322 44994 44334
rect 30482 44270 30494 44322
rect 30546 44270 30558 44322
rect 35298 44270 35310 44322
rect 35362 44270 35374 44322
rect 28366 44258 28418 44270
rect 44942 44258 44994 44270
rect 48414 44322 48466 44334
rect 48414 44258 48466 44270
rect 48526 44322 48578 44334
rect 48526 44258 48578 44270
rect 49086 44322 49138 44334
rect 49086 44258 49138 44270
rect 49422 44322 49474 44334
rect 49422 44258 49474 44270
rect 49646 44322 49698 44334
rect 55570 44270 55582 44322
rect 55634 44270 55646 44322
rect 49646 44258 49698 44270
rect 1710 44210 1762 44222
rect 1710 44146 1762 44158
rect 8990 44210 9042 44222
rect 20190 44210 20242 44222
rect 14018 44158 14030 44210
rect 14082 44158 14094 44210
rect 8990 44146 9042 44158
rect 20190 44146 20242 44158
rect 20750 44210 20802 44222
rect 20750 44146 20802 44158
rect 24222 44210 24274 44222
rect 24222 44146 24274 44158
rect 24558 44210 24610 44222
rect 26686 44210 26738 44222
rect 41582 44210 41634 44222
rect 24882 44158 24894 44210
rect 24946 44158 24958 44210
rect 35074 44158 35086 44210
rect 35138 44158 35150 44210
rect 38658 44158 38670 44210
rect 38722 44158 38734 44210
rect 24558 44146 24610 44158
rect 26686 44146 26738 44158
rect 41582 44146 41634 44158
rect 48862 44210 48914 44222
rect 48862 44146 48914 44158
rect 2046 44098 2098 44110
rect 2046 44034 2098 44046
rect 2494 44098 2546 44110
rect 2494 44034 2546 44046
rect 11566 44098 11618 44110
rect 11566 44034 11618 44046
rect 12014 44098 12066 44110
rect 12014 44034 12066 44046
rect 20078 44098 20130 44110
rect 20078 44034 20130 44046
rect 21534 44098 21586 44110
rect 21534 44034 21586 44046
rect 23998 44098 24050 44110
rect 23998 44034 24050 44046
rect 26462 44098 26514 44110
rect 26462 44034 26514 44046
rect 29262 44098 29314 44110
rect 29262 44034 29314 44046
rect 34078 44098 34130 44110
rect 34078 44034 34130 44046
rect 38334 44098 38386 44110
rect 38334 44034 38386 44046
rect 43374 44098 43426 44110
rect 43374 44034 43426 44046
rect 48750 44098 48802 44110
rect 48750 44034 48802 44046
rect 49310 44098 49362 44110
rect 49310 44034 49362 44046
rect 1344 43930 58576 43964
rect 1344 43878 19838 43930
rect 19890 43878 19942 43930
rect 19994 43878 20046 43930
rect 20098 43878 50558 43930
rect 50610 43878 50662 43930
rect 50714 43878 50766 43930
rect 50818 43878 58576 43930
rect 1344 43844 58576 43878
rect 11454 43762 11506 43774
rect 11454 43698 11506 43710
rect 12574 43762 12626 43774
rect 12574 43698 12626 43710
rect 7646 43650 7698 43662
rect 7646 43586 7698 43598
rect 7758 43650 7810 43662
rect 7758 43586 7810 43598
rect 11790 43650 11842 43662
rect 11790 43586 11842 43598
rect 12350 43650 12402 43662
rect 24110 43650 24162 43662
rect 14466 43598 14478 43650
rect 14530 43598 14542 43650
rect 21522 43598 21534 43650
rect 21586 43598 21598 43650
rect 12350 43586 12402 43598
rect 24110 43586 24162 43598
rect 24334 43650 24386 43662
rect 24334 43586 24386 43598
rect 28926 43650 28978 43662
rect 28926 43586 28978 43598
rect 29150 43650 29202 43662
rect 29150 43586 29202 43598
rect 32286 43650 32338 43662
rect 37998 43650 38050 43662
rect 39566 43650 39618 43662
rect 33954 43598 33966 43650
rect 34018 43598 34030 43650
rect 35970 43598 35982 43650
rect 36034 43598 36046 43650
rect 38770 43598 38782 43650
rect 38834 43598 38846 43650
rect 32286 43586 32338 43598
rect 37998 43586 38050 43598
rect 39566 43586 39618 43598
rect 41358 43650 41410 43662
rect 41358 43586 41410 43598
rect 42142 43650 42194 43662
rect 47966 43650 48018 43662
rect 43810 43598 43822 43650
rect 43874 43598 43886 43650
rect 42142 43586 42194 43598
rect 47966 43586 48018 43598
rect 11678 43538 11730 43550
rect 4274 43486 4286 43538
rect 4338 43486 4350 43538
rect 11678 43474 11730 43486
rect 12238 43538 12290 43550
rect 12238 43474 12290 43486
rect 12910 43538 12962 43550
rect 12910 43474 12962 43486
rect 13246 43538 13298 43550
rect 19182 43538 19234 43550
rect 22878 43538 22930 43550
rect 13682 43486 13694 43538
rect 13746 43486 13758 43538
rect 18162 43486 18174 43538
rect 18226 43486 18238 43538
rect 18386 43486 18398 43538
rect 18450 43486 18462 43538
rect 22194 43486 22206 43538
rect 22258 43486 22270 43538
rect 22642 43486 22654 43538
rect 22706 43486 22718 43538
rect 13246 43474 13298 43486
rect 19182 43474 19234 43486
rect 22878 43474 22930 43486
rect 23102 43538 23154 43550
rect 23774 43538 23826 43550
rect 23314 43486 23326 43538
rect 23378 43486 23390 43538
rect 23102 43474 23154 43486
rect 23774 43474 23826 43486
rect 23886 43538 23938 43550
rect 29486 43538 29538 43550
rect 34750 43538 34802 43550
rect 39118 43538 39170 43550
rect 25554 43486 25566 43538
rect 25618 43486 25630 43538
rect 29922 43486 29934 43538
rect 29986 43486 29998 43538
rect 33730 43486 33742 43538
rect 33794 43486 33806 43538
rect 35746 43486 35758 43538
rect 35810 43486 35822 43538
rect 37762 43486 37774 43538
rect 37826 43486 37838 43538
rect 23886 43474 23938 43486
rect 29486 43474 29538 43486
rect 34750 43474 34802 43486
rect 39118 43474 39170 43486
rect 40910 43538 40962 43550
rect 40910 43474 40962 43486
rect 41582 43538 41634 43550
rect 41582 43474 41634 43486
rect 41918 43538 41970 43550
rect 41918 43474 41970 43486
rect 42590 43538 42642 43550
rect 46846 43538 46898 43550
rect 43026 43486 43038 43538
rect 43090 43486 43102 43538
rect 42590 43474 42642 43486
rect 46846 43474 46898 43486
rect 47070 43538 47122 43550
rect 47070 43474 47122 43486
rect 47406 43538 47458 43550
rect 47406 43474 47458 43486
rect 47518 43538 47570 43550
rect 47518 43474 47570 43486
rect 48190 43538 48242 43550
rect 48850 43486 48862 43538
rect 48914 43486 48926 43538
rect 48190 43474 48242 43486
rect 4846 43426 4898 43438
rect 4846 43362 4898 43374
rect 10446 43426 10498 43438
rect 17502 43426 17554 43438
rect 22990 43426 23042 43438
rect 29374 43426 29426 43438
rect 16594 43374 16606 43426
rect 16658 43374 16670 43426
rect 18498 43374 18510 43426
rect 18562 43374 18574 43426
rect 19394 43374 19406 43426
rect 19458 43374 19470 43426
rect 26338 43374 26350 43426
rect 26402 43374 26414 43426
rect 28466 43374 28478 43426
rect 28530 43374 28542 43426
rect 10446 43362 10498 43374
rect 17502 43362 17554 43374
rect 22990 43362 23042 43374
rect 29374 43362 29426 43374
rect 30382 43426 30434 43438
rect 30382 43362 30434 43374
rect 34414 43426 34466 43438
rect 36430 43426 36482 43438
rect 35186 43374 35198 43426
rect 35250 43374 35262 43426
rect 34414 43362 34466 43374
rect 36430 43362 36482 43374
rect 41134 43426 41186 43438
rect 41134 43362 41186 43374
rect 42366 43426 42418 43438
rect 46398 43426 46450 43438
rect 45938 43374 45950 43426
rect 46002 43374 46014 43426
rect 42366 43362 42418 43374
rect 46398 43362 46450 43374
rect 47182 43426 47234 43438
rect 47182 43362 47234 43374
rect 47742 43426 47794 43438
rect 49522 43374 49534 43426
rect 49586 43374 49598 43426
rect 51650 43374 51662 43426
rect 51714 43374 51726 43426
rect 47742 43362 47794 43374
rect 1934 43314 1986 43326
rect 1934 43250 1986 43262
rect 10334 43314 10386 43326
rect 10334 43250 10386 43262
rect 11790 43314 11842 43326
rect 11790 43250 11842 43262
rect 13022 43314 13074 43326
rect 13022 43250 13074 43262
rect 13358 43314 13410 43326
rect 36194 43262 36206 43314
rect 36258 43311 36270 43314
rect 36418 43311 36430 43314
rect 36258 43265 36430 43311
rect 36258 43262 36270 43265
rect 36418 43262 36430 43265
rect 36482 43262 36494 43314
rect 13358 43250 13410 43262
rect 1344 43146 58576 43180
rect 1344 43094 4478 43146
rect 4530 43094 4582 43146
rect 4634 43094 4686 43146
rect 4738 43094 35198 43146
rect 35250 43094 35302 43146
rect 35354 43094 35406 43146
rect 35458 43094 58576 43146
rect 1344 43060 58576 43094
rect 9662 42978 9714 42990
rect 9662 42914 9714 42926
rect 9886 42978 9938 42990
rect 9886 42914 9938 42926
rect 10110 42978 10162 42990
rect 17950 42978 18002 42990
rect 11442 42926 11454 42978
rect 11506 42926 11518 42978
rect 10110 42914 10162 42926
rect 17950 42914 18002 42926
rect 18174 42978 18226 42990
rect 19742 42978 19794 42990
rect 19394 42926 19406 42978
rect 19458 42926 19470 42978
rect 18174 42914 18226 42926
rect 19742 42914 19794 42926
rect 22094 42978 22146 42990
rect 22094 42914 22146 42926
rect 57934 42978 57986 42990
rect 57934 42914 57986 42926
rect 9326 42866 9378 42878
rect 9326 42802 9378 42814
rect 10222 42866 10274 42878
rect 10222 42802 10274 42814
rect 17726 42866 17778 42878
rect 17726 42802 17778 42814
rect 19182 42866 19234 42878
rect 19182 42802 19234 42814
rect 20750 42866 20802 42878
rect 20750 42802 20802 42814
rect 21982 42866 22034 42878
rect 21982 42802 22034 42814
rect 25790 42866 25842 42878
rect 32510 42866 32562 42878
rect 50206 42866 50258 42878
rect 27906 42814 27918 42866
rect 27970 42814 27982 42866
rect 49522 42814 49534 42866
rect 49586 42814 49598 42866
rect 25790 42802 25842 42814
rect 32510 42802 32562 42814
rect 50206 42802 50258 42814
rect 50654 42866 50706 42878
rect 50654 42802 50706 42814
rect 13694 42754 13746 42766
rect 10658 42702 10670 42754
rect 10722 42702 10734 42754
rect 13694 42690 13746 42702
rect 14030 42754 14082 42766
rect 14030 42690 14082 42702
rect 19966 42754 20018 42766
rect 19966 42690 20018 42702
rect 23774 42754 23826 42766
rect 23774 42690 23826 42702
rect 23998 42754 24050 42766
rect 23998 42690 24050 42702
rect 24334 42754 24386 42766
rect 24334 42690 24386 42702
rect 24558 42754 24610 42766
rect 24558 42690 24610 42702
rect 25006 42754 25058 42766
rect 25006 42690 25058 42702
rect 26238 42754 26290 42766
rect 26238 42690 26290 42702
rect 26686 42754 26738 42766
rect 26686 42690 26738 42702
rect 26798 42754 26850 42766
rect 26798 42690 26850 42702
rect 27134 42754 27186 42766
rect 29598 42754 29650 42766
rect 27570 42702 27582 42754
rect 27634 42702 27646 42754
rect 27134 42690 27186 42702
rect 29598 42690 29650 42702
rect 30158 42754 30210 42766
rect 30158 42690 30210 42702
rect 30718 42754 30770 42766
rect 30718 42690 30770 42702
rect 31054 42754 31106 42766
rect 31054 42690 31106 42702
rect 31390 42754 31442 42766
rect 31390 42690 31442 42702
rect 32734 42754 32786 42766
rect 32734 42690 32786 42702
rect 33182 42754 33234 42766
rect 33182 42690 33234 42702
rect 33630 42754 33682 42766
rect 33630 42690 33682 42702
rect 34078 42754 34130 42766
rect 34078 42690 34130 42702
rect 34190 42754 34242 42766
rect 34190 42690 34242 42702
rect 34638 42754 34690 42766
rect 34638 42690 34690 42702
rect 34974 42754 35026 42766
rect 34974 42690 35026 42702
rect 35086 42754 35138 42766
rect 35086 42690 35138 42702
rect 36206 42754 36258 42766
rect 36206 42690 36258 42702
rect 37662 42754 37714 42766
rect 37662 42690 37714 42702
rect 38110 42754 38162 42766
rect 38110 42690 38162 42702
rect 38334 42754 38386 42766
rect 38334 42690 38386 42702
rect 38670 42754 38722 42766
rect 38670 42690 38722 42702
rect 38894 42754 38946 42766
rect 38894 42690 38946 42702
rect 39678 42754 39730 42766
rect 39678 42690 39730 42702
rect 39902 42754 39954 42766
rect 39902 42690 39954 42702
rect 40238 42754 40290 42766
rect 40238 42690 40290 42702
rect 40574 42754 40626 42766
rect 40574 42690 40626 42702
rect 40686 42754 40738 42766
rect 40686 42690 40738 42702
rect 41358 42754 41410 42766
rect 41358 42690 41410 42702
rect 41582 42754 41634 42766
rect 41582 42690 41634 42702
rect 42478 42754 42530 42766
rect 42478 42690 42530 42702
rect 42702 42754 42754 42766
rect 42702 42690 42754 42702
rect 45390 42754 45442 42766
rect 45390 42690 45442 42702
rect 45838 42754 45890 42766
rect 45838 42690 45890 42702
rect 46062 42754 46114 42766
rect 46062 42690 46114 42702
rect 46398 42754 46450 42766
rect 46398 42690 46450 42702
rect 46622 42754 46674 42766
rect 46622 42690 46674 42702
rect 46958 42754 47010 42766
rect 46958 42690 47010 42702
rect 47294 42754 47346 42766
rect 47294 42690 47346 42702
rect 47630 42754 47682 42766
rect 47630 42690 47682 42702
rect 47854 42754 47906 42766
rect 47854 42690 47906 42702
rect 48190 42754 48242 42766
rect 48190 42690 48242 42702
rect 48414 42754 48466 42766
rect 48414 42690 48466 42702
rect 48750 42754 48802 42766
rect 49074 42702 49086 42754
rect 49138 42702 49150 42754
rect 49746 42702 49758 42754
rect 49810 42702 49822 42754
rect 55570 42702 55582 42754
rect 55634 42702 55646 42754
rect 48750 42690 48802 42702
rect 1710 42642 1762 42654
rect 1710 42578 1762 42590
rect 10894 42642 10946 42654
rect 10894 42578 10946 42590
rect 11006 42642 11058 42654
rect 11006 42578 11058 42590
rect 13918 42642 13970 42654
rect 13918 42578 13970 42590
rect 22430 42642 22482 42654
rect 22430 42578 22482 42590
rect 25230 42642 25282 42654
rect 25230 42578 25282 42590
rect 26014 42642 26066 42654
rect 26014 42578 26066 42590
rect 29710 42642 29762 42654
rect 29710 42578 29762 42590
rect 31614 42642 31666 42654
rect 31614 42578 31666 42590
rect 31950 42642 32002 42654
rect 31950 42578 32002 42590
rect 33406 42642 33458 42654
rect 33406 42578 33458 42590
rect 35870 42642 35922 42654
rect 35870 42578 35922 42590
rect 36430 42642 36482 42654
rect 39230 42642 39282 42654
rect 37314 42590 37326 42642
rect 37378 42590 37390 42642
rect 36430 42578 36482 42590
rect 39230 42578 39282 42590
rect 41022 42642 41074 42654
rect 41022 42578 41074 42590
rect 41918 42642 41970 42654
rect 41918 42578 41970 42590
rect 42254 42642 42306 42654
rect 44818 42590 44830 42642
rect 44882 42590 44894 42642
rect 42254 42578 42306 42590
rect 2046 42530 2098 42542
rect 2046 42466 2098 42478
rect 2494 42530 2546 42542
rect 2494 42466 2546 42478
rect 10222 42530 10274 42542
rect 10222 42466 10274 42478
rect 18622 42530 18674 42542
rect 18622 42466 18674 42478
rect 21646 42530 21698 42542
rect 21646 42466 21698 42478
rect 22766 42530 22818 42542
rect 22766 42466 22818 42478
rect 23102 42530 23154 42542
rect 23886 42530 23938 42542
rect 23426 42478 23438 42530
rect 23490 42478 23502 42530
rect 23102 42466 23154 42478
rect 23886 42466 23938 42478
rect 24782 42530 24834 42542
rect 24782 42466 24834 42478
rect 26350 42530 26402 42542
rect 26350 42466 26402 42478
rect 27022 42530 27074 42542
rect 27022 42466 27074 42478
rect 29934 42530 29986 42542
rect 29934 42466 29986 42478
rect 31166 42530 31218 42542
rect 31166 42466 31218 42478
rect 32958 42530 33010 42542
rect 32958 42466 33010 42478
rect 33854 42530 33906 42542
rect 33854 42466 33906 42478
rect 34750 42530 34802 42542
rect 34750 42466 34802 42478
rect 36318 42530 36370 42542
rect 36318 42466 36370 42478
rect 36990 42530 37042 42542
rect 36990 42466 37042 42478
rect 37998 42530 38050 42542
rect 37998 42466 38050 42478
rect 39118 42530 39170 42542
rect 39118 42466 39170 42478
rect 40014 42530 40066 42542
rect 40014 42466 40066 42478
rect 40910 42530 40962 42542
rect 40910 42466 40962 42478
rect 41806 42530 41858 42542
rect 41806 42466 41858 42478
rect 42366 42530 42418 42542
rect 42366 42466 42418 42478
rect 45166 42530 45218 42542
rect 45166 42466 45218 42478
rect 45726 42530 45778 42542
rect 45726 42466 45778 42478
rect 46622 42530 46674 42542
rect 46622 42466 46674 42478
rect 47406 42530 47458 42542
rect 47406 42466 47458 42478
rect 48526 42530 48578 42542
rect 48526 42466 48578 42478
rect 49310 42530 49362 42542
rect 49310 42466 49362 42478
rect 49534 42530 49586 42542
rect 49534 42466 49586 42478
rect 50542 42530 50594 42542
rect 50542 42466 50594 42478
rect 1344 42362 58576 42396
rect 1344 42310 19838 42362
rect 19890 42310 19942 42362
rect 19994 42310 20046 42362
rect 20098 42310 50558 42362
rect 50610 42310 50662 42362
rect 50714 42310 50766 42362
rect 50818 42310 58576 42362
rect 1344 42276 58576 42310
rect 10894 42194 10946 42206
rect 10894 42130 10946 42142
rect 25230 42194 25282 42206
rect 26910 42194 26962 42206
rect 26674 42142 26686 42194
rect 26738 42142 26750 42194
rect 25230 42130 25282 42142
rect 26910 42130 26962 42142
rect 35422 42194 35474 42206
rect 35422 42130 35474 42142
rect 37886 42194 37938 42206
rect 37886 42130 37938 42142
rect 39342 42194 39394 42206
rect 39342 42130 39394 42142
rect 42254 42194 42306 42206
rect 46510 42194 46562 42206
rect 45826 42142 45838 42194
rect 45890 42142 45902 42194
rect 42254 42130 42306 42142
rect 46510 42130 46562 42142
rect 48078 42194 48130 42206
rect 48078 42130 48130 42142
rect 2046 42082 2098 42094
rect 2046 42018 2098 42030
rect 9886 42082 9938 42094
rect 24558 42082 24610 42094
rect 13234 42030 13246 42082
rect 13298 42030 13310 42082
rect 18834 42030 18846 42082
rect 18898 42030 18910 42082
rect 22306 42030 22318 42082
rect 22370 42030 22382 42082
rect 9886 42018 9938 42030
rect 24558 42018 24610 42030
rect 27134 42082 27186 42094
rect 27134 42018 27186 42030
rect 27246 42082 27298 42094
rect 41022 42082 41074 42094
rect 30818 42030 30830 42082
rect 30882 42030 30894 42082
rect 27246 42018 27298 42030
rect 41022 42018 41074 42030
rect 47518 42082 47570 42094
rect 47518 42018 47570 42030
rect 49310 42082 49362 42094
rect 49310 42018 49362 42030
rect 49534 42082 49586 42094
rect 49534 42018 49586 42030
rect 1710 41970 1762 41982
rect 1710 41906 1762 41918
rect 9774 41970 9826 41982
rect 10782 41970 10834 41982
rect 10322 41918 10334 41970
rect 10386 41918 10398 41970
rect 9774 41906 9826 41918
rect 10782 41906 10834 41918
rect 11006 41970 11058 41982
rect 23886 41970 23938 41982
rect 12562 41918 12574 41970
rect 12626 41918 12638 41970
rect 19058 41918 19070 41970
rect 19122 41918 19134 41970
rect 23090 41918 23102 41970
rect 23154 41918 23166 41970
rect 11006 41906 11058 41918
rect 23886 41906 23938 41918
rect 24334 41970 24386 41982
rect 26126 41970 26178 41982
rect 27694 41970 27746 41982
rect 25442 41918 25454 41970
rect 25506 41918 25518 41970
rect 26450 41918 26462 41970
rect 26514 41918 26526 41970
rect 24334 41906 24386 41918
rect 26126 41906 26178 41918
rect 27694 41906 27746 41918
rect 29150 41970 29202 41982
rect 29150 41906 29202 41918
rect 29262 41970 29314 41982
rect 29262 41906 29314 41918
rect 29486 41970 29538 41982
rect 29486 41906 29538 41918
rect 29598 41970 29650 41982
rect 29598 41906 29650 41918
rect 30494 41970 30546 41982
rect 30494 41906 30546 41918
rect 33406 41970 33458 41982
rect 33406 41906 33458 41918
rect 34302 41970 34354 41982
rect 34302 41906 34354 41918
rect 34862 41970 34914 41982
rect 36766 41970 36818 41982
rect 35634 41918 35646 41970
rect 35698 41918 35710 41970
rect 34862 41906 34914 41918
rect 36766 41906 36818 41918
rect 37326 41970 37378 41982
rect 37326 41906 37378 41918
rect 37550 41970 37602 41982
rect 39006 41970 39058 41982
rect 38546 41918 38558 41970
rect 38610 41918 38622 41970
rect 37550 41906 37602 41918
rect 39006 41906 39058 41918
rect 39678 41970 39730 41982
rect 39678 41906 39730 41918
rect 41246 41970 41298 41982
rect 41246 41906 41298 41918
rect 41470 41970 41522 41982
rect 41470 41906 41522 41918
rect 41582 41970 41634 41982
rect 41582 41906 41634 41918
rect 46174 41970 46226 41982
rect 47182 41970 47234 41982
rect 46722 41918 46734 41970
rect 46786 41918 46798 41970
rect 49074 41918 49086 41970
rect 49138 41918 49150 41970
rect 49746 41918 49758 41970
rect 49810 41918 49822 41970
rect 53442 41918 53454 41970
rect 53506 41918 53518 41970
rect 46174 41906 46226 41918
rect 47182 41906 47234 41918
rect 2494 41858 2546 41870
rect 2494 41794 2546 41806
rect 10558 41858 10610 41870
rect 23774 41858 23826 41870
rect 15362 41806 15374 41858
rect 15426 41806 15438 41858
rect 20178 41806 20190 41858
rect 20242 41806 20254 41858
rect 10558 41794 10610 41806
rect 23774 41794 23826 41806
rect 24110 41858 24162 41870
rect 24110 41794 24162 41806
rect 29374 41858 29426 41870
rect 29374 41794 29426 41806
rect 33966 41858 34018 41870
rect 33966 41794 34018 41806
rect 36318 41858 36370 41870
rect 36318 41794 36370 41806
rect 41358 41858 41410 41870
rect 41358 41794 41410 41806
rect 49422 41858 49474 41870
rect 49422 41794 49474 41806
rect 53230 41858 53282 41870
rect 53230 41794 53282 41806
rect 9886 41746 9938 41758
rect 55346 41694 55358 41746
rect 55410 41694 55422 41746
rect 9886 41682 9938 41694
rect 1344 41578 58576 41612
rect 1344 41526 4478 41578
rect 4530 41526 4582 41578
rect 4634 41526 4686 41578
rect 4738 41526 35198 41578
rect 35250 41526 35302 41578
rect 35354 41526 35406 41578
rect 35458 41526 58576 41578
rect 1344 41492 58576 41526
rect 10782 41410 10834 41422
rect 10782 41346 10834 41358
rect 11006 41410 11058 41422
rect 11006 41346 11058 41358
rect 11678 41410 11730 41422
rect 50990 41410 51042 41422
rect 34402 41358 34414 41410
rect 34466 41407 34478 41410
rect 34962 41407 34974 41410
rect 34466 41361 34974 41407
rect 34466 41358 34478 41361
rect 34962 41358 34974 41361
rect 35026 41358 35038 41410
rect 11678 41346 11730 41358
rect 50990 41346 51042 41358
rect 57934 41410 57986 41422
rect 57934 41346 57986 41358
rect 10110 41298 10162 41310
rect 10110 41234 10162 41246
rect 15486 41298 15538 41310
rect 15486 41234 15538 41246
rect 16046 41298 16098 41310
rect 16046 41234 16098 41246
rect 21982 41298 22034 41310
rect 28030 41298 28082 41310
rect 26562 41246 26574 41298
rect 26626 41246 26638 41298
rect 27458 41246 27470 41298
rect 27522 41246 27534 41298
rect 21982 41234 22034 41246
rect 28030 41234 28082 41246
rect 28702 41298 28754 41310
rect 28702 41234 28754 41246
rect 29150 41298 29202 41310
rect 34414 41298 34466 41310
rect 32498 41246 32510 41298
rect 32562 41246 32574 41298
rect 29150 41234 29202 41246
rect 34414 41234 34466 41246
rect 38110 41298 38162 41310
rect 51102 41298 51154 41310
rect 41794 41246 41806 41298
rect 41858 41246 41870 41298
rect 43922 41246 43934 41298
rect 43986 41246 43998 41298
rect 48626 41246 48638 41298
rect 48690 41246 48702 41298
rect 38110 41234 38162 41246
rect 51102 41234 51154 41246
rect 55022 41298 55074 41310
rect 55022 41234 55074 41246
rect 10558 41186 10610 41198
rect 15710 41186 15762 41198
rect 19406 41186 19458 41198
rect 11218 41134 11230 41186
rect 11282 41134 11294 41186
rect 16594 41134 16606 41186
rect 16658 41134 16670 41186
rect 10558 41122 10610 41134
rect 15710 41122 15762 41134
rect 19406 41122 19458 41134
rect 19966 41186 20018 41198
rect 19966 41122 20018 41134
rect 24110 41186 24162 41198
rect 29262 41186 29314 41198
rect 35198 41186 35250 41198
rect 45166 41186 45218 41198
rect 51550 41186 51602 41198
rect 25554 41134 25566 41186
rect 25618 41134 25630 41186
rect 29698 41134 29710 41186
rect 29762 41134 29774 41186
rect 41122 41134 41134 41186
rect 41186 41134 41198 41186
rect 49186 41134 49198 41186
rect 49250 41134 49262 41186
rect 52658 41134 52670 41186
rect 52722 41134 52734 41186
rect 55570 41134 55582 41186
rect 55634 41134 55646 41186
rect 24110 41122 24162 41134
rect 29262 41122 29314 41134
rect 35198 41122 35250 41134
rect 45166 41122 45218 41134
rect 51550 41122 51602 41134
rect 1710 41074 1762 41086
rect 1710 41010 1762 41022
rect 2382 41074 2434 41086
rect 2382 41010 2434 41022
rect 2718 41074 2770 41086
rect 2718 41010 2770 41022
rect 11566 41074 11618 41086
rect 11566 41010 11618 41022
rect 12238 41074 12290 41086
rect 12238 41010 12290 41022
rect 18734 41074 18786 41086
rect 18734 41010 18786 41022
rect 21870 41074 21922 41086
rect 22990 41074 23042 41086
rect 25790 41074 25842 41086
rect 22642 41022 22654 41074
rect 22706 41022 22718 41074
rect 24770 41022 24782 41074
rect 24834 41022 24846 41074
rect 21870 41010 21922 41022
rect 22990 41010 23042 41022
rect 25790 41010 25842 41022
rect 27022 41074 27074 41086
rect 30370 41022 30382 41074
rect 30434 41022 30446 41074
rect 27022 41010 27074 41022
rect 2046 40962 2098 40974
rect 2046 40898 2098 40910
rect 3166 40962 3218 40974
rect 3166 40898 3218 40910
rect 10670 40962 10722 40974
rect 10670 40898 10722 40910
rect 11790 40962 11842 40974
rect 11790 40898 11842 40910
rect 12014 40962 12066 40974
rect 12014 40898 12066 40910
rect 12686 40962 12738 40974
rect 12686 40898 12738 40910
rect 16382 40962 16434 40974
rect 16382 40898 16434 40910
rect 18622 40962 18674 40974
rect 19630 40962 19682 40974
rect 19058 40910 19070 40962
rect 19122 40910 19134 40962
rect 18622 40898 18674 40910
rect 19630 40898 19682 40910
rect 19854 40962 19906 40974
rect 19854 40898 19906 40910
rect 23550 40962 23602 40974
rect 23550 40898 23602 40910
rect 25118 40962 25170 40974
rect 25118 40898 25170 40910
rect 26126 40962 26178 40974
rect 26126 40898 26178 40910
rect 34750 40962 34802 40974
rect 34750 40898 34802 40910
rect 51438 40962 51490 40974
rect 51438 40898 51490 40910
rect 1344 40794 58576 40828
rect 1344 40742 19838 40794
rect 19890 40742 19942 40794
rect 19994 40742 20046 40794
rect 20098 40742 50558 40794
rect 50610 40742 50662 40794
rect 50714 40742 50766 40794
rect 50818 40742 58576 40794
rect 1344 40708 58576 40742
rect 2494 40626 2546 40638
rect 21422 40626 21474 40638
rect 21074 40574 21086 40626
rect 21138 40574 21150 40626
rect 2494 40562 2546 40574
rect 21422 40562 21474 40574
rect 23102 40626 23154 40638
rect 23102 40562 23154 40574
rect 23886 40626 23938 40638
rect 23886 40562 23938 40574
rect 24446 40626 24498 40638
rect 24446 40562 24498 40574
rect 24670 40626 24722 40638
rect 24670 40562 24722 40574
rect 25342 40626 25394 40638
rect 25342 40562 25394 40574
rect 26910 40626 26962 40638
rect 26910 40562 26962 40574
rect 35310 40626 35362 40638
rect 35310 40562 35362 40574
rect 37214 40626 37266 40638
rect 37214 40562 37266 40574
rect 22094 40514 22146 40526
rect 2034 40462 2046 40514
rect 2098 40462 2110 40514
rect 16034 40462 16046 40514
rect 16098 40462 16110 40514
rect 18610 40462 18622 40514
rect 18674 40462 18686 40514
rect 22094 40450 22146 40462
rect 22766 40514 22818 40526
rect 22766 40450 22818 40462
rect 23438 40514 23490 40526
rect 23438 40450 23490 40462
rect 24334 40514 24386 40526
rect 24334 40450 24386 40462
rect 25790 40514 25842 40526
rect 34190 40514 34242 40526
rect 30594 40462 30606 40514
rect 30658 40462 30670 40514
rect 25790 40450 25842 40462
rect 34190 40450 34242 40462
rect 35758 40514 35810 40526
rect 35758 40450 35810 40462
rect 36318 40514 36370 40526
rect 36318 40450 36370 40462
rect 38446 40514 38498 40526
rect 49522 40462 49534 40514
rect 49586 40462 49598 40514
rect 38446 40450 38498 40462
rect 1710 40402 1762 40414
rect 1710 40338 1762 40350
rect 2942 40402 2994 40414
rect 2942 40338 2994 40350
rect 11230 40402 11282 40414
rect 23998 40402 24050 40414
rect 16818 40350 16830 40402
rect 16882 40350 16894 40402
rect 17826 40350 17838 40402
rect 17890 40350 17902 40402
rect 21858 40350 21870 40402
rect 21922 40350 21934 40402
rect 11230 40338 11282 40350
rect 23998 40338 24050 40350
rect 26462 40402 26514 40414
rect 33854 40402 33906 40414
rect 27234 40350 27246 40402
rect 27298 40350 27310 40402
rect 26462 40338 26514 40350
rect 33854 40338 33906 40350
rect 33966 40402 34018 40414
rect 34862 40402 34914 40414
rect 34402 40350 34414 40402
rect 34466 40350 34478 40402
rect 33966 40338 34018 40350
rect 34862 40338 34914 40350
rect 34974 40402 35026 40414
rect 34974 40338 35026 40350
rect 35198 40402 35250 40414
rect 35198 40338 35250 40350
rect 36206 40402 36258 40414
rect 36206 40338 36258 40350
rect 38670 40402 38722 40414
rect 38670 40338 38722 40350
rect 38894 40402 38946 40414
rect 38894 40338 38946 40350
rect 39006 40402 39058 40414
rect 39006 40338 39058 40350
rect 39566 40402 39618 40414
rect 39566 40338 39618 40350
rect 39678 40402 39730 40414
rect 39678 40338 39730 40350
rect 39902 40402 39954 40414
rect 39902 40338 39954 40350
rect 40014 40402 40066 40414
rect 41234 40350 41246 40402
rect 41298 40350 41310 40402
rect 42018 40350 42030 40402
rect 42082 40350 42094 40402
rect 44930 40350 44942 40402
rect 44994 40350 45006 40402
rect 48738 40350 48750 40402
rect 48802 40350 48814 40402
rect 53442 40350 53454 40402
rect 53506 40350 53518 40402
rect 40014 40338 40066 40350
rect 17390 40290 17442 40302
rect 34078 40290 34130 40302
rect 13906 40238 13918 40290
rect 13970 40238 13982 40290
rect 20738 40238 20750 40290
rect 20802 40238 20814 40290
rect 17390 40226 17442 40238
rect 34078 40226 34130 40238
rect 35086 40290 35138 40302
rect 35086 40226 35138 40238
rect 35870 40290 35922 40302
rect 35870 40226 35922 40238
rect 36878 40290 36930 40302
rect 36878 40226 36930 40238
rect 38782 40290 38834 40302
rect 38782 40226 38834 40238
rect 39790 40290 39842 40302
rect 44146 40238 44158 40290
rect 44210 40238 44222 40290
rect 45602 40238 45614 40290
rect 45666 40238 45678 40290
rect 47730 40238 47742 40290
rect 47794 40238 47806 40290
rect 51650 40238 51662 40290
rect 51714 40238 51726 40290
rect 39790 40226 39842 40238
rect 17502 40178 17554 40190
rect 17502 40114 17554 40126
rect 23886 40178 23938 40190
rect 55346 40126 55358 40178
rect 55410 40126 55422 40178
rect 23886 40114 23938 40126
rect 1344 40010 58576 40044
rect 1344 39958 4478 40010
rect 4530 39958 4582 40010
rect 4634 39958 4686 40010
rect 4738 39958 35198 40010
rect 35250 39958 35302 40010
rect 35354 39958 35406 40010
rect 35458 39958 58576 40010
rect 1344 39924 58576 39958
rect 42926 39842 42978 39854
rect 12898 39790 12910 39842
rect 12962 39790 12974 39842
rect 42926 39778 42978 39790
rect 57934 39842 57986 39854
rect 57934 39778 57986 39790
rect 13582 39730 13634 39742
rect 19742 39730 19794 39742
rect 20750 39730 20802 39742
rect 11106 39678 11118 39730
rect 11170 39678 11182 39730
rect 16818 39678 16830 39730
rect 16882 39678 16894 39730
rect 18946 39678 18958 39730
rect 19010 39678 19022 39730
rect 19954 39678 19966 39730
rect 20018 39678 20030 39730
rect 13582 39666 13634 39678
rect 19742 39666 19794 39678
rect 20750 39666 20802 39678
rect 21422 39730 21474 39742
rect 32398 39730 32450 39742
rect 41582 39730 41634 39742
rect 23202 39678 23214 39730
rect 23266 39678 23278 39730
rect 31266 39678 31278 39730
rect 31330 39678 31342 39730
rect 33954 39678 33966 39730
rect 34018 39678 34030 39730
rect 36082 39678 36094 39730
rect 36146 39678 36158 39730
rect 37874 39678 37886 39730
rect 37938 39678 37950 39730
rect 40002 39678 40014 39730
rect 40066 39678 40078 39730
rect 21422 39666 21474 39678
rect 32398 39666 32450 39678
rect 41582 39666 41634 39678
rect 43374 39730 43426 39742
rect 43374 39666 43426 39678
rect 43486 39730 43538 39742
rect 43486 39666 43538 39678
rect 47742 39730 47794 39742
rect 51426 39678 51438 39730
rect 51490 39678 51502 39730
rect 47742 39666 47794 39678
rect 19294 39618 19346 39630
rect 10434 39566 10446 39618
rect 10498 39566 10510 39618
rect 10994 39566 11006 39618
rect 11058 39566 11070 39618
rect 11666 39566 11678 39618
rect 11730 39566 11742 39618
rect 12674 39566 12686 39618
rect 12738 39566 12750 39618
rect 16034 39566 16046 39618
rect 16098 39566 16110 39618
rect 19294 39554 19346 39566
rect 19518 39618 19570 39630
rect 41470 39618 41522 39630
rect 43038 39618 43090 39630
rect 46286 39618 46338 39630
rect 26786 39566 26798 39618
rect 26850 39566 26862 39618
rect 30706 39566 30718 39618
rect 30770 39566 30782 39618
rect 31378 39566 31390 39618
rect 31442 39566 31454 39618
rect 33282 39566 33294 39618
rect 33346 39566 33358 39618
rect 37202 39566 37214 39618
rect 37266 39566 37278 39618
rect 40674 39566 40686 39618
rect 40738 39566 40750 39618
rect 41906 39566 41918 39618
rect 41970 39566 41982 39618
rect 45378 39566 45390 39618
rect 45442 39566 45454 39618
rect 45938 39566 45950 39618
rect 46002 39566 46014 39618
rect 19518 39554 19570 39566
rect 41470 39554 41522 39566
rect 43038 39554 43090 39566
rect 46286 39554 46338 39566
rect 46958 39618 47010 39630
rect 48626 39566 48638 39618
rect 48690 39566 48702 39618
rect 55570 39566 55582 39618
rect 55634 39566 55646 39618
rect 46958 39554 47010 39566
rect 1710 39506 1762 39518
rect 1710 39442 1762 39454
rect 2046 39506 2098 39518
rect 2046 39442 2098 39454
rect 12910 39506 12962 39518
rect 12910 39442 12962 39454
rect 15710 39506 15762 39518
rect 15710 39442 15762 39454
rect 19966 39506 20018 39518
rect 19966 39442 20018 39454
rect 29822 39506 29874 39518
rect 29822 39442 29874 39454
rect 31838 39506 31890 39518
rect 55358 39506 55410 39518
rect 40898 39454 40910 39506
rect 40962 39454 40974 39506
rect 47282 39454 47294 39506
rect 47346 39454 47358 39506
rect 49298 39454 49310 39506
rect 49362 39454 49374 39506
rect 31838 39442 31890 39454
rect 55358 39442 55410 39454
rect 2494 39394 2546 39406
rect 2494 39330 2546 39342
rect 13470 39394 13522 39406
rect 13470 39330 13522 39342
rect 14030 39394 14082 39406
rect 14030 39330 14082 39342
rect 15374 39394 15426 39406
rect 15374 39330 15426 39342
rect 15598 39394 15650 39406
rect 15598 39330 15650 39342
rect 20190 39394 20242 39406
rect 20190 39330 20242 39342
rect 27470 39394 27522 39406
rect 30942 39394 30994 39406
rect 30146 39342 30158 39394
rect 30210 39342 30222 39394
rect 27470 39330 27522 39342
rect 30942 39330 30994 39342
rect 31166 39394 31218 39406
rect 31166 39330 31218 39342
rect 31726 39394 31778 39406
rect 31726 39330 31778 39342
rect 41358 39394 41410 39406
rect 41358 39330 41410 39342
rect 41694 39394 41746 39406
rect 46174 39394 46226 39406
rect 45602 39342 45614 39394
rect 45666 39342 45678 39394
rect 41694 39330 41746 39342
rect 46174 39330 46226 39342
rect 46398 39394 46450 39406
rect 46398 39330 46450 39342
rect 46510 39394 46562 39406
rect 46510 39330 46562 39342
rect 47630 39394 47682 39406
rect 47630 39330 47682 39342
rect 1344 39226 58576 39260
rect 1344 39174 19838 39226
rect 19890 39174 19942 39226
rect 19994 39174 20046 39226
rect 20098 39174 50558 39226
rect 50610 39174 50662 39226
rect 50714 39174 50766 39226
rect 50818 39174 58576 39226
rect 1344 39140 58576 39174
rect 14590 39058 14642 39070
rect 16046 39058 16098 39070
rect 15250 39006 15262 39058
rect 15314 39006 15326 39058
rect 14590 38994 14642 39006
rect 16046 38994 16098 39006
rect 17502 39058 17554 39070
rect 17502 38994 17554 39006
rect 18062 39058 18114 39070
rect 18062 38994 18114 39006
rect 18510 39058 18562 39070
rect 18510 38994 18562 39006
rect 25454 39058 25506 39070
rect 25454 38994 25506 39006
rect 31726 39058 31778 39070
rect 32510 39058 32562 39070
rect 32162 39006 32174 39058
rect 32226 39006 32238 39058
rect 31726 38994 31778 39006
rect 32510 38994 32562 39006
rect 39342 39058 39394 39070
rect 39342 38994 39394 39006
rect 49086 39058 49138 39070
rect 49086 38994 49138 39006
rect 49198 39058 49250 39070
rect 49198 38994 49250 39006
rect 49310 39058 49362 39070
rect 49310 38994 49362 39006
rect 24670 38946 24722 38958
rect 31166 38946 31218 38958
rect 11890 38894 11902 38946
rect 11954 38894 11966 38946
rect 22082 38894 22094 38946
rect 22146 38894 22158 38946
rect 29586 38894 29598 38946
rect 29650 38894 29662 38946
rect 24670 38882 24722 38894
rect 31166 38882 31218 38894
rect 39454 38946 39506 38958
rect 39454 38882 39506 38894
rect 49646 38946 49698 38958
rect 49646 38882 49698 38894
rect 31390 38834 31442 38846
rect 4274 38782 4286 38834
rect 4338 38782 4350 38834
rect 11218 38782 11230 38834
rect 11282 38782 11294 38834
rect 15026 38782 15038 38834
rect 15090 38782 15102 38834
rect 20402 38782 20414 38834
rect 20466 38782 20478 38834
rect 20850 38782 20862 38834
rect 20914 38782 20926 38834
rect 21298 38782 21310 38834
rect 21362 38782 21374 38834
rect 30258 38782 30270 38834
rect 30322 38782 30334 38834
rect 31390 38770 31442 38782
rect 31614 38834 31666 38846
rect 41022 38834 41074 38846
rect 38322 38782 38334 38834
rect 38386 38782 38398 38834
rect 31614 38770 31666 38782
rect 41022 38770 41074 38782
rect 49422 38834 49474 38846
rect 53442 38782 53454 38834
rect 53506 38782 53518 38834
rect 49422 38770 49474 38782
rect 10670 38722 10722 38734
rect 10670 38658 10722 38670
rect 10782 38722 10834 38734
rect 15710 38722 15762 38734
rect 14018 38670 14030 38722
rect 14082 38670 14094 38722
rect 10782 38658 10834 38670
rect 15710 38658 15762 38670
rect 16606 38722 16658 38734
rect 24558 38722 24610 38734
rect 24210 38670 24222 38722
rect 24274 38670 24286 38722
rect 16606 38658 16658 38670
rect 24558 38658 24610 38670
rect 27246 38722 27298 38734
rect 30830 38722 30882 38734
rect 27458 38670 27470 38722
rect 27522 38670 27534 38722
rect 27246 38658 27298 38670
rect 30830 38658 30882 38670
rect 31502 38722 31554 38734
rect 38894 38722 38946 38734
rect 33282 38670 33294 38722
rect 33346 38670 33358 38722
rect 31502 38658 31554 38670
rect 38894 38658 38946 38670
rect 53230 38722 53282 38734
rect 53230 38658 53282 38670
rect 1934 38610 1986 38622
rect 1934 38546 1986 38558
rect 15598 38610 15650 38622
rect 40910 38610 40962 38622
rect 20850 38558 20862 38610
rect 20914 38558 20926 38610
rect 55346 38558 55358 38610
rect 55410 38558 55422 38610
rect 15598 38546 15650 38558
rect 40910 38546 40962 38558
rect 1344 38442 58576 38476
rect 1344 38390 4478 38442
rect 4530 38390 4582 38442
rect 4634 38390 4686 38442
rect 4738 38390 35198 38442
rect 35250 38390 35302 38442
rect 35354 38390 35406 38442
rect 35458 38390 58576 38442
rect 1344 38356 58576 38390
rect 22094 38274 22146 38286
rect 13458 38222 13470 38274
rect 13522 38222 13534 38274
rect 20738 38222 20750 38274
rect 20802 38222 20814 38274
rect 22094 38210 22146 38222
rect 27582 38274 27634 38286
rect 27582 38210 27634 38222
rect 33854 38274 33906 38286
rect 33854 38210 33906 38222
rect 57934 38274 57986 38286
rect 57934 38210 57986 38222
rect 18286 38162 18338 38174
rect 9762 38110 9774 38162
rect 9826 38110 9838 38162
rect 11890 38110 11902 38162
rect 11954 38110 11966 38162
rect 18286 38098 18338 38110
rect 21758 38162 21810 38174
rect 21758 38098 21810 38110
rect 23886 38162 23938 38174
rect 33966 38162 34018 38174
rect 43262 38162 43314 38174
rect 27122 38110 27134 38162
rect 27186 38110 27198 38162
rect 27906 38110 27918 38162
rect 27970 38110 27982 38162
rect 31378 38110 31390 38162
rect 31442 38110 31454 38162
rect 33506 38110 33518 38162
rect 33570 38110 33582 38162
rect 38210 38110 38222 38162
rect 38274 38110 38286 38162
rect 40338 38110 40350 38162
rect 40402 38110 40414 38162
rect 23886 38098 23938 38110
rect 33966 38098 34018 38110
rect 43262 38098 43314 38110
rect 14478 38050 14530 38062
rect 16158 38050 16210 38062
rect 17502 38050 17554 38062
rect 9090 37998 9102 38050
rect 9154 37998 9166 38050
rect 13682 37998 13694 38050
rect 13746 37998 13758 38050
rect 14578 37998 14590 38050
rect 14642 37998 14654 38050
rect 15698 37998 15710 38050
rect 15762 37998 15774 38050
rect 16706 37998 16718 38050
rect 16770 37998 16782 38050
rect 14478 37986 14530 37998
rect 16158 37986 16210 37998
rect 17502 37986 17554 37998
rect 17950 38050 18002 38062
rect 17950 37986 18002 37998
rect 18062 38050 18114 38062
rect 18062 37986 18114 37998
rect 18398 38050 18450 38062
rect 18398 37986 18450 37998
rect 18622 38050 18674 38062
rect 18622 37986 18674 37998
rect 19854 38050 19906 38062
rect 19854 37986 19906 37998
rect 20190 38050 20242 38062
rect 20190 37986 20242 37998
rect 20414 38050 20466 38062
rect 20414 37986 20466 37998
rect 22990 38050 23042 38062
rect 28478 38050 28530 38062
rect 24322 37998 24334 38050
rect 24386 37998 24398 38050
rect 22990 37986 23042 37998
rect 28478 37986 28530 37998
rect 29374 38050 29426 38062
rect 29374 37986 29426 37998
rect 30270 38050 30322 38062
rect 42254 38050 42306 38062
rect 47518 38050 47570 38062
rect 30594 37998 30606 38050
rect 30658 37998 30670 38050
rect 37426 37998 37438 38050
rect 37490 37998 37502 38050
rect 47170 37998 47182 38050
rect 47234 37998 47246 38050
rect 30270 37986 30322 37998
rect 42254 37986 42306 37998
rect 47518 37986 47570 37998
rect 55358 38050 55410 38062
rect 55570 37998 55582 38050
rect 55634 37998 55646 38050
rect 55358 37986 55410 37998
rect 1710 37938 1762 37950
rect 1710 37874 1762 37886
rect 13470 37938 13522 37950
rect 13470 37874 13522 37886
rect 17390 37938 17442 37950
rect 22206 37938 22258 37950
rect 30158 37938 30210 37950
rect 19506 37886 19518 37938
rect 19570 37886 19582 37938
rect 24994 37886 25006 37938
rect 25058 37886 25070 37938
rect 17390 37874 17442 37886
rect 22206 37874 22258 37886
rect 30158 37874 30210 37886
rect 43822 37938 43874 37950
rect 43822 37874 43874 37886
rect 46846 37938 46898 37950
rect 46846 37874 46898 37886
rect 48526 37938 48578 37950
rect 48526 37874 48578 37886
rect 2046 37826 2098 37838
rect 2046 37762 2098 37774
rect 2494 37826 2546 37838
rect 17278 37826 17330 37838
rect 16482 37774 16494 37826
rect 16546 37774 16558 37826
rect 2494 37762 2546 37774
rect 17278 37762 17330 37774
rect 19294 37826 19346 37838
rect 19294 37762 19346 37774
rect 22094 37826 22146 37838
rect 23326 37826 23378 37838
rect 22642 37774 22654 37826
rect 22706 37774 22718 37826
rect 22094 37762 22146 37774
rect 23326 37762 23378 37774
rect 27806 37826 27858 37838
rect 27806 37762 27858 37774
rect 28142 37826 28194 37838
rect 28142 37762 28194 37774
rect 28366 37826 28418 37838
rect 28366 37762 28418 37774
rect 29150 37826 29202 37838
rect 29150 37762 29202 37774
rect 29262 37826 29314 37838
rect 29262 37762 29314 37774
rect 29598 37826 29650 37838
rect 29598 37762 29650 37774
rect 29934 37826 29986 37838
rect 29934 37762 29986 37774
rect 34526 37826 34578 37838
rect 35422 37826 35474 37838
rect 34850 37774 34862 37826
rect 34914 37774 34926 37826
rect 34526 37762 34578 37774
rect 35422 37762 35474 37774
rect 42366 37826 42418 37838
rect 42366 37762 42418 37774
rect 42478 37826 42530 37838
rect 42478 37762 42530 37774
rect 42590 37826 42642 37838
rect 42590 37762 42642 37774
rect 42702 37826 42754 37838
rect 42702 37762 42754 37774
rect 43710 37826 43762 37838
rect 43710 37762 43762 37774
rect 46734 37826 46786 37838
rect 46734 37762 46786 37774
rect 47406 37826 47458 37838
rect 47406 37762 47458 37774
rect 47630 37826 47682 37838
rect 47630 37762 47682 37774
rect 47742 37826 47794 37838
rect 47742 37762 47794 37774
rect 48414 37826 48466 37838
rect 48414 37762 48466 37774
rect 1344 37658 58576 37692
rect 1344 37606 19838 37658
rect 19890 37606 19942 37658
rect 19994 37606 20046 37658
rect 20098 37606 50558 37658
rect 50610 37606 50662 37658
rect 50714 37606 50766 37658
rect 50818 37606 58576 37658
rect 1344 37572 58576 37606
rect 17614 37490 17666 37502
rect 17614 37426 17666 37438
rect 17838 37490 17890 37502
rect 17838 37426 17890 37438
rect 18958 37490 19010 37502
rect 18958 37426 19010 37438
rect 21870 37490 21922 37502
rect 21870 37426 21922 37438
rect 22990 37490 23042 37502
rect 22990 37426 23042 37438
rect 24334 37490 24386 37502
rect 24334 37426 24386 37438
rect 26126 37490 26178 37502
rect 26126 37426 26178 37438
rect 26238 37490 26290 37502
rect 26238 37426 26290 37438
rect 33630 37490 33682 37502
rect 33630 37426 33682 37438
rect 41470 37490 41522 37502
rect 41470 37426 41522 37438
rect 49310 37490 49362 37502
rect 49310 37426 49362 37438
rect 2046 37378 2098 37390
rect 20974 37378 21026 37390
rect 11778 37326 11790 37378
rect 11842 37326 11854 37378
rect 2046 37314 2098 37326
rect 20974 37314 21026 37326
rect 21198 37378 21250 37390
rect 21198 37314 21250 37326
rect 22094 37378 22146 37390
rect 22094 37314 22146 37326
rect 22766 37378 22818 37390
rect 22766 37314 22818 37326
rect 24558 37378 24610 37390
rect 24558 37314 24610 37326
rect 25342 37378 25394 37390
rect 30382 37378 30434 37390
rect 29138 37326 29150 37378
rect 29202 37326 29214 37378
rect 25342 37314 25394 37326
rect 30382 37314 30434 37326
rect 30494 37378 30546 37390
rect 30494 37314 30546 37326
rect 30942 37378 30994 37390
rect 30942 37314 30994 37326
rect 31390 37378 31442 37390
rect 31390 37314 31442 37326
rect 31502 37378 31554 37390
rect 34962 37326 34974 37378
rect 35026 37326 35038 37378
rect 42578 37326 42590 37378
rect 42642 37326 42654 37378
rect 31502 37314 31554 37326
rect 1710 37266 1762 37278
rect 18062 37266 18114 37278
rect 18622 37266 18674 37278
rect 16706 37214 16718 37266
rect 16770 37214 16782 37266
rect 18386 37214 18398 37266
rect 18450 37214 18462 37266
rect 1710 37202 1762 37214
rect 18062 37202 18114 37214
rect 18622 37202 18674 37214
rect 18846 37266 18898 37278
rect 20526 37266 20578 37278
rect 20066 37214 20078 37266
rect 20130 37214 20142 37266
rect 18846 37202 18898 37214
rect 20526 37202 20578 37214
rect 22206 37266 22258 37278
rect 22206 37202 22258 37214
rect 22654 37266 22706 37278
rect 24110 37266 24162 37278
rect 23650 37214 23662 37266
rect 23714 37214 23726 37266
rect 22654 37202 22706 37214
rect 24110 37202 24162 37214
rect 24670 37266 24722 37278
rect 24670 37202 24722 37214
rect 25454 37266 25506 37278
rect 25454 37202 25506 37214
rect 25678 37266 25730 37278
rect 25678 37202 25730 37214
rect 26350 37266 26402 37278
rect 30158 37266 30210 37278
rect 48862 37266 48914 37278
rect 29810 37214 29822 37266
rect 29874 37214 29886 37266
rect 34290 37214 34302 37266
rect 34354 37214 34366 37266
rect 37426 37214 37438 37266
rect 37490 37214 37502 37266
rect 41906 37214 41918 37266
rect 41970 37214 41982 37266
rect 45154 37214 45166 37266
rect 45218 37214 45230 37266
rect 26350 37202 26402 37214
rect 30158 37202 30210 37214
rect 48862 37202 48914 37214
rect 48974 37266 49026 37278
rect 48974 37202 49026 37214
rect 49198 37266 49250 37278
rect 53442 37214 53454 37266
rect 53506 37214 53518 37266
rect 49198 37202 49250 37214
rect 2494 37154 2546 37166
rect 2494 37090 2546 37102
rect 10334 37154 10386 37166
rect 10334 37090 10386 37102
rect 17950 37154 18002 37166
rect 19406 37154 19458 37166
rect 21646 37154 21698 37166
rect 41134 37154 41186 37166
rect 49086 37154 49138 37166
rect 18946 37102 18958 37154
rect 19010 37102 19022 37154
rect 20850 37102 20862 37154
rect 20914 37102 20926 37154
rect 27010 37102 27022 37154
rect 27074 37102 27086 37154
rect 37090 37102 37102 37154
rect 37154 37102 37166 37154
rect 38210 37102 38222 37154
rect 38274 37102 38286 37154
rect 40338 37102 40350 37154
rect 40402 37102 40414 37154
rect 44706 37102 44718 37154
rect 44770 37102 44782 37154
rect 45826 37102 45838 37154
rect 45890 37102 45902 37154
rect 47954 37102 47966 37154
rect 48018 37102 48030 37154
rect 17950 37090 18002 37102
rect 19406 37090 19458 37102
rect 21646 37090 21698 37102
rect 41134 37090 41186 37102
rect 49086 37090 49138 37102
rect 10222 37042 10274 37054
rect 10222 36978 10274 36990
rect 19518 37042 19570 37054
rect 19518 36978 19570 36990
rect 25342 37042 25394 37054
rect 25342 36978 25394 36990
rect 30830 37042 30882 37054
rect 30830 36978 30882 36990
rect 31502 37042 31554 37054
rect 55346 36990 55358 37042
rect 55410 36990 55422 37042
rect 31502 36978 31554 36990
rect 1344 36874 58576 36908
rect 1344 36822 4478 36874
rect 4530 36822 4582 36874
rect 4634 36822 4686 36874
rect 4738 36822 35198 36874
rect 35250 36822 35302 36874
rect 35354 36822 35406 36874
rect 35458 36822 58576 36874
rect 1344 36788 58576 36822
rect 16830 36706 16882 36718
rect 16830 36642 16882 36654
rect 50430 36706 50482 36718
rect 50430 36642 50482 36654
rect 57934 36706 57986 36718
rect 57934 36642 57986 36654
rect 1934 36594 1986 36606
rect 1934 36530 1986 36542
rect 4846 36594 4898 36606
rect 23662 36594 23714 36606
rect 9202 36542 9214 36594
rect 9266 36542 9278 36594
rect 11330 36542 11342 36594
rect 11394 36542 11406 36594
rect 14242 36542 14254 36594
rect 14306 36542 14318 36594
rect 16370 36542 16382 36594
rect 16434 36542 16446 36594
rect 17490 36542 17502 36594
rect 17554 36542 17566 36594
rect 19618 36542 19630 36594
rect 19682 36542 19694 36594
rect 4846 36530 4898 36542
rect 23662 36530 23714 36542
rect 24446 36594 24498 36606
rect 24446 36530 24498 36542
rect 27470 36594 27522 36606
rect 27470 36530 27522 36542
rect 29262 36594 29314 36606
rect 43486 36594 43538 36606
rect 35074 36542 35086 36594
rect 35138 36542 35150 36594
rect 29262 36530 29314 36542
rect 43486 36530 43538 36542
rect 55022 36594 55074 36606
rect 55022 36530 55074 36542
rect 21310 36482 21362 36494
rect 29374 36482 29426 36494
rect 4162 36430 4174 36482
rect 4226 36430 4238 36482
rect 8418 36430 8430 36482
rect 8482 36430 8494 36482
rect 13458 36430 13470 36482
rect 13522 36430 13534 36482
rect 20402 36430 20414 36482
rect 20466 36430 20478 36482
rect 25890 36430 25902 36482
rect 25954 36430 25966 36482
rect 21310 36418 21362 36430
rect 29374 36418 29426 36430
rect 29822 36482 29874 36494
rect 30718 36482 30770 36494
rect 30146 36430 30158 36482
rect 30210 36430 30222 36482
rect 29822 36418 29874 36430
rect 30718 36418 30770 36430
rect 31054 36482 31106 36494
rect 32162 36430 32174 36482
rect 32226 36430 32238 36482
rect 35634 36430 35646 36482
rect 35698 36430 35710 36482
rect 36306 36430 36318 36482
rect 36370 36430 36382 36482
rect 42242 36430 42254 36482
rect 42306 36430 42318 36482
rect 42802 36430 42814 36482
rect 42866 36430 42878 36482
rect 46162 36430 46174 36482
rect 46226 36430 46238 36482
rect 52770 36430 52782 36482
rect 52834 36430 52846 36482
rect 55570 36430 55582 36482
rect 55634 36430 55646 36482
rect 31054 36418 31106 36430
rect 16718 36370 16770 36382
rect 16718 36306 16770 36318
rect 21870 36370 21922 36382
rect 21870 36306 21922 36318
rect 22206 36370 22258 36382
rect 22206 36306 22258 36318
rect 22654 36370 22706 36382
rect 22654 36306 22706 36318
rect 22766 36370 22818 36382
rect 44270 36370 44322 36382
rect 50542 36370 50594 36382
rect 25666 36318 25678 36370
rect 25730 36318 25742 36370
rect 27234 36318 27246 36370
rect 27298 36318 27310 36370
rect 32946 36318 32958 36370
rect 33010 36318 33022 36370
rect 37202 36318 37214 36370
rect 37266 36318 37278 36370
rect 42578 36318 42590 36370
rect 42642 36318 42654 36370
rect 48738 36318 48750 36370
rect 48802 36318 48814 36370
rect 22766 36306 22818 36318
rect 44270 36306 44322 36318
rect 50542 36306 50594 36318
rect 50990 36370 51042 36382
rect 50990 36306 51042 36318
rect 12910 36258 12962 36270
rect 12910 36194 12962 36206
rect 16830 36258 16882 36270
rect 16830 36194 16882 36206
rect 21422 36258 21474 36270
rect 21422 36194 21474 36206
rect 21646 36258 21698 36270
rect 21646 36194 21698 36206
rect 22430 36258 22482 36270
rect 22430 36194 22482 36206
rect 23214 36258 23266 36270
rect 23214 36194 23266 36206
rect 24894 36258 24946 36270
rect 24894 36194 24946 36206
rect 28590 36258 28642 36270
rect 28590 36194 28642 36206
rect 29150 36258 29202 36270
rect 29150 36194 29202 36206
rect 30382 36258 30434 36270
rect 30382 36194 30434 36206
rect 30830 36258 30882 36270
rect 30830 36194 30882 36206
rect 35870 36258 35922 36270
rect 35870 36194 35922 36206
rect 35982 36258 36034 36270
rect 35982 36194 36034 36206
rect 36094 36258 36146 36270
rect 36094 36194 36146 36206
rect 43374 36258 43426 36270
rect 43374 36194 43426 36206
rect 44158 36258 44210 36270
rect 44158 36194 44210 36206
rect 50878 36258 50930 36270
rect 50878 36194 50930 36206
rect 52110 36258 52162 36270
rect 52110 36194 52162 36206
rect 1344 36090 58576 36124
rect 1344 36038 19838 36090
rect 19890 36038 19942 36090
rect 19994 36038 20046 36090
rect 20098 36038 50558 36090
rect 50610 36038 50662 36090
rect 50714 36038 50766 36090
rect 50818 36038 58576 36090
rect 1344 36004 58576 36038
rect 2718 35922 2770 35934
rect 20750 35922 20802 35934
rect 18050 35870 18062 35922
rect 18114 35870 18126 35922
rect 2718 35858 2770 35870
rect 20750 35858 20802 35870
rect 23550 35922 23602 35934
rect 23550 35858 23602 35870
rect 23998 35922 24050 35934
rect 23998 35858 24050 35870
rect 26014 35922 26066 35934
rect 26014 35858 26066 35870
rect 26462 35922 26514 35934
rect 26462 35858 26514 35870
rect 26910 35922 26962 35934
rect 26910 35858 26962 35870
rect 27358 35922 27410 35934
rect 27358 35858 27410 35870
rect 33518 35922 33570 35934
rect 33518 35858 33570 35870
rect 33630 35922 33682 35934
rect 33630 35858 33682 35870
rect 33742 35922 33794 35934
rect 33742 35858 33794 35870
rect 34414 35922 34466 35934
rect 34414 35858 34466 35870
rect 39790 35922 39842 35934
rect 39790 35858 39842 35870
rect 45166 35922 45218 35934
rect 45166 35858 45218 35870
rect 45502 35922 45554 35934
rect 46286 35922 46338 35934
rect 45826 35870 45838 35922
rect 45890 35870 45902 35922
rect 45502 35858 45554 35870
rect 46286 35858 46338 35870
rect 46398 35922 46450 35934
rect 46398 35858 46450 35870
rect 46510 35922 46562 35934
rect 46510 35858 46562 35870
rect 47966 35922 48018 35934
rect 47966 35858 48018 35870
rect 48078 35922 48130 35934
rect 48078 35858 48130 35870
rect 2046 35810 2098 35822
rect 19406 35810 19458 35822
rect 14354 35758 14366 35810
rect 14418 35758 14430 35810
rect 17490 35758 17502 35810
rect 17554 35758 17566 35810
rect 18946 35758 18958 35810
rect 19010 35758 19022 35810
rect 2046 35746 2098 35758
rect 19406 35746 19458 35758
rect 19742 35810 19794 35822
rect 22990 35810 23042 35822
rect 33182 35810 33234 35822
rect 20402 35758 20414 35810
rect 20466 35758 20478 35810
rect 30370 35758 30382 35810
rect 30434 35758 30446 35810
rect 19742 35746 19794 35758
rect 22990 35746 23042 35758
rect 33182 35746 33234 35758
rect 34526 35810 34578 35822
rect 38446 35810 38498 35822
rect 35970 35758 35982 35810
rect 36034 35758 36046 35810
rect 34526 35746 34578 35758
rect 38446 35746 38498 35758
rect 38782 35810 38834 35822
rect 38782 35746 38834 35758
rect 39454 35810 39506 35822
rect 39454 35746 39506 35758
rect 41022 35810 41074 35822
rect 41022 35746 41074 35758
rect 46846 35810 46898 35822
rect 49522 35758 49534 35810
rect 49586 35758 49598 35810
rect 46846 35746 46898 35758
rect 1710 35698 1762 35710
rect 1710 35634 1762 35646
rect 2382 35698 2434 35710
rect 2382 35634 2434 35646
rect 10558 35698 10610 35710
rect 12238 35698 12290 35710
rect 22318 35698 22370 35710
rect 10770 35646 10782 35698
rect 10834 35646 10846 35698
rect 11778 35646 11790 35698
rect 11842 35646 11854 35698
rect 12674 35646 12686 35698
rect 12738 35646 12750 35698
rect 13570 35646 13582 35698
rect 13634 35646 13646 35698
rect 17378 35646 17390 35698
rect 17442 35646 17454 35698
rect 18386 35646 18398 35698
rect 18450 35646 18462 35698
rect 21410 35646 21422 35698
rect 21474 35646 21486 35698
rect 10558 35634 10610 35646
rect 12238 35634 12290 35646
rect 22318 35634 22370 35646
rect 22654 35698 22706 35710
rect 33406 35698 33458 35710
rect 39678 35698 39730 35710
rect 25778 35646 25790 35698
rect 25842 35646 25854 35698
rect 29586 35646 29598 35698
rect 29650 35646 29662 35698
rect 35298 35646 35310 35698
rect 35362 35646 35374 35698
rect 22654 35634 22706 35646
rect 33406 35634 33458 35646
rect 39678 35634 39730 35646
rect 39902 35698 39954 35710
rect 40910 35698 40962 35710
rect 46622 35698 46674 35710
rect 40114 35646 40126 35698
rect 40178 35646 40190 35698
rect 41346 35646 41358 35698
rect 41410 35646 41422 35698
rect 39902 35634 39954 35646
rect 40910 35634 40962 35646
rect 46622 35634 46674 35646
rect 47630 35698 47682 35710
rect 47630 35634 47682 35646
rect 47742 35698 47794 35710
rect 48738 35646 48750 35698
rect 48802 35646 48814 35698
rect 53442 35646 53454 35698
rect 53506 35646 53518 35698
rect 47742 35634 47794 35646
rect 3166 35586 3218 35598
rect 3166 35522 3218 35534
rect 10222 35586 10274 35598
rect 22094 35586 22146 35598
rect 13122 35534 13134 35586
rect 13186 35534 13198 35586
rect 16482 35534 16494 35586
rect 16546 35534 16558 35586
rect 21634 35534 21646 35586
rect 21698 35534 21710 35586
rect 10222 35522 10274 35534
rect 22094 35522 22146 35534
rect 22542 35586 22594 35598
rect 44718 35586 44770 35598
rect 53230 35586 53282 35598
rect 32498 35534 32510 35586
rect 32562 35534 32574 35586
rect 38098 35534 38110 35586
rect 38162 35534 38174 35586
rect 42130 35534 42142 35586
rect 42194 35534 42206 35586
rect 44258 35534 44270 35586
rect 44322 35534 44334 35586
rect 47954 35534 47966 35586
rect 48018 35534 48030 35586
rect 51650 35534 51662 35586
rect 51714 35534 51726 35586
rect 22542 35522 22594 35534
rect 44718 35522 44770 35534
rect 53230 35522 53282 35534
rect 10110 35474 10162 35486
rect 11106 35422 11118 35474
rect 11170 35422 11182 35474
rect 55346 35422 55358 35474
rect 55410 35422 55422 35474
rect 10110 35410 10162 35422
rect 1344 35306 58576 35340
rect 1344 35254 4478 35306
rect 4530 35254 4582 35306
rect 4634 35254 4686 35306
rect 4738 35254 35198 35306
rect 35250 35254 35302 35306
rect 35354 35254 35406 35306
rect 35458 35254 58576 35306
rect 1344 35220 58576 35254
rect 16830 35138 16882 35150
rect 16830 35074 16882 35086
rect 16942 35138 16994 35150
rect 16942 35074 16994 35086
rect 17278 35138 17330 35150
rect 17278 35074 17330 35086
rect 32062 35138 32114 35150
rect 32062 35074 32114 35086
rect 33294 35138 33346 35150
rect 33294 35074 33346 35086
rect 37102 35138 37154 35150
rect 43262 35138 43314 35150
rect 37426 35086 37438 35138
rect 37490 35135 37502 35138
rect 38098 35135 38110 35138
rect 37490 35089 38110 35135
rect 37490 35086 37502 35089
rect 38098 35086 38110 35089
rect 38162 35086 38174 35138
rect 37102 35074 37154 35086
rect 43262 35074 43314 35086
rect 44942 35138 44994 35150
rect 44942 35074 44994 35086
rect 56590 35138 56642 35150
rect 56590 35074 56642 35086
rect 2494 35026 2546 35038
rect 17726 35026 17778 35038
rect 9090 34974 9102 35026
rect 9154 34974 9166 35026
rect 11218 34974 11230 35026
rect 11282 34974 11294 35026
rect 12450 34974 12462 35026
rect 12514 34974 12526 35026
rect 16370 34974 16382 35026
rect 16434 34974 16446 35026
rect 2494 34962 2546 34974
rect 17726 34962 17778 34974
rect 18510 35026 18562 35038
rect 18510 34962 18562 34974
rect 19070 35026 19122 35038
rect 30606 35026 30658 35038
rect 22642 34974 22654 35026
rect 22706 34974 22718 35026
rect 19070 34962 19122 34974
rect 30606 34962 30658 34974
rect 36542 35026 36594 35038
rect 36542 34962 36594 34974
rect 37214 35026 37266 35038
rect 41682 34974 41694 35026
rect 41746 34974 41758 35026
rect 47058 34974 47070 35026
rect 47122 34974 47134 35026
rect 49186 34974 49198 35026
rect 49250 34974 49262 35026
rect 37214 34962 37266 34974
rect 17166 34914 17218 34926
rect 8418 34862 8430 34914
rect 8482 34862 8494 34914
rect 13458 34862 13470 34914
rect 13522 34862 13534 34914
rect 17166 34850 17218 34862
rect 18062 34914 18114 34926
rect 18062 34850 18114 34862
rect 18734 34914 18786 34926
rect 18734 34850 18786 34862
rect 21646 34914 21698 34926
rect 21646 34850 21698 34862
rect 22318 34914 22370 34926
rect 26238 34914 26290 34926
rect 25554 34862 25566 34914
rect 25618 34862 25630 34914
rect 22318 34850 22370 34862
rect 26238 34850 26290 34862
rect 26910 34914 26962 34926
rect 26910 34850 26962 34862
rect 27022 34914 27074 34926
rect 27022 34850 27074 34862
rect 27470 34914 27522 34926
rect 27918 34914 27970 34926
rect 27682 34862 27694 34914
rect 27746 34862 27758 34914
rect 27470 34850 27522 34862
rect 27918 34850 27970 34862
rect 31278 34914 31330 34926
rect 31278 34850 31330 34862
rect 32510 34914 32562 34926
rect 32510 34850 32562 34862
rect 34302 34914 34354 34926
rect 35086 34914 35138 34926
rect 34738 34862 34750 34914
rect 34802 34862 34814 34914
rect 34302 34850 34354 34862
rect 35086 34850 35138 34862
rect 36094 34914 36146 34926
rect 36094 34850 36146 34862
rect 38446 34914 38498 34926
rect 38446 34850 38498 34862
rect 41246 34914 41298 34926
rect 41246 34850 41298 34862
rect 41582 34914 41634 34926
rect 41582 34850 41634 34862
rect 42254 34914 42306 34926
rect 42254 34850 42306 34862
rect 42590 34914 42642 34926
rect 42590 34850 42642 34862
rect 42702 34914 42754 34926
rect 45714 34862 45726 34914
rect 45778 34862 45790 34914
rect 46386 34862 46398 34914
rect 46450 34862 46462 34914
rect 55570 34862 55582 34914
rect 55634 34862 55646 34914
rect 42702 34850 42754 34862
rect 1710 34802 1762 34814
rect 18286 34802 18338 34814
rect 14242 34750 14254 34802
rect 14306 34750 14318 34802
rect 1710 34738 1762 34750
rect 18286 34738 18338 34750
rect 20638 34802 20690 34814
rect 20638 34738 20690 34750
rect 20750 34802 20802 34814
rect 20750 34738 20802 34750
rect 21758 34802 21810 34814
rect 28030 34802 28082 34814
rect 31950 34802 32002 34814
rect 24770 34750 24782 34802
rect 24834 34750 24846 34802
rect 31602 34750 31614 34802
rect 31666 34750 31678 34802
rect 21758 34738 21810 34750
rect 28030 34738 28082 34750
rect 31950 34738 32002 34750
rect 33182 34802 33234 34814
rect 33182 34738 33234 34750
rect 35422 34802 35474 34814
rect 35422 34738 35474 34750
rect 35758 34802 35810 34814
rect 35758 34738 35810 34750
rect 38782 34802 38834 34814
rect 38782 34738 38834 34750
rect 39678 34802 39730 34814
rect 43150 34802 43202 34814
rect 40450 34750 40462 34802
rect 40514 34750 40526 34802
rect 39678 34738 39730 34750
rect 43150 34738 43202 34750
rect 43934 34802 43986 34814
rect 43934 34738 43986 34750
rect 44830 34802 44882 34814
rect 44830 34738 44882 34750
rect 2046 34690 2098 34702
rect 2046 34626 2098 34638
rect 2942 34690 2994 34702
rect 2942 34626 2994 34638
rect 12126 34690 12178 34702
rect 12126 34626 12178 34638
rect 12910 34690 12962 34702
rect 12910 34626 12962 34638
rect 20414 34690 20466 34702
rect 20414 34626 20466 34638
rect 21870 34690 21922 34702
rect 27246 34690 27298 34702
rect 29262 34690 29314 34702
rect 25890 34638 25902 34690
rect 25954 34638 25966 34690
rect 28466 34638 28478 34690
rect 28530 34638 28542 34690
rect 21870 34626 21922 34638
rect 27246 34626 27298 34638
rect 29262 34626 29314 34638
rect 32062 34690 32114 34702
rect 33294 34690 33346 34702
rect 32834 34638 32846 34690
rect 32898 34638 32910 34690
rect 32062 34626 32114 34638
rect 33294 34626 33346 34638
rect 33854 34690 33906 34702
rect 33854 34626 33906 34638
rect 35310 34690 35362 34702
rect 35310 34626 35362 34638
rect 35870 34690 35922 34702
rect 35870 34626 35922 34638
rect 37662 34690 37714 34702
rect 37662 34626 37714 34638
rect 38222 34690 38274 34702
rect 38222 34626 38274 34638
rect 38670 34690 38722 34702
rect 38670 34626 38722 34638
rect 39342 34690 39394 34702
rect 39342 34626 39394 34638
rect 40126 34690 40178 34702
rect 40126 34626 40178 34638
rect 41358 34690 41410 34702
rect 41358 34626 41410 34638
rect 41694 34690 41746 34702
rect 41694 34626 41746 34638
rect 42366 34690 42418 34702
rect 42366 34626 42418 34638
rect 42478 34690 42530 34702
rect 42478 34626 42530 34638
rect 43262 34690 43314 34702
rect 43262 34626 43314 34638
rect 43598 34690 43650 34702
rect 43598 34626 43650 34638
rect 43822 34690 43874 34702
rect 43822 34626 43874 34638
rect 44942 34690 44994 34702
rect 44942 34626 44994 34638
rect 45950 34690 46002 34702
rect 45950 34626 46002 34638
rect 1344 34522 58576 34556
rect 1344 34470 19838 34522
rect 19890 34470 19942 34522
rect 19994 34470 20046 34522
rect 20098 34470 50558 34522
rect 50610 34470 50662 34522
rect 50714 34470 50766 34522
rect 50818 34470 58576 34522
rect 1344 34436 58576 34470
rect 16158 34354 16210 34366
rect 15138 34302 15150 34354
rect 15202 34302 15214 34354
rect 16158 34290 16210 34302
rect 24334 34354 24386 34366
rect 24334 34290 24386 34302
rect 26574 34354 26626 34366
rect 26574 34290 26626 34302
rect 27694 34354 27746 34366
rect 27694 34290 27746 34302
rect 30942 34354 30994 34366
rect 30942 34290 30994 34302
rect 31726 34354 31778 34366
rect 31726 34290 31778 34302
rect 33854 34354 33906 34366
rect 33854 34290 33906 34302
rect 34302 34354 34354 34366
rect 34302 34290 34354 34302
rect 38782 34354 38834 34366
rect 38782 34290 38834 34302
rect 39678 34354 39730 34366
rect 39678 34290 39730 34302
rect 39790 34354 39842 34366
rect 39790 34290 39842 34302
rect 41246 34354 41298 34366
rect 41246 34290 41298 34302
rect 45950 34354 46002 34366
rect 45950 34290 46002 34302
rect 46510 34354 46562 34366
rect 46510 34290 46562 34302
rect 47406 34354 47458 34366
rect 47406 34290 47458 34302
rect 47630 34354 47682 34366
rect 47630 34290 47682 34302
rect 15710 34242 15762 34254
rect 15710 34178 15762 34190
rect 23998 34242 24050 34254
rect 23998 34178 24050 34190
rect 25230 34242 25282 34254
rect 29486 34242 29538 34254
rect 39342 34242 39394 34254
rect 26226 34190 26238 34242
rect 26290 34190 26302 34242
rect 28018 34190 28030 34242
rect 28082 34190 28094 34242
rect 31266 34190 31278 34242
rect 31330 34190 31342 34242
rect 25230 34178 25282 34190
rect 29486 34178 29538 34190
rect 39342 34178 39394 34190
rect 39454 34242 39506 34254
rect 39454 34178 39506 34190
rect 40014 34242 40066 34254
rect 40014 34178 40066 34190
rect 40126 34242 40178 34254
rect 40126 34178 40178 34190
rect 40910 34242 40962 34254
rect 40910 34178 40962 34190
rect 41022 34242 41074 34254
rect 45614 34242 45666 34254
rect 46734 34242 46786 34254
rect 42242 34190 42254 34242
rect 42306 34190 42318 34242
rect 46274 34190 46286 34242
rect 46338 34190 46350 34242
rect 41022 34178 41074 34190
rect 45614 34178 45666 34190
rect 46734 34178 46786 34190
rect 46846 34242 46898 34254
rect 49522 34190 49534 34242
rect 49586 34190 49598 34242
rect 46846 34178 46898 34190
rect 10558 34130 10610 34142
rect 12238 34130 12290 34142
rect 13582 34130 13634 34142
rect 16270 34130 16322 34142
rect 4274 34078 4286 34130
rect 4338 34078 4350 34130
rect 10994 34078 11006 34130
rect 11058 34078 11070 34130
rect 11778 34078 11790 34130
rect 11842 34078 11854 34130
rect 13010 34078 13022 34130
rect 13074 34078 13086 34130
rect 14018 34078 14030 34130
rect 14082 34078 14094 34130
rect 10558 34066 10610 34078
rect 12238 34066 12290 34078
rect 13582 34066 13634 34078
rect 16270 34066 16322 34078
rect 23662 34130 23714 34142
rect 23662 34066 23714 34078
rect 24222 34130 24274 34142
rect 24222 34066 24274 34078
rect 24446 34130 24498 34142
rect 25454 34130 25506 34142
rect 24658 34078 24670 34130
rect 24722 34078 24734 34130
rect 24446 34066 24498 34078
rect 25454 34066 25506 34078
rect 25678 34130 25730 34142
rect 25678 34066 25730 34078
rect 25790 34130 25842 34142
rect 25790 34066 25842 34078
rect 26910 34130 26962 34142
rect 29822 34130 29874 34142
rect 28354 34078 28366 34130
rect 28418 34078 28430 34130
rect 28914 34078 28926 34130
rect 28978 34078 28990 34130
rect 29586 34078 29598 34130
rect 29650 34078 29662 34130
rect 26910 34066 26962 34078
rect 29822 34066 29874 34078
rect 34414 34130 34466 34142
rect 34414 34066 34466 34078
rect 34750 34130 34802 34142
rect 34750 34066 34802 34078
rect 35086 34130 35138 34142
rect 47742 34130 47794 34142
rect 35522 34078 35534 34130
rect 35586 34078 35598 34130
rect 41458 34078 41470 34130
rect 41522 34078 41534 34130
rect 48738 34078 48750 34130
rect 48802 34078 48814 34130
rect 53442 34078 53454 34130
rect 53506 34078 53518 34130
rect 35086 34066 35138 34078
rect 47742 34066 47794 34078
rect 4734 34018 4786 34030
rect 23214 34018 23266 34030
rect 13234 33966 13246 34018
rect 13298 33966 13310 34018
rect 4734 33954 4786 33966
rect 23214 33954 23266 33966
rect 23550 34018 23602 34030
rect 23550 33954 23602 33966
rect 25566 34018 25618 34030
rect 25566 33954 25618 33966
rect 27022 34018 27074 34030
rect 32398 34018 32450 34030
rect 28578 33966 28590 34018
rect 28642 33966 28654 34018
rect 27022 33954 27074 33966
rect 32398 33954 32450 33966
rect 33294 34018 33346 34030
rect 33294 33954 33346 33966
rect 34638 34018 34690 34030
rect 44830 34018 44882 34030
rect 36194 33966 36206 34018
rect 36258 33966 36270 34018
rect 38322 33966 38334 34018
rect 38386 33966 38398 34018
rect 44370 33966 44382 34018
rect 44434 33966 44446 34018
rect 34638 33954 34690 33966
rect 44830 33954 44882 33966
rect 48190 34018 48242 34030
rect 51650 33966 51662 34018
rect 51714 33966 51726 34018
rect 48190 33954 48242 33966
rect 1934 33906 1986 33918
rect 15486 33906 15538 33918
rect 11106 33854 11118 33906
rect 11170 33854 11182 33906
rect 1934 33842 1986 33854
rect 15486 33842 15538 33854
rect 16158 33906 16210 33918
rect 55346 33854 55358 33906
rect 55410 33854 55422 33906
rect 16158 33842 16210 33854
rect 1344 33738 58576 33772
rect 1344 33686 4478 33738
rect 4530 33686 4582 33738
rect 4634 33686 4686 33738
rect 4738 33686 35198 33738
rect 35250 33686 35302 33738
rect 35354 33686 35406 33738
rect 35458 33686 58576 33738
rect 1344 33652 58576 33686
rect 14590 33570 14642 33582
rect 14590 33506 14642 33518
rect 27470 33570 27522 33582
rect 27470 33506 27522 33518
rect 34414 33570 34466 33582
rect 34414 33506 34466 33518
rect 48078 33570 48130 33582
rect 48078 33506 48130 33518
rect 48862 33570 48914 33582
rect 48862 33506 48914 33518
rect 49422 33570 49474 33582
rect 49422 33506 49474 33518
rect 50542 33570 50594 33582
rect 50542 33506 50594 33518
rect 57934 33570 57986 33582
rect 57934 33506 57986 33518
rect 18062 33458 18114 33470
rect 11106 33406 11118 33458
rect 11170 33406 11182 33458
rect 18062 33394 18114 33406
rect 18510 33458 18562 33470
rect 18510 33394 18562 33406
rect 21982 33458 22034 33470
rect 32622 33458 32674 33470
rect 23090 33406 23102 33458
rect 23154 33406 23166 33458
rect 25218 33406 25230 33458
rect 25282 33406 25294 33458
rect 21982 33394 22034 33406
rect 32622 33394 32674 33406
rect 35982 33458 36034 33470
rect 35982 33394 36034 33406
rect 18846 33346 18898 33358
rect 8194 33294 8206 33346
rect 8258 33294 8270 33346
rect 14914 33294 14926 33346
rect 14978 33294 14990 33346
rect 15138 33294 15150 33346
rect 15202 33294 15214 33346
rect 18846 33282 18898 33294
rect 19630 33346 19682 33358
rect 27694 33346 27746 33358
rect 25890 33294 25902 33346
rect 25954 33294 25966 33346
rect 19630 33282 19682 33294
rect 27694 33282 27746 33294
rect 27918 33346 27970 33358
rect 27918 33282 27970 33294
rect 28590 33346 28642 33358
rect 28590 33282 28642 33294
rect 30046 33346 30098 33358
rect 30046 33282 30098 33294
rect 31502 33346 31554 33358
rect 31502 33282 31554 33294
rect 34862 33346 34914 33358
rect 34862 33282 34914 33294
rect 35086 33346 35138 33358
rect 35086 33282 35138 33294
rect 36542 33346 36594 33358
rect 36542 33282 36594 33294
rect 36878 33346 36930 33358
rect 36878 33282 36930 33294
rect 37214 33346 37266 33358
rect 37214 33282 37266 33294
rect 37662 33346 37714 33358
rect 37662 33282 37714 33294
rect 40910 33346 40962 33358
rect 40910 33282 40962 33294
rect 41246 33346 41298 33358
rect 41246 33282 41298 33294
rect 46062 33346 46114 33358
rect 46062 33282 46114 33294
rect 46398 33346 46450 33358
rect 46398 33282 46450 33294
rect 47966 33346 48018 33358
rect 47966 33282 48018 33294
rect 48750 33346 48802 33358
rect 48750 33282 48802 33294
rect 49534 33346 49586 33358
rect 49534 33282 49586 33294
rect 49758 33346 49810 33358
rect 49758 33282 49810 33294
rect 50094 33346 50146 33358
rect 50094 33282 50146 33294
rect 50654 33346 50706 33358
rect 55570 33294 55582 33346
rect 55634 33294 55646 33346
rect 50654 33282 50706 33294
rect 1710 33234 1762 33246
rect 14702 33234 14754 33246
rect 8978 33182 8990 33234
rect 9042 33182 9054 33234
rect 1710 33170 1762 33182
rect 14702 33170 14754 33182
rect 16942 33234 16994 33246
rect 29374 33234 29426 33246
rect 34974 33234 35026 33246
rect 27122 33182 27134 33234
rect 27186 33182 27198 33234
rect 32162 33182 32174 33234
rect 32226 33182 32238 33234
rect 16942 33170 16994 33182
rect 29374 33170 29426 33182
rect 34974 33170 35026 33182
rect 55358 33234 55410 33246
rect 55358 33170 55410 33182
rect 2046 33122 2098 33134
rect 2046 33058 2098 33070
rect 2494 33122 2546 33134
rect 26574 33122 26626 33134
rect 19170 33070 19182 33122
rect 19234 33070 19246 33122
rect 2494 33058 2546 33070
rect 26574 33058 26626 33070
rect 28366 33122 28418 33134
rect 28366 33058 28418 33070
rect 28478 33122 28530 33134
rect 28478 33058 28530 33070
rect 29150 33122 29202 33134
rect 29150 33058 29202 33070
rect 29262 33122 29314 33134
rect 29262 33058 29314 33070
rect 29598 33122 29650 33134
rect 29598 33058 29650 33070
rect 30158 33122 30210 33134
rect 30158 33058 30210 33070
rect 30382 33122 30434 33134
rect 30382 33058 30434 33070
rect 30830 33122 30882 33134
rect 31838 33122 31890 33134
rect 31154 33070 31166 33122
rect 31218 33070 31230 33122
rect 30830 33058 30882 33070
rect 31838 33058 31890 33070
rect 34190 33122 34242 33134
rect 34190 33058 34242 33070
rect 34302 33122 34354 33134
rect 35870 33122 35922 33134
rect 35522 33070 35534 33122
rect 35586 33070 35598 33122
rect 34302 33058 34354 33070
rect 35870 33058 35922 33070
rect 36094 33122 36146 33134
rect 36094 33058 36146 33070
rect 37102 33122 37154 33134
rect 37102 33058 37154 33070
rect 38110 33122 38162 33134
rect 38110 33058 38162 33070
rect 39566 33122 39618 33134
rect 39566 33058 39618 33070
rect 40686 33122 40738 33134
rect 40686 33058 40738 33070
rect 41022 33122 41074 33134
rect 41022 33058 41074 33070
rect 43374 33122 43426 33134
rect 43374 33058 43426 33070
rect 46286 33122 46338 33134
rect 46286 33058 46338 33070
rect 47742 33122 47794 33134
rect 47742 33058 47794 33070
rect 48078 33122 48130 33134
rect 48078 33058 48130 33070
rect 48862 33122 48914 33134
rect 48862 33058 48914 33070
rect 49422 33122 49474 33134
rect 49422 33058 49474 33070
rect 49982 33122 50034 33134
rect 49982 33058 50034 33070
rect 50542 33122 50594 33134
rect 50542 33058 50594 33070
rect 1344 32954 58576 32988
rect 1344 32902 19838 32954
rect 19890 32902 19942 32954
rect 19994 32902 20046 32954
rect 20098 32902 50558 32954
rect 50610 32902 50662 32954
rect 50714 32902 50766 32954
rect 50818 32902 58576 32954
rect 1344 32868 58576 32902
rect 9886 32786 9938 32798
rect 9426 32734 9438 32786
rect 9490 32783 9502 32786
rect 9650 32783 9662 32786
rect 9490 32737 9662 32783
rect 9490 32734 9502 32737
rect 9650 32734 9662 32737
rect 9714 32734 9726 32786
rect 9886 32722 9938 32734
rect 14926 32786 14978 32798
rect 18734 32786 18786 32798
rect 16146 32734 16158 32786
rect 16210 32734 16222 32786
rect 14926 32722 14978 32734
rect 18734 32722 18786 32734
rect 22430 32786 22482 32798
rect 22430 32722 22482 32734
rect 24782 32786 24834 32798
rect 24782 32722 24834 32734
rect 25118 32786 25170 32798
rect 25118 32722 25170 32734
rect 30942 32786 30994 32798
rect 30942 32722 30994 32734
rect 34190 32786 34242 32798
rect 34190 32722 34242 32734
rect 34414 32786 34466 32798
rect 34414 32722 34466 32734
rect 35198 32786 35250 32798
rect 35198 32722 35250 32734
rect 35534 32786 35586 32798
rect 35534 32722 35586 32734
rect 43038 32786 43090 32798
rect 43038 32722 43090 32734
rect 2046 32674 2098 32686
rect 2046 32610 2098 32622
rect 15150 32674 15202 32686
rect 15150 32610 15202 32622
rect 16718 32674 16770 32686
rect 16718 32610 16770 32622
rect 17614 32674 17666 32686
rect 17614 32610 17666 32622
rect 17726 32674 17778 32686
rect 17726 32610 17778 32622
rect 17950 32674 18002 32686
rect 22542 32674 22594 32686
rect 19842 32622 19854 32674
rect 19906 32622 19918 32674
rect 17950 32610 18002 32622
rect 22542 32610 22594 32622
rect 24558 32674 24610 32686
rect 24558 32610 24610 32622
rect 25342 32674 25394 32686
rect 25342 32610 25394 32622
rect 26238 32674 26290 32686
rect 33630 32674 33682 32686
rect 35982 32674 36034 32686
rect 26562 32622 26574 32674
rect 26626 32622 26638 32674
rect 29026 32622 29038 32674
rect 29090 32622 29102 32674
rect 31266 32622 31278 32674
rect 31330 32622 31342 32674
rect 34738 32622 34750 32674
rect 34802 32622 34814 32674
rect 26238 32610 26290 32622
rect 33630 32610 33682 32622
rect 35982 32610 36034 32622
rect 1710 32562 1762 32574
rect 13134 32562 13186 32574
rect 11778 32510 11790 32562
rect 11842 32510 11854 32562
rect 12114 32510 12126 32562
rect 12178 32510 12190 32562
rect 12674 32510 12686 32562
rect 12738 32510 12750 32562
rect 1710 32498 1762 32510
rect 13134 32498 13186 32510
rect 13470 32562 13522 32574
rect 14590 32562 14642 32574
rect 13570 32510 13582 32562
rect 13634 32510 13646 32562
rect 13470 32498 13522 32510
rect 14590 32498 14642 32510
rect 16494 32562 16546 32574
rect 16494 32498 16546 32510
rect 18062 32562 18114 32574
rect 18062 32498 18114 32510
rect 18510 32562 18562 32574
rect 22766 32562 22818 32574
rect 24446 32562 24498 32574
rect 19170 32510 19182 32562
rect 19234 32510 19246 32562
rect 22978 32510 22990 32562
rect 23042 32510 23054 32562
rect 18510 32498 18562 32510
rect 22766 32498 22818 32510
rect 24446 32498 24498 32510
rect 25454 32562 25506 32574
rect 31614 32562 31666 32574
rect 29810 32510 29822 32562
rect 29874 32510 29886 32562
rect 25454 32498 25506 32510
rect 31614 32498 31666 32510
rect 32174 32562 32226 32574
rect 35422 32562 35474 32574
rect 33170 32510 33182 32562
rect 33234 32510 33246 32562
rect 32174 32498 32226 32510
rect 35422 32498 35474 32510
rect 35646 32562 35698 32574
rect 35646 32498 35698 32510
rect 36318 32562 36370 32574
rect 36318 32498 36370 32510
rect 36542 32562 36594 32574
rect 37426 32510 37438 32562
rect 37490 32510 37502 32562
rect 43698 32510 43710 32562
rect 43762 32510 43774 32562
rect 47058 32510 47070 32562
rect 47122 32510 47134 32562
rect 53442 32510 53454 32562
rect 53506 32510 53518 32562
rect 36542 32498 36594 32510
rect 2494 32450 2546 32462
rect 2494 32386 2546 32398
rect 8990 32450 9042 32462
rect 8990 32386 9042 32398
rect 9998 32450 10050 32462
rect 9998 32386 10050 32398
rect 15598 32450 15650 32462
rect 15598 32386 15650 32398
rect 18622 32450 18674 32462
rect 23438 32450 23490 32462
rect 21970 32398 21982 32450
rect 22034 32398 22046 32450
rect 22418 32398 22430 32450
rect 22482 32398 22494 32450
rect 18622 32386 18674 32398
rect 23438 32386 23490 32398
rect 24222 32450 24274 32462
rect 24222 32386 24274 32398
rect 26014 32450 26066 32462
rect 30718 32450 30770 32462
rect 26898 32398 26910 32450
rect 26962 32398 26974 32450
rect 26014 32386 26066 32398
rect 30718 32386 30770 32398
rect 36430 32450 36482 32462
rect 43262 32450 43314 32462
rect 49198 32450 49250 32462
rect 38210 32398 38222 32450
rect 38274 32398 38286 32450
rect 40338 32398 40350 32450
rect 40402 32398 40414 32450
rect 44146 32398 44158 32450
rect 44210 32398 44222 32450
rect 46274 32398 46286 32450
rect 46338 32398 46350 32450
rect 36430 32386 36482 32398
rect 43262 32386 43314 32398
rect 49198 32386 49250 32398
rect 8878 32338 8930 32350
rect 14814 32338 14866 32350
rect 12002 32286 12014 32338
rect 12066 32286 12078 32338
rect 55346 32286 55358 32338
rect 55410 32286 55422 32338
rect 8878 32274 8930 32286
rect 14814 32274 14866 32286
rect 1344 32170 58576 32204
rect 1344 32118 4478 32170
rect 4530 32118 4582 32170
rect 4634 32118 4686 32170
rect 4738 32118 35198 32170
rect 35250 32118 35302 32170
rect 35354 32118 35406 32170
rect 35458 32118 58576 32170
rect 1344 32084 58576 32118
rect 14030 32002 14082 32014
rect 14030 31938 14082 31950
rect 16270 32002 16322 32014
rect 16270 31938 16322 31950
rect 21646 32002 21698 32014
rect 21646 31938 21698 31950
rect 21982 32002 22034 32014
rect 24434 31950 24446 32002
rect 24498 31999 24510 32002
rect 24770 31999 24782 32002
rect 24498 31953 24782 31999
rect 24498 31950 24510 31953
rect 24770 31950 24782 31953
rect 24834 31950 24846 32002
rect 36978 31950 36990 32002
rect 37042 31950 37054 32002
rect 21982 31938 22034 31950
rect 1934 31890 1986 31902
rect 1934 31826 1986 31838
rect 4846 31890 4898 31902
rect 14702 31890 14754 31902
rect 23102 31890 23154 31902
rect 8642 31838 8654 31890
rect 8706 31838 8718 31890
rect 10770 31838 10782 31890
rect 10834 31838 10846 31890
rect 11666 31838 11678 31890
rect 11730 31838 11742 31890
rect 16706 31838 16718 31890
rect 16770 31838 16782 31890
rect 18834 31838 18846 31890
rect 18898 31838 18910 31890
rect 4846 31826 4898 31838
rect 14702 31826 14754 31838
rect 23102 31826 23154 31838
rect 24894 31890 24946 31902
rect 37326 31890 37378 31902
rect 25666 31838 25678 31890
rect 25730 31838 25742 31890
rect 24894 31826 24946 31838
rect 37326 31826 37378 31838
rect 39006 31890 39058 31902
rect 45502 31890 45554 31902
rect 55022 31890 55074 31902
rect 44034 31838 44046 31890
rect 44098 31838 44110 31890
rect 50530 31838 50542 31890
rect 50594 31838 50606 31890
rect 39006 31826 39058 31838
rect 45502 31826 45554 31838
rect 55022 31826 55074 31838
rect 57934 31890 57986 31902
rect 57934 31826 57986 31838
rect 12126 31778 12178 31790
rect 4162 31726 4174 31778
rect 4226 31726 4238 31778
rect 7970 31726 7982 31778
rect 8034 31726 8046 31778
rect 11330 31726 11342 31778
rect 11394 31726 11406 31778
rect 12126 31714 12178 31726
rect 14478 31778 14530 31790
rect 14478 31714 14530 31726
rect 15374 31778 15426 31790
rect 15374 31714 15426 31726
rect 15598 31778 15650 31790
rect 15598 31714 15650 31726
rect 15822 31778 15874 31790
rect 27134 31778 27186 31790
rect 19618 31726 19630 31778
rect 19682 31726 19694 31778
rect 15822 31714 15874 31726
rect 27134 31714 27186 31726
rect 29374 31778 29426 31790
rect 35310 31778 35362 31790
rect 34962 31726 34974 31778
rect 35026 31726 35038 31778
rect 29374 31714 29426 31726
rect 35310 31714 35362 31726
rect 37550 31778 37602 31790
rect 39678 31778 39730 31790
rect 39442 31726 39454 31778
rect 39506 31726 39518 31778
rect 37550 31714 37602 31726
rect 39678 31714 39730 31726
rect 40014 31778 40066 31790
rect 45614 31778 45666 31790
rect 41122 31726 41134 31778
rect 41186 31726 41198 31778
rect 46498 31726 46510 31778
rect 46562 31726 46574 31778
rect 47618 31726 47630 31778
rect 47682 31726 47694 31778
rect 52658 31726 52670 31778
rect 52722 31726 52734 31778
rect 55570 31726 55582 31778
rect 55634 31726 55646 31778
rect 40014 31714 40066 31726
rect 45614 31714 45666 31726
rect 14142 31666 14194 31678
rect 25230 31666 25282 31678
rect 22642 31614 22654 31666
rect 22706 31614 22718 31666
rect 14142 31602 14194 31614
rect 25230 31602 25282 31614
rect 26350 31666 26402 31678
rect 26350 31602 26402 31614
rect 26910 31666 26962 31678
rect 26910 31602 26962 31614
rect 28590 31666 28642 31678
rect 39902 31666 39954 31678
rect 29922 31614 29934 31666
rect 29986 31614 29998 31666
rect 41906 31614 41918 31666
rect 41970 31614 41982 31666
rect 48402 31614 48414 31666
rect 48466 31614 48478 31666
rect 28590 31602 28642 31614
rect 39902 31602 39954 31614
rect 12686 31554 12738 31566
rect 12686 31490 12738 31502
rect 13694 31554 13746 31566
rect 13694 31490 13746 31502
rect 14030 31554 14082 31566
rect 21758 31554 21810 31566
rect 15026 31502 15038 31554
rect 15090 31502 15102 31554
rect 14030 31490 14082 31502
rect 21758 31490 21810 31502
rect 22318 31554 22370 31566
rect 22318 31490 22370 31502
rect 23550 31554 23602 31566
rect 23550 31490 23602 31502
rect 23998 31554 24050 31566
rect 23998 31490 24050 31502
rect 24558 31554 24610 31566
rect 24558 31490 24610 31502
rect 25454 31554 25506 31566
rect 25454 31490 25506 31502
rect 25678 31554 25730 31566
rect 25678 31490 25730 31502
rect 25790 31554 25842 31566
rect 25790 31490 25842 31502
rect 26238 31554 26290 31566
rect 26238 31490 26290 31502
rect 26798 31554 26850 31566
rect 26798 31490 26850 31502
rect 27470 31554 27522 31566
rect 27470 31490 27522 31502
rect 27694 31554 27746 31566
rect 27694 31490 27746 31502
rect 27806 31554 27858 31566
rect 27806 31490 27858 31502
rect 28142 31554 28194 31566
rect 28142 31490 28194 31502
rect 35422 31554 35474 31566
rect 35422 31490 35474 31502
rect 35534 31554 35586 31566
rect 35534 31490 35586 31502
rect 35758 31554 35810 31566
rect 35758 31490 35810 31502
rect 36318 31554 36370 31566
rect 36318 31490 36370 31502
rect 38894 31554 38946 31566
rect 38894 31490 38946 31502
rect 39118 31554 39170 31566
rect 39118 31490 39170 31502
rect 45166 31554 45218 31566
rect 45166 31490 45218 31502
rect 45390 31554 45442 31566
rect 45390 31490 45442 31502
rect 45838 31554 45890 31566
rect 46958 31554 47010 31566
rect 46274 31502 46286 31554
rect 46338 31502 46350 31554
rect 47282 31502 47294 31554
rect 47346 31502 47358 31554
rect 45838 31490 45890 31502
rect 46958 31490 47010 31502
rect 1344 31386 58576 31420
rect 1344 31334 19838 31386
rect 19890 31334 19942 31386
rect 19994 31334 20046 31386
rect 20098 31334 50558 31386
rect 50610 31334 50662 31386
rect 50714 31334 50766 31386
rect 50818 31334 58576 31386
rect 1344 31300 58576 31334
rect 2046 31218 2098 31230
rect 31502 31218 31554 31230
rect 16034 31166 16046 31218
rect 16098 31166 16110 31218
rect 2046 31154 2098 31166
rect 31502 31154 31554 31166
rect 32174 31218 32226 31230
rect 32174 31154 32226 31166
rect 38222 31218 38274 31230
rect 41246 31218 41298 31230
rect 38994 31166 39006 31218
rect 39058 31166 39070 31218
rect 38222 31154 38274 31166
rect 41246 31154 41298 31166
rect 42142 31218 42194 31230
rect 42142 31154 42194 31166
rect 42254 31218 42306 31230
rect 42254 31154 42306 31166
rect 42702 31218 42754 31230
rect 42702 31154 42754 31166
rect 45726 31218 45778 31230
rect 46162 31166 46174 31218
rect 46226 31166 46238 31218
rect 45726 31154 45778 31166
rect 2718 31106 2770 31118
rect 16606 31106 16658 31118
rect 14914 31054 14926 31106
rect 14978 31054 14990 31106
rect 2718 31042 2770 31054
rect 16606 31042 16658 31054
rect 17502 31106 17554 31118
rect 17502 31042 17554 31054
rect 17614 31106 17666 31118
rect 30830 31106 30882 31118
rect 20850 31054 20862 31106
rect 20914 31054 20926 31106
rect 23538 31054 23550 31106
rect 23602 31054 23614 31106
rect 24098 31054 24110 31106
rect 24162 31054 24174 31106
rect 17614 31042 17666 31054
rect 30830 31042 30882 31054
rect 30942 31106 30994 31118
rect 36318 31106 36370 31118
rect 31826 31054 31838 31106
rect 31890 31054 31902 31106
rect 32498 31054 32510 31106
rect 32562 31054 32574 31106
rect 33842 31054 33854 31106
rect 33906 31054 33918 31106
rect 30942 31042 30994 31054
rect 36318 31042 36370 31054
rect 36430 31106 36482 31118
rect 50754 31054 50766 31106
rect 50818 31054 50830 31106
rect 36430 31042 36482 31054
rect 1710 30994 1762 31006
rect 1710 30930 1762 30942
rect 2382 30994 2434 31006
rect 16382 30994 16434 31006
rect 31166 30994 31218 31006
rect 38110 30994 38162 31006
rect 10098 30942 10110 30994
rect 10162 30942 10174 30994
rect 10546 30942 10558 30994
rect 10610 30942 10622 30994
rect 11218 30942 11230 30994
rect 11282 30942 11294 30994
rect 11890 30942 11902 30994
rect 11954 30942 11966 30994
rect 15586 30942 15598 30994
rect 15650 30942 15662 30994
rect 20066 30942 20078 30994
rect 20130 30942 20142 30994
rect 24434 30942 24446 30994
rect 24498 30942 24510 30994
rect 25218 30942 25230 30994
rect 25282 30942 25294 30994
rect 33058 30942 33070 30994
rect 33122 30942 33134 30994
rect 2382 30930 2434 30942
rect 16382 30930 16434 30942
rect 31166 30930 31218 30942
rect 38110 30930 38162 30942
rect 38334 30994 38386 31006
rect 39342 30994 39394 31006
rect 38658 30942 38670 30994
rect 38722 30942 38734 30994
rect 38334 30930 38386 30942
rect 39342 30930 39394 30942
rect 41358 30994 41410 31006
rect 41358 30930 41410 30942
rect 41582 30994 41634 31006
rect 41582 30930 41634 30942
rect 42030 30994 42082 31006
rect 42030 30930 42082 30942
rect 42590 30994 42642 31006
rect 42590 30930 42642 30942
rect 42814 30994 42866 31006
rect 45166 30994 45218 31006
rect 43138 30942 43150 30994
rect 43202 30942 43214 30994
rect 42814 30930 42866 30942
rect 45166 30930 45218 30942
rect 45614 30994 45666 31006
rect 45614 30930 45666 30942
rect 45838 30994 45890 31006
rect 45838 30930 45890 30942
rect 47406 30994 47458 31006
rect 47406 30930 47458 30942
rect 47854 30994 47906 31006
rect 47854 30930 47906 30942
rect 48078 30994 48130 31006
rect 49074 30942 49086 30994
rect 49138 30942 49150 30994
rect 48078 30930 48130 30942
rect 3166 30882 3218 30894
rect 23214 30882 23266 30894
rect 36990 30882 37042 30894
rect 10882 30830 10894 30882
rect 10946 30830 10958 30882
rect 12450 30830 12462 30882
rect 12514 30830 12526 30882
rect 12786 30830 12798 30882
rect 12850 30830 12862 30882
rect 22978 30830 22990 30882
rect 23042 30830 23054 30882
rect 27234 30830 27246 30882
rect 27298 30830 27310 30882
rect 35970 30830 35982 30882
rect 36034 30830 36046 30882
rect 3166 30818 3218 30830
rect 23214 30818 23266 30830
rect 36990 30818 37042 30830
rect 39566 30882 39618 30894
rect 39566 30818 39618 30830
rect 46510 30882 46562 30894
rect 46510 30818 46562 30830
rect 46734 30882 46786 30894
rect 46734 30818 46786 30830
rect 47182 30882 47234 30894
rect 47182 30818 47234 30830
rect 47966 30882 48018 30894
rect 47966 30818 48018 30830
rect 17502 30770 17554 30782
rect 10322 30718 10334 30770
rect 10386 30718 10398 30770
rect 17502 30706 17554 30718
rect 36430 30770 36482 30782
rect 36430 30706 36482 30718
rect 41246 30770 41298 30782
rect 41246 30706 41298 30718
rect 1344 30602 58576 30636
rect 1344 30550 4478 30602
rect 4530 30550 4582 30602
rect 4634 30550 4686 30602
rect 4738 30550 35198 30602
rect 35250 30550 35302 30602
rect 35354 30550 35406 30602
rect 35458 30550 58576 30602
rect 1344 30516 58576 30550
rect 46734 30434 46786 30446
rect 42690 30382 42702 30434
rect 42754 30382 42766 30434
rect 46734 30370 46786 30382
rect 2494 30322 2546 30334
rect 19406 30322 19458 30334
rect 10770 30270 10782 30322
rect 10834 30270 10846 30322
rect 16370 30270 16382 30322
rect 16434 30270 16446 30322
rect 2494 30258 2546 30270
rect 19406 30258 19458 30270
rect 23774 30322 23826 30334
rect 35198 30322 35250 30334
rect 25890 30270 25902 30322
rect 25954 30270 25966 30322
rect 29474 30270 29486 30322
rect 29538 30270 29550 30322
rect 29810 30270 29822 30322
rect 29874 30270 29886 30322
rect 31154 30270 31166 30322
rect 31218 30270 31230 30322
rect 23774 30258 23826 30270
rect 35198 30258 35250 30270
rect 35758 30322 35810 30334
rect 35758 30258 35810 30270
rect 38782 30322 38834 30334
rect 48862 30322 48914 30334
rect 42130 30270 42142 30322
rect 42194 30270 42206 30322
rect 47618 30270 47630 30322
rect 47682 30270 47694 30322
rect 38782 30258 38834 30270
rect 48862 30258 48914 30270
rect 49870 30322 49922 30334
rect 55346 30270 55358 30322
rect 55410 30270 55422 30322
rect 49870 30258 49922 30270
rect 11342 30210 11394 30222
rect 19742 30210 19794 30222
rect 7970 30158 7982 30210
rect 8034 30158 8046 30210
rect 13570 30158 13582 30210
rect 13634 30158 13646 30210
rect 11342 30146 11394 30158
rect 19742 30146 19794 30158
rect 20302 30210 20354 30222
rect 20302 30146 20354 30158
rect 21534 30210 21586 30222
rect 22318 30210 22370 30222
rect 21858 30158 21870 30210
rect 21922 30158 21934 30210
rect 21534 30146 21586 30158
rect 22318 30146 22370 30158
rect 22542 30210 22594 30222
rect 22542 30146 22594 30158
rect 22766 30210 22818 30222
rect 27470 30210 27522 30222
rect 26562 30158 26574 30210
rect 26626 30158 26638 30210
rect 22766 30146 22818 30158
rect 27470 30146 27522 30158
rect 27582 30210 27634 30222
rect 27582 30146 27634 30158
rect 28030 30210 28082 30222
rect 28030 30146 28082 30158
rect 28702 30210 28754 30222
rect 32958 30210 33010 30222
rect 34078 30210 34130 30222
rect 29138 30158 29150 30210
rect 29202 30158 29214 30210
rect 30258 30158 30270 30210
rect 30322 30158 30334 30210
rect 31266 30158 31278 30210
rect 31330 30158 31342 30210
rect 32050 30158 32062 30210
rect 32114 30158 32126 30210
rect 32498 30158 32510 30210
rect 32562 30158 32574 30210
rect 33394 30158 33406 30210
rect 33458 30158 33470 30210
rect 28702 30146 28754 30158
rect 32958 30146 33010 30158
rect 34078 30146 34130 30158
rect 37326 30210 37378 30222
rect 37326 30146 37378 30158
rect 37886 30210 37938 30222
rect 39230 30210 39282 30222
rect 43262 30210 43314 30222
rect 38322 30158 38334 30210
rect 38386 30158 38398 30210
rect 40562 30158 40574 30210
rect 40626 30158 40638 30210
rect 41458 30158 41470 30210
rect 41522 30158 41534 30210
rect 42242 30158 42254 30210
rect 42306 30158 42318 30210
rect 37886 30146 37938 30158
rect 39230 30146 39282 30158
rect 43262 30146 43314 30158
rect 44942 30210 44994 30222
rect 44942 30146 44994 30158
rect 45614 30210 45666 30222
rect 45614 30146 45666 30158
rect 45950 30210 46002 30222
rect 45950 30146 46002 30158
rect 46846 30210 46898 30222
rect 48750 30210 48802 30222
rect 47842 30158 47854 30210
rect 47906 30158 47918 30210
rect 46846 30146 46898 30158
rect 48750 30146 48802 30158
rect 49422 30210 49474 30222
rect 49422 30146 49474 30158
rect 49646 30210 49698 30222
rect 49646 30146 49698 30158
rect 50430 30210 50482 30222
rect 50430 30146 50482 30158
rect 53230 30210 53282 30222
rect 53442 30158 53454 30210
rect 53506 30158 53518 30210
rect 53230 30146 53282 30158
rect 1710 30098 1762 30110
rect 1710 30034 1762 30046
rect 2046 30098 2098 30110
rect 18398 30098 18450 30110
rect 8642 30046 8654 30098
rect 8706 30046 8718 30098
rect 14242 30046 14254 30098
rect 14306 30046 14318 30098
rect 2046 30034 2098 30046
rect 18398 30034 18450 30046
rect 22206 30098 22258 30110
rect 22206 30034 22258 30046
rect 23326 30098 23378 30110
rect 23326 30034 23378 30046
rect 27246 30098 27298 30110
rect 36990 30098 37042 30110
rect 31378 30046 31390 30098
rect 31442 30046 31454 30098
rect 33618 30046 33630 30098
rect 33682 30046 33694 30098
rect 27246 30034 27298 30046
rect 36990 30034 37042 30046
rect 39118 30098 39170 30110
rect 39118 30034 39170 30046
rect 39566 30098 39618 30110
rect 43374 30098 43426 30110
rect 41346 30046 41358 30098
rect 41410 30046 41422 30098
rect 39566 30034 39618 30046
rect 43374 30034 43426 30046
rect 45054 30098 45106 30110
rect 45054 30034 45106 30046
rect 45390 30098 45442 30110
rect 45390 30034 45442 30046
rect 46286 30098 46338 30110
rect 46286 30034 46338 30046
rect 46734 30098 46786 30110
rect 46734 30034 46786 30046
rect 48414 30098 48466 30110
rect 48414 30034 48466 30046
rect 50766 30098 50818 30110
rect 50766 30034 50818 30046
rect 2942 29986 2994 29998
rect 2942 29922 2994 29934
rect 11902 29986 11954 29998
rect 11902 29922 11954 29934
rect 12350 29986 12402 29998
rect 12350 29922 12402 29934
rect 18286 29986 18338 29998
rect 18286 29922 18338 29934
rect 20862 29986 20914 29998
rect 20862 29922 20914 29934
rect 21310 29986 21362 29998
rect 21310 29922 21362 29934
rect 21422 29986 21474 29998
rect 21422 29922 21474 29934
rect 27694 29986 27746 29998
rect 27694 29922 27746 29934
rect 28142 29986 28194 29998
rect 28142 29922 28194 29934
rect 28254 29986 28306 29998
rect 28254 29922 28306 29934
rect 37102 29986 37154 29998
rect 37102 29922 37154 29934
rect 39342 29986 39394 29998
rect 44382 29986 44434 29998
rect 40450 29934 40462 29986
rect 40514 29934 40526 29986
rect 39342 29922 39394 29934
rect 44382 29922 44434 29934
rect 45278 29986 45330 29998
rect 45278 29922 45330 29934
rect 45838 29986 45890 29998
rect 45838 29922 45890 29934
rect 48974 29986 49026 29998
rect 50654 29986 50706 29998
rect 50194 29934 50206 29986
rect 50258 29934 50270 29986
rect 48974 29922 49026 29934
rect 50654 29922 50706 29934
rect 1344 29818 58576 29852
rect 1344 29766 19838 29818
rect 19890 29766 19942 29818
rect 19994 29766 20046 29818
rect 20098 29766 50558 29818
rect 50610 29766 50662 29818
rect 50714 29766 50766 29818
rect 50818 29766 58576 29818
rect 1344 29732 58576 29766
rect 8878 29650 8930 29662
rect 8878 29586 8930 29598
rect 16046 29650 16098 29662
rect 16046 29586 16098 29598
rect 16270 29650 16322 29662
rect 25454 29650 25506 29662
rect 22642 29598 22654 29650
rect 22706 29647 22718 29650
rect 23090 29647 23102 29650
rect 22706 29601 23102 29647
rect 22706 29598 22718 29601
rect 23090 29598 23102 29601
rect 23154 29598 23166 29650
rect 16270 29586 16322 29598
rect 25454 29586 25506 29598
rect 25566 29650 25618 29662
rect 25566 29586 25618 29598
rect 31278 29650 31330 29662
rect 31278 29586 31330 29598
rect 32286 29650 32338 29662
rect 32286 29586 32338 29598
rect 33182 29650 33234 29662
rect 33182 29586 33234 29598
rect 33630 29650 33682 29662
rect 33630 29586 33682 29598
rect 38782 29650 38834 29662
rect 38782 29586 38834 29598
rect 39342 29650 39394 29662
rect 39342 29586 39394 29598
rect 40462 29650 40514 29662
rect 40462 29586 40514 29598
rect 46510 29650 46562 29662
rect 46510 29586 46562 29598
rect 46622 29650 46674 29662
rect 46622 29586 46674 29598
rect 46734 29650 46786 29662
rect 46734 29586 46786 29598
rect 47854 29650 47906 29662
rect 47854 29586 47906 29598
rect 2046 29538 2098 29550
rect 2046 29474 2098 29486
rect 12462 29538 12514 29550
rect 12462 29474 12514 29486
rect 15822 29538 15874 29550
rect 15822 29474 15874 29486
rect 16718 29538 16770 29550
rect 16718 29474 16770 29486
rect 24558 29538 24610 29550
rect 24558 29474 24610 29486
rect 29822 29538 29874 29550
rect 29822 29474 29874 29486
rect 31502 29538 31554 29550
rect 40238 29538 40290 29550
rect 47406 29538 47458 29550
rect 34402 29486 34414 29538
rect 34466 29486 34478 29538
rect 37538 29486 37550 29538
rect 37602 29486 37614 29538
rect 41122 29486 41134 29538
rect 41186 29486 41198 29538
rect 31502 29474 31554 29486
rect 40238 29474 40290 29486
rect 47406 29474 47458 29486
rect 1710 29426 1762 29438
rect 11454 29426 11506 29438
rect 12798 29426 12850 29438
rect 23550 29426 23602 29438
rect 10098 29374 10110 29426
rect 10162 29374 10174 29426
rect 10546 29374 10558 29426
rect 10610 29374 10622 29426
rect 11218 29374 11230 29426
rect 11282 29374 11294 29426
rect 12226 29374 12238 29426
rect 12290 29374 12302 29426
rect 13010 29374 13022 29426
rect 13074 29374 13086 29426
rect 14018 29374 14030 29426
rect 14082 29374 14094 29426
rect 15138 29374 15150 29426
rect 15202 29374 15214 29426
rect 22642 29374 22654 29426
rect 22706 29374 22718 29426
rect 1710 29362 1762 29374
rect 11454 29362 11506 29374
rect 12798 29362 12850 29374
rect 23550 29362 23602 29374
rect 24446 29426 24498 29438
rect 24446 29362 24498 29374
rect 24782 29426 24834 29438
rect 24782 29362 24834 29374
rect 25790 29426 25842 29438
rect 25790 29362 25842 29374
rect 25902 29426 25954 29438
rect 32174 29426 32226 29438
rect 36094 29426 36146 29438
rect 26674 29374 26686 29426
rect 26738 29374 26750 29426
rect 30034 29374 30046 29426
rect 30098 29374 30110 29426
rect 30482 29374 30494 29426
rect 30546 29374 30558 29426
rect 31826 29374 31838 29426
rect 31890 29374 31902 29426
rect 34962 29374 34974 29426
rect 35026 29374 35038 29426
rect 35746 29374 35758 29426
rect 35810 29374 35822 29426
rect 25902 29362 25954 29374
rect 32174 29362 32226 29374
rect 36094 29362 36146 29374
rect 37214 29426 37266 29438
rect 39118 29426 39170 29438
rect 38322 29374 38334 29426
rect 38386 29374 38398 29426
rect 38546 29374 38558 29426
rect 38610 29374 38622 29426
rect 37214 29362 37266 29374
rect 39118 29362 39170 29374
rect 39454 29426 39506 29438
rect 39454 29362 39506 29374
rect 40126 29426 40178 29438
rect 47182 29426 47234 29438
rect 46162 29374 46174 29426
rect 46226 29374 46238 29426
rect 47618 29374 47630 29426
rect 47682 29374 47694 29426
rect 40126 29362 40178 29374
rect 47182 29362 47234 29374
rect 2494 29314 2546 29326
rect 2494 29250 2546 29262
rect 8990 29314 9042 29326
rect 15934 29314 15986 29326
rect 23326 29314 23378 29326
rect 13682 29262 13694 29314
rect 13746 29262 13758 29314
rect 15474 29262 15486 29314
rect 15538 29262 15550 29314
rect 17602 29262 17614 29314
rect 17666 29262 17678 29314
rect 8990 29250 9042 29262
rect 15934 29250 15986 29262
rect 23326 29250 23378 29262
rect 24110 29314 24162 29326
rect 24110 29250 24162 29262
rect 25678 29314 25730 29326
rect 31390 29314 31442 29326
rect 27346 29262 27358 29314
rect 27410 29262 27422 29314
rect 29474 29262 29486 29314
rect 29538 29262 29550 29314
rect 25678 29250 25730 29262
rect 31390 29250 31442 29262
rect 34638 29314 34690 29326
rect 34638 29250 34690 29262
rect 36654 29314 36706 29326
rect 36654 29250 36706 29262
rect 38110 29314 38162 29326
rect 48862 29314 48914 29326
rect 38658 29262 38670 29314
rect 38722 29262 38734 29314
rect 38110 29250 38162 29262
rect 48862 29250 48914 29262
rect 16606 29202 16658 29214
rect 10322 29150 10334 29202
rect 10386 29150 10398 29202
rect 13458 29150 13470 29202
rect 13522 29150 13534 29202
rect 16606 29138 16658 29150
rect 32286 29202 32338 29214
rect 32286 29138 32338 29150
rect 47518 29202 47570 29214
rect 47518 29138 47570 29150
rect 1344 29034 58576 29068
rect 1344 28982 4478 29034
rect 4530 28982 4582 29034
rect 4634 28982 4686 29034
rect 4738 28982 35198 29034
rect 35250 28982 35302 29034
rect 35354 28982 35406 29034
rect 35458 28982 58576 29034
rect 1344 28948 58576 28982
rect 22542 28866 22594 28878
rect 22542 28802 22594 28814
rect 22878 28866 22930 28878
rect 28366 28866 28418 28878
rect 28018 28814 28030 28866
rect 28082 28814 28094 28866
rect 22878 28802 22930 28814
rect 28366 28802 28418 28814
rect 29262 28866 29314 28878
rect 33742 28866 33794 28878
rect 42702 28866 42754 28878
rect 31378 28814 31390 28866
rect 31442 28814 31454 28866
rect 39778 28814 39790 28866
rect 39842 28863 39854 28866
rect 40114 28863 40126 28866
rect 39842 28817 40126 28863
rect 39842 28814 39854 28817
rect 40114 28814 40126 28817
rect 40178 28814 40190 28866
rect 41346 28814 41358 28866
rect 41410 28814 41422 28866
rect 42354 28814 42366 28866
rect 42418 28814 42430 28866
rect 29262 28802 29314 28814
rect 33742 28802 33794 28814
rect 42702 28802 42754 28814
rect 45950 28866 46002 28878
rect 45950 28802 46002 28814
rect 57934 28866 57986 28878
rect 57934 28802 57986 28814
rect 21646 28754 21698 28766
rect 27134 28754 27186 28766
rect 17154 28702 17166 28754
rect 17218 28702 17230 28754
rect 18274 28702 18286 28754
rect 18338 28702 18350 28754
rect 20402 28702 20414 28754
rect 20466 28702 20478 28754
rect 24658 28702 24670 28754
rect 24722 28702 24734 28754
rect 26786 28702 26798 28754
rect 26850 28702 26862 28754
rect 21646 28690 21698 28702
rect 27134 28690 27186 28702
rect 28590 28754 28642 28766
rect 35646 28754 35698 28766
rect 31154 28702 31166 28754
rect 31218 28702 31230 28754
rect 28590 28690 28642 28702
rect 35646 28690 35698 28702
rect 37550 28754 37602 28766
rect 37550 28690 37602 28702
rect 38670 28754 38722 28766
rect 38670 28690 38722 28702
rect 40350 28754 40402 28766
rect 40350 28690 40402 28702
rect 42926 28754 42978 28766
rect 42926 28690 42978 28702
rect 47854 28754 47906 28766
rect 47854 28690 47906 28702
rect 55358 28754 55410 28766
rect 55358 28690 55410 28702
rect 1710 28642 1762 28654
rect 1710 28578 1762 28590
rect 2494 28642 2546 28654
rect 13470 28642 13522 28654
rect 21422 28642 21474 28654
rect 12786 28590 12798 28642
rect 12850 28590 12862 28642
rect 14242 28590 14254 28642
rect 14306 28590 14318 28642
rect 17490 28590 17502 28642
rect 17554 28590 17566 28642
rect 2494 28578 2546 28590
rect 13470 28578 13522 28590
rect 21422 28578 21474 28590
rect 21870 28642 21922 28654
rect 21870 28578 21922 28590
rect 21982 28642 22034 28654
rect 21982 28578 22034 28590
rect 22654 28642 22706 28654
rect 30606 28642 30658 28654
rect 35534 28642 35586 28654
rect 36094 28642 36146 28654
rect 23986 28590 23998 28642
rect 24050 28590 24062 28642
rect 31042 28590 31054 28642
rect 31106 28590 31118 28642
rect 34514 28590 34526 28642
rect 34578 28590 34590 28642
rect 34962 28590 34974 28642
rect 35026 28590 35038 28642
rect 35858 28590 35870 28642
rect 35922 28590 35934 28642
rect 22654 28578 22706 28590
rect 30606 28578 30658 28590
rect 35534 28578 35586 28590
rect 36094 28578 36146 28590
rect 36430 28642 36482 28654
rect 36430 28578 36482 28590
rect 36990 28642 37042 28654
rect 36990 28578 37042 28590
rect 39790 28642 39842 28654
rect 43486 28642 43538 28654
rect 40786 28590 40798 28642
rect 40850 28590 40862 28642
rect 41346 28590 41358 28642
rect 41410 28590 41422 28642
rect 41794 28590 41806 28642
rect 41858 28590 41870 28642
rect 39790 28578 39842 28590
rect 43486 28578 43538 28590
rect 43598 28642 43650 28654
rect 43598 28578 43650 28590
rect 44942 28642 44994 28654
rect 44942 28578 44994 28590
rect 45054 28642 45106 28654
rect 46958 28642 47010 28654
rect 45602 28590 45614 28642
rect 45666 28590 45678 28642
rect 46274 28590 46286 28642
rect 46338 28590 46350 28642
rect 45054 28578 45106 28590
rect 46958 28578 47010 28590
rect 47518 28642 47570 28654
rect 55570 28590 55582 28642
rect 55634 28590 55646 28642
rect 47518 28578 47570 28590
rect 13582 28530 13634 28542
rect 22990 28530 23042 28542
rect 8418 28478 8430 28530
rect 8482 28478 8494 28530
rect 15026 28478 15038 28530
rect 15090 28478 15102 28530
rect 13582 28466 13634 28478
rect 22990 28466 23042 28478
rect 23214 28530 23266 28542
rect 23214 28466 23266 28478
rect 23438 28530 23490 28542
rect 23438 28466 23490 28478
rect 29150 28530 29202 28542
rect 29150 28466 29202 28478
rect 29934 28530 29986 28542
rect 29934 28466 29986 28478
rect 32398 28530 32450 28542
rect 32398 28466 32450 28478
rect 32734 28530 32786 28542
rect 32734 28466 32786 28478
rect 32846 28530 32898 28542
rect 32846 28466 32898 28478
rect 33854 28530 33906 28542
rect 33854 28466 33906 28478
rect 35198 28530 35250 28542
rect 35198 28466 35250 28478
rect 36318 28530 36370 28542
rect 36318 28466 36370 28478
rect 37998 28530 38050 28542
rect 37998 28466 38050 28478
rect 39118 28530 39170 28542
rect 39118 28466 39170 28478
rect 44270 28530 44322 28542
rect 44270 28466 44322 28478
rect 45166 28530 45218 28542
rect 45166 28466 45218 28478
rect 47182 28530 47234 28542
rect 47182 28466 47234 28478
rect 2046 28418 2098 28430
rect 2046 28354 2098 28366
rect 22542 28418 22594 28430
rect 22542 28354 22594 28366
rect 27694 28418 27746 28430
rect 27694 28354 27746 28366
rect 29262 28418 29314 28430
rect 29262 28354 29314 28366
rect 30046 28418 30098 28430
rect 30046 28354 30098 28366
rect 30158 28418 30210 28430
rect 30158 28354 30210 28366
rect 32286 28418 32338 28430
rect 32286 28354 32338 28366
rect 33070 28418 33122 28430
rect 33070 28354 33122 28366
rect 33742 28418 33794 28430
rect 33742 28354 33794 28366
rect 38110 28418 38162 28430
rect 38110 28354 38162 28366
rect 38334 28418 38386 28430
rect 38334 28354 38386 28366
rect 44046 28418 44098 28430
rect 44046 28354 44098 28366
rect 44158 28418 44210 28430
rect 44158 28354 44210 28366
rect 46062 28418 46114 28430
rect 46062 28354 46114 28366
rect 47294 28418 47346 28430
rect 47294 28354 47346 28366
rect 1344 28250 58576 28284
rect 1344 28198 19838 28250
rect 19890 28198 19942 28250
rect 19994 28198 20046 28250
rect 20098 28198 50558 28250
rect 50610 28198 50662 28250
rect 50714 28198 50766 28250
rect 50818 28198 58576 28250
rect 1344 28164 58576 28198
rect 14366 28082 14418 28094
rect 14366 28018 14418 28030
rect 15710 28082 15762 28094
rect 15710 28018 15762 28030
rect 15822 28082 15874 28094
rect 15822 28018 15874 28030
rect 15934 28082 15986 28094
rect 15934 28018 15986 28030
rect 16718 28082 16770 28094
rect 16718 28018 16770 28030
rect 17502 28082 17554 28094
rect 17502 28018 17554 28030
rect 22542 28082 22594 28094
rect 22542 28018 22594 28030
rect 23326 28082 23378 28094
rect 23326 28018 23378 28030
rect 24670 28082 24722 28094
rect 24670 28018 24722 28030
rect 25342 28082 25394 28094
rect 25342 28018 25394 28030
rect 26798 28082 26850 28094
rect 26798 28018 26850 28030
rect 27918 28082 27970 28094
rect 27918 28018 27970 28030
rect 30270 28082 30322 28094
rect 32062 28082 32114 28094
rect 45726 28082 45778 28094
rect 30594 28030 30606 28082
rect 30658 28030 30670 28082
rect 31154 28030 31166 28082
rect 31218 28030 31230 28082
rect 40898 28030 40910 28082
rect 40962 28030 40974 28082
rect 30270 28018 30322 28030
rect 32062 28018 32114 28030
rect 45726 28018 45778 28030
rect 46510 28082 46562 28094
rect 46510 28018 46562 28030
rect 2046 27970 2098 27982
rect 2046 27906 2098 27918
rect 9998 27970 10050 27982
rect 16494 27970 16546 27982
rect 11778 27918 11790 27970
rect 11842 27918 11854 27970
rect 9998 27906 10050 27918
rect 16494 27906 16546 27918
rect 16830 27970 16882 27982
rect 16830 27906 16882 27918
rect 24110 27970 24162 27982
rect 24110 27906 24162 27918
rect 29374 27970 29426 27982
rect 29374 27906 29426 27918
rect 29710 27970 29762 27982
rect 29710 27906 29762 27918
rect 29822 27970 29874 27982
rect 29822 27906 29874 27918
rect 32286 27970 32338 27982
rect 32286 27906 32338 27918
rect 41694 27970 41746 27982
rect 50318 27970 50370 27982
rect 44482 27918 44494 27970
rect 44546 27918 44558 27970
rect 49522 27918 49534 27970
rect 49586 27918 49598 27970
rect 41694 27906 41746 27918
rect 50318 27906 50370 27918
rect 50430 27970 50482 27982
rect 50430 27906 50482 27918
rect 1710 27858 1762 27870
rect 16382 27858 16434 27870
rect 22318 27858 22370 27870
rect 11106 27806 11118 27858
rect 11170 27806 11182 27858
rect 19058 27806 19070 27858
rect 19122 27806 19134 27858
rect 1710 27794 1762 27806
rect 16382 27794 16434 27806
rect 22318 27794 22370 27806
rect 22990 27858 23042 27870
rect 24222 27858 24274 27870
rect 23538 27806 23550 27858
rect 23602 27806 23614 27858
rect 22990 27794 23042 27806
rect 24222 27794 24274 27806
rect 25230 27858 25282 27870
rect 25230 27794 25282 27806
rect 25566 27858 25618 27870
rect 29038 27858 29090 27870
rect 25890 27806 25902 27858
rect 25954 27806 25966 27858
rect 25566 27794 25618 27806
rect 29038 27794 29090 27806
rect 31502 27858 31554 27870
rect 31502 27794 31554 27806
rect 31726 27858 31778 27870
rect 41246 27858 41298 27870
rect 48078 27858 48130 27870
rect 50094 27858 50146 27870
rect 32498 27806 32510 27858
rect 32562 27806 32574 27858
rect 33058 27806 33070 27858
rect 33122 27806 33134 27858
rect 37426 27806 37438 27858
rect 37490 27806 37502 27858
rect 45266 27806 45278 27858
rect 45330 27806 45342 27858
rect 48738 27806 48750 27858
rect 48802 27806 48814 27858
rect 49298 27806 49310 27858
rect 49362 27806 49374 27858
rect 31726 27794 31778 27806
rect 41246 27794 41298 27806
rect 48078 27794 48130 27806
rect 50094 27794 50146 27806
rect 2494 27746 2546 27758
rect 18286 27746 18338 27758
rect 13906 27694 13918 27746
rect 13970 27694 13982 27746
rect 2494 27682 2546 27694
rect 18286 27682 18338 27694
rect 18846 27746 18898 27758
rect 22430 27746 22482 27758
rect 28478 27746 28530 27758
rect 19842 27694 19854 27746
rect 19906 27694 19918 27746
rect 21970 27694 21982 27746
rect 22034 27694 22046 27746
rect 26226 27694 26238 27746
rect 26290 27694 26302 27746
rect 18846 27682 18898 27694
rect 22430 27682 22482 27694
rect 28478 27682 28530 27694
rect 32398 27746 32450 27758
rect 47966 27746 48018 27758
rect 33842 27694 33854 27746
rect 33906 27694 33918 27746
rect 35970 27694 35982 27746
rect 36034 27694 36046 27746
rect 38210 27694 38222 27746
rect 38274 27694 38286 27746
rect 40338 27694 40350 27746
rect 40402 27694 40414 27746
rect 41570 27694 41582 27746
rect 41634 27694 41646 27746
rect 42354 27694 42366 27746
rect 42418 27694 42430 27746
rect 49634 27694 49646 27746
rect 49698 27694 49710 27746
rect 32398 27682 32450 27694
rect 47966 27682 48018 27694
rect 9886 27634 9938 27646
rect 23214 27634 23266 27646
rect 18498 27582 18510 27634
rect 18562 27631 18574 27634
rect 18834 27631 18846 27634
rect 18562 27585 18846 27631
rect 18562 27582 18574 27585
rect 18834 27582 18846 27585
rect 18898 27582 18910 27634
rect 9886 27570 9938 27582
rect 23214 27570 23266 27582
rect 24110 27634 24162 27646
rect 24110 27570 24162 27582
rect 29822 27634 29874 27646
rect 29822 27570 29874 27582
rect 41918 27634 41970 27646
rect 41918 27570 41970 27582
rect 1344 27466 58576 27500
rect 1344 27414 4478 27466
rect 4530 27414 4582 27466
rect 4634 27414 4686 27466
rect 4738 27414 35198 27466
rect 35250 27414 35302 27466
rect 35354 27414 35406 27466
rect 35458 27414 58576 27466
rect 1344 27380 58576 27414
rect 35198 27298 35250 27310
rect 14018 27246 14030 27298
rect 14082 27246 14094 27298
rect 18386 27246 18398 27298
rect 18450 27246 18462 27298
rect 22530 27246 22542 27298
rect 22594 27246 22606 27298
rect 35198 27234 35250 27246
rect 43038 27298 43090 27310
rect 43038 27234 43090 27246
rect 46846 27298 46898 27310
rect 46846 27234 46898 27246
rect 16606 27186 16658 27198
rect 20862 27186 20914 27198
rect 25902 27186 25954 27198
rect 9090 27134 9102 27186
rect 9154 27134 9166 27186
rect 11218 27134 11230 27186
rect 11282 27134 11294 27186
rect 14354 27134 14366 27186
rect 14418 27134 14430 27186
rect 18498 27134 18510 27186
rect 18562 27134 18574 27186
rect 22642 27134 22654 27186
rect 22706 27134 22718 27186
rect 24658 27134 24670 27186
rect 24722 27134 24734 27186
rect 16606 27122 16658 27134
rect 20862 27122 20914 27134
rect 25902 27122 25954 27134
rect 26350 27186 26402 27198
rect 26350 27122 26402 27134
rect 27134 27186 27186 27198
rect 32510 27186 32562 27198
rect 29922 27134 29934 27186
rect 29986 27134 29998 27186
rect 32050 27134 32062 27186
rect 32114 27134 32126 27186
rect 27134 27122 27186 27134
rect 32510 27122 32562 27134
rect 33966 27186 34018 27198
rect 41582 27186 41634 27198
rect 37986 27134 37998 27186
rect 38050 27134 38062 27186
rect 33966 27122 34018 27134
rect 41582 27122 41634 27134
rect 43934 27186 43986 27198
rect 47394 27134 47406 27186
rect 47458 27134 47470 27186
rect 48514 27134 48526 27186
rect 48578 27134 48590 27186
rect 43934 27122 43986 27134
rect 15486 27074 15538 27086
rect 21646 27074 21698 27086
rect 23326 27074 23378 27086
rect 8418 27022 8430 27074
rect 8482 27022 8494 27074
rect 13682 27022 13694 27074
rect 13746 27022 13758 27074
rect 14130 27022 14142 27074
rect 14194 27022 14206 27074
rect 14690 27022 14702 27074
rect 14754 27022 14766 27074
rect 15810 27022 15822 27074
rect 15874 27022 15886 27074
rect 17602 27022 17614 27074
rect 17666 27022 17678 27074
rect 18834 27022 18846 27074
rect 18898 27022 18910 27074
rect 19618 27022 19630 27074
rect 19682 27022 19694 27074
rect 22418 27022 22430 27074
rect 22482 27022 22494 27074
rect 15486 27010 15538 27022
rect 21646 27010 21698 27022
rect 23326 27010 23378 27022
rect 23998 27074 24050 27086
rect 23998 27010 24050 27022
rect 24222 27074 24274 27086
rect 24222 27010 24274 27022
rect 25118 27074 25170 27086
rect 25118 27010 25170 27022
rect 27470 27074 27522 27086
rect 27470 27010 27522 27022
rect 28030 27074 28082 27086
rect 33294 27074 33346 27086
rect 29250 27022 29262 27074
rect 29314 27022 29326 27074
rect 28030 27010 28082 27022
rect 33294 27010 33346 27022
rect 33406 27074 33458 27086
rect 33406 27010 33458 27022
rect 34078 27074 34130 27086
rect 34078 27010 34130 27022
rect 34414 27074 34466 27086
rect 34414 27010 34466 27022
rect 34526 27074 34578 27086
rect 34526 27010 34578 27022
rect 34862 27074 34914 27086
rect 38334 27074 38386 27086
rect 35746 27022 35758 27074
rect 35810 27022 35822 27074
rect 37762 27022 37774 27074
rect 37826 27022 37838 27074
rect 34862 27010 34914 27022
rect 38334 27010 38386 27022
rect 39006 27074 39058 27086
rect 40350 27074 40402 27086
rect 40002 27022 40014 27074
rect 40066 27022 40078 27074
rect 39006 27010 39058 27022
rect 40350 27010 40402 27022
rect 41806 27074 41858 27086
rect 41806 27010 41858 27022
rect 42142 27074 42194 27086
rect 43262 27074 43314 27086
rect 42466 27022 42478 27074
rect 42530 27022 42542 27074
rect 42690 27022 42702 27074
rect 42754 27022 42766 27074
rect 42142 27010 42194 27022
rect 43262 27010 43314 27022
rect 43598 27074 43650 27086
rect 43598 27010 43650 27022
rect 45390 27074 45442 27086
rect 45390 27010 45442 27022
rect 45726 27074 45778 27086
rect 45726 27010 45778 27022
rect 46062 27074 46114 27086
rect 46062 27010 46114 27022
rect 46174 27074 46226 27086
rect 46498 27022 46510 27074
rect 46562 27022 46574 27074
rect 47730 27022 47742 27074
rect 47794 27022 47806 27074
rect 51314 27022 51326 27074
rect 51378 27022 51390 27074
rect 46174 27010 46226 27022
rect 1710 26962 1762 26974
rect 1710 26898 1762 26910
rect 2382 26962 2434 26974
rect 2382 26898 2434 26910
rect 2718 26962 2770 26974
rect 2718 26898 2770 26910
rect 3166 26962 3218 26974
rect 3166 26898 3218 26910
rect 16942 26962 16994 26974
rect 16942 26898 16994 26910
rect 17054 26962 17106 26974
rect 20078 26962 20130 26974
rect 17378 26910 17390 26962
rect 17442 26910 17454 26962
rect 17054 26898 17106 26910
rect 20078 26898 20130 26910
rect 21310 26962 21362 26974
rect 21310 26898 21362 26910
rect 21534 26962 21586 26974
rect 21534 26898 21586 26910
rect 24558 26962 24610 26974
rect 33854 26962 33906 26974
rect 25442 26910 25454 26962
rect 25506 26910 25518 26962
rect 24558 26898 24610 26910
rect 33854 26898 33906 26910
rect 34750 26962 34802 26974
rect 34750 26898 34802 26910
rect 35310 26962 35362 26974
rect 35310 26898 35362 26910
rect 35534 26962 35586 26974
rect 35534 26898 35586 26910
rect 36318 26962 36370 26974
rect 36318 26898 36370 26910
rect 37326 26962 37378 26974
rect 37326 26898 37378 26910
rect 37550 26962 37602 26974
rect 37550 26898 37602 26910
rect 38446 26962 38498 26974
rect 38446 26898 38498 26910
rect 39454 26962 39506 26974
rect 39454 26898 39506 26910
rect 42926 26962 42978 26974
rect 42926 26898 42978 26910
rect 43374 26962 43426 26974
rect 43374 26898 43426 26910
rect 44830 26962 44882 26974
rect 44830 26898 44882 26910
rect 45838 26962 45890 26974
rect 45838 26898 45890 26910
rect 46734 26962 46786 26974
rect 46734 26898 46786 26910
rect 48190 26962 48242 26974
rect 50642 26910 50654 26962
rect 50706 26910 50718 26962
rect 48190 26898 48242 26910
rect 2046 26850 2098 26862
rect 2046 26786 2098 26798
rect 23774 26850 23826 26862
rect 23774 26786 23826 26798
rect 23886 26850 23938 26862
rect 23886 26786 23938 26798
rect 24782 26850 24834 26862
rect 24782 26786 24834 26798
rect 37998 26850 38050 26862
rect 37998 26786 38050 26798
rect 38558 26850 38610 26862
rect 38558 26786 38610 26798
rect 42030 26850 42082 26862
rect 42030 26786 42082 26798
rect 44942 26850 44994 26862
rect 44942 26786 44994 26798
rect 1344 26682 58576 26716
rect 1344 26630 19838 26682
rect 19890 26630 19942 26682
rect 19994 26630 20046 26682
rect 20098 26630 50558 26682
rect 50610 26630 50662 26682
rect 50714 26630 50766 26682
rect 50818 26630 58576 26682
rect 1344 26596 58576 26630
rect 2046 26514 2098 26526
rect 2046 26450 2098 26462
rect 2494 26514 2546 26526
rect 2494 26450 2546 26462
rect 25118 26514 25170 26526
rect 25118 26450 25170 26462
rect 25230 26514 25282 26526
rect 25230 26450 25282 26462
rect 26014 26514 26066 26526
rect 38334 26514 38386 26526
rect 28914 26462 28926 26514
rect 28978 26462 28990 26514
rect 26014 26450 26066 26462
rect 38334 26450 38386 26462
rect 38782 26514 38834 26526
rect 38782 26450 38834 26462
rect 46174 26514 46226 26526
rect 46174 26450 46226 26462
rect 46846 26514 46898 26526
rect 47742 26514 47794 26526
rect 47170 26462 47182 26514
rect 47234 26462 47246 26514
rect 46846 26450 46898 26462
rect 47742 26450 47794 26462
rect 48078 26514 48130 26526
rect 48078 26450 48130 26462
rect 48190 26514 48242 26526
rect 48190 26450 48242 26462
rect 49646 26514 49698 26526
rect 49646 26450 49698 26462
rect 49758 26514 49810 26526
rect 49758 26450 49810 26462
rect 50094 26514 50146 26526
rect 50094 26450 50146 26462
rect 20078 26402 20130 26414
rect 15586 26350 15598 26402
rect 15650 26350 15662 26402
rect 16818 26350 16830 26402
rect 16882 26350 16894 26402
rect 20078 26338 20130 26350
rect 23662 26402 23714 26414
rect 23662 26338 23714 26350
rect 23998 26402 24050 26414
rect 23998 26338 24050 26350
rect 24446 26402 24498 26414
rect 24446 26338 24498 26350
rect 24558 26402 24610 26414
rect 24558 26338 24610 26350
rect 25454 26402 25506 26414
rect 39006 26402 39058 26414
rect 26338 26350 26350 26402
rect 26402 26350 26414 26402
rect 25454 26338 25506 26350
rect 39006 26338 39058 26350
rect 47966 26402 48018 26414
rect 47966 26338 48018 26350
rect 1710 26290 1762 26302
rect 1710 26226 1762 26238
rect 11118 26290 11170 26302
rect 11118 26226 11170 26238
rect 11678 26290 11730 26302
rect 16494 26290 16546 26302
rect 19070 26290 19122 26302
rect 20414 26290 20466 26302
rect 23438 26290 23490 26302
rect 12002 26238 12014 26290
rect 12066 26238 12078 26290
rect 15362 26238 15374 26290
rect 15426 26238 15438 26290
rect 17602 26238 17614 26290
rect 17666 26238 17678 26290
rect 18050 26238 18062 26290
rect 18114 26238 18126 26290
rect 18834 26238 18846 26290
rect 18898 26238 18910 26290
rect 19506 26238 19518 26290
rect 19570 26238 19582 26290
rect 20626 26238 20638 26290
rect 20690 26238 20702 26290
rect 21634 26238 21646 26290
rect 21698 26238 21710 26290
rect 22530 26238 22542 26290
rect 22594 26238 22606 26290
rect 11678 26226 11730 26238
rect 16494 26226 16546 26238
rect 19070 26226 19122 26238
rect 20414 26226 20466 26238
rect 23438 26226 23490 26238
rect 24222 26290 24274 26302
rect 24222 26226 24274 26238
rect 25790 26290 25842 26302
rect 25790 26226 25842 26238
rect 28590 26290 28642 26302
rect 34750 26290 34802 26302
rect 36430 26290 36482 26302
rect 34290 26238 34302 26290
rect 34354 26238 34366 26290
rect 35186 26238 35198 26290
rect 35250 26238 35262 26290
rect 36082 26238 36094 26290
rect 36146 26238 36158 26290
rect 28590 26226 28642 26238
rect 34750 26226 34802 26238
rect 36430 26226 36482 26238
rect 37886 26290 37938 26302
rect 37886 26226 37938 26238
rect 38558 26290 38610 26302
rect 38558 26226 38610 26238
rect 39118 26290 39170 26302
rect 43934 26290 43986 26302
rect 48974 26290 49026 26302
rect 43138 26238 43150 26290
rect 43202 26238 43214 26290
rect 44370 26238 44382 26290
rect 44434 26238 44446 26290
rect 44930 26238 44942 26290
rect 44994 26238 45006 26290
rect 45266 26238 45278 26290
rect 45330 26238 45342 26290
rect 39118 26226 39170 26238
rect 43934 26226 43986 26238
rect 48974 26226 49026 26238
rect 49870 26290 49922 26302
rect 49870 26226 49922 26238
rect 2942 26178 2994 26190
rect 2942 26114 2994 26126
rect 8318 26178 8370 26190
rect 16158 26178 16210 26190
rect 23886 26178 23938 26190
rect 12786 26126 12798 26178
rect 12850 26126 12862 26178
rect 14914 26126 14926 26178
rect 14978 26126 14990 26178
rect 21522 26126 21534 26178
rect 21586 26126 21598 26178
rect 23090 26126 23102 26178
rect 23154 26126 23166 26178
rect 8318 26114 8370 26126
rect 16158 26114 16210 26126
rect 23886 26114 23938 26126
rect 26798 26178 26850 26190
rect 26798 26114 26850 26126
rect 27246 26178 27298 26190
rect 27246 26114 27298 26126
rect 27694 26178 27746 26190
rect 27694 26114 27746 26126
rect 28142 26178 28194 26190
rect 36878 26178 36930 26190
rect 33730 26126 33742 26178
rect 33794 26126 33806 26178
rect 28142 26114 28194 26126
rect 36878 26114 36930 26126
rect 37326 26178 37378 26190
rect 46622 26178 46674 26190
rect 42914 26126 42926 26178
rect 42978 26126 42990 26178
rect 37326 26114 37378 26126
rect 46622 26114 46674 26126
rect 48750 26178 48802 26190
rect 48750 26114 48802 26126
rect 8206 26066 8258 26078
rect 36766 26066 36818 26078
rect 17938 26014 17950 26066
rect 18002 26014 18014 26066
rect 20962 26014 20974 26066
rect 21026 26014 21038 26066
rect 35858 26014 35870 26066
rect 35922 26014 35934 26066
rect 8206 26002 8258 26014
rect 36766 26002 36818 26014
rect 37438 26066 37490 26078
rect 44818 26014 44830 26066
rect 44882 26014 44894 26066
rect 49298 26014 49310 26066
rect 49362 26014 49374 26066
rect 37438 26002 37490 26014
rect 1344 25898 58576 25932
rect 1344 25846 4478 25898
rect 4530 25846 4582 25898
rect 4634 25846 4686 25898
rect 4738 25846 35198 25898
rect 35250 25846 35302 25898
rect 35354 25846 35406 25898
rect 35458 25846 58576 25898
rect 1344 25812 58576 25846
rect 13470 25730 13522 25742
rect 11106 25678 11118 25730
rect 11170 25678 11182 25730
rect 13470 25666 13522 25678
rect 20638 25730 20690 25742
rect 33506 25678 33518 25730
rect 33570 25678 33582 25730
rect 20638 25666 20690 25678
rect 13582 25618 13634 25630
rect 19070 25618 19122 25630
rect 7186 25566 7198 25618
rect 7250 25566 7262 25618
rect 9314 25566 9326 25618
rect 9378 25566 9390 25618
rect 11330 25566 11342 25618
rect 11394 25566 11406 25618
rect 14690 25566 14702 25618
rect 14754 25566 14766 25618
rect 16258 25566 16270 25618
rect 16322 25566 16334 25618
rect 18386 25566 18398 25618
rect 18450 25566 18462 25618
rect 19730 25566 19742 25618
rect 19794 25566 19806 25618
rect 35186 25566 35198 25618
rect 35250 25566 35262 25618
rect 37762 25566 37774 25618
rect 37826 25566 37838 25618
rect 39890 25566 39902 25618
rect 39954 25566 39966 25618
rect 41234 25566 41246 25618
rect 41298 25566 41310 25618
rect 45602 25566 45614 25618
rect 45666 25566 45678 25618
rect 47730 25566 47742 25618
rect 47794 25566 47806 25618
rect 13582 25554 13634 25566
rect 19070 25554 19122 25566
rect 14254 25506 14306 25518
rect 6514 25454 6526 25506
rect 6578 25454 6590 25506
rect 10434 25454 10446 25506
rect 10498 25454 10510 25506
rect 11666 25454 11678 25506
rect 11730 25454 11742 25506
rect 12338 25454 12350 25506
rect 12402 25454 12414 25506
rect 14254 25442 14306 25454
rect 15150 25506 15202 25518
rect 27134 25506 27186 25518
rect 33406 25506 33458 25518
rect 15474 25454 15486 25506
rect 15538 25454 15550 25506
rect 19394 25454 19406 25506
rect 19458 25454 19470 25506
rect 26562 25454 26574 25506
rect 26626 25454 26638 25506
rect 28130 25454 28142 25506
rect 28194 25454 28206 25506
rect 31266 25454 31278 25506
rect 31330 25454 31342 25506
rect 32162 25454 32174 25506
rect 32226 25454 32238 25506
rect 33282 25454 33294 25506
rect 33346 25454 33358 25506
rect 15150 25442 15202 25454
rect 27134 25442 27186 25454
rect 33406 25442 33458 25454
rect 33742 25506 33794 25518
rect 40574 25506 40626 25518
rect 33954 25454 33966 25506
rect 34018 25454 34030 25506
rect 34850 25454 34862 25506
rect 34914 25454 34926 25506
rect 37090 25454 37102 25506
rect 37154 25454 37166 25506
rect 44146 25454 44158 25506
rect 44210 25454 44222 25506
rect 44818 25454 44830 25506
rect 44882 25454 44894 25506
rect 33742 25442 33794 25454
rect 40574 25442 40626 25454
rect 1710 25394 1762 25406
rect 1710 25330 1762 25342
rect 2046 25394 2098 25406
rect 12910 25394 12962 25406
rect 10210 25342 10222 25394
rect 10274 25342 10286 25394
rect 2046 25330 2098 25342
rect 12910 25330 12962 25342
rect 20750 25394 20802 25406
rect 40238 25394 40290 25406
rect 57598 25394 57650 25406
rect 21858 25342 21870 25394
rect 21922 25342 21934 25394
rect 27458 25342 27470 25394
rect 27522 25342 27534 25394
rect 28354 25342 28366 25394
rect 28418 25342 28430 25394
rect 31714 25342 31726 25394
rect 31778 25342 31790 25394
rect 43362 25342 43374 25394
rect 43426 25342 43438 25394
rect 20750 25330 20802 25342
rect 40238 25330 40290 25342
rect 57598 25330 57650 25342
rect 58158 25394 58210 25406
rect 58158 25330 58210 25342
rect 2494 25282 2546 25294
rect 20638 25282 20690 25294
rect 35870 25282 35922 25294
rect 13906 25230 13918 25282
rect 13970 25230 13982 25282
rect 31042 25230 31054 25282
rect 31106 25230 31118 25282
rect 2494 25218 2546 25230
rect 20638 25218 20690 25230
rect 35870 25218 35922 25230
rect 40350 25282 40402 25294
rect 40350 25218 40402 25230
rect 41022 25282 41074 25294
rect 41022 25218 41074 25230
rect 57822 25282 57874 25294
rect 57822 25218 57874 25230
rect 1344 25114 58576 25148
rect 1344 25062 19838 25114
rect 19890 25062 19942 25114
rect 19994 25062 20046 25114
rect 20098 25062 50558 25114
rect 50610 25062 50662 25114
rect 50714 25062 50766 25114
rect 50818 25062 58576 25114
rect 1344 25028 58576 25062
rect 10222 24946 10274 24958
rect 14926 24946 14978 24958
rect 14578 24894 14590 24946
rect 14642 24894 14654 24946
rect 10222 24882 10274 24894
rect 14926 24882 14978 24894
rect 15486 24946 15538 24958
rect 15486 24882 15538 24894
rect 18734 24946 18786 24958
rect 18734 24882 18786 24894
rect 19182 24946 19234 24958
rect 19182 24882 19234 24894
rect 19966 24946 20018 24958
rect 19966 24882 20018 24894
rect 23774 24946 23826 24958
rect 23774 24882 23826 24894
rect 24334 24946 24386 24958
rect 24334 24882 24386 24894
rect 24558 24946 24610 24958
rect 24558 24882 24610 24894
rect 34190 24946 34242 24958
rect 34190 24882 34242 24894
rect 48078 24946 48130 24958
rect 48078 24882 48130 24894
rect 57822 24946 57874 24958
rect 57822 24882 57874 24894
rect 2046 24834 2098 24846
rect 2046 24770 2098 24782
rect 11118 24834 11170 24846
rect 11118 24770 11170 24782
rect 14254 24834 14306 24846
rect 14254 24770 14306 24782
rect 18062 24834 18114 24846
rect 23886 24834 23938 24846
rect 22418 24782 22430 24834
rect 22482 24782 22494 24834
rect 18062 24770 18114 24782
rect 23886 24770 23938 24782
rect 24670 24834 24722 24846
rect 24670 24770 24722 24782
rect 25342 24834 25394 24846
rect 25342 24770 25394 24782
rect 25454 24834 25506 24846
rect 33406 24834 33458 24846
rect 25778 24782 25790 24834
rect 25842 24782 25854 24834
rect 26786 24782 26798 24834
rect 26850 24782 26862 24834
rect 25454 24770 25506 24782
rect 33406 24770 33458 24782
rect 33854 24834 33906 24846
rect 33854 24770 33906 24782
rect 33966 24834 34018 24846
rect 48190 24834 48242 24846
rect 50654 24834 50706 24846
rect 43586 24782 43598 24834
rect 43650 24782 43662 24834
rect 48738 24782 48750 24834
rect 48802 24782 48814 24834
rect 33966 24770 34018 24782
rect 48190 24770 48242 24782
rect 50654 24770 50706 24782
rect 1710 24722 1762 24734
rect 23550 24722 23602 24734
rect 5618 24670 5630 24722
rect 5682 24670 5694 24722
rect 11778 24670 11790 24722
rect 11842 24670 11854 24722
rect 12226 24670 12238 24722
rect 12290 24670 12302 24722
rect 13010 24670 13022 24722
rect 13074 24670 13086 24722
rect 14018 24670 14030 24722
rect 14082 24670 14094 24722
rect 23202 24670 23214 24722
rect 23266 24670 23278 24722
rect 1710 24658 1762 24670
rect 23550 24658 23602 24670
rect 23998 24722 24050 24734
rect 23998 24658 24050 24670
rect 25118 24722 25170 24734
rect 25118 24658 25170 24670
rect 26126 24722 26178 24734
rect 41582 24722 41634 24734
rect 47854 24722 47906 24734
rect 50542 24722 50594 24734
rect 26562 24670 26574 24722
rect 26626 24670 26638 24722
rect 30258 24670 30270 24722
rect 30322 24670 30334 24722
rect 31154 24670 31166 24722
rect 31218 24670 31230 24722
rect 32050 24670 32062 24722
rect 32114 24670 32126 24722
rect 36194 24670 36206 24722
rect 36258 24670 36270 24722
rect 41458 24670 41470 24722
rect 41522 24670 41534 24722
rect 42354 24670 42366 24722
rect 42418 24670 42430 24722
rect 43362 24670 43374 24722
rect 43426 24670 43438 24722
rect 44034 24670 44046 24722
rect 44098 24670 44110 24722
rect 49410 24670 49422 24722
rect 49474 24670 49486 24722
rect 49970 24670 49982 24722
rect 50034 24670 50046 24722
rect 26126 24658 26178 24670
rect 41582 24658 41634 24670
rect 47854 24658 47906 24670
rect 50542 24658 50594 24670
rect 58158 24722 58210 24734
rect 58158 24658 58210 24670
rect 2494 24610 2546 24622
rect 8766 24610 8818 24622
rect 6290 24558 6302 24610
rect 6354 24558 6366 24610
rect 8418 24558 8430 24610
rect 8482 24558 8494 24610
rect 2494 24546 2546 24558
rect 8766 24546 8818 24558
rect 8878 24610 8930 24622
rect 8878 24546 8930 24558
rect 9662 24610 9714 24622
rect 17726 24610 17778 24622
rect 12562 24558 12574 24610
rect 12626 24558 12638 24610
rect 9662 24546 9714 24558
rect 17726 24546 17778 24558
rect 19630 24610 19682 24622
rect 33294 24610 33346 24622
rect 20290 24558 20302 24610
rect 20354 24558 20366 24610
rect 27234 24558 27246 24610
rect 27298 24558 27310 24610
rect 29474 24558 29486 24610
rect 29538 24558 29550 24610
rect 31490 24558 31502 24610
rect 31554 24558 31566 24610
rect 32386 24558 32398 24610
rect 32450 24558 32462 24610
rect 19630 24546 19682 24558
rect 33294 24546 33346 24558
rect 34638 24610 34690 24622
rect 47294 24610 47346 24622
rect 37090 24558 37102 24610
rect 37154 24558 37166 24610
rect 42690 24558 42702 24610
rect 42754 24558 42766 24610
rect 44706 24558 44718 24610
rect 44770 24558 44782 24610
rect 46834 24558 46846 24610
rect 46898 24558 46910 24610
rect 34638 24546 34690 24558
rect 47294 24546 47346 24558
rect 48974 24610 49026 24622
rect 48974 24546 49026 24558
rect 57598 24610 57650 24622
rect 57598 24546 57650 24558
rect 11230 24498 11282 24510
rect 18174 24498 18226 24510
rect 50430 24498 50482 24510
rect 13346 24446 13358 24498
rect 13410 24446 13422 24498
rect 18498 24446 18510 24498
rect 18562 24495 18574 24498
rect 19282 24495 19294 24498
rect 18562 24449 19294 24495
rect 18562 24446 18574 24449
rect 19282 24446 19294 24449
rect 19346 24495 19358 24498
rect 19842 24495 19854 24498
rect 19346 24449 19854 24495
rect 19346 24446 19358 24449
rect 19842 24446 19854 24449
rect 19906 24446 19918 24498
rect 43026 24446 43038 24498
rect 43090 24446 43102 24498
rect 11230 24434 11282 24446
rect 18174 24434 18226 24446
rect 50430 24434 50482 24446
rect 1344 24330 58576 24364
rect 1344 24278 4478 24330
rect 4530 24278 4582 24330
rect 4634 24278 4686 24330
rect 4738 24278 35198 24330
rect 35250 24278 35302 24330
rect 35354 24278 35406 24330
rect 35458 24278 58576 24330
rect 1344 24244 58576 24278
rect 23550 24162 23602 24174
rect 8306 24110 8318 24162
rect 8370 24110 8382 24162
rect 23550 24098 23602 24110
rect 29262 24162 29314 24174
rect 29262 24098 29314 24110
rect 43486 24162 43538 24174
rect 43486 24098 43538 24110
rect 19854 24050 19906 24062
rect 9986 23998 9998 24050
rect 10050 23998 10062 24050
rect 12114 23998 12126 24050
rect 12178 23998 12190 24050
rect 19854 23986 19906 23998
rect 21534 24050 21586 24062
rect 21534 23986 21586 23998
rect 23214 24050 23266 24062
rect 23214 23986 23266 23998
rect 23662 24050 23714 24062
rect 28254 24050 28306 24062
rect 27682 23998 27694 24050
rect 27746 23998 27758 24050
rect 23662 23986 23714 23998
rect 28254 23986 28306 23998
rect 28590 24050 28642 24062
rect 36206 24050 36258 24062
rect 32722 23998 32734 24050
rect 32786 23998 32798 24050
rect 34850 23998 34862 24050
rect 34914 23998 34926 24050
rect 28590 23986 28642 23998
rect 36206 23986 36258 23998
rect 38782 24050 38834 24062
rect 43598 24050 43650 24062
rect 39106 23998 39118 24050
rect 39170 23998 39182 24050
rect 38782 23986 38834 23998
rect 43598 23986 43650 23998
rect 7198 23938 7250 23950
rect 7198 23874 7250 23886
rect 7646 23938 7698 23950
rect 7646 23874 7698 23886
rect 7758 23938 7810 23950
rect 7758 23874 7810 23886
rect 8094 23938 8146 23950
rect 35758 23938 35810 23950
rect 37998 23938 38050 23950
rect 43150 23938 43202 23950
rect 12898 23886 12910 23938
rect 12962 23886 12974 23938
rect 17266 23886 17278 23938
rect 17330 23886 17342 23938
rect 19282 23886 19294 23938
rect 19346 23886 19358 23938
rect 22642 23886 22654 23938
rect 22706 23886 22718 23938
rect 22978 23886 22990 23938
rect 23042 23886 23054 23938
rect 24882 23886 24894 23938
rect 24946 23886 24958 23938
rect 31938 23886 31950 23938
rect 32002 23886 32014 23938
rect 37426 23886 37438 23938
rect 37490 23886 37502 23938
rect 42018 23886 42030 23938
rect 42082 23886 42094 23938
rect 50082 23886 50094 23938
rect 50146 23886 50158 23938
rect 50642 23886 50654 23938
rect 50706 23886 50718 23938
rect 8094 23874 8146 23886
rect 35758 23874 35810 23886
rect 37998 23874 38050 23886
rect 43150 23874 43202 23886
rect 1710 23826 1762 23838
rect 1710 23762 1762 23774
rect 2046 23826 2098 23838
rect 2046 23762 2098 23774
rect 6974 23826 7026 23838
rect 6974 23762 7026 23774
rect 8318 23826 8370 23838
rect 20750 23826 20802 23838
rect 13682 23774 13694 23826
rect 13746 23774 13758 23826
rect 19058 23774 19070 23826
rect 19122 23774 19134 23826
rect 8318 23762 8370 23774
rect 20750 23762 20802 23774
rect 24334 23826 24386 23838
rect 24334 23762 24386 23774
rect 24446 23826 24498 23838
rect 29150 23826 29202 23838
rect 25554 23774 25566 23826
rect 25618 23774 25630 23826
rect 24446 23762 24498 23774
rect 29150 23762 29202 23774
rect 29598 23826 29650 23838
rect 29598 23762 29650 23774
rect 36990 23826 37042 23838
rect 43934 23826 43986 23838
rect 41234 23774 41246 23826
rect 41298 23774 41310 23826
rect 36990 23762 37042 23774
rect 43934 23762 43986 23774
rect 44046 23826 44098 23838
rect 58158 23826 58210 23838
rect 46946 23774 46958 23826
rect 47010 23774 47022 23826
rect 50418 23774 50430 23826
rect 50482 23774 50494 23826
rect 44046 23762 44098 23774
rect 58158 23762 58210 23774
rect 2494 23714 2546 23726
rect 2494 23650 2546 23662
rect 20302 23714 20354 23726
rect 20302 23650 20354 23662
rect 21870 23714 21922 23726
rect 21870 23650 21922 23662
rect 29934 23714 29986 23726
rect 29934 23650 29986 23662
rect 35198 23714 35250 23726
rect 35198 23650 35250 23662
rect 42590 23714 42642 23726
rect 42590 23650 42642 23662
rect 57598 23714 57650 23726
rect 57598 23650 57650 23662
rect 57822 23714 57874 23726
rect 57822 23650 57874 23662
rect 1344 23546 58576 23580
rect 1344 23494 19838 23546
rect 19890 23494 19942 23546
rect 19994 23494 20046 23546
rect 20098 23494 50558 23546
rect 50610 23494 50662 23546
rect 50714 23494 50766 23546
rect 50818 23494 58576 23546
rect 1344 23460 58576 23494
rect 14366 23378 14418 23390
rect 14366 23314 14418 23326
rect 15150 23378 15202 23390
rect 15150 23314 15202 23326
rect 22206 23378 22258 23390
rect 22206 23314 22258 23326
rect 39230 23378 39282 23390
rect 39230 23314 39282 23326
rect 40238 23378 40290 23390
rect 40238 23314 40290 23326
rect 49982 23378 50034 23390
rect 49982 23314 50034 23326
rect 50206 23378 50258 23390
rect 50206 23314 50258 23326
rect 2046 23266 2098 23278
rect 2046 23202 2098 23214
rect 13470 23266 13522 23278
rect 13470 23202 13522 23214
rect 13806 23266 13858 23278
rect 22654 23266 22706 23278
rect 18162 23214 18174 23266
rect 18226 23214 18238 23266
rect 20962 23214 20974 23266
rect 21026 23214 21038 23266
rect 13806 23202 13858 23214
rect 22654 23202 22706 23214
rect 27470 23266 27522 23278
rect 28366 23266 28418 23278
rect 47854 23266 47906 23278
rect 27794 23214 27806 23266
rect 27858 23214 27870 23266
rect 35634 23214 35646 23266
rect 35698 23214 35710 23266
rect 27470 23202 27522 23214
rect 28366 23202 28418 23214
rect 47854 23202 47906 23214
rect 47966 23266 48018 23278
rect 47966 23202 48018 23214
rect 50318 23266 50370 23278
rect 50318 23202 50370 23214
rect 1710 23154 1762 23166
rect 11230 23154 11282 23166
rect 20638 23154 20690 23166
rect 5394 23102 5406 23154
rect 5458 23102 5470 23154
rect 9762 23102 9774 23154
rect 9826 23102 9838 23154
rect 10322 23102 10334 23154
rect 10386 23102 10398 23154
rect 11106 23102 11118 23154
rect 11170 23102 11182 23154
rect 11778 23102 11790 23154
rect 11842 23102 11854 23154
rect 13010 23102 13022 23154
rect 13074 23102 13086 23154
rect 17490 23102 17502 23154
rect 17554 23102 17566 23154
rect 1710 23090 1762 23102
rect 11230 23090 11282 23102
rect 20638 23090 20690 23102
rect 23550 23154 23602 23166
rect 25342 23154 25394 23166
rect 24546 23102 24558 23154
rect 24610 23102 24622 23154
rect 23550 23090 23602 23102
rect 25342 23090 25394 23102
rect 25678 23154 25730 23166
rect 25678 23090 25730 23102
rect 26014 23154 26066 23166
rect 26014 23090 26066 23102
rect 26350 23154 26402 23166
rect 26350 23090 26402 23102
rect 27134 23154 27186 23166
rect 39790 23154 39842 23166
rect 31826 23102 31838 23154
rect 31890 23102 31902 23154
rect 34626 23102 34638 23154
rect 34690 23102 34702 23154
rect 27134 23090 27186 23102
rect 39790 23090 39842 23102
rect 40910 23154 40962 23166
rect 42590 23154 42642 23166
rect 41346 23102 41358 23154
rect 41410 23102 41422 23154
rect 42130 23102 42142 23154
rect 42194 23102 42206 23154
rect 40910 23090 40962 23102
rect 42590 23090 42642 23102
rect 42926 23154 42978 23166
rect 44606 23154 44658 23166
rect 43026 23102 43038 23154
rect 43090 23102 43102 23154
rect 44370 23102 44382 23154
rect 44434 23102 44446 23154
rect 42926 23090 42978 23102
rect 44606 23090 44658 23102
rect 44942 23154 44994 23166
rect 46846 23154 46898 23166
rect 45154 23102 45166 23154
rect 45218 23102 45230 23154
rect 45938 23102 45950 23154
rect 46002 23102 46014 23154
rect 46386 23102 46398 23154
rect 46450 23102 46462 23154
rect 44942 23090 44994 23102
rect 46846 23090 46898 23102
rect 47294 23154 47346 23166
rect 47294 23090 47346 23102
rect 47518 23154 47570 23166
rect 49646 23154 49698 23166
rect 49410 23102 49422 23154
rect 49474 23102 49486 23154
rect 47518 23090 47570 23102
rect 49646 23090 49698 23102
rect 2494 23042 2546 23054
rect 14702 23042 14754 23054
rect 6066 22990 6078 23042
rect 6130 22990 6142 23042
rect 8194 22990 8206 23042
rect 8258 22990 8270 23042
rect 12114 22990 12126 23042
rect 12178 22990 12190 23042
rect 12674 22990 12686 23042
rect 12738 22990 12750 23042
rect 2494 22978 2546 22990
rect 14702 22978 14754 22990
rect 16718 23042 16770 23054
rect 21422 23042 21474 23054
rect 20290 22990 20302 23042
rect 20354 22990 20366 23042
rect 16718 22978 16770 22990
rect 21422 22978 21474 22990
rect 23102 23042 23154 23054
rect 23102 22978 23154 22990
rect 24110 23042 24162 23054
rect 24110 22978 24162 22990
rect 26126 23042 26178 23054
rect 26126 22978 26178 22990
rect 26574 23042 26626 23054
rect 33182 23042 33234 23054
rect 28914 22990 28926 23042
rect 28978 22990 28990 23042
rect 31042 22990 31054 23042
rect 31106 22990 31118 23042
rect 26574 22978 26626 22990
rect 33182 22978 33234 22990
rect 47406 23042 47458 23054
rect 47406 22978 47458 22990
rect 48750 23042 48802 23054
rect 48750 22978 48802 22990
rect 14590 22930 14642 22942
rect 10098 22878 10110 22930
rect 10162 22878 10174 22930
rect 14590 22866 14642 22878
rect 16830 22930 16882 22942
rect 47966 22930 48018 22942
rect 22082 22878 22094 22930
rect 22146 22927 22158 22930
rect 23090 22927 23102 22930
rect 22146 22881 23102 22927
rect 22146 22878 22158 22881
rect 23090 22878 23102 22881
rect 23154 22878 23166 22930
rect 42802 22878 42814 22930
rect 42866 22878 42878 22930
rect 43922 22878 43934 22930
rect 43986 22878 43998 22930
rect 16830 22866 16882 22878
rect 47966 22866 48018 22878
rect 1344 22762 58576 22796
rect 1344 22710 4478 22762
rect 4530 22710 4582 22762
rect 4634 22710 4686 22762
rect 4738 22710 35198 22762
rect 35250 22710 35302 22762
rect 35354 22710 35406 22762
rect 35458 22710 58576 22762
rect 1344 22676 58576 22710
rect 6974 22594 7026 22606
rect 26910 22594 26962 22606
rect 7746 22542 7758 22594
rect 7810 22542 7822 22594
rect 20514 22542 20526 22594
rect 20578 22542 20590 22594
rect 30930 22542 30942 22594
rect 30994 22542 31006 22594
rect 6974 22530 7026 22542
rect 26910 22530 26962 22542
rect 7086 22482 7138 22494
rect 7086 22418 7138 22430
rect 10782 22482 10834 22494
rect 28142 22482 28194 22494
rect 43150 22482 43202 22494
rect 11778 22430 11790 22482
rect 11842 22430 11854 22482
rect 14354 22430 14366 22482
rect 14418 22430 14430 22482
rect 14802 22430 14814 22482
rect 14866 22430 14878 22482
rect 16930 22430 16942 22482
rect 16994 22430 17006 22482
rect 23314 22430 23326 22482
rect 23378 22430 23390 22482
rect 31154 22430 31166 22482
rect 31218 22430 31230 22482
rect 33506 22430 33518 22482
rect 33570 22430 33582 22482
rect 35634 22430 35646 22482
rect 35698 22430 35710 22482
rect 40450 22430 40462 22482
rect 40514 22430 40526 22482
rect 41234 22430 41246 22482
rect 41298 22430 41310 22482
rect 42130 22430 42142 22482
rect 42194 22430 42206 22482
rect 10782 22418 10834 22430
rect 28142 22418 28194 22430
rect 43150 22418 43202 22430
rect 43486 22482 43538 22494
rect 45266 22430 45278 22482
rect 45330 22430 45342 22482
rect 47842 22430 47854 22482
rect 47906 22430 47918 22482
rect 49970 22430 49982 22482
rect 50034 22430 50046 22482
rect 43486 22418 43538 22430
rect 8430 22370 8482 22382
rect 7970 22318 7982 22370
rect 8034 22318 8046 22370
rect 8430 22306 8482 22318
rect 8766 22370 8818 22382
rect 10446 22370 10498 22382
rect 19742 22370 19794 22382
rect 27694 22370 27746 22382
rect 9202 22318 9214 22370
rect 9266 22318 9278 22370
rect 10098 22318 10110 22370
rect 10162 22318 10174 22370
rect 11218 22318 11230 22370
rect 11282 22318 11294 22370
rect 17714 22318 17726 22370
rect 17778 22318 17790 22370
rect 18386 22318 18398 22370
rect 18450 22318 18462 22370
rect 18834 22318 18846 22370
rect 18898 22318 18910 22370
rect 19506 22318 19518 22370
rect 19570 22318 19582 22370
rect 20402 22318 20414 22370
rect 20466 22318 20478 22370
rect 25218 22318 25230 22370
rect 25282 22318 25294 22370
rect 8766 22306 8818 22318
rect 10446 22306 10498 22318
rect 19742 22306 19794 22318
rect 27694 22306 27746 22318
rect 30270 22370 30322 22382
rect 32286 22370 32338 22382
rect 40798 22370 40850 22382
rect 30706 22318 30718 22370
rect 30770 22318 30782 22370
rect 31714 22318 31726 22370
rect 31778 22318 31790 22370
rect 32386 22318 32398 22370
rect 32450 22318 32462 22370
rect 36306 22318 36318 22370
rect 36370 22318 36382 22370
rect 37538 22318 37550 22370
rect 37602 22318 37614 22370
rect 30270 22306 30322 22318
rect 32286 22306 32338 22318
rect 40798 22306 40850 22318
rect 41694 22370 41746 22382
rect 41694 22306 41746 22318
rect 43598 22370 43650 22382
rect 45502 22370 45554 22382
rect 44818 22318 44830 22370
rect 44882 22318 44894 22370
rect 43598 22306 43650 22318
rect 45502 22306 45554 22318
rect 46174 22370 46226 22382
rect 47058 22318 47070 22370
rect 47122 22318 47134 22370
rect 46174 22306 46226 22318
rect 1710 22258 1762 22270
rect 1710 22194 1762 22206
rect 2382 22258 2434 22270
rect 2382 22194 2434 22206
rect 13582 22258 13634 22270
rect 13582 22194 13634 22206
rect 20750 22258 20802 22270
rect 20750 22194 20802 22206
rect 27134 22258 27186 22270
rect 44158 22258 44210 22270
rect 38322 22206 38334 22258
rect 38386 22206 38398 22258
rect 27134 22194 27186 22206
rect 44158 22194 44210 22206
rect 45950 22258 46002 22270
rect 45950 22194 46002 22206
rect 57598 22258 57650 22270
rect 57598 22194 57650 22206
rect 58158 22258 58210 22270
rect 58158 22194 58210 22206
rect 2046 22146 2098 22158
rect 2046 22082 2098 22094
rect 2718 22146 2770 22158
rect 2718 22082 2770 22094
rect 3166 22146 3218 22158
rect 3166 22082 3218 22094
rect 12238 22146 12290 22158
rect 12238 22082 12290 22094
rect 13470 22146 13522 22158
rect 13470 22082 13522 22094
rect 13918 22146 13970 22158
rect 13918 22082 13970 22094
rect 27022 22146 27074 22158
rect 27022 22082 27074 22094
rect 28590 22146 28642 22158
rect 28590 22082 28642 22094
rect 42590 22146 42642 22158
rect 42590 22082 42642 22094
rect 44046 22146 44098 22158
rect 44046 22082 44098 22094
rect 45054 22146 45106 22158
rect 45054 22082 45106 22094
rect 45278 22146 45330 22158
rect 45278 22082 45330 22094
rect 45838 22146 45890 22158
rect 45838 22082 45890 22094
rect 46622 22146 46674 22158
rect 46622 22082 46674 22094
rect 57822 22146 57874 22158
rect 57822 22082 57874 22094
rect 1344 21978 58576 22012
rect 1344 21926 19838 21978
rect 19890 21926 19942 21978
rect 19994 21926 20046 21978
rect 20098 21926 50558 21978
rect 50610 21926 50662 21978
rect 50714 21926 50766 21978
rect 50818 21926 58576 21978
rect 1344 21892 58576 21926
rect 2494 21810 2546 21822
rect 2494 21746 2546 21758
rect 18174 21810 18226 21822
rect 18174 21746 18226 21758
rect 22878 21810 22930 21822
rect 22878 21746 22930 21758
rect 23102 21810 23154 21822
rect 23102 21746 23154 21758
rect 25342 21810 25394 21822
rect 25342 21746 25394 21758
rect 31054 21810 31106 21822
rect 31054 21746 31106 21758
rect 32510 21810 32562 21822
rect 32510 21746 32562 21758
rect 33070 21810 33122 21822
rect 33070 21746 33122 21758
rect 34526 21810 34578 21822
rect 34526 21746 34578 21758
rect 40126 21810 40178 21822
rect 40126 21746 40178 21758
rect 41022 21810 41074 21822
rect 41022 21746 41074 21758
rect 41470 21810 41522 21822
rect 41470 21746 41522 21758
rect 41918 21810 41970 21822
rect 47518 21810 47570 21822
rect 46498 21758 46510 21810
rect 46562 21758 46574 21810
rect 41918 21746 41970 21758
rect 47518 21746 47570 21758
rect 47854 21810 47906 21822
rect 47854 21746 47906 21758
rect 2046 21698 2098 21710
rect 2046 21634 2098 21646
rect 8990 21698 9042 21710
rect 24558 21698 24610 21710
rect 10994 21646 11006 21698
rect 11058 21646 11070 21698
rect 14242 21646 14254 21698
rect 14306 21646 14318 21698
rect 23762 21646 23774 21698
rect 23826 21646 23838 21698
rect 8990 21634 9042 21646
rect 24558 21634 24610 21646
rect 25454 21698 25506 21710
rect 25454 21634 25506 21646
rect 26350 21698 26402 21710
rect 26350 21634 26402 21646
rect 30494 21698 30546 21710
rect 30494 21634 30546 21646
rect 30942 21698 30994 21710
rect 35870 21698 35922 21710
rect 35522 21646 35534 21698
rect 35586 21646 35598 21698
rect 30942 21634 30994 21646
rect 35870 21634 35922 21646
rect 36430 21698 36482 21710
rect 39790 21698 39842 21710
rect 37090 21646 37102 21698
rect 37154 21646 37166 21698
rect 36430 21634 36482 21646
rect 39790 21634 39842 21646
rect 42254 21698 42306 21710
rect 47294 21698 47346 21710
rect 44034 21646 44046 21698
rect 44098 21646 44110 21698
rect 42254 21634 42306 21646
rect 47294 21634 47346 21646
rect 1710 21586 1762 21598
rect 1710 21522 1762 21534
rect 6302 21586 6354 21598
rect 7982 21586 8034 21598
rect 18510 21586 18562 21598
rect 23550 21586 23602 21598
rect 6514 21534 6526 21586
rect 6578 21534 6590 21586
rect 7858 21534 7870 21586
rect 7922 21534 7934 21586
rect 8754 21534 8766 21586
rect 8818 21534 8830 21586
rect 10210 21534 10222 21586
rect 10274 21534 10286 21586
rect 13458 21534 13470 21586
rect 13522 21534 13534 21586
rect 19506 21534 19518 21586
rect 19570 21534 19582 21586
rect 6302 21522 6354 21534
rect 7982 21522 8034 21534
rect 18510 21522 18562 21534
rect 23550 21522 23602 21534
rect 24110 21586 24162 21598
rect 24110 21522 24162 21534
rect 24334 21586 24386 21598
rect 24334 21522 24386 21534
rect 24670 21586 24722 21598
rect 24670 21522 24722 21534
rect 25118 21586 25170 21598
rect 26238 21586 26290 21598
rect 30606 21586 30658 21598
rect 26002 21534 26014 21586
rect 26066 21534 26078 21586
rect 27234 21534 27246 21586
rect 27298 21534 27310 21586
rect 25118 21522 25170 21534
rect 26238 21522 26290 21534
rect 30606 21522 30658 21534
rect 33966 21586 34018 21598
rect 33966 21522 34018 21534
rect 35198 21586 35250 21598
rect 46846 21586 46898 21598
rect 37538 21534 37550 21586
rect 37602 21534 37614 21586
rect 38546 21534 38558 21586
rect 38610 21534 38622 21586
rect 39554 21534 39566 21586
rect 39618 21534 39630 21586
rect 43362 21534 43374 21586
rect 43426 21534 43438 21586
rect 35198 21522 35250 21534
rect 46846 21522 46898 21534
rect 47182 21586 47234 21598
rect 47182 21522 47234 21534
rect 2942 21474 2994 21486
rect 2942 21410 2994 21422
rect 9662 21474 9714 21486
rect 16718 21474 16770 21486
rect 13122 21422 13134 21474
rect 13186 21422 13198 21474
rect 16370 21422 16382 21474
rect 16434 21422 16446 21474
rect 9662 21410 9714 21422
rect 16718 21410 16770 21422
rect 17614 21474 17666 21486
rect 22990 21474 23042 21486
rect 31502 21474 31554 21486
rect 18946 21422 18958 21474
rect 19010 21422 19022 21474
rect 20178 21422 20190 21474
rect 20242 21422 20254 21474
rect 22306 21422 22318 21474
rect 22370 21422 22382 21474
rect 27906 21422 27918 21474
rect 27970 21422 27982 21474
rect 30034 21422 30046 21474
rect 30098 21422 30110 21474
rect 17614 21410 17666 21422
rect 22990 21410 23042 21422
rect 31502 21410 31554 21422
rect 31950 21474 32002 21486
rect 40238 21474 40290 21486
rect 33506 21422 33518 21474
rect 33570 21422 33582 21474
rect 37986 21422 37998 21474
rect 38050 21422 38062 21474
rect 42690 21422 42702 21474
rect 42754 21422 42766 21474
rect 46162 21422 46174 21474
rect 46226 21422 46238 21474
rect 31950 21410 32002 21422
rect 40238 21410 40290 21422
rect 9550 21362 9602 21374
rect 8978 21310 8990 21362
rect 9042 21310 9054 21362
rect 9550 21298 9602 21310
rect 16830 21362 16882 21374
rect 30494 21362 30546 21374
rect 26786 21310 26798 21362
rect 26850 21310 26862 21362
rect 38658 21310 38670 21362
rect 38722 21310 38734 21362
rect 16830 21298 16882 21310
rect 30494 21298 30546 21310
rect 1344 21194 58576 21228
rect 1344 21142 4478 21194
rect 4530 21142 4582 21194
rect 4634 21142 4686 21194
rect 4738 21142 35198 21194
rect 35250 21142 35302 21194
rect 35354 21142 35406 21194
rect 35458 21142 58576 21194
rect 1344 21108 58576 21142
rect 20302 21026 20354 21038
rect 10098 20974 10110 21026
rect 10162 20974 10174 21026
rect 16594 20974 16606 21026
rect 16658 20974 16670 21026
rect 23426 20974 23438 21026
rect 23490 20974 23502 21026
rect 30258 20974 30270 21026
rect 30322 20974 30334 21026
rect 40226 20974 40238 21026
rect 40290 20974 40302 21026
rect 20302 20962 20354 20974
rect 20414 20914 20466 20926
rect 28142 20914 28194 20926
rect 44046 20914 44098 20926
rect 6850 20862 6862 20914
rect 6914 20862 6926 20914
rect 8978 20862 8990 20914
rect 9042 20862 9054 20914
rect 10322 20862 10334 20914
rect 10386 20862 10398 20914
rect 11890 20862 11902 20914
rect 11954 20862 11966 20914
rect 19954 20862 19966 20914
rect 20018 20862 20030 20914
rect 21298 20862 21310 20914
rect 21362 20862 21374 20914
rect 23090 20862 23102 20914
rect 23154 20862 23166 20914
rect 24322 20862 24334 20914
rect 24386 20862 24398 20914
rect 32050 20862 32062 20914
rect 32114 20862 32126 20914
rect 38434 20862 38446 20914
rect 38498 20862 38510 20914
rect 20414 20850 20466 20862
rect 28142 20850 28194 20862
rect 44046 20850 44098 20862
rect 45278 20914 45330 20926
rect 45278 20850 45330 20862
rect 48302 20914 48354 20926
rect 48302 20850 48354 20862
rect 12910 20802 12962 20814
rect 15710 20802 15762 20814
rect 6066 20750 6078 20802
rect 6130 20750 6142 20802
rect 9538 20750 9550 20802
rect 9602 20750 9614 20802
rect 10546 20750 10558 20802
rect 10610 20750 10622 20802
rect 11442 20750 11454 20802
rect 11506 20750 11518 20802
rect 14242 20750 14254 20802
rect 14306 20750 14318 20802
rect 15362 20750 15374 20802
rect 15426 20750 15438 20802
rect 12910 20738 12962 20750
rect 15710 20738 15762 20750
rect 16046 20802 16098 20814
rect 23998 20802 24050 20814
rect 28254 20802 28306 20814
rect 16146 20750 16158 20802
rect 16210 20750 16222 20802
rect 17154 20750 17166 20802
rect 17218 20750 17230 20802
rect 17826 20750 17838 20802
rect 17890 20750 17902 20802
rect 21522 20750 21534 20802
rect 21586 20750 21598 20802
rect 22418 20750 22430 20802
rect 22482 20750 22494 20802
rect 23762 20750 23774 20802
rect 23826 20750 23838 20802
rect 27234 20750 27246 20802
rect 27298 20750 27310 20802
rect 16046 20738 16098 20750
rect 23998 20738 24050 20750
rect 28254 20738 28306 20750
rect 28702 20802 28754 20814
rect 31054 20802 31106 20814
rect 36206 20802 36258 20814
rect 29586 20750 29598 20802
rect 29650 20750 29662 20802
rect 30146 20750 30158 20802
rect 30210 20750 30222 20802
rect 30818 20750 30830 20802
rect 30882 20750 30894 20802
rect 31490 20750 31502 20802
rect 31554 20750 31566 20802
rect 28702 20738 28754 20750
rect 31054 20738 31106 20750
rect 36206 20738 36258 20750
rect 37550 20802 37602 20814
rect 39566 20802 39618 20814
rect 41582 20802 41634 20814
rect 37986 20750 37998 20802
rect 38050 20750 38062 20802
rect 38994 20750 39006 20802
rect 39058 20750 39070 20802
rect 40002 20750 40014 20802
rect 40066 20750 40078 20802
rect 37550 20738 37602 20750
rect 39566 20738 39618 20750
rect 41582 20738 41634 20750
rect 42926 20802 42978 20814
rect 42926 20738 42978 20750
rect 47854 20802 47906 20814
rect 47854 20738 47906 20750
rect 1710 20690 1762 20702
rect 34302 20690 34354 20702
rect 9314 20638 9326 20690
rect 9378 20638 9390 20690
rect 14018 20638 14030 20690
rect 14082 20638 14094 20690
rect 26450 20638 26462 20690
rect 26514 20638 26526 20690
rect 1710 20626 1762 20638
rect 34302 20626 34354 20638
rect 34974 20690 35026 20702
rect 34974 20626 35026 20638
rect 41470 20690 41522 20702
rect 41470 20626 41522 20638
rect 41694 20690 41746 20702
rect 41694 20626 41746 20638
rect 42366 20690 42418 20702
rect 42366 20626 42418 20638
rect 42590 20690 42642 20702
rect 42590 20626 42642 20638
rect 47742 20690 47794 20702
rect 47742 20626 47794 20638
rect 2046 20578 2098 20590
rect 2046 20514 2098 20526
rect 2494 20578 2546 20590
rect 2494 20514 2546 20526
rect 12350 20578 12402 20590
rect 12350 20514 12402 20526
rect 13694 20578 13746 20590
rect 13694 20514 13746 20526
rect 27806 20578 27858 20590
rect 27806 20514 27858 20526
rect 28030 20578 28082 20590
rect 28030 20514 28082 20526
rect 34750 20578 34802 20590
rect 34750 20514 34802 20526
rect 34862 20578 34914 20590
rect 34862 20514 34914 20526
rect 35534 20578 35586 20590
rect 35534 20514 35586 20526
rect 35646 20578 35698 20590
rect 35646 20514 35698 20526
rect 35758 20578 35810 20590
rect 35758 20514 35810 20526
rect 37102 20578 37154 20590
rect 37102 20514 37154 20526
rect 40686 20578 40738 20590
rect 40686 20514 40738 20526
rect 42814 20578 42866 20590
rect 42814 20514 42866 20526
rect 43598 20578 43650 20590
rect 43598 20514 43650 20526
rect 45838 20578 45890 20590
rect 45838 20514 45890 20526
rect 46286 20578 46338 20590
rect 46286 20514 46338 20526
rect 46846 20578 46898 20590
rect 46846 20514 46898 20526
rect 47294 20578 47346 20590
rect 47294 20514 47346 20526
rect 47518 20578 47570 20590
rect 47518 20514 47570 20526
rect 1344 20410 58576 20444
rect 1344 20358 19838 20410
rect 19890 20358 19942 20410
rect 19994 20358 20046 20410
rect 20098 20358 50558 20410
rect 50610 20358 50662 20410
rect 50714 20358 50766 20410
rect 50818 20358 58576 20410
rect 1344 20324 58576 20358
rect 15150 20242 15202 20254
rect 15150 20178 15202 20190
rect 17950 20242 18002 20254
rect 17950 20178 18002 20190
rect 18510 20242 18562 20254
rect 18510 20178 18562 20190
rect 38670 20242 38722 20254
rect 42478 20242 42530 20254
rect 41234 20190 41246 20242
rect 41298 20190 41310 20242
rect 38670 20178 38722 20190
rect 42478 20178 42530 20190
rect 47406 20242 47458 20254
rect 47406 20178 47458 20190
rect 2046 20130 2098 20142
rect 2046 20066 2098 20078
rect 16046 20130 16098 20142
rect 25342 20130 25394 20142
rect 22530 20078 22542 20130
rect 22594 20078 22606 20130
rect 16046 20066 16098 20078
rect 25342 20066 25394 20078
rect 31390 20130 31442 20142
rect 33406 20130 33458 20142
rect 33058 20078 33070 20130
rect 33122 20078 33134 20130
rect 31390 20066 31442 20078
rect 33406 20066 33458 20078
rect 33966 20130 34018 20142
rect 33966 20066 34018 20078
rect 34190 20130 34242 20142
rect 39454 20130 39506 20142
rect 36082 20078 36094 20130
rect 36146 20078 36158 20130
rect 34190 20066 34242 20078
rect 39454 20066 39506 20078
rect 39678 20130 39730 20142
rect 45614 20130 45666 20142
rect 40002 20078 40014 20130
rect 40066 20078 40078 20130
rect 42914 20078 42926 20130
rect 42978 20078 42990 20130
rect 39678 20066 39730 20078
rect 45614 20066 45666 20078
rect 46846 20130 46898 20142
rect 46846 20066 46898 20078
rect 47742 20130 47794 20142
rect 47742 20066 47794 20078
rect 1710 20018 1762 20030
rect 18734 20018 18786 20030
rect 31166 20018 31218 20030
rect 6066 19966 6078 20018
rect 6130 19966 6142 20018
rect 14802 19966 14814 20018
rect 14866 19966 14878 20018
rect 19170 19966 19182 20018
rect 19234 19966 19246 20018
rect 19954 19966 19966 20018
rect 20018 19966 20030 20018
rect 20850 19966 20862 20018
rect 20914 19966 20926 20018
rect 21858 19966 21870 20018
rect 21922 19966 21934 20018
rect 25666 19966 25678 20018
rect 25730 19966 25742 20018
rect 1710 19954 1762 19966
rect 18734 19954 18786 19966
rect 31166 19954 31218 19966
rect 31502 20018 31554 20030
rect 31502 19954 31554 19966
rect 34414 20018 34466 20030
rect 34414 19954 34466 19966
rect 34862 20018 34914 20030
rect 41694 20018 41746 20030
rect 35410 19966 35422 20018
rect 35474 19966 35486 20018
rect 34862 19954 34914 19966
rect 41694 19954 41746 19966
rect 41806 20018 41858 20030
rect 47630 20018 47682 20030
rect 42018 19966 42030 20018
rect 42082 19966 42094 20018
rect 43362 19966 43374 20018
rect 43426 19966 43438 20018
rect 44482 19966 44494 20018
rect 44546 19966 44558 20018
rect 45154 19966 45166 20018
rect 45218 19966 45230 20018
rect 41806 19954 41858 19966
rect 47630 19954 47682 19966
rect 47854 20018 47906 20030
rect 47854 19954 47906 19966
rect 2494 19906 2546 19918
rect 15710 19906 15762 19918
rect 6850 19854 6862 19906
rect 6914 19854 6926 19906
rect 8978 19854 8990 19906
rect 9042 19854 9054 19906
rect 10210 19854 10222 19906
rect 10274 19854 10286 19906
rect 2494 19842 2546 19854
rect 15710 19842 15762 19854
rect 16606 19906 16658 19918
rect 16606 19842 16658 19854
rect 17502 19906 17554 19918
rect 31950 19906 32002 19918
rect 19618 19854 19630 19906
rect 19682 19854 19694 19906
rect 21298 19854 21310 19906
rect 21362 19854 21374 19906
rect 24658 19854 24670 19906
rect 24722 19854 24734 19906
rect 27682 19854 27694 19906
rect 27746 19854 27758 19906
rect 17502 19842 17554 19854
rect 31950 19842 32002 19854
rect 34302 19906 34354 19918
rect 46062 19906 46114 19918
rect 38210 19854 38222 19906
rect 38274 19854 38286 19906
rect 43810 19854 43822 19906
rect 43874 19854 43886 19906
rect 34302 19842 34354 19854
rect 46062 19842 46114 19854
rect 48862 19906 48914 19918
rect 48862 19842 48914 19854
rect 17390 19794 17442 19806
rect 46622 19794 46674 19806
rect 19282 19742 19294 19794
rect 19346 19742 19358 19794
rect 44034 19742 44046 19794
rect 44098 19742 44110 19794
rect 45826 19742 45838 19794
rect 45890 19791 45902 19794
rect 46386 19791 46398 19794
rect 45890 19745 46398 19791
rect 45890 19742 45902 19745
rect 46386 19742 46398 19745
rect 46450 19742 46462 19794
rect 17390 19730 17442 19742
rect 46622 19730 46674 19742
rect 46958 19794 47010 19806
rect 46958 19730 47010 19742
rect 1344 19626 58576 19660
rect 1344 19574 4478 19626
rect 4530 19574 4582 19626
rect 4634 19574 4686 19626
rect 4738 19574 35198 19626
rect 35250 19574 35302 19626
rect 35354 19574 35406 19626
rect 35458 19574 58576 19626
rect 1344 19540 58576 19574
rect 6862 19458 6914 19470
rect 22318 19458 22370 19470
rect 9762 19406 9774 19458
rect 9826 19406 9838 19458
rect 12786 19406 12798 19458
rect 12850 19406 12862 19458
rect 14690 19406 14702 19458
rect 14754 19406 14766 19458
rect 16818 19406 16830 19458
rect 16882 19406 16894 19458
rect 6862 19394 6914 19406
rect 22318 19394 22370 19406
rect 27246 19458 27298 19470
rect 37102 19458 37154 19470
rect 35298 19406 35310 19458
rect 35362 19406 35374 19458
rect 37426 19406 37438 19458
rect 37490 19455 37502 19458
rect 37874 19455 37886 19458
rect 37490 19409 37886 19455
rect 37490 19406 37502 19409
rect 37874 19406 37886 19409
rect 37938 19455 37950 19458
rect 38210 19455 38222 19458
rect 37938 19409 38222 19455
rect 37938 19406 37950 19409
rect 38210 19406 38222 19409
rect 38274 19406 38286 19458
rect 27246 19394 27298 19406
rect 37102 19394 37154 19406
rect 6750 19346 6802 19358
rect 19854 19346 19906 19358
rect 14578 19294 14590 19346
rect 14642 19294 14654 19346
rect 6750 19282 6802 19294
rect 19854 19282 19906 19294
rect 20414 19346 20466 19358
rect 20414 19282 20466 19294
rect 21310 19346 21362 19358
rect 21310 19282 21362 19294
rect 24782 19346 24834 19358
rect 37662 19346 37714 19358
rect 34962 19294 34974 19346
rect 35026 19294 35038 19346
rect 24782 19282 24834 19294
rect 37662 19282 37714 19294
rect 38110 19346 38162 19358
rect 42702 19346 42754 19358
rect 42242 19294 42254 19346
rect 42306 19294 42318 19346
rect 47954 19294 47966 19346
rect 48018 19294 48030 19346
rect 50082 19294 50094 19346
rect 50146 19294 50158 19346
rect 38110 19282 38162 19294
rect 42702 19282 42754 19294
rect 7198 19234 7250 19246
rect 8878 19234 8930 19246
rect 11902 19234 11954 19246
rect 17726 19234 17778 19246
rect 22766 19234 22818 19246
rect 25566 19234 25618 19246
rect 7410 19182 7422 19234
rect 7474 19182 7486 19234
rect 8754 19182 8766 19234
rect 8818 19182 8830 19234
rect 9650 19182 9662 19234
rect 9714 19182 9726 19234
rect 10434 19182 10446 19234
rect 10498 19182 10510 19234
rect 10994 19182 11006 19234
rect 11058 19182 11070 19234
rect 11442 19182 11454 19234
rect 11506 19182 11518 19234
rect 12338 19182 12350 19234
rect 12402 19182 12414 19234
rect 13906 19182 13918 19234
rect 13970 19182 13982 19234
rect 14354 19182 14366 19234
rect 14418 19182 14430 19234
rect 14914 19182 14926 19234
rect 14978 19182 14990 19234
rect 15810 19182 15822 19234
rect 15874 19182 15886 19234
rect 16930 19182 16942 19234
rect 16994 19182 17006 19234
rect 17826 19182 17838 19234
rect 17890 19182 17902 19234
rect 18610 19182 18622 19234
rect 18674 19182 18686 19234
rect 19058 19182 19070 19234
rect 19122 19182 19134 19234
rect 21746 19182 21758 19234
rect 21810 19182 21822 19234
rect 23314 19182 23326 19234
rect 23378 19182 23390 19234
rect 25106 19182 25118 19234
rect 25170 19182 25182 19234
rect 7198 19170 7250 19182
rect 8878 19170 8930 19182
rect 11902 19170 11954 19182
rect 17726 19170 17778 19182
rect 22766 19170 22818 19182
rect 25566 19170 25618 19182
rect 26014 19234 26066 19246
rect 26014 19170 26066 19182
rect 27470 19234 27522 19246
rect 27470 19170 27522 19182
rect 27694 19234 27746 19246
rect 27694 19170 27746 19182
rect 28142 19234 28194 19246
rect 28142 19170 28194 19182
rect 28254 19234 28306 19246
rect 28254 19170 28306 19182
rect 29262 19234 29314 19246
rect 29262 19170 29314 19182
rect 30270 19234 30322 19246
rect 30270 19170 30322 19182
rect 30942 19234 30994 19246
rect 30942 19170 30994 19182
rect 31166 19234 31218 19246
rect 31166 19170 31218 19182
rect 31502 19234 31554 19246
rect 35758 19234 35810 19246
rect 37214 19234 37266 19246
rect 42590 19234 42642 19246
rect 32162 19182 32174 19234
rect 32226 19182 32238 19234
rect 36082 19182 36094 19234
rect 36146 19182 36158 19234
rect 39330 19182 39342 19234
rect 39394 19182 39406 19234
rect 31502 19170 31554 19182
rect 35758 19170 35810 19182
rect 37214 19170 37266 19182
rect 42590 19170 42642 19182
rect 43710 19234 43762 19246
rect 43710 19170 43762 19182
rect 45502 19234 45554 19246
rect 45502 19170 45554 19182
rect 46398 19234 46450 19246
rect 47170 19182 47182 19234
rect 47234 19182 47246 19234
rect 46398 19170 46450 19182
rect 9886 19122 9938 19134
rect 9886 19058 9938 19070
rect 12910 19122 12962 19134
rect 12910 19058 12962 19070
rect 16382 19122 16434 19134
rect 16382 19058 16434 19070
rect 16718 19122 16770 19134
rect 16718 19058 16770 19070
rect 20750 19122 20802 19134
rect 20750 19058 20802 19070
rect 22430 19122 22482 19134
rect 22430 19058 22482 19070
rect 23550 19122 23602 19134
rect 23550 19058 23602 19070
rect 24110 19122 24162 19134
rect 24110 19058 24162 19070
rect 25454 19122 25506 19134
rect 29710 19122 29762 19134
rect 26898 19070 26910 19122
rect 26962 19070 26974 19122
rect 25454 19058 25506 19070
rect 29710 19058 29762 19070
rect 29934 19122 29986 19134
rect 35870 19122 35922 19134
rect 32834 19070 32846 19122
rect 32898 19070 32910 19122
rect 29934 19058 29986 19070
rect 35870 19058 35922 19070
rect 37102 19122 37154 19134
rect 37102 19058 37154 19070
rect 38558 19122 38610 19134
rect 42926 19122 42978 19134
rect 40114 19070 40126 19122
rect 40178 19070 40190 19122
rect 38558 19058 38610 19070
rect 42926 19058 42978 19070
rect 43150 19122 43202 19134
rect 43150 19058 43202 19070
rect 44942 19122 44994 19134
rect 44942 19058 44994 19070
rect 45054 19122 45106 19134
rect 45054 19058 45106 19070
rect 46174 19122 46226 19134
rect 46174 19058 46226 19070
rect 46286 19122 46338 19134
rect 46286 19058 46338 19070
rect 22318 19010 22370 19022
rect 22318 18946 22370 18958
rect 22878 19010 22930 19022
rect 22878 18946 22930 18958
rect 22990 19010 23042 19022
rect 22990 18946 23042 18958
rect 23662 19010 23714 19022
rect 23662 18946 23714 18958
rect 23886 19010 23938 19022
rect 23886 18946 23938 18958
rect 25678 19010 25730 19022
rect 25678 18946 25730 18958
rect 26126 19010 26178 19022
rect 26126 18946 26178 18958
rect 26238 19010 26290 19022
rect 26238 18946 26290 18958
rect 26462 19010 26514 19022
rect 26462 18946 26514 18958
rect 28030 19010 28082 19022
rect 28030 18946 28082 18958
rect 29598 19010 29650 19022
rect 29598 18946 29650 18958
rect 30382 19010 30434 19022
rect 30382 18946 30434 18958
rect 30494 19010 30546 19022
rect 30494 18946 30546 18958
rect 31390 19010 31442 19022
rect 31390 18946 31442 18958
rect 39006 19010 39058 19022
rect 39006 18946 39058 18958
rect 43486 19010 43538 19022
rect 43486 18946 43538 18958
rect 43598 19010 43650 19022
rect 43598 18946 43650 18958
rect 43934 19010 43986 19022
rect 43934 18946 43986 18958
rect 44718 19010 44770 19022
rect 46834 18958 46846 19010
rect 46898 18958 46910 19010
rect 44718 18946 44770 18958
rect 1344 18842 58576 18876
rect 1344 18790 19838 18842
rect 19890 18790 19942 18842
rect 19994 18790 20046 18842
rect 20098 18790 50558 18842
rect 50610 18790 50662 18842
rect 50714 18790 50766 18842
rect 50818 18790 58576 18842
rect 1344 18756 58576 18790
rect 11790 18674 11842 18686
rect 11790 18610 11842 18622
rect 22430 18674 22482 18686
rect 22430 18610 22482 18622
rect 24558 18674 24610 18686
rect 24558 18610 24610 18622
rect 33630 18674 33682 18686
rect 33630 18610 33682 18622
rect 40126 18674 40178 18686
rect 40126 18610 40178 18622
rect 40350 18674 40402 18686
rect 40350 18610 40402 18622
rect 47854 18674 47906 18686
rect 47854 18610 47906 18622
rect 2046 18562 2098 18574
rect 2046 18498 2098 18510
rect 24670 18562 24722 18574
rect 24670 18498 24722 18510
rect 34078 18562 34130 18574
rect 34078 18498 34130 18510
rect 36318 18562 36370 18574
rect 36318 18498 36370 18510
rect 37326 18562 37378 18574
rect 39902 18562 39954 18574
rect 39442 18510 39454 18562
rect 39506 18510 39518 18562
rect 37326 18498 37378 18510
rect 39902 18498 39954 18510
rect 40910 18562 40962 18574
rect 46846 18562 46898 18574
rect 45938 18510 45950 18562
rect 46002 18510 46014 18562
rect 40910 18498 40962 18510
rect 46846 18498 46898 18510
rect 1710 18450 1762 18462
rect 7982 18450 8034 18462
rect 10110 18450 10162 18462
rect 16046 18450 16098 18462
rect 6514 18398 6526 18450
rect 6578 18398 6590 18450
rect 6962 18398 6974 18450
rect 7026 18398 7038 18450
rect 7858 18398 7870 18450
rect 7922 18398 7934 18450
rect 8754 18398 8766 18450
rect 8818 18398 8830 18450
rect 12226 18398 12238 18450
rect 12290 18398 12302 18450
rect 1710 18386 1762 18398
rect 7982 18386 8034 18398
rect 10110 18386 10162 18398
rect 16046 18386 16098 18398
rect 16270 18450 16322 18462
rect 16270 18386 16322 18398
rect 16494 18450 16546 18462
rect 18958 18450 19010 18462
rect 20638 18450 20690 18462
rect 16706 18398 16718 18450
rect 16770 18398 16782 18450
rect 17714 18398 17726 18450
rect 17778 18398 17790 18450
rect 19170 18398 19182 18450
rect 19234 18398 19246 18450
rect 20178 18398 20190 18450
rect 20242 18398 20254 18450
rect 16494 18386 16546 18398
rect 18958 18386 19010 18398
rect 20638 18386 20690 18398
rect 20974 18450 21026 18462
rect 22206 18450 22258 18462
rect 21074 18398 21086 18450
rect 21138 18398 21150 18450
rect 20974 18386 21026 18398
rect 22206 18386 22258 18398
rect 22542 18450 22594 18462
rect 22542 18386 22594 18398
rect 22766 18450 22818 18462
rect 23998 18450 24050 18462
rect 23650 18398 23662 18450
rect 23714 18398 23726 18450
rect 22766 18386 22818 18398
rect 23998 18386 24050 18398
rect 24334 18450 24386 18462
rect 24334 18386 24386 18398
rect 25790 18450 25842 18462
rect 32286 18450 32338 18462
rect 29026 18398 29038 18450
rect 29090 18398 29102 18450
rect 29698 18398 29710 18450
rect 29762 18398 29774 18450
rect 25790 18386 25842 18398
rect 32286 18386 32338 18398
rect 33742 18450 33794 18462
rect 33742 18386 33794 18398
rect 33854 18450 33906 18462
rect 34862 18450 34914 18462
rect 34514 18398 34526 18450
rect 34578 18398 34590 18450
rect 33854 18386 33906 18398
rect 34862 18386 34914 18398
rect 35310 18450 35362 18462
rect 35310 18386 35362 18398
rect 35534 18450 35586 18462
rect 35534 18386 35586 18398
rect 35758 18450 35810 18462
rect 35758 18386 35810 18398
rect 35870 18450 35922 18462
rect 37102 18450 37154 18462
rect 36530 18398 36542 18450
rect 36594 18398 36606 18450
rect 36754 18398 36766 18450
rect 36818 18398 36830 18450
rect 35870 18386 35922 18398
rect 37102 18386 37154 18398
rect 37774 18450 37826 18462
rect 39118 18450 39170 18462
rect 38658 18398 38670 18450
rect 38722 18398 38734 18450
rect 37774 18386 37826 18398
rect 39118 18386 39170 18398
rect 40238 18450 40290 18462
rect 40238 18386 40290 18398
rect 41134 18450 41186 18462
rect 46286 18450 46338 18462
rect 41458 18398 41470 18450
rect 41522 18398 41534 18450
rect 42130 18398 42142 18450
rect 42194 18398 42206 18450
rect 42914 18398 42926 18450
rect 42978 18398 42990 18450
rect 45714 18398 45726 18450
rect 45778 18398 45790 18450
rect 41134 18386 41186 18398
rect 46286 18386 46338 18398
rect 46622 18450 46674 18462
rect 46622 18386 46674 18398
rect 47406 18450 47458 18462
rect 47406 18386 47458 18398
rect 47742 18450 47794 18462
rect 47742 18386 47794 18398
rect 48078 18450 48130 18462
rect 51650 18398 51662 18450
rect 51714 18398 51726 18450
rect 48078 18386 48130 18398
rect 2494 18338 2546 18350
rect 9550 18338 9602 18350
rect 8866 18286 8878 18338
rect 8930 18286 8942 18338
rect 2494 18274 2546 18286
rect 9550 18274 9602 18286
rect 10558 18338 10610 18350
rect 15374 18338 15426 18350
rect 18622 18338 18674 18350
rect 11330 18286 11342 18338
rect 11394 18286 11406 18338
rect 12898 18286 12910 18338
rect 12962 18286 12974 18338
rect 15026 18286 15038 18338
rect 15090 18286 15102 18338
rect 18050 18286 18062 18338
rect 18114 18286 18126 18338
rect 10558 18274 10610 18286
rect 15374 18274 15426 18286
rect 18622 18274 18674 18286
rect 24110 18338 24162 18350
rect 24110 18274 24162 18286
rect 25342 18338 25394 18350
rect 25342 18274 25394 18286
rect 28590 18338 28642 18350
rect 33406 18338 33458 18350
rect 31826 18286 31838 18338
rect 31890 18286 31902 18338
rect 28590 18274 28642 18286
rect 33406 18274 33458 18286
rect 35086 18338 35138 18350
rect 37214 18338 37266 18350
rect 41022 18338 41074 18350
rect 46734 18338 46786 18350
rect 36306 18286 36318 18338
rect 36370 18286 36382 18338
rect 38322 18286 38334 18338
rect 38386 18286 38398 18338
rect 45042 18286 45054 18338
rect 45106 18286 45118 18338
rect 48738 18286 48750 18338
rect 48802 18286 48814 18338
rect 50866 18286 50878 18338
rect 50930 18286 50942 18338
rect 35086 18274 35138 18286
rect 37214 18274 37266 18286
rect 41022 18274 41074 18286
rect 46734 18274 46786 18286
rect 10446 18226 10498 18238
rect 8194 18174 8206 18226
rect 8258 18174 8270 18226
rect 10446 18162 10498 18174
rect 15598 18226 15650 18238
rect 18510 18226 18562 18238
rect 16706 18174 16718 18226
rect 16770 18174 16782 18226
rect 19618 18174 19630 18226
rect 19682 18174 19694 18226
rect 15598 18162 15650 18174
rect 18510 18162 18562 18174
rect 1344 18058 58576 18092
rect 1344 18006 4478 18058
rect 4530 18006 4582 18058
rect 4634 18006 4686 18058
rect 4738 18006 35198 18058
rect 35250 18006 35302 18058
rect 35354 18006 35406 18058
rect 35458 18006 58576 18058
rect 1344 17972 58576 18006
rect 34078 17890 34130 17902
rect 14018 17838 14030 17890
rect 14082 17838 14094 17890
rect 17042 17838 17054 17890
rect 17106 17838 17118 17890
rect 28242 17838 28254 17890
rect 28306 17887 28318 17890
rect 28578 17887 28590 17890
rect 28306 17841 28590 17887
rect 28306 17838 28318 17841
rect 28578 17838 28590 17841
rect 28642 17838 28654 17890
rect 34078 17826 34130 17838
rect 40910 17890 40962 17902
rect 48974 17890 49026 17902
rect 41234 17838 41246 17890
rect 41298 17838 41310 17890
rect 40910 17826 40962 17838
rect 48974 17826 49026 17838
rect 11118 17778 11170 17790
rect 7858 17726 7870 17778
rect 7922 17726 7934 17778
rect 9986 17726 9998 17778
rect 10050 17726 10062 17778
rect 11118 17714 11170 17726
rect 12126 17778 12178 17790
rect 19630 17778 19682 17790
rect 16146 17726 16158 17778
rect 16210 17726 16222 17778
rect 17378 17726 17390 17778
rect 17442 17726 17454 17778
rect 12126 17714 12178 17726
rect 19630 17714 19682 17726
rect 20078 17778 20130 17790
rect 25342 17778 25394 17790
rect 22082 17726 22094 17778
rect 22146 17726 22158 17778
rect 24210 17726 24222 17778
rect 24274 17726 24286 17778
rect 20078 17714 20130 17726
rect 25342 17714 25394 17726
rect 28254 17778 28306 17790
rect 30830 17778 30882 17790
rect 33630 17778 33682 17790
rect 30034 17726 30046 17778
rect 30098 17726 30110 17778
rect 31602 17726 31614 17778
rect 31666 17726 31678 17778
rect 32386 17726 32398 17778
rect 32450 17726 32462 17778
rect 28254 17714 28306 17726
rect 30830 17714 30882 17726
rect 33630 17714 33682 17726
rect 34862 17778 34914 17790
rect 34862 17714 34914 17726
rect 35982 17778 36034 17790
rect 40686 17778 40738 17790
rect 37762 17726 37774 17778
rect 37826 17726 37838 17778
rect 39890 17726 39902 17778
rect 39954 17726 39966 17778
rect 35982 17714 36034 17726
rect 40686 17714 40738 17726
rect 43038 17778 43090 17790
rect 43038 17714 43090 17726
rect 43598 17778 43650 17790
rect 43598 17714 43650 17726
rect 43934 17778 43986 17790
rect 43934 17714 43986 17726
rect 46398 17778 46450 17790
rect 46398 17714 46450 17726
rect 49758 17778 49810 17790
rect 49758 17714 49810 17726
rect 50206 17778 50258 17790
rect 50206 17714 50258 17726
rect 12350 17666 12402 17678
rect 7074 17614 7086 17666
rect 7138 17614 7150 17666
rect 12350 17602 12402 17614
rect 12910 17666 12962 17678
rect 15150 17666 15202 17678
rect 16494 17666 16546 17678
rect 18510 17666 18562 17678
rect 31054 17666 31106 17678
rect 13682 17614 13694 17666
rect 13746 17614 13758 17666
rect 14242 17614 14254 17666
rect 14306 17614 14318 17666
rect 14802 17614 14814 17666
rect 14866 17614 14878 17666
rect 15586 17614 15598 17666
rect 15650 17614 15662 17666
rect 16930 17614 16942 17666
rect 16994 17614 17006 17666
rect 18050 17614 18062 17666
rect 18114 17614 18126 17666
rect 18946 17614 18958 17666
rect 19010 17614 19022 17666
rect 21410 17614 21422 17666
rect 21474 17614 21486 17666
rect 24770 17614 24782 17666
rect 24834 17614 24846 17666
rect 30258 17614 30270 17666
rect 30322 17614 30334 17666
rect 12910 17602 12962 17614
rect 15150 17602 15202 17614
rect 16494 17602 16546 17614
rect 18510 17602 18562 17614
rect 31054 17602 31106 17614
rect 33182 17666 33234 17678
rect 33182 17602 33234 17614
rect 33966 17666 34018 17678
rect 33966 17602 34018 17614
rect 34974 17666 35026 17678
rect 34974 17602 35026 17614
rect 35310 17666 35362 17678
rect 35310 17602 35362 17614
rect 35870 17666 35922 17678
rect 35870 17602 35922 17614
rect 36206 17666 36258 17678
rect 41470 17666 41522 17678
rect 37090 17614 37102 17666
rect 37154 17614 37166 17666
rect 36206 17602 36258 17614
rect 41470 17602 41522 17614
rect 41806 17666 41858 17678
rect 41806 17602 41858 17614
rect 44718 17666 44770 17678
rect 44718 17602 44770 17614
rect 47294 17666 47346 17678
rect 47294 17602 47346 17614
rect 48190 17666 48242 17678
rect 48190 17602 48242 17614
rect 48414 17666 48466 17678
rect 48414 17602 48466 17614
rect 48750 17666 48802 17678
rect 48750 17602 48802 17614
rect 1710 17554 1762 17566
rect 1710 17490 1762 17502
rect 2382 17554 2434 17566
rect 2382 17490 2434 17502
rect 2718 17554 2770 17566
rect 2718 17490 2770 17502
rect 19518 17554 19570 17566
rect 19518 17490 19570 17502
rect 31614 17554 31666 17566
rect 34078 17554 34130 17566
rect 32834 17502 32846 17554
rect 32898 17502 32910 17554
rect 31614 17490 31666 17502
rect 34078 17490 34130 17502
rect 34750 17554 34802 17566
rect 34750 17490 34802 17502
rect 36430 17554 36482 17566
rect 36430 17490 36482 17502
rect 45726 17554 45778 17566
rect 45726 17490 45778 17502
rect 45838 17554 45890 17566
rect 45838 17490 45890 17502
rect 47406 17554 47458 17566
rect 47406 17490 47458 17502
rect 2046 17442 2098 17454
rect 2046 17378 2098 17390
rect 3166 17442 3218 17454
rect 3166 17378 3218 17390
rect 11006 17442 11058 17454
rect 31390 17442 31442 17454
rect 24546 17390 24558 17442
rect 24610 17390 24622 17442
rect 11006 17378 11058 17390
rect 31390 17378 31442 17390
rect 31950 17442 32002 17454
rect 31950 17378 32002 17390
rect 40350 17442 40402 17454
rect 40350 17378 40402 17390
rect 41694 17442 41746 17454
rect 41694 17378 41746 17390
rect 42590 17442 42642 17454
rect 42590 17378 42642 17390
rect 45054 17442 45106 17454
rect 45054 17378 45106 17390
rect 45278 17442 45330 17454
rect 45278 17378 45330 17390
rect 45390 17442 45442 17454
rect 45390 17378 45442 17390
rect 45502 17442 45554 17454
rect 45502 17378 45554 17390
rect 46734 17442 46786 17454
rect 46734 17378 46786 17390
rect 47630 17442 47682 17454
rect 47630 17378 47682 17390
rect 47966 17442 48018 17454
rect 47966 17378 48018 17390
rect 48302 17442 48354 17454
rect 49298 17390 49310 17442
rect 49362 17390 49374 17442
rect 48302 17378 48354 17390
rect 1344 17274 58576 17308
rect 1344 17222 19838 17274
rect 19890 17222 19942 17274
rect 19994 17222 20046 17274
rect 20098 17222 50558 17274
rect 50610 17222 50662 17274
rect 50714 17222 50766 17274
rect 50818 17222 58576 17274
rect 1344 17188 58576 17222
rect 2494 17106 2546 17118
rect 2494 17042 2546 17054
rect 13358 17106 13410 17118
rect 13358 17042 13410 17054
rect 23214 17106 23266 17118
rect 23214 17042 23266 17054
rect 24334 17106 24386 17118
rect 24334 17042 24386 17054
rect 25342 17106 25394 17118
rect 25342 17042 25394 17054
rect 26910 17106 26962 17118
rect 26910 17042 26962 17054
rect 28142 17106 28194 17118
rect 28142 17042 28194 17054
rect 28590 17106 28642 17118
rect 30270 17106 30322 17118
rect 28914 17054 28926 17106
rect 28978 17054 28990 17106
rect 28590 17042 28642 17054
rect 30270 17042 30322 17054
rect 30830 17106 30882 17118
rect 30830 17042 30882 17054
rect 31502 17106 31554 17118
rect 31502 17042 31554 17054
rect 32062 17106 32114 17118
rect 32062 17042 32114 17054
rect 33182 17106 33234 17118
rect 33182 17042 33234 17054
rect 33966 17106 34018 17118
rect 33966 17042 34018 17054
rect 34190 17106 34242 17118
rect 34190 17042 34242 17054
rect 35198 17106 35250 17118
rect 35198 17042 35250 17054
rect 35758 17106 35810 17118
rect 35758 17042 35810 17054
rect 36542 17106 36594 17118
rect 36542 17042 36594 17054
rect 38894 17106 38946 17118
rect 38894 17042 38946 17054
rect 39678 17106 39730 17118
rect 39678 17042 39730 17054
rect 40126 17106 40178 17118
rect 40126 17042 40178 17054
rect 41358 17106 41410 17118
rect 41358 17042 41410 17054
rect 42814 17106 42866 17118
rect 42814 17042 42866 17054
rect 46398 17106 46450 17118
rect 46398 17042 46450 17054
rect 46958 17106 47010 17118
rect 46958 17042 47010 17054
rect 47406 17106 47458 17118
rect 47406 17042 47458 17054
rect 48862 17106 48914 17118
rect 48862 17042 48914 17054
rect 49086 17106 49138 17118
rect 49086 17042 49138 17054
rect 49310 17106 49362 17118
rect 49310 17042 49362 17054
rect 49758 17106 49810 17118
rect 49758 17042 49810 17054
rect 2046 16994 2098 17006
rect 13470 16994 13522 17006
rect 23550 16994 23602 17006
rect 10546 16942 10558 16994
rect 10610 16942 10622 16994
rect 14690 16942 14702 16994
rect 14754 16942 14766 16994
rect 2046 16930 2098 16942
rect 13470 16930 13522 16942
rect 23550 16930 23602 16942
rect 24446 16994 24498 17006
rect 24446 16930 24498 16942
rect 25454 16994 25506 17006
rect 25454 16930 25506 16942
rect 36430 16994 36482 17006
rect 36430 16930 36482 16942
rect 36990 16994 37042 17006
rect 36990 16930 37042 16942
rect 39118 16994 39170 17006
rect 39118 16930 39170 16942
rect 39230 16994 39282 17006
rect 39230 16930 39282 16942
rect 43374 16994 43426 17006
rect 43374 16930 43426 16942
rect 43710 16994 43762 17006
rect 43710 16930 43762 16942
rect 43934 16994 43986 17006
rect 43934 16930 43986 16942
rect 44270 16994 44322 17006
rect 44270 16930 44322 16942
rect 45838 16994 45890 17006
rect 45838 16930 45890 16942
rect 46286 16994 46338 17006
rect 46286 16930 46338 16942
rect 49198 16994 49250 17006
rect 49198 16930 49250 16942
rect 26798 16882 26850 16894
rect 1810 16830 1822 16882
rect 1874 16830 1886 16882
rect 9874 16830 9886 16882
rect 9938 16830 9950 16882
rect 14018 16830 14030 16882
rect 14082 16830 14094 16882
rect 21858 16830 21870 16882
rect 21922 16830 21934 16882
rect 23874 16830 23886 16882
rect 23938 16830 23950 16882
rect 26798 16818 26850 16830
rect 27022 16882 27074 16894
rect 27022 16818 27074 16830
rect 27470 16882 27522 16894
rect 27470 16818 27522 16830
rect 27694 16882 27746 16894
rect 27694 16818 27746 16830
rect 27918 16882 27970 16894
rect 27918 16818 27970 16830
rect 31950 16882 32002 16894
rect 31950 16818 32002 16830
rect 34750 16882 34802 16894
rect 34750 16818 34802 16830
rect 34974 16882 35026 16894
rect 34974 16818 35026 16830
rect 35310 16882 35362 16894
rect 40798 16882 40850 16894
rect 41806 16882 41858 16894
rect 37650 16830 37662 16882
rect 37714 16830 37726 16882
rect 38658 16830 38670 16882
rect 38722 16830 38734 16882
rect 41122 16830 41134 16882
rect 41186 16830 41198 16882
rect 35310 16818 35362 16830
rect 40798 16818 40850 16830
rect 41806 16818 41858 16830
rect 42030 16882 42082 16894
rect 46622 16882 46674 16894
rect 42354 16830 42366 16882
rect 42418 16830 42430 16882
rect 44930 16830 44942 16882
rect 44994 16830 45006 16882
rect 42030 16818 42082 16830
rect 46622 16818 46674 16830
rect 8878 16770 8930 16782
rect 26462 16770 26514 16782
rect 12674 16718 12686 16770
rect 12738 16718 12750 16770
rect 16818 16718 16830 16770
rect 16882 16718 16894 16770
rect 17602 16718 17614 16770
rect 17666 16718 17678 16770
rect 8878 16706 8930 16718
rect 26462 16706 26514 16718
rect 27806 16770 27858 16782
rect 27806 16706 27858 16718
rect 30606 16770 30658 16782
rect 38334 16770 38386 16782
rect 37874 16718 37886 16770
rect 37938 16718 37950 16770
rect 30606 16706 30658 16718
rect 38334 16706 38386 16718
rect 41918 16770 41970 16782
rect 41918 16706 41970 16718
rect 43486 16770 43538 16782
rect 47854 16770 47906 16782
rect 45154 16718 45166 16770
rect 45218 16718 45230 16770
rect 43486 16706 43538 16718
rect 47854 16706 47906 16718
rect 8990 16658 9042 16670
rect 8990 16594 9042 16606
rect 23886 16658 23938 16670
rect 23886 16594 23938 16606
rect 24334 16658 24386 16670
rect 24334 16594 24386 16606
rect 25342 16658 25394 16670
rect 26238 16658 26290 16670
rect 25890 16606 25902 16658
rect 25954 16606 25966 16658
rect 25342 16594 25394 16606
rect 26238 16594 26290 16606
rect 30942 16658 30994 16670
rect 30942 16594 30994 16606
rect 32062 16658 32114 16670
rect 32062 16594 32114 16606
rect 36542 16658 36594 16670
rect 36542 16594 36594 16606
rect 38670 16658 38722 16670
rect 38670 16594 38722 16606
rect 41022 16658 41074 16670
rect 41022 16594 41074 16606
rect 45614 16658 45666 16670
rect 45614 16594 45666 16606
rect 45950 16658 46002 16670
rect 45950 16594 46002 16606
rect 1344 16490 58576 16524
rect 1344 16438 4478 16490
rect 4530 16438 4582 16490
rect 4634 16438 4686 16490
rect 4738 16438 35198 16490
rect 35250 16438 35302 16490
rect 35354 16438 35406 16490
rect 35458 16438 58576 16490
rect 1344 16404 58576 16438
rect 49086 16322 49138 16334
rect 38322 16270 38334 16322
rect 38386 16319 38398 16322
rect 38658 16319 38670 16322
rect 38386 16273 38670 16319
rect 38386 16270 38398 16273
rect 38658 16270 38670 16273
rect 38722 16270 38734 16322
rect 49086 16258 49138 16270
rect 1822 16210 1874 16222
rect 12686 16210 12738 16222
rect 22878 16210 22930 16222
rect 9090 16158 9102 16210
rect 9154 16158 9166 16210
rect 11218 16158 11230 16210
rect 11282 16158 11294 16210
rect 17266 16158 17278 16210
rect 17330 16158 17342 16210
rect 18610 16158 18622 16210
rect 18674 16158 18686 16210
rect 20738 16158 20750 16210
rect 20802 16158 20814 16210
rect 1822 16146 1874 16158
rect 12686 16146 12738 16158
rect 22878 16146 22930 16158
rect 25342 16210 25394 16222
rect 30046 16210 30098 16222
rect 37102 16210 37154 16222
rect 28578 16158 28590 16210
rect 28642 16158 28654 16210
rect 30594 16158 30606 16210
rect 30658 16158 30670 16210
rect 25342 16146 25394 16158
rect 30046 16146 30098 16158
rect 37102 16146 37154 16158
rect 46286 16210 46338 16222
rect 46286 16146 46338 16158
rect 47294 16210 47346 16222
rect 47294 16146 47346 16158
rect 49982 16210 50034 16222
rect 49982 16146 50034 16158
rect 37998 16098 38050 16110
rect 44830 16098 44882 16110
rect 8418 16046 8430 16098
rect 8482 16046 8494 16098
rect 14466 16046 14478 16098
rect 14530 16046 14542 16098
rect 17826 16046 17838 16098
rect 17890 16046 17902 16098
rect 23650 16046 23662 16098
rect 23714 16046 23726 16098
rect 23874 16046 23886 16098
rect 23938 16046 23950 16098
rect 24546 16046 24558 16098
rect 24610 16046 24622 16098
rect 25778 16046 25790 16098
rect 25842 16046 25854 16098
rect 35634 16046 35646 16098
rect 35698 16046 35710 16098
rect 42802 16046 42814 16098
rect 42866 16046 42878 16098
rect 37998 16034 38050 16046
rect 44830 16034 44882 16046
rect 45054 16098 45106 16110
rect 45054 16034 45106 16046
rect 45502 16098 45554 16110
rect 46622 16098 46674 16110
rect 45826 16046 45838 16098
rect 45890 16046 45902 16098
rect 45502 16034 45554 16046
rect 46622 16034 46674 16046
rect 47630 16098 47682 16110
rect 47630 16034 47682 16046
rect 47854 16098 47906 16110
rect 47854 16034 47906 16046
rect 48414 16098 48466 16110
rect 48414 16034 48466 16046
rect 49534 16098 49586 16110
rect 49534 16034 49586 16046
rect 50430 16098 50482 16110
rect 50430 16034 50482 16046
rect 29374 15986 29426 15998
rect 15138 15934 15150 15986
rect 15202 15934 15214 15986
rect 23762 15934 23774 15986
rect 23826 15934 23838 15986
rect 26450 15934 26462 15986
rect 26514 15934 26526 15986
rect 29374 15922 29426 15934
rect 37886 15986 37938 15998
rect 46734 15986 46786 15998
rect 39218 15934 39230 15986
rect 39282 15934 39294 15986
rect 37886 15922 37938 15934
rect 46734 15922 46786 15934
rect 49422 15986 49474 15998
rect 49422 15922 49474 15934
rect 12798 15874 12850 15886
rect 12798 15810 12850 15822
rect 29038 15874 29090 15886
rect 29038 15810 29090 15822
rect 29262 15874 29314 15886
rect 29262 15810 29314 15822
rect 36206 15874 36258 15886
rect 36206 15810 36258 15822
rect 37662 15874 37714 15886
rect 37662 15810 37714 15822
rect 38446 15874 38498 15886
rect 38446 15810 38498 15822
rect 44942 15874 44994 15886
rect 44942 15810 44994 15822
rect 46958 15874 47010 15886
rect 48750 15874 48802 15886
rect 48178 15822 48190 15874
rect 48242 15822 48254 15874
rect 46958 15810 47010 15822
rect 48750 15810 48802 15822
rect 48974 15874 49026 15886
rect 48974 15810 49026 15822
rect 49198 15874 49250 15886
rect 49198 15810 49250 15822
rect 1344 15706 58576 15740
rect 1344 15654 19838 15706
rect 19890 15654 19942 15706
rect 19994 15654 20046 15706
rect 20098 15654 50558 15706
rect 50610 15654 50662 15706
rect 50714 15654 50766 15706
rect 50818 15654 58576 15706
rect 1344 15620 58576 15654
rect 16382 15538 16434 15550
rect 16382 15474 16434 15486
rect 16718 15538 16770 15550
rect 16718 15474 16770 15486
rect 22990 15538 23042 15550
rect 22990 15474 23042 15486
rect 25342 15538 25394 15550
rect 25342 15474 25394 15486
rect 26238 15538 26290 15550
rect 26238 15474 26290 15486
rect 26350 15538 26402 15550
rect 26350 15474 26402 15486
rect 26462 15538 26514 15550
rect 26462 15474 26514 15486
rect 28030 15538 28082 15550
rect 28030 15474 28082 15486
rect 29598 15538 29650 15550
rect 29598 15474 29650 15486
rect 32286 15538 32338 15550
rect 32286 15474 32338 15486
rect 33294 15538 33346 15550
rect 33294 15474 33346 15486
rect 35198 15538 35250 15550
rect 35198 15474 35250 15486
rect 35870 15538 35922 15550
rect 35870 15474 35922 15486
rect 35982 15538 36034 15550
rect 35982 15474 36034 15486
rect 36878 15538 36930 15550
rect 36878 15474 36930 15486
rect 39118 15538 39170 15550
rect 42702 15538 42754 15550
rect 40338 15486 40350 15538
rect 40402 15486 40414 15538
rect 39118 15474 39170 15486
rect 42702 15474 42754 15486
rect 48750 15538 48802 15550
rect 48750 15474 48802 15486
rect 48862 15538 48914 15550
rect 48862 15474 48914 15486
rect 49758 15538 49810 15550
rect 49758 15474 49810 15486
rect 50430 15538 50482 15550
rect 50430 15474 50482 15486
rect 16830 15426 16882 15438
rect 13682 15374 13694 15426
rect 13746 15374 13758 15426
rect 16830 15362 16882 15374
rect 22318 15426 22370 15438
rect 22318 15362 22370 15374
rect 22654 15426 22706 15438
rect 22654 15362 22706 15374
rect 22766 15426 22818 15438
rect 22766 15362 22818 15374
rect 26798 15426 26850 15438
rect 26798 15362 26850 15374
rect 28142 15426 28194 15438
rect 28142 15362 28194 15374
rect 29822 15426 29874 15438
rect 29822 15362 29874 15374
rect 29934 15426 29986 15438
rect 29934 15362 29986 15374
rect 32174 15426 32226 15438
rect 32174 15362 32226 15374
rect 33518 15426 33570 15438
rect 33518 15362 33570 15374
rect 39006 15426 39058 15438
rect 48078 15426 48130 15438
rect 42018 15374 42030 15426
rect 42082 15374 42094 15426
rect 39006 15362 39058 15374
rect 48078 15362 48130 15374
rect 21870 15314 21922 15326
rect 14466 15262 14478 15314
rect 14530 15262 14542 15314
rect 17714 15262 17726 15314
rect 17778 15262 17790 15314
rect 21870 15250 21922 15262
rect 23774 15314 23826 15326
rect 23774 15250 23826 15262
rect 24110 15314 24162 15326
rect 24110 15250 24162 15262
rect 24334 15314 24386 15326
rect 25230 15314 25282 15326
rect 24658 15262 24670 15314
rect 24722 15262 24734 15314
rect 24334 15250 24386 15262
rect 25230 15250 25282 15262
rect 25566 15314 25618 15326
rect 25566 15250 25618 15262
rect 25790 15314 25842 15326
rect 27694 15314 27746 15326
rect 28702 15314 28754 15326
rect 27234 15262 27246 15314
rect 27298 15262 27310 15314
rect 28354 15262 28366 15314
rect 28418 15262 28430 15314
rect 25790 15250 25842 15262
rect 27694 15250 27746 15262
rect 28702 15250 28754 15262
rect 29150 15314 29202 15326
rect 29150 15250 29202 15262
rect 30158 15314 30210 15326
rect 32510 15314 32562 15326
rect 30482 15262 30494 15314
rect 30546 15262 30558 15314
rect 30930 15262 30942 15314
rect 30994 15262 31006 15314
rect 31826 15262 31838 15314
rect 31890 15262 31902 15314
rect 30158 15250 30210 15262
rect 32510 15250 32562 15262
rect 33070 15314 33122 15326
rect 33070 15250 33122 15262
rect 33966 15314 34018 15326
rect 33966 15250 34018 15262
rect 34190 15314 34242 15326
rect 34190 15250 34242 15262
rect 34638 15314 34690 15326
rect 34638 15250 34690 15262
rect 34750 15314 34802 15326
rect 34750 15250 34802 15262
rect 35310 15314 35362 15326
rect 35310 15250 35362 15262
rect 35422 15314 35474 15326
rect 35422 15250 35474 15262
rect 35758 15314 35810 15326
rect 35758 15250 35810 15262
rect 36430 15314 36482 15326
rect 39790 15314 39842 15326
rect 37650 15262 37662 15314
rect 37714 15262 37726 15314
rect 38322 15262 38334 15314
rect 38386 15262 38398 15314
rect 36430 15250 36482 15262
rect 39790 15250 39842 15262
rect 40014 15314 40066 15326
rect 48974 15314 49026 15326
rect 41010 15262 41022 15314
rect 41074 15262 41086 15314
rect 41570 15262 41582 15314
rect 41634 15262 41646 15314
rect 43026 15262 43038 15314
rect 43090 15262 43102 15314
rect 43810 15262 43822 15314
rect 43874 15262 43886 15314
rect 46610 15262 46622 15314
rect 46674 15262 46686 15314
rect 47282 15262 47294 15314
rect 47346 15262 47358 15314
rect 49298 15262 49310 15314
rect 49362 15262 49374 15314
rect 50978 15262 50990 15314
rect 51042 15262 51054 15314
rect 40014 15250 40066 15262
rect 48974 15250 49026 15262
rect 23550 15202 23602 15214
rect 11554 15150 11566 15202
rect 11618 15150 11630 15202
rect 18386 15150 18398 15202
rect 18450 15150 18462 15202
rect 20514 15150 20526 15202
rect 20578 15150 20590 15202
rect 23550 15138 23602 15150
rect 24222 15202 24274 15214
rect 24222 15138 24274 15150
rect 33182 15202 33234 15214
rect 33182 15138 33234 15150
rect 34078 15202 34130 15214
rect 46510 15202 46562 15214
rect 37874 15150 37886 15202
rect 37938 15150 37950 15202
rect 41906 15150 41918 15202
rect 41970 15150 41982 15202
rect 45938 15150 45950 15202
rect 46002 15150 46014 15202
rect 52770 15150 52782 15202
rect 52834 15150 52846 15202
rect 34078 15138 34130 15150
rect 46510 15138 46562 15150
rect 31278 15090 31330 15102
rect 39118 15090 39170 15102
rect 21858 15038 21870 15090
rect 21922 15087 21934 15090
rect 22306 15087 22318 15090
rect 21922 15041 22318 15087
rect 21922 15038 21934 15041
rect 22306 15038 22318 15041
rect 22370 15038 22382 15090
rect 23202 15038 23214 15090
rect 23266 15038 23278 15090
rect 38098 15038 38110 15090
rect 38162 15038 38174 15090
rect 46722 15038 46734 15090
rect 46786 15038 46798 15090
rect 31278 15026 31330 15038
rect 39118 15026 39170 15038
rect 1344 14922 58576 14956
rect 1344 14870 4478 14922
rect 4530 14870 4582 14922
rect 4634 14870 4686 14922
rect 4738 14870 35198 14922
rect 35250 14870 35302 14922
rect 35354 14870 35406 14922
rect 35458 14870 58576 14922
rect 1344 14836 58576 14870
rect 36318 14754 36370 14766
rect 10098 14702 10110 14754
rect 10162 14702 10174 14754
rect 18722 14702 18734 14754
rect 18786 14702 18798 14754
rect 27906 14702 27918 14754
rect 27970 14751 27982 14754
rect 28466 14751 28478 14754
rect 27970 14705 28478 14751
rect 27970 14702 27982 14705
rect 28466 14702 28478 14705
rect 28530 14702 28542 14754
rect 29362 14702 29374 14754
rect 29426 14702 29438 14754
rect 36318 14690 36370 14702
rect 36878 14754 36930 14766
rect 36878 14690 36930 14702
rect 23886 14642 23938 14654
rect 27134 14642 27186 14654
rect 10434 14590 10446 14642
rect 10498 14590 10510 14642
rect 12114 14590 12126 14642
rect 12178 14590 12190 14642
rect 21858 14590 21870 14642
rect 21922 14590 21934 14642
rect 23090 14590 23102 14642
rect 23154 14590 23166 14642
rect 25442 14590 25454 14642
rect 25506 14590 25518 14642
rect 23886 14578 23938 14590
rect 27134 14578 27186 14590
rect 27806 14642 27858 14654
rect 27806 14578 27858 14590
rect 28142 14642 28194 14654
rect 28142 14578 28194 14590
rect 28590 14642 28642 14654
rect 28590 14578 28642 14590
rect 30718 14642 30770 14654
rect 44046 14642 44098 14654
rect 31826 14590 31838 14642
rect 31890 14590 31902 14642
rect 33394 14590 33406 14642
rect 33458 14590 33470 14642
rect 35522 14590 35534 14642
rect 35586 14590 35598 14642
rect 40898 14590 40910 14642
rect 40962 14590 40974 14642
rect 43026 14590 43038 14642
rect 43090 14590 43102 14642
rect 30718 14578 30770 14590
rect 44046 14578 44098 14590
rect 45502 14642 45554 14654
rect 45502 14578 45554 14590
rect 47518 14642 47570 14654
rect 50754 14590 50766 14642
rect 50818 14590 50830 14642
rect 47518 14578 47570 14590
rect 9550 14530 9602 14542
rect 17950 14530 18002 14542
rect 19630 14530 19682 14542
rect 9762 14478 9774 14530
rect 9826 14478 9838 14530
rect 11106 14478 11118 14530
rect 11170 14478 11182 14530
rect 11890 14478 11902 14530
rect 11954 14478 11966 14530
rect 18162 14478 18174 14530
rect 18226 14478 18238 14530
rect 19282 14478 19294 14530
rect 19346 14478 19358 14530
rect 9550 14466 9602 14478
rect 17950 14466 18002 14478
rect 19630 14466 19682 14478
rect 19966 14530 20018 14542
rect 24110 14530 24162 14542
rect 20402 14478 20414 14530
rect 20466 14478 20478 14530
rect 19966 14466 20018 14478
rect 24110 14466 24162 14478
rect 24334 14530 24386 14542
rect 24334 14466 24386 14478
rect 24782 14530 24834 14542
rect 26462 14530 26514 14542
rect 25218 14478 25230 14530
rect 25282 14478 25294 14530
rect 26114 14478 26126 14530
rect 26178 14478 26190 14530
rect 24782 14466 24834 14478
rect 26462 14466 26514 14478
rect 29710 14530 29762 14542
rect 29710 14466 29762 14478
rect 29934 14530 29986 14542
rect 30606 14530 30658 14542
rect 36206 14530 36258 14542
rect 30258 14478 30270 14530
rect 30322 14478 30334 14530
rect 31154 14478 31166 14530
rect 31218 14478 31230 14530
rect 32162 14478 32174 14530
rect 32226 14478 32238 14530
rect 32610 14478 32622 14530
rect 32674 14478 32686 14530
rect 29934 14466 29986 14478
rect 30606 14466 30658 14478
rect 36206 14466 36258 14478
rect 38110 14530 38162 14542
rect 38110 14466 38162 14478
rect 38334 14530 38386 14542
rect 44830 14530 44882 14542
rect 38658 14478 38670 14530
rect 38722 14478 38734 14530
rect 39778 14478 39790 14530
rect 39842 14478 39854 14530
rect 40226 14478 40238 14530
rect 40290 14478 40302 14530
rect 38334 14466 38386 14478
rect 44830 14466 44882 14478
rect 45166 14530 45218 14542
rect 45166 14466 45218 14478
rect 46286 14530 46338 14542
rect 46286 14466 46338 14478
rect 46622 14530 46674 14542
rect 47058 14478 47070 14530
rect 47122 14478 47134 14530
rect 47954 14478 47966 14530
rect 48018 14478 48030 14530
rect 46622 14466 46674 14478
rect 21422 14418 21474 14430
rect 26574 14418 26626 14430
rect 25106 14366 25118 14418
rect 25170 14366 25182 14418
rect 21422 14354 21474 14366
rect 26574 14354 26626 14366
rect 30830 14418 30882 14430
rect 36990 14418 37042 14430
rect 31266 14366 31278 14418
rect 31330 14366 31342 14418
rect 30830 14354 30882 14366
rect 36990 14354 37042 14366
rect 37438 14418 37490 14430
rect 37438 14354 37490 14366
rect 37886 14418 37938 14430
rect 45950 14418 46002 14430
rect 38770 14366 38782 14418
rect 38834 14366 38846 14418
rect 37886 14354 37938 14366
rect 45950 14354 46002 14366
rect 46062 14418 46114 14430
rect 48626 14366 48638 14418
rect 48690 14366 48702 14418
rect 46062 14354 46114 14366
rect 21310 14306 21362 14318
rect 21310 14242 21362 14254
rect 22318 14306 22370 14318
rect 22318 14242 22370 14254
rect 22654 14306 22706 14318
rect 22654 14242 22706 14254
rect 24222 14306 24274 14318
rect 24222 14242 24274 14254
rect 36318 14306 36370 14318
rect 36318 14242 36370 14254
rect 37214 14306 37266 14318
rect 37214 14242 37266 14254
rect 38222 14306 38274 14318
rect 43486 14306 43538 14318
rect 39666 14254 39678 14306
rect 39730 14254 39742 14306
rect 38222 14242 38274 14254
rect 43486 14242 43538 14254
rect 44942 14306 44994 14318
rect 44942 14242 44994 14254
rect 1344 14138 58576 14172
rect 1344 14086 19838 14138
rect 19890 14086 19942 14138
rect 19994 14086 20046 14138
rect 20098 14086 50558 14138
rect 50610 14086 50662 14138
rect 50714 14086 50766 14138
rect 50818 14086 58576 14138
rect 1344 14052 58576 14086
rect 28254 13970 28306 13982
rect 27570 13918 27582 13970
rect 27634 13918 27646 13970
rect 28254 13906 28306 13918
rect 35086 13970 35138 13982
rect 35086 13906 35138 13918
rect 36318 13970 36370 13982
rect 36318 13906 36370 13918
rect 38782 13970 38834 13982
rect 38782 13906 38834 13918
rect 39230 13970 39282 13982
rect 39230 13906 39282 13918
rect 40126 13970 40178 13982
rect 40126 13906 40178 13918
rect 40238 13970 40290 13982
rect 40238 13906 40290 13918
rect 40350 13970 40402 13982
rect 40350 13906 40402 13918
rect 42142 13970 42194 13982
rect 42142 13906 42194 13918
rect 42366 13970 42418 13982
rect 42366 13906 42418 13918
rect 43038 13970 43090 13982
rect 43038 13906 43090 13918
rect 43486 13970 43538 13982
rect 43486 13906 43538 13918
rect 44494 13970 44546 13982
rect 44494 13906 44546 13918
rect 47854 13970 47906 13982
rect 47854 13906 47906 13918
rect 48750 13970 48802 13982
rect 48750 13906 48802 13918
rect 49198 13970 49250 13982
rect 49198 13906 49250 13918
rect 49870 13970 49922 13982
rect 49870 13906 49922 13918
rect 25230 13858 25282 13870
rect 27246 13858 27298 13870
rect 19282 13806 19294 13858
rect 19346 13806 19358 13858
rect 22530 13806 22542 13858
rect 22594 13806 22606 13858
rect 26898 13806 26910 13858
rect 26962 13806 26974 13858
rect 25230 13794 25282 13806
rect 27246 13794 27298 13806
rect 27918 13858 27970 13870
rect 33406 13858 33458 13870
rect 28578 13806 28590 13858
rect 28642 13806 28654 13858
rect 31154 13806 31166 13858
rect 31218 13806 31230 13858
rect 27918 13794 27970 13806
rect 33406 13794 33458 13806
rect 35198 13858 35250 13870
rect 35198 13794 35250 13806
rect 36766 13858 36818 13870
rect 36766 13794 36818 13806
rect 37438 13858 37490 13870
rect 37438 13794 37490 13806
rect 41918 13858 41970 13870
rect 41918 13794 41970 13806
rect 42478 13858 42530 13870
rect 47630 13858 47682 13870
rect 46722 13806 46734 13858
rect 46786 13806 46798 13858
rect 42478 13794 42530 13806
rect 47630 13794 47682 13806
rect 34526 13746 34578 13758
rect 18498 13694 18510 13746
rect 18562 13694 18574 13746
rect 21858 13694 21870 13746
rect 21922 13694 21934 13746
rect 25890 13694 25902 13746
rect 25954 13694 25966 13746
rect 31938 13694 31950 13746
rect 32002 13694 32014 13746
rect 34290 13694 34302 13746
rect 34354 13694 34366 13746
rect 34526 13682 34578 13694
rect 34862 13746 34914 13758
rect 34862 13682 34914 13694
rect 37326 13746 37378 13758
rect 37326 13682 37378 13694
rect 37886 13746 37938 13758
rect 39006 13746 39058 13758
rect 38434 13694 38446 13746
rect 38498 13694 38510 13746
rect 37886 13682 37938 13694
rect 39006 13682 39058 13694
rect 39678 13746 39730 13758
rect 45614 13746 45666 13758
rect 47406 13746 47458 13758
rect 41458 13694 41470 13746
rect 41522 13694 41534 13746
rect 46162 13694 46174 13746
rect 46226 13694 46238 13746
rect 47058 13694 47070 13746
rect 47122 13694 47134 13746
rect 39678 13682 39730 13694
rect 45614 13682 45666 13694
rect 47406 13682 47458 13694
rect 48974 13746 49026 13758
rect 48974 13682 49026 13694
rect 32398 13634 32450 13646
rect 21410 13582 21422 13634
rect 21474 13582 21486 13634
rect 24658 13582 24670 13634
rect 24722 13582 24734 13634
rect 26002 13582 26014 13634
rect 26066 13582 26078 13634
rect 29026 13582 29038 13634
rect 29090 13582 29102 13634
rect 32398 13570 32450 13582
rect 33630 13634 33682 13646
rect 33630 13570 33682 13582
rect 35870 13634 35922 13646
rect 35870 13570 35922 13582
rect 38894 13634 38946 13646
rect 43934 13634 43986 13646
rect 47518 13634 47570 13646
rect 41122 13582 41134 13634
rect 41186 13582 41198 13634
rect 46722 13582 46734 13634
rect 46786 13582 46798 13634
rect 38894 13570 38946 13582
rect 43934 13570 43986 13582
rect 47518 13570 47570 13582
rect 48862 13634 48914 13646
rect 48862 13570 48914 13582
rect 32286 13522 32338 13534
rect 32286 13458 32338 13470
rect 37438 13522 37490 13534
rect 37438 13458 37490 13470
rect 38110 13522 38162 13534
rect 38110 13458 38162 13470
rect 1344 13354 58576 13388
rect 1344 13302 4478 13354
rect 4530 13302 4582 13354
rect 4634 13302 4686 13354
rect 4738 13302 35198 13354
rect 35250 13302 35302 13354
rect 35354 13302 35406 13354
rect 35458 13302 58576 13354
rect 1344 13268 58576 13302
rect 33406 13186 33458 13198
rect 40350 13186 40402 13198
rect 24434 13134 24446 13186
rect 24498 13134 24510 13186
rect 30818 13134 30830 13186
rect 30882 13134 30894 13186
rect 33730 13134 33742 13186
rect 33794 13134 33806 13186
rect 33406 13122 33458 13134
rect 40350 13122 40402 13134
rect 46846 13186 46898 13198
rect 46846 13122 46898 13134
rect 20750 13074 20802 13086
rect 20750 13010 20802 13022
rect 27582 13074 27634 13086
rect 27582 13010 27634 13022
rect 28254 13074 28306 13086
rect 28254 13010 28306 13022
rect 29374 13074 29426 13086
rect 29374 13010 29426 13022
rect 30270 13074 30322 13086
rect 33182 13074 33234 13086
rect 31042 13022 31054 13074
rect 31106 13022 31118 13074
rect 32386 13022 32398 13074
rect 32450 13022 32462 13074
rect 30270 13010 30322 13022
rect 33182 13010 33234 13022
rect 35310 13074 35362 13086
rect 35310 13010 35362 13022
rect 35870 13074 35922 13086
rect 48526 13074 48578 13086
rect 37874 13022 37886 13074
rect 37938 13022 37950 13074
rect 40002 13022 40014 13074
rect 40066 13022 40078 13074
rect 44258 13022 44270 13074
rect 44322 13022 44334 13074
rect 45490 13022 45502 13074
rect 45554 13022 45566 13074
rect 35870 13010 35922 13022
rect 48526 13010 48578 13022
rect 49422 13074 49474 13086
rect 49422 13010 49474 13022
rect 22990 12962 23042 12974
rect 25006 12962 25058 12974
rect 23650 12910 23662 12962
rect 23714 12910 23726 12962
rect 24098 12910 24110 12962
rect 24162 12910 24174 12962
rect 24658 12910 24670 12962
rect 24722 12910 24734 12962
rect 22990 12898 23042 12910
rect 25006 12898 25058 12910
rect 25342 12962 25394 12974
rect 26238 12962 26290 12974
rect 25442 12910 25454 12962
rect 25506 12910 25518 12962
rect 25342 12898 25394 12910
rect 26238 12898 26290 12910
rect 26574 12962 26626 12974
rect 31950 12962 32002 12974
rect 31490 12910 31502 12962
rect 31554 12910 31566 12962
rect 26574 12898 26626 12910
rect 31950 12898 32002 12910
rect 36430 12962 36482 12974
rect 40798 12962 40850 12974
rect 37090 12910 37102 12962
rect 37154 12910 37166 12962
rect 36430 12898 36482 12910
rect 40798 12898 40850 12910
rect 41134 12962 41186 12974
rect 46286 12962 46338 12974
rect 41458 12910 41470 12962
rect 41522 12910 41534 12962
rect 45826 12910 45838 12962
rect 45890 12910 45902 12962
rect 41134 12898 41186 12910
rect 46286 12898 46338 12910
rect 46622 12962 46674 12974
rect 46622 12898 46674 12910
rect 47518 12962 47570 12974
rect 47518 12898 47570 12910
rect 48190 12962 48242 12974
rect 48190 12898 48242 12910
rect 48414 12962 48466 12974
rect 48414 12898 48466 12910
rect 49086 12962 49138 12974
rect 49086 12898 49138 12910
rect 32510 12850 32562 12862
rect 32510 12786 32562 12798
rect 34190 12850 34242 12862
rect 34190 12786 34242 12798
rect 34750 12850 34802 12862
rect 34750 12786 34802 12798
rect 40462 12850 40514 12862
rect 47742 12850 47794 12862
rect 42130 12798 42142 12850
rect 42194 12798 42206 12850
rect 47170 12798 47182 12850
rect 47234 12798 47246 12850
rect 40462 12786 40514 12798
rect 47742 12786 47794 12798
rect 26462 12738 26514 12750
rect 26462 12674 26514 12686
rect 27022 12738 27074 12750
rect 27022 12674 27074 12686
rect 32286 12738 32338 12750
rect 32286 12674 32338 12686
rect 34638 12738 34690 12750
rect 34638 12674 34690 12686
rect 40910 12738 40962 12750
rect 40910 12674 40962 12686
rect 47630 12738 47682 12750
rect 47630 12674 47682 12686
rect 48638 12738 48690 12750
rect 48638 12674 48690 12686
rect 1344 12570 58576 12604
rect 1344 12518 19838 12570
rect 19890 12518 19942 12570
rect 19994 12518 20046 12570
rect 20098 12518 50558 12570
rect 50610 12518 50662 12570
rect 50714 12518 50766 12570
rect 50818 12518 58576 12570
rect 1344 12484 58576 12518
rect 19966 12402 20018 12414
rect 19966 12338 20018 12350
rect 24782 12402 24834 12414
rect 24782 12338 24834 12350
rect 25230 12402 25282 12414
rect 25230 12338 25282 12350
rect 30270 12402 30322 12414
rect 30270 12338 30322 12350
rect 31054 12402 31106 12414
rect 31054 12338 31106 12350
rect 32398 12402 32450 12414
rect 32398 12338 32450 12350
rect 33294 12402 33346 12414
rect 33294 12338 33346 12350
rect 40238 12402 40290 12414
rect 40238 12338 40290 12350
rect 41134 12402 41186 12414
rect 41134 12338 41186 12350
rect 42590 12402 42642 12414
rect 42590 12338 42642 12350
rect 43934 12402 43986 12414
rect 43934 12338 43986 12350
rect 44606 12402 44658 12414
rect 44606 12338 44658 12350
rect 47966 12402 48018 12414
rect 47966 12338 48018 12350
rect 48190 12402 48242 12414
rect 48190 12338 48242 12350
rect 48862 12402 48914 12414
rect 48862 12338 48914 12350
rect 23998 12290 24050 12302
rect 20962 12238 20974 12290
rect 21026 12238 21038 12290
rect 23998 12226 24050 12238
rect 31278 12290 31330 12302
rect 31278 12226 31330 12238
rect 31390 12290 31442 12302
rect 31390 12226 31442 12238
rect 38670 12290 38722 12302
rect 38670 12226 38722 12238
rect 44270 12290 44322 12302
rect 44270 12226 44322 12238
rect 44382 12290 44434 12302
rect 44382 12226 44434 12238
rect 47854 12290 47906 12302
rect 47854 12226 47906 12238
rect 20302 12178 20354 12190
rect 25790 12178 25842 12190
rect 29262 12178 29314 12190
rect 30830 12178 30882 12190
rect 34750 12178 34802 12190
rect 38334 12178 38386 12190
rect 20738 12126 20750 12178
rect 20802 12126 20814 12178
rect 21522 12126 21534 12178
rect 21586 12126 21598 12178
rect 21970 12126 21982 12178
rect 22034 12126 22046 12178
rect 22530 12126 22542 12178
rect 22594 12126 22606 12178
rect 23762 12126 23774 12178
rect 23826 12126 23838 12178
rect 25442 12126 25454 12178
rect 25506 12126 25518 12178
rect 27682 12126 27694 12178
rect 27746 12126 27758 12178
rect 28018 12126 28030 12178
rect 28082 12126 28094 12178
rect 28690 12126 28702 12178
rect 28754 12126 28766 12178
rect 29698 12126 29710 12178
rect 29762 12126 29774 12178
rect 33954 12126 33966 12178
rect 34018 12126 34030 12178
rect 36194 12126 36206 12178
rect 36258 12126 36270 12178
rect 36754 12126 36766 12178
rect 36818 12126 36830 12178
rect 37874 12126 37886 12178
rect 37938 12126 37950 12178
rect 20302 12114 20354 12126
rect 25790 12114 25842 12126
rect 29262 12114 29314 12126
rect 30830 12114 30882 12126
rect 34750 12114 34802 12126
rect 38334 12114 38386 12126
rect 38894 12178 38946 12190
rect 41470 12178 41522 12190
rect 39554 12126 39566 12178
rect 39618 12126 39630 12178
rect 38894 12114 38946 12126
rect 41470 12114 41522 12126
rect 42814 12178 42866 12190
rect 45042 12126 45054 12178
rect 45106 12126 45118 12178
rect 45490 12126 45502 12178
rect 45554 12126 45566 12178
rect 46050 12126 46062 12178
rect 46114 12126 46126 12178
rect 47282 12126 47294 12178
rect 47346 12126 47358 12178
rect 42814 12114 42866 12126
rect 25566 12066 25618 12078
rect 22194 12014 22206 12066
rect 22258 12014 22270 12066
rect 25566 12002 25618 12014
rect 26126 12066 26178 12078
rect 26126 12002 26178 12014
rect 26574 12066 26626 12078
rect 31838 12066 31890 12078
rect 35310 12066 35362 12078
rect 28130 12014 28142 12066
rect 28194 12014 28206 12066
rect 33618 12014 33630 12066
rect 33682 12014 33694 12066
rect 35746 12014 35758 12066
rect 35810 12014 35822 12066
rect 37314 12014 37326 12066
rect 37378 12014 37390 12066
rect 43250 12014 43262 12066
rect 43314 12014 43326 12066
rect 45714 12014 45726 12066
rect 45778 12014 45790 12066
rect 47394 12014 47406 12066
rect 47458 12014 47470 12066
rect 26574 12002 26626 12014
rect 31838 12002 31890 12014
rect 35310 12002 35362 12014
rect 22082 11902 22094 11954
rect 22146 11902 22158 11954
rect 28802 11902 28814 11954
rect 28866 11902 28878 11954
rect 36530 11902 36542 11954
rect 36594 11902 36606 11954
rect 45378 11902 45390 11954
rect 45442 11902 45454 11954
rect 1344 11786 58576 11820
rect 1344 11734 4478 11786
rect 4530 11734 4582 11786
rect 4634 11734 4686 11786
rect 4738 11734 35198 11786
rect 35250 11734 35302 11786
rect 35354 11734 35406 11786
rect 35458 11734 58576 11786
rect 1344 11700 58576 11734
rect 19730 11566 19742 11618
rect 19794 11566 19806 11618
rect 21186 11566 21198 11618
rect 21250 11615 21262 11618
rect 21410 11615 21422 11618
rect 21250 11569 21422 11615
rect 21250 11566 21262 11569
rect 21410 11566 21422 11569
rect 21474 11566 21486 11618
rect 32050 11566 32062 11618
rect 32114 11566 32126 11618
rect 38658 11566 38670 11618
rect 38722 11566 38734 11618
rect 41458 11566 41470 11618
rect 41522 11566 41534 11618
rect 21534 11506 21586 11518
rect 19842 11454 19854 11506
rect 19906 11454 19918 11506
rect 21534 11442 21586 11454
rect 22654 11506 22706 11518
rect 32510 11506 32562 11518
rect 46174 11506 46226 11518
rect 31938 11454 31950 11506
rect 32002 11454 32014 11506
rect 34290 11454 34302 11506
rect 34354 11454 34366 11506
rect 36418 11454 36430 11506
rect 36482 11454 36494 11506
rect 40450 11454 40462 11506
rect 40514 11454 40526 11506
rect 46498 11454 46510 11506
rect 46562 11454 46574 11506
rect 48626 11454 48638 11506
rect 48690 11454 48702 11506
rect 22654 11442 22706 11454
rect 32510 11442 32562 11454
rect 46174 11442 46226 11454
rect 18734 11394 18786 11406
rect 29374 11394 29426 11406
rect 31054 11394 31106 11406
rect 37998 11394 38050 11406
rect 39902 11394 39954 11406
rect 42590 11394 42642 11406
rect 18386 11342 18398 11394
rect 18450 11342 18462 11394
rect 19506 11342 19518 11394
rect 19570 11342 19582 11394
rect 20514 11342 20526 11394
rect 20578 11342 20590 11394
rect 23314 11342 23326 11394
rect 23378 11342 23390 11394
rect 29810 11342 29822 11394
rect 29874 11342 29886 11394
rect 30818 11342 30830 11394
rect 30882 11342 30894 11394
rect 31490 11342 31502 11394
rect 31554 11342 31566 11394
rect 32946 11342 32958 11394
rect 33010 11342 33022 11394
rect 33618 11342 33630 11394
rect 33682 11342 33694 11394
rect 37202 11342 37214 11394
rect 37266 11342 37278 11394
rect 38098 11342 38110 11394
rect 38162 11342 38174 11394
rect 39218 11342 39230 11394
rect 39282 11342 39294 11394
rect 41346 11342 41358 11394
rect 41410 11342 41422 11394
rect 42130 11342 42142 11394
rect 42194 11342 42206 11394
rect 18734 11330 18786 11342
rect 29374 11330 29426 11342
rect 31054 11330 31106 11342
rect 37998 11330 38050 11342
rect 39902 11330 39954 11342
rect 42590 11330 42642 11342
rect 42926 11394 42978 11406
rect 44830 11394 44882 11406
rect 43026 11342 43038 11394
rect 43090 11342 43102 11394
rect 45154 11342 45166 11394
rect 45218 11342 45230 11394
rect 49298 11342 49310 11394
rect 49362 11342 49374 11394
rect 42926 11330 42978 11342
rect 44830 11330 44882 11342
rect 36990 11282 37042 11294
rect 40462 11282 40514 11294
rect 45502 11282 45554 11294
rect 20738 11230 20750 11282
rect 20802 11230 20814 11282
rect 25330 11230 25342 11282
rect 25394 11230 25406 11282
rect 33170 11230 33182 11282
rect 33234 11230 33246 11282
rect 39666 11230 39678 11282
rect 39730 11230 39742 11282
rect 40898 11230 40910 11282
rect 40962 11230 40974 11282
rect 36990 11218 37042 11230
rect 40462 11218 40514 11230
rect 45502 11218 45554 11230
rect 46062 11282 46114 11294
rect 46062 11218 46114 11230
rect 23102 11170 23154 11182
rect 23102 11106 23154 11118
rect 32398 11170 32450 11182
rect 32398 11106 32450 11118
rect 40238 11170 40290 11182
rect 40238 11106 40290 11118
rect 44382 11170 44434 11182
rect 44382 11106 44434 11118
rect 45390 11170 45442 11182
rect 45390 11106 45442 11118
rect 1344 11002 58576 11036
rect 1344 10950 19838 11002
rect 19890 10950 19942 11002
rect 19994 10950 20046 11002
rect 20098 10950 50558 11002
rect 50610 10950 50662 11002
rect 50714 10950 50766 11002
rect 50818 10950 58576 11002
rect 1344 10916 58576 10950
rect 32510 10834 32562 10846
rect 32510 10770 32562 10782
rect 39678 10834 39730 10846
rect 39678 10770 39730 10782
rect 41134 10834 41186 10846
rect 41134 10770 41186 10782
rect 42254 10834 42306 10846
rect 42254 10770 42306 10782
rect 31950 10722 32002 10734
rect 35758 10722 35810 10734
rect 33058 10670 33070 10722
rect 33122 10670 33134 10722
rect 38770 10670 38782 10722
rect 38834 10670 38846 10722
rect 31950 10658 32002 10670
rect 35758 10658 35810 10670
rect 21422 10610 21474 10622
rect 34750 10610 34802 10622
rect 36766 10610 36818 10622
rect 21858 10558 21870 10610
rect 21922 10558 21934 10610
rect 27010 10558 27022 10610
rect 27074 10558 27086 10610
rect 30370 10558 30382 10610
rect 30434 10558 30446 10610
rect 33394 10558 33406 10610
rect 33458 10558 33470 10610
rect 34290 10558 34302 10610
rect 34354 10558 34366 10610
rect 35522 10558 35534 10610
rect 35586 10558 35598 10610
rect 36642 10558 36654 10610
rect 36706 10558 36718 10610
rect 37202 10558 37214 10610
rect 37266 10558 37278 10610
rect 38322 10558 38334 10610
rect 38386 10558 38398 10610
rect 46498 10558 46510 10610
rect 46562 10558 46574 10610
rect 21422 10546 21474 10558
rect 34750 10546 34802 10558
rect 36766 10546 36818 10558
rect 31614 10498 31666 10510
rect 41918 10498 41970 10510
rect 20962 10446 20974 10498
rect 21026 10446 21038 10498
rect 22530 10446 22542 10498
rect 22594 10446 22606 10498
rect 24658 10446 24670 10498
rect 24722 10446 24734 10498
rect 27794 10446 27806 10498
rect 27858 10446 27870 10498
rect 29922 10446 29934 10498
rect 29986 10446 29998 10498
rect 30706 10446 30718 10498
rect 30770 10446 30782 10498
rect 37650 10446 37662 10498
rect 37714 10446 37726 10498
rect 31614 10434 31666 10446
rect 41918 10434 41970 10446
rect 42366 10498 42418 10510
rect 44818 10446 44830 10498
rect 44882 10446 44894 10498
rect 42366 10434 42418 10446
rect 31502 10386 31554 10398
rect 34066 10334 34078 10386
rect 34130 10334 34142 10386
rect 36194 10334 36206 10386
rect 36258 10334 36270 10386
rect 31502 10322 31554 10334
rect 1344 10218 58576 10252
rect 1344 10166 4478 10218
rect 4530 10166 4582 10218
rect 4634 10166 4686 10218
rect 4738 10166 35198 10218
rect 35250 10166 35302 10218
rect 35354 10166 35406 10218
rect 35458 10166 58576 10218
rect 1344 10132 58576 10166
rect 31602 9998 31614 10050
rect 31666 9998 31678 10050
rect 36430 9938 36482 9950
rect 44382 9938 44434 9950
rect 25106 9886 25118 9938
rect 25170 9886 25182 9938
rect 28354 9886 28366 9938
rect 28418 9886 28430 9938
rect 31042 9886 31054 9938
rect 31106 9886 31118 9938
rect 35970 9886 35982 9938
rect 36034 9886 36046 9938
rect 37426 9886 37438 9938
rect 37490 9886 37502 9938
rect 38546 9886 38558 9938
rect 38610 9886 38622 9938
rect 42242 9886 42254 9938
rect 42306 9886 42318 9938
rect 43026 9886 43038 9938
rect 43090 9886 43102 9938
rect 47730 9886 47742 9938
rect 47794 9886 47806 9938
rect 36430 9874 36482 9886
rect 44382 9874 44434 9886
rect 32062 9826 32114 9838
rect 36990 9826 37042 9838
rect 42590 9826 42642 9838
rect 22194 9774 22206 9826
rect 22258 9774 22270 9826
rect 25442 9774 25454 9826
rect 25506 9774 25518 9826
rect 30482 9774 30494 9826
rect 30546 9774 30558 9826
rect 30706 9774 30718 9826
rect 30770 9774 30782 9826
rect 31266 9774 31278 9826
rect 31330 9774 31342 9826
rect 32498 9774 32510 9826
rect 32562 9774 32574 9826
rect 33170 9774 33182 9826
rect 33234 9774 33246 9826
rect 38882 9774 38894 9826
rect 38946 9774 38958 9826
rect 39330 9774 39342 9826
rect 39394 9774 39406 9826
rect 44818 9774 44830 9826
rect 44882 9774 44894 9826
rect 32062 9762 32114 9774
rect 36990 9762 37042 9774
rect 42590 9762 42642 9774
rect 22978 9662 22990 9714
rect 23042 9662 23054 9714
rect 26226 9662 26238 9714
rect 26290 9662 26302 9714
rect 33842 9662 33854 9714
rect 33906 9662 33918 9714
rect 40114 9662 40126 9714
rect 40178 9662 40190 9714
rect 45602 9662 45614 9714
rect 45666 9662 45678 9714
rect 21646 9602 21698 9614
rect 21646 9538 21698 9550
rect 29710 9602 29762 9614
rect 29710 9538 29762 9550
rect 38110 9602 38162 9614
rect 38110 9538 38162 9550
rect 1344 9434 58576 9468
rect 1344 9382 19838 9434
rect 19890 9382 19942 9434
rect 19994 9382 20046 9434
rect 20098 9382 50558 9434
rect 50610 9382 50662 9434
rect 50714 9382 50766 9434
rect 50818 9382 58576 9434
rect 1344 9348 58576 9382
rect 22878 9266 22930 9278
rect 22878 9202 22930 9214
rect 24446 9266 24498 9278
rect 24446 9202 24498 9214
rect 32622 9266 32674 9278
rect 32622 9202 32674 9214
rect 38782 9266 38834 9278
rect 38782 9202 38834 9214
rect 39230 9266 39282 9278
rect 39230 9202 39282 9214
rect 40238 9266 40290 9278
rect 40238 9202 40290 9214
rect 40910 9266 40962 9278
rect 40910 9202 40962 9214
rect 45614 9266 45666 9278
rect 45614 9202 45666 9214
rect 46622 9266 46674 9278
rect 46622 9202 46674 9214
rect 22990 9154 23042 9166
rect 22990 9090 23042 9102
rect 24558 9154 24610 9166
rect 39678 9154 39730 9166
rect 25330 9102 25342 9154
rect 25394 9102 25406 9154
rect 30818 9102 30830 9154
rect 30882 9102 30894 9154
rect 24558 9090 24610 9102
rect 39678 9090 39730 9102
rect 40350 9154 40402 9166
rect 40350 9090 40402 9102
rect 45502 9154 45554 9166
rect 45502 9090 45554 9102
rect 23886 9042 23938 9054
rect 23426 8990 23438 9042
rect 23490 8990 23502 9042
rect 25778 8990 25790 9042
rect 25842 8990 25854 9042
rect 26562 8990 26574 9042
rect 26626 8990 26638 9042
rect 27794 8990 27806 9042
rect 27858 8990 27870 9042
rect 31602 8990 31614 9042
rect 31666 8990 31678 9042
rect 38322 8990 38334 9042
rect 38386 8990 38398 9042
rect 42354 8990 42366 9042
rect 42418 8990 42430 9042
rect 23886 8978 23938 8990
rect 41470 8930 41522 8942
rect 46062 8930 46114 8942
rect 26226 8878 26238 8930
rect 26290 8878 26302 8930
rect 27906 8878 27918 8930
rect 27970 8878 27982 8930
rect 28690 8878 28702 8930
rect 28754 8878 28766 8930
rect 36306 8878 36318 8930
rect 36370 8878 36382 8930
rect 43026 8878 43038 8930
rect 43090 8878 43102 8930
rect 45154 8878 45166 8930
rect 45218 8878 45230 8930
rect 41470 8866 41522 8878
rect 46062 8866 46114 8878
rect 39566 8818 39618 8830
rect 26562 8766 26574 8818
rect 26626 8766 26638 8818
rect 39566 8754 39618 8766
rect 45950 8818 46002 8830
rect 45950 8754 46002 8766
rect 1344 8650 58576 8684
rect 1344 8598 4478 8650
rect 4530 8598 4582 8650
rect 4634 8598 4686 8650
rect 4738 8598 35198 8650
rect 35250 8598 35302 8650
rect 35354 8598 35406 8650
rect 35458 8598 58576 8650
rect 1344 8564 58576 8598
rect 26462 8482 26514 8494
rect 26462 8418 26514 8430
rect 33966 8482 34018 8494
rect 42466 8430 42478 8482
rect 42530 8430 42542 8482
rect 33966 8418 34018 8430
rect 24222 8370 24274 8382
rect 24222 8306 24274 8318
rect 26574 8370 26626 8382
rect 26574 8306 26626 8318
rect 28030 8370 28082 8382
rect 28030 8306 28082 8318
rect 28142 8370 28194 8382
rect 34078 8370 34130 8382
rect 31490 8318 31502 8370
rect 31554 8318 31566 8370
rect 33618 8318 33630 8370
rect 33682 8318 33694 8370
rect 28142 8306 28194 8318
rect 34078 8306 34130 8318
rect 36318 8370 36370 8382
rect 40686 8370 40738 8382
rect 39890 8318 39902 8370
rect 39954 8318 39966 8370
rect 42690 8318 42702 8370
rect 42754 8318 42766 8370
rect 45714 8318 45726 8370
rect 45778 8318 45790 8370
rect 47842 8318 47854 8370
rect 47906 8318 47918 8370
rect 36318 8306 36370 8318
rect 40686 8306 40738 8318
rect 30818 8206 30830 8258
rect 30882 8206 30894 8258
rect 36978 8206 36990 8258
rect 37042 8206 37054 8258
rect 41794 8206 41806 8258
rect 41858 8206 41870 8258
rect 42354 8206 42366 8258
rect 42418 8206 42430 8258
rect 42914 8206 42926 8258
rect 42978 8206 42990 8258
rect 43810 8206 43822 8258
rect 43874 8206 43886 8258
rect 44930 8206 44942 8258
rect 44994 8206 45006 8258
rect 36430 8146 36482 8158
rect 44270 8146 44322 8158
rect 37762 8094 37774 8146
rect 37826 8094 37838 8146
rect 36430 8082 36482 8094
rect 44270 8082 44322 8094
rect 1344 7866 58576 7900
rect 1344 7814 19838 7866
rect 19890 7814 19942 7866
rect 19994 7814 20046 7866
rect 20098 7814 50558 7866
rect 50610 7814 50662 7866
rect 50714 7814 50766 7866
rect 50818 7814 58576 7866
rect 1344 7780 58576 7814
rect 42254 7698 42306 7710
rect 42254 7634 42306 7646
rect 45726 7698 45778 7710
rect 45726 7634 45778 7646
rect 39554 7534 39566 7586
rect 39618 7534 39630 7586
rect 40338 7422 40350 7474
rect 40402 7422 40414 7474
rect 42914 7422 42926 7474
rect 42978 7422 42990 7474
rect 43362 7422 43374 7474
rect 43426 7422 43438 7474
rect 43810 7422 43822 7474
rect 43874 7422 43886 7474
rect 44706 7422 44718 7474
rect 44770 7422 44782 7474
rect 42142 7362 42194 7374
rect 37426 7310 37438 7362
rect 37490 7310 37502 7362
rect 43698 7310 43710 7362
rect 43762 7310 43774 7362
rect 45154 7310 45166 7362
rect 45218 7310 45230 7362
rect 42142 7298 42194 7310
rect 43138 7198 43150 7250
rect 43202 7198 43214 7250
rect 1344 7082 58576 7116
rect 1344 7030 4478 7082
rect 4530 7030 4582 7082
rect 4634 7030 4686 7082
rect 4738 7030 35198 7082
rect 35250 7030 35302 7082
rect 35354 7030 35406 7082
rect 35458 7030 58576 7082
rect 1344 6996 58576 7030
rect 1344 6298 58576 6332
rect 1344 6246 19838 6298
rect 19890 6246 19942 6298
rect 19994 6246 20046 6298
rect 20098 6246 50558 6298
rect 50610 6246 50662 6298
rect 50714 6246 50766 6298
rect 50818 6246 58576 6298
rect 1344 6212 58576 6246
rect 42590 6130 42642 6142
rect 42590 6066 42642 6078
rect 45614 6018 45666 6030
rect 45614 5954 45666 5966
rect 43362 5854 43374 5906
rect 43426 5854 43438 5906
rect 43586 5854 43598 5906
rect 43650 5854 43662 5906
rect 44482 5854 44494 5906
rect 44546 5854 44558 5906
rect 45266 5854 45278 5906
rect 45330 5854 45342 5906
rect 29598 5794 29650 5806
rect 43810 5742 43822 5794
rect 43874 5742 43886 5794
rect 29598 5730 29650 5742
rect 45042 5630 45054 5682
rect 45106 5630 45118 5682
rect 1344 5514 58576 5548
rect 1344 5462 4478 5514
rect 4530 5462 4582 5514
rect 4634 5462 4686 5514
rect 4738 5462 35198 5514
rect 35250 5462 35302 5514
rect 35354 5462 35406 5514
rect 35458 5462 58576 5514
rect 1344 5428 58576 5462
rect 28702 5122 28754 5134
rect 28702 5058 28754 5070
rect 29150 5122 29202 5134
rect 30034 5070 30046 5122
rect 30098 5070 30110 5122
rect 29150 5058 29202 5070
rect 29486 5010 29538 5022
rect 29486 4946 29538 4958
rect 29822 5010 29874 5022
rect 29822 4946 29874 4958
rect 1344 4730 58576 4764
rect 1344 4678 19838 4730
rect 19890 4678 19942 4730
rect 19994 4678 20046 4730
rect 20098 4678 50558 4730
rect 50610 4678 50662 4730
rect 50714 4678 50766 4730
rect 50818 4678 58576 4730
rect 1344 4644 58576 4678
rect 26910 4562 26962 4574
rect 26910 4498 26962 4510
rect 30830 4562 30882 4574
rect 30830 4498 30882 4510
rect 30494 4338 30546 4350
rect 27346 4286 27358 4338
rect 27410 4286 27422 4338
rect 30494 4274 30546 4286
rect 16830 4226 16882 4238
rect 16830 4162 16882 4174
rect 18398 4226 18450 4238
rect 18398 4162 18450 4174
rect 19070 4226 19122 4238
rect 19070 4162 19122 4174
rect 19742 4226 19794 4238
rect 19742 4162 19794 4174
rect 20862 4226 20914 4238
rect 20862 4162 20914 4174
rect 23550 4226 23602 4238
rect 23550 4162 23602 4174
rect 24334 4226 24386 4238
rect 24334 4162 24386 4174
rect 24670 4226 24722 4238
rect 24670 4162 24722 4174
rect 30270 4226 30322 4238
rect 30270 4162 30322 4174
rect 31390 4226 31442 4238
rect 31390 4162 31442 4174
rect 33630 4226 33682 4238
rect 33630 4162 33682 4174
rect 34302 4226 34354 4238
rect 34302 4162 34354 4174
rect 36430 4226 36482 4238
rect 36430 4162 36482 4174
rect 37102 4226 37154 4238
rect 37102 4162 37154 4174
rect 37774 4226 37826 4238
rect 37774 4162 37826 4174
rect 38446 4226 38498 4238
rect 38446 4162 38498 4174
rect 39678 4226 39730 4238
rect 39678 4162 39730 4174
rect 40350 4226 40402 4238
rect 40350 4162 40402 4174
rect 41134 4226 41186 4238
rect 41134 4162 41186 4174
rect 43374 4226 43426 4238
rect 43374 4162 43426 4174
rect 44046 4226 44098 4238
rect 44046 4162 44098 4174
rect 28142 4114 28194 4126
rect 24210 4062 24222 4114
rect 24274 4111 24286 4114
rect 24658 4111 24670 4114
rect 24274 4065 24670 4111
rect 24274 4062 24286 4065
rect 24658 4062 24670 4065
rect 24722 4062 24734 4114
rect 28142 4050 28194 4062
rect 1344 3946 58576 3980
rect 1344 3894 4478 3946
rect 4530 3894 4582 3946
rect 4634 3894 4686 3946
rect 4738 3894 35198 3946
rect 35250 3894 35302 3946
rect 35354 3894 35406 3946
rect 35458 3894 58576 3946
rect 1344 3860 58576 3894
rect 29374 3666 29426 3678
rect 29374 3602 29426 3614
rect 27246 3554 27298 3566
rect 33854 3554 33906 3566
rect 16258 3502 16270 3554
rect 16322 3502 16334 3554
rect 17266 3502 17278 3554
rect 17330 3502 17342 3554
rect 17938 3502 17950 3554
rect 18002 3502 18014 3554
rect 18610 3502 18622 3554
rect 18674 3502 18686 3554
rect 23202 3502 23214 3554
rect 23266 3502 23278 3554
rect 23874 3502 23886 3554
rect 23938 3502 23950 3554
rect 26002 3502 26014 3554
rect 26066 3502 26078 3554
rect 27570 3502 27582 3554
rect 27634 3502 27646 3554
rect 28354 3502 28366 3554
rect 28418 3502 28430 3554
rect 31490 3502 31502 3554
rect 31554 3502 31566 3554
rect 27246 3490 27298 3502
rect 33854 3490 33906 3502
rect 34526 3554 34578 3566
rect 34526 3490 34578 3502
rect 36654 3554 36706 3566
rect 36654 3490 36706 3502
rect 37326 3554 37378 3566
rect 38210 3502 38222 3554
rect 38274 3502 38286 3554
rect 37326 3490 37378 3502
rect 12686 3442 12738 3454
rect 12686 3378 12738 3390
rect 13134 3442 13186 3454
rect 13134 3378 13186 3390
rect 13470 3442 13522 3454
rect 13470 3378 13522 3390
rect 15822 3442 15874 3454
rect 15822 3378 15874 3390
rect 16046 3442 16098 3454
rect 16046 3378 16098 3390
rect 17054 3442 17106 3454
rect 17054 3378 17106 3390
rect 18174 3442 18226 3454
rect 18174 3378 18226 3390
rect 18846 3442 18898 3454
rect 18846 3378 18898 3390
rect 19182 3442 19234 3454
rect 19182 3378 19234 3390
rect 19518 3442 19570 3454
rect 19518 3378 19570 3390
rect 19854 3442 19906 3454
rect 19854 3378 19906 3390
rect 20190 3442 20242 3454
rect 20190 3378 20242 3390
rect 21086 3442 21138 3454
rect 21086 3378 21138 3390
rect 21422 3442 21474 3454
rect 21422 3378 21474 3390
rect 21870 3442 21922 3454
rect 21870 3378 21922 3390
rect 22990 3442 23042 3454
rect 22990 3378 23042 3390
rect 23662 3442 23714 3454
rect 23662 3378 23714 3390
rect 24558 3442 24610 3454
rect 24558 3378 24610 3390
rect 24894 3442 24946 3454
rect 24894 3378 24946 3390
rect 25566 3442 25618 3454
rect 25566 3378 25618 3390
rect 25790 3442 25842 3454
rect 25790 3378 25842 3390
rect 26798 3442 26850 3454
rect 26798 3378 26850 3390
rect 27806 3442 27858 3454
rect 27806 3378 27858 3390
rect 31278 3442 31330 3454
rect 31278 3378 31330 3390
rect 32958 3442 33010 3454
rect 32958 3378 33010 3390
rect 33182 3442 33234 3454
rect 33182 3378 33234 3390
rect 33518 3442 33570 3454
rect 33518 3378 33570 3390
rect 34190 3442 34242 3454
rect 34190 3378 34242 3390
rect 34862 3442 34914 3454
rect 34862 3378 34914 3390
rect 35534 3442 35586 3454
rect 35534 3378 35586 3390
rect 35982 3442 36034 3454
rect 35982 3378 36034 3390
rect 36318 3442 36370 3454
rect 36318 3378 36370 3390
rect 36990 3442 37042 3454
rect 36990 3378 37042 3390
rect 37662 3442 37714 3454
rect 37662 3378 37714 3390
rect 37998 3442 38050 3454
rect 37998 3378 38050 3390
rect 38670 3442 38722 3454
rect 38670 3378 38722 3390
rect 39006 3442 39058 3454
rect 39006 3378 39058 3390
rect 39902 3442 39954 3454
rect 39902 3378 39954 3390
rect 40238 3442 40290 3454
rect 40238 3378 40290 3390
rect 40574 3442 40626 3454
rect 40574 3378 40626 3390
rect 40910 3442 40962 3454
rect 40910 3378 40962 3390
rect 41246 3442 41298 3454
rect 41246 3378 41298 3390
rect 41582 3442 41634 3454
rect 41582 3378 41634 3390
rect 42366 3442 42418 3454
rect 42366 3378 42418 3390
rect 42590 3442 42642 3454
rect 42590 3378 42642 3390
rect 42926 3442 42978 3454
rect 42926 3378 42978 3390
rect 43598 3442 43650 3454
rect 43598 3378 43650 3390
rect 43934 3442 43986 3454
rect 43934 3378 43986 3390
rect 44270 3442 44322 3454
rect 44270 3378 44322 3390
rect 44606 3442 44658 3454
rect 44606 3378 44658 3390
rect 1344 3162 58576 3196
rect 1344 3110 19838 3162
rect 19890 3110 19942 3162
rect 19994 3110 20046 3162
rect 20098 3110 50558 3162
rect 50610 3110 50662 3162
rect 50714 3110 50766 3162
rect 50818 3110 58576 3162
rect 1344 3076 58576 3110
<< via1 >>
rect 19838 76806 19890 76858
rect 19942 76806 19994 76858
rect 20046 76806 20098 76858
rect 50558 76806 50610 76858
rect 50662 76806 50714 76858
rect 50766 76806 50818 76858
rect 4478 76022 4530 76074
rect 4582 76022 4634 76074
rect 4686 76022 4738 76074
rect 35198 76022 35250 76074
rect 35302 76022 35354 76074
rect 35406 76022 35458 76074
rect 19838 75238 19890 75290
rect 19942 75238 19994 75290
rect 20046 75238 20098 75290
rect 50558 75238 50610 75290
rect 50662 75238 50714 75290
rect 50766 75238 50818 75290
rect 4478 74454 4530 74506
rect 4582 74454 4634 74506
rect 4686 74454 4738 74506
rect 35198 74454 35250 74506
rect 35302 74454 35354 74506
rect 35406 74454 35458 74506
rect 19838 73670 19890 73722
rect 19942 73670 19994 73722
rect 20046 73670 20098 73722
rect 50558 73670 50610 73722
rect 50662 73670 50714 73722
rect 50766 73670 50818 73722
rect 4478 72886 4530 72938
rect 4582 72886 4634 72938
rect 4686 72886 4738 72938
rect 35198 72886 35250 72938
rect 35302 72886 35354 72938
rect 35406 72886 35458 72938
rect 19838 72102 19890 72154
rect 19942 72102 19994 72154
rect 20046 72102 20098 72154
rect 50558 72102 50610 72154
rect 50662 72102 50714 72154
rect 50766 72102 50818 72154
rect 40238 71934 40290 71986
rect 39118 71822 39170 71874
rect 39902 71710 39954 71762
rect 36990 71598 37042 71650
rect 40350 71598 40402 71650
rect 40910 71598 40962 71650
rect 41022 71486 41074 71538
rect 4478 71318 4530 71370
rect 4582 71318 4634 71370
rect 4686 71318 4738 71370
rect 35198 71318 35250 71370
rect 35302 71318 35354 71370
rect 35406 71318 35458 71370
rect 34414 71038 34466 71090
rect 31614 70926 31666 70978
rect 41918 70926 41970 70978
rect 32286 70814 32338 70866
rect 34862 70814 34914 70866
rect 37214 70814 37266 70866
rect 34750 70702 34802 70754
rect 42702 70702 42754 70754
rect 19838 70534 19890 70586
rect 19942 70534 19994 70586
rect 20046 70534 20098 70586
rect 50558 70534 50610 70586
rect 50662 70534 50714 70586
rect 50766 70534 50818 70586
rect 31054 70366 31106 70418
rect 32398 70366 32450 70418
rect 40238 70366 40290 70418
rect 33966 70254 34018 70306
rect 41694 70254 41746 70306
rect 27806 70142 27858 70194
rect 31166 70142 31218 70194
rect 33182 70142 33234 70194
rect 36430 70142 36482 70194
rect 39790 70142 39842 70194
rect 40126 70142 40178 70194
rect 40350 70142 40402 70194
rect 40910 70142 40962 70194
rect 23998 70030 24050 70082
rect 25454 70030 25506 70082
rect 25790 70030 25842 70082
rect 28590 70030 28642 70082
rect 30718 70030 30770 70082
rect 32510 70030 32562 70082
rect 36094 70030 36146 70082
rect 37214 70030 37266 70082
rect 39342 70030 39394 70082
rect 43822 70030 43874 70082
rect 23886 69918 23938 69970
rect 25902 69918 25954 69970
rect 4478 69750 4530 69802
rect 4582 69750 4634 69802
rect 4686 69750 4738 69802
rect 35198 69750 35250 69802
rect 35302 69750 35354 69802
rect 35406 69750 35458 69802
rect 31278 69582 31330 69634
rect 35646 69582 35698 69634
rect 36430 69582 36482 69634
rect 22878 69470 22930 69522
rect 25006 69470 25058 69522
rect 26126 69470 26178 69522
rect 28254 69470 28306 69522
rect 30942 69470 30994 69522
rect 32958 69470 33010 69522
rect 34302 69470 34354 69522
rect 38446 69470 38498 69522
rect 42590 69470 42642 69522
rect 22206 69358 22258 69410
rect 25342 69358 25394 69410
rect 30382 69358 30434 69410
rect 33406 69358 33458 69410
rect 34414 69358 34466 69410
rect 35310 69358 35362 69410
rect 39678 69358 39730 69410
rect 29038 69246 29090 69298
rect 29374 69246 29426 69298
rect 30606 69246 30658 69298
rect 31390 69246 31442 69298
rect 31838 69246 31890 69298
rect 34974 69246 35026 69298
rect 35534 69246 35586 69298
rect 36318 69246 36370 69298
rect 37550 69246 37602 69298
rect 39230 69246 39282 69298
rect 39342 69246 39394 69298
rect 40462 69246 40514 69298
rect 43710 69246 43762 69298
rect 45278 69246 45330 69298
rect 29262 69134 29314 69186
rect 29710 69134 29762 69186
rect 29822 69134 29874 69186
rect 29934 69134 29986 69186
rect 30830 69134 30882 69186
rect 31054 69134 31106 69186
rect 31614 69134 31666 69186
rect 32846 69134 32898 69186
rect 33070 69134 33122 69186
rect 33966 69134 34018 69186
rect 34190 69134 34242 69186
rect 34638 69134 34690 69186
rect 34750 69134 34802 69186
rect 35646 69134 35698 69186
rect 37214 69134 37266 69186
rect 37438 69134 37490 69186
rect 37662 69134 37714 69186
rect 38110 69134 38162 69186
rect 38334 69134 38386 69186
rect 38558 69134 38610 69186
rect 42926 69134 42978 69186
rect 43262 69134 43314 69186
rect 43598 69134 43650 69186
rect 44158 69134 44210 69186
rect 45390 69134 45442 69186
rect 19838 68966 19890 69018
rect 19942 68966 19994 69018
rect 20046 68966 20098 69018
rect 50558 68966 50610 69018
rect 50662 68966 50714 69018
rect 50766 68966 50818 69018
rect 24558 68798 24610 68850
rect 24670 68798 24722 68850
rect 33294 68798 33346 68850
rect 33518 68798 33570 68850
rect 37326 68798 37378 68850
rect 38110 68798 38162 68850
rect 38222 68798 38274 68850
rect 41358 68798 41410 68850
rect 41470 68798 41522 68850
rect 23774 68686 23826 68738
rect 27806 68686 27858 68738
rect 34414 68686 34466 68738
rect 35982 68686 36034 68738
rect 36430 68686 36482 68738
rect 36654 68686 36706 68738
rect 38782 68686 38834 68738
rect 39230 68686 39282 68738
rect 40350 68686 40402 68738
rect 41246 68686 41298 68738
rect 42366 68686 42418 68738
rect 22766 68574 22818 68626
rect 23326 68574 23378 68626
rect 23550 68574 23602 68626
rect 23998 68574 24050 68626
rect 24446 68574 24498 68626
rect 25454 68574 25506 68626
rect 32958 68574 33010 68626
rect 34750 68574 34802 68626
rect 35646 68574 35698 68626
rect 36318 68574 36370 68626
rect 36766 68574 36818 68626
rect 37102 68574 37154 68626
rect 37550 68574 37602 68626
rect 37886 68574 37938 68626
rect 38558 68574 38610 68626
rect 39118 68574 39170 68626
rect 39454 68574 39506 68626
rect 39790 68574 39842 68626
rect 40126 68574 40178 68626
rect 40910 68574 40962 68626
rect 45838 68574 45890 68626
rect 19854 68462 19906 68514
rect 21982 68462 22034 68514
rect 23886 68462 23938 68514
rect 33406 68462 33458 68514
rect 35310 68462 35362 68514
rect 37214 68462 37266 68514
rect 40014 68462 40066 68514
rect 4478 68182 4530 68234
rect 4582 68182 4634 68234
rect 4686 68182 4738 68234
rect 35198 68182 35250 68234
rect 35302 68182 35354 68234
rect 35406 68182 35458 68234
rect 21422 68014 21474 68066
rect 37438 68014 37490 68066
rect 40910 68014 40962 68066
rect 20750 67902 20802 67954
rect 24782 67902 24834 67954
rect 25678 67902 25730 67954
rect 29150 67902 29202 67954
rect 29262 67902 29314 67954
rect 30382 67902 30434 67954
rect 32510 67902 32562 67954
rect 41358 67902 41410 67954
rect 43486 67902 43538 67954
rect 44830 67902 44882 67954
rect 46958 67902 47010 67954
rect 21870 67790 21922 67842
rect 22542 67790 22594 67842
rect 22878 67790 22930 67842
rect 23438 67790 23490 67842
rect 25118 67790 25170 67842
rect 26126 67790 26178 67842
rect 28030 67790 28082 67842
rect 28254 67790 28306 67842
rect 29710 67790 29762 67842
rect 37550 67790 37602 67842
rect 40798 67790 40850 67842
rect 44158 67790 44210 67842
rect 47630 67790 47682 67842
rect 21310 67678 21362 67730
rect 21982 67678 22034 67730
rect 24894 67678 24946 67730
rect 36206 67678 36258 67730
rect 37438 67678 37490 67730
rect 38446 67678 38498 67730
rect 41022 67678 41074 67730
rect 22094 67566 22146 67618
rect 23102 67566 23154 67618
rect 23774 67566 23826 67618
rect 24446 67566 24498 67618
rect 24670 67566 24722 67618
rect 25566 67566 25618 67618
rect 25790 67566 25842 67618
rect 26238 67566 26290 67618
rect 26462 67566 26514 67618
rect 28590 67566 28642 67618
rect 33070 67566 33122 67618
rect 33406 67566 33458 67618
rect 35646 67566 35698 67618
rect 35870 67566 35922 67618
rect 38110 67566 38162 67618
rect 38782 67566 38834 67618
rect 40238 67566 40290 67618
rect 40574 67566 40626 67618
rect 19838 67398 19890 67450
rect 19942 67398 19994 67450
rect 20046 67398 20098 67450
rect 50558 67398 50610 67450
rect 50662 67398 50714 67450
rect 50766 67398 50818 67450
rect 20526 67230 20578 67282
rect 21982 67230 22034 67282
rect 22542 67230 22594 67282
rect 22878 67230 22930 67282
rect 29262 67230 29314 67282
rect 39678 67230 39730 67282
rect 21310 67118 21362 67170
rect 22654 67118 22706 67170
rect 23550 67118 23602 67170
rect 23998 67118 24050 67170
rect 24222 67118 24274 67170
rect 29150 67118 29202 67170
rect 29486 67118 29538 67170
rect 29710 67118 29762 67170
rect 30382 67118 30434 67170
rect 30494 67118 30546 67170
rect 31278 67118 31330 67170
rect 32062 67118 32114 67170
rect 41470 67118 41522 67170
rect 41806 67118 41858 67170
rect 42478 67118 42530 67170
rect 43262 67118 43314 67170
rect 43486 67118 43538 67170
rect 44494 67118 44546 67170
rect 45502 67118 45554 67170
rect 20302 67006 20354 67058
rect 21086 67006 21138 67058
rect 21422 67006 21474 67058
rect 21758 67006 21810 67058
rect 22318 67006 22370 67058
rect 23102 67006 23154 67058
rect 24334 67006 24386 67058
rect 30046 67006 30098 67058
rect 30606 67006 30658 67058
rect 30942 67006 30994 67058
rect 31502 67006 31554 67058
rect 41134 67006 41186 67058
rect 42030 67006 42082 67058
rect 42702 67006 42754 67058
rect 43038 67006 43090 67058
rect 43934 67006 43986 67058
rect 44046 67006 44098 67058
rect 44718 67006 44770 67058
rect 44942 67006 44994 67058
rect 45390 67006 45442 67058
rect 45614 67006 45666 67058
rect 15374 66894 15426 66946
rect 19854 66894 19906 66946
rect 21870 66894 21922 66946
rect 25678 66894 25730 66946
rect 26126 66894 26178 66946
rect 26462 66894 26514 66946
rect 27022 66894 27074 66946
rect 28702 66894 28754 66946
rect 34414 66894 34466 66946
rect 36766 66894 36818 66946
rect 40238 66894 40290 66946
rect 42814 66894 42866 66946
rect 43374 66894 43426 66946
rect 44606 66894 44658 66946
rect 15262 66782 15314 66834
rect 25678 66782 25730 66834
rect 26462 66782 26514 66834
rect 4478 66614 4530 66666
rect 4582 66614 4634 66666
rect 4686 66614 4738 66666
rect 35198 66614 35250 66666
rect 35302 66614 35354 66666
rect 35406 66614 35458 66666
rect 14030 66446 14082 66498
rect 22318 66446 22370 66498
rect 26126 66446 26178 66498
rect 31054 66446 31106 66498
rect 41134 66446 41186 66498
rect 43374 66446 43426 66498
rect 43934 66446 43986 66498
rect 17390 66334 17442 66386
rect 21422 66334 21474 66386
rect 25566 66334 25618 66386
rect 34526 66334 34578 66386
rect 48078 66334 48130 66386
rect 14478 66222 14530 66274
rect 19966 66222 20018 66274
rect 21646 66222 21698 66274
rect 21982 66222 22034 66274
rect 25790 66222 25842 66274
rect 26238 66222 26290 66274
rect 27806 66222 27858 66274
rect 28142 66222 28194 66274
rect 35198 66222 35250 66274
rect 35422 66222 35474 66274
rect 37326 66222 37378 66274
rect 37662 66222 37714 66274
rect 38670 66222 38722 66274
rect 41246 66222 41298 66274
rect 41582 66222 41634 66274
rect 42254 66222 42306 66274
rect 42702 66222 42754 66274
rect 44158 66222 44210 66274
rect 45166 66222 45218 66274
rect 13918 66110 13970 66162
rect 15262 66110 15314 66162
rect 24670 66110 24722 66162
rect 25454 66110 25506 66162
rect 26126 66110 26178 66162
rect 28366 66110 28418 66162
rect 30270 66110 30322 66162
rect 30606 66110 30658 66162
rect 30942 66110 30994 66162
rect 31054 66110 31106 66162
rect 33630 66110 33682 66162
rect 34078 66110 34130 66162
rect 36206 66110 36258 66162
rect 36430 66110 36482 66162
rect 36990 66110 37042 66162
rect 39902 66110 39954 66162
rect 41918 66110 41970 66162
rect 42478 66110 42530 66162
rect 43262 66110 43314 66162
rect 43598 66110 43650 66162
rect 45950 66110 46002 66162
rect 14030 65998 14082 66050
rect 20190 65998 20242 66050
rect 20638 65998 20690 66050
rect 21310 65998 21362 66050
rect 22206 65998 22258 66050
rect 24446 65998 24498 66050
rect 24782 65998 24834 66050
rect 25006 65998 25058 66050
rect 25230 65998 25282 66050
rect 27022 65998 27074 66050
rect 27246 65998 27298 66050
rect 27358 65998 27410 66050
rect 27470 65998 27522 66050
rect 27918 65998 27970 66050
rect 29374 65998 29426 66050
rect 30046 65998 30098 66050
rect 32734 65998 32786 66050
rect 33294 65998 33346 66050
rect 33518 65998 33570 66050
rect 33966 65998 34018 66050
rect 35758 65998 35810 66050
rect 36318 65998 36370 66050
rect 37326 65998 37378 66050
rect 39118 65998 39170 66050
rect 39230 65998 39282 66050
rect 39342 65998 39394 66050
rect 39566 65998 39618 66050
rect 39790 65998 39842 66050
rect 40350 65998 40402 66050
rect 41134 65998 41186 66050
rect 41694 65998 41746 66050
rect 43038 65998 43090 66050
rect 43822 65998 43874 66050
rect 19838 65830 19890 65882
rect 19942 65830 19994 65882
rect 20046 65830 20098 65882
rect 50558 65830 50610 65882
rect 50662 65830 50714 65882
rect 50766 65830 50818 65882
rect 16382 65662 16434 65714
rect 25790 65662 25842 65714
rect 43598 65662 43650 65714
rect 43822 65662 43874 65714
rect 44158 65662 44210 65714
rect 44382 65662 44434 65714
rect 45390 65662 45442 65714
rect 16494 65550 16546 65602
rect 18510 65550 18562 65602
rect 20750 65550 20802 65602
rect 23214 65550 23266 65602
rect 24222 65550 24274 65602
rect 27358 65550 27410 65602
rect 30270 65550 30322 65602
rect 32174 65550 32226 65602
rect 34190 65550 34242 65602
rect 43934 65550 43986 65602
rect 44494 65550 44546 65602
rect 45278 65550 45330 65602
rect 47518 65550 47570 65602
rect 9886 65438 9938 65490
rect 13134 65438 13186 65490
rect 16158 65438 16210 65490
rect 17390 65438 17442 65490
rect 17614 65438 17666 65490
rect 17726 65438 17778 65490
rect 17838 65438 17890 65490
rect 18062 65438 18114 65490
rect 18398 65438 18450 65490
rect 19966 65438 20018 65490
rect 23438 65438 23490 65490
rect 24446 65438 24498 65490
rect 25230 65438 25282 65490
rect 25566 65438 25618 65490
rect 26574 65438 26626 65490
rect 30046 65438 30098 65490
rect 30158 65438 30210 65490
rect 30718 65438 30770 65490
rect 31950 65438 32002 65490
rect 32510 65438 32562 65490
rect 32958 65438 33010 65490
rect 33406 65438 33458 65490
rect 33630 65438 33682 65490
rect 33966 65438 34018 65490
rect 34526 65438 34578 65490
rect 40238 65438 40290 65490
rect 41246 65438 41298 65490
rect 47854 65438 47906 65490
rect 10558 65326 10610 65378
rect 12686 65326 12738 65378
rect 13806 65326 13858 65378
rect 15934 65326 15986 65378
rect 22878 65326 22930 65378
rect 25678 65326 25730 65378
rect 26126 65326 26178 65378
rect 26238 65326 26290 65378
rect 29486 65326 29538 65378
rect 33518 65326 33570 65378
rect 34078 65326 34130 65378
rect 37438 65326 37490 65378
rect 41022 65326 41074 65378
rect 41806 65326 41858 65378
rect 42142 65326 42194 65378
rect 42590 65326 42642 65378
rect 43038 65326 43090 65378
rect 40910 65214 40962 65266
rect 41470 65214 41522 65266
rect 41806 65214 41858 65266
rect 42366 65214 42418 65266
rect 42590 65214 42642 65266
rect 4478 65046 4530 65098
rect 4582 65046 4634 65098
rect 4686 65046 4738 65098
rect 35198 65046 35250 65098
rect 35302 65046 35354 65098
rect 35406 65046 35458 65098
rect 26574 64878 26626 64930
rect 26910 64878 26962 64930
rect 29934 64878 29986 64930
rect 30942 64878 30994 64930
rect 34974 64878 35026 64930
rect 36430 64878 36482 64930
rect 41694 64878 41746 64930
rect 43038 64878 43090 64930
rect 43598 64878 43650 64930
rect 12910 64766 12962 64818
rect 13918 64766 13970 64818
rect 17502 64766 17554 64818
rect 20750 64766 20802 64818
rect 23774 64766 23826 64818
rect 25902 64766 25954 64818
rect 31950 64766 32002 64818
rect 34078 64766 34130 64818
rect 10110 64654 10162 64706
rect 13694 64654 13746 64706
rect 14254 64654 14306 64706
rect 14590 64654 14642 64706
rect 17950 64654 18002 64706
rect 21646 64654 21698 64706
rect 22990 64654 23042 64706
rect 27246 64654 27298 64706
rect 27470 64654 27522 64706
rect 27806 64654 27858 64706
rect 28030 64654 28082 64706
rect 29374 64654 29426 64706
rect 29822 64654 29874 64706
rect 31166 64654 31218 64706
rect 34638 64654 34690 64706
rect 35758 64654 35810 64706
rect 35870 64654 35922 64706
rect 37438 64654 37490 64706
rect 41134 64654 41186 64706
rect 42030 64654 42082 64706
rect 42702 64654 42754 64706
rect 44718 64654 44770 64706
rect 45166 64654 45218 64706
rect 10782 64542 10834 64594
rect 15374 64542 15426 64594
rect 18622 64542 18674 64594
rect 21310 64542 21362 64594
rect 21422 64542 21474 64594
rect 28142 64542 28194 64594
rect 28590 64542 28642 64594
rect 29150 64542 29202 64594
rect 34414 64542 34466 64594
rect 35982 64542 36034 64594
rect 37214 64542 37266 64594
rect 38222 64542 38274 64594
rect 41022 64542 41074 64594
rect 41246 64542 41298 64594
rect 42254 64542 42306 64594
rect 43038 64542 43090 64594
rect 44046 64542 44098 64594
rect 13806 64430 13858 64482
rect 14030 64430 14082 64482
rect 22766 64430 22818 64482
rect 26350 64430 26402 64482
rect 26462 64430 26514 64482
rect 29598 64430 29650 64482
rect 30158 64430 30210 64482
rect 30606 64430 30658 64482
rect 40462 64430 40514 64482
rect 42478 64430 42530 64482
rect 43598 64430 43650 64482
rect 43934 64430 43986 64482
rect 45278 64430 45330 64482
rect 45390 64430 45442 64482
rect 45950 64430 46002 64482
rect 46846 64430 46898 64482
rect 19838 64262 19890 64314
rect 19942 64262 19994 64314
rect 20046 64262 20098 64314
rect 50558 64262 50610 64314
rect 50662 64262 50714 64314
rect 50766 64262 50818 64314
rect 11678 64094 11730 64146
rect 11790 64094 11842 64146
rect 12798 64094 12850 64146
rect 14814 64094 14866 64146
rect 15598 64094 15650 64146
rect 16158 64094 16210 64146
rect 16270 64094 16322 64146
rect 16382 64094 16434 64146
rect 17950 64094 18002 64146
rect 19294 64094 19346 64146
rect 20302 64094 20354 64146
rect 22542 64094 22594 64146
rect 22990 64094 23042 64146
rect 26126 64094 26178 64146
rect 26574 64094 26626 64146
rect 28590 64094 28642 64146
rect 30382 64094 30434 64146
rect 31726 64094 31778 64146
rect 33518 64094 33570 64146
rect 33854 64094 33906 64146
rect 37774 64094 37826 64146
rect 37998 64094 38050 64146
rect 38670 64094 38722 64146
rect 38894 64094 38946 64146
rect 39566 64094 39618 64146
rect 41022 64094 41074 64146
rect 42478 64094 42530 64146
rect 47182 64094 47234 64146
rect 12462 63982 12514 64034
rect 13470 63982 13522 64034
rect 13918 63982 13970 64034
rect 14030 63982 14082 64034
rect 14926 63982 14978 64034
rect 15262 63982 15314 64034
rect 23550 63982 23602 64034
rect 26686 63982 26738 64034
rect 28814 63982 28866 64034
rect 28926 63982 28978 64034
rect 29374 63982 29426 64034
rect 31614 63982 31666 64034
rect 31950 63982 32002 64034
rect 32510 63982 32562 64034
rect 33630 63982 33682 64034
rect 34078 63982 34130 64034
rect 34190 63982 34242 64034
rect 41918 63982 41970 64034
rect 42590 63982 42642 64034
rect 43822 63982 43874 64034
rect 47630 63982 47682 64034
rect 48974 63982 49026 64034
rect 11454 63870 11506 63922
rect 11566 63870 11618 63922
rect 12014 63870 12066 63922
rect 12574 63870 12626 63922
rect 13022 63870 13074 63922
rect 13358 63870 13410 63922
rect 13694 63870 13746 63922
rect 16046 63870 16098 63922
rect 16606 63870 16658 63922
rect 17390 63870 17442 63922
rect 20190 63870 20242 63922
rect 20526 63870 20578 63922
rect 22318 63870 22370 63922
rect 22654 63870 22706 63922
rect 23774 63870 23826 63922
rect 24222 63870 24274 63922
rect 24446 63870 24498 63922
rect 25454 63870 25506 63922
rect 25902 63870 25954 63922
rect 26014 63870 26066 63922
rect 27694 63870 27746 63922
rect 28366 63870 28418 63922
rect 29598 63870 29650 63922
rect 30046 63870 30098 63922
rect 30494 63870 30546 63922
rect 32174 63870 32226 63922
rect 33182 63870 33234 63922
rect 33294 63870 33346 63922
rect 37438 63870 37490 63922
rect 38334 63870 38386 63922
rect 39342 63870 39394 63922
rect 40126 63870 40178 63922
rect 40798 63870 40850 63922
rect 41134 63870 41186 63922
rect 41358 63870 41410 63922
rect 42030 63870 42082 63922
rect 42254 63870 42306 63922
rect 43150 63870 43202 63922
rect 47070 63870 47122 63922
rect 47854 63870 47906 63922
rect 48302 63870 48354 63922
rect 49422 63870 49474 63922
rect 12462 63758 12514 63810
rect 17502 63758 17554 63810
rect 19406 63758 19458 63810
rect 22206 63758 22258 63810
rect 24334 63758 24386 63810
rect 27582 63758 27634 63810
rect 29486 63758 29538 63810
rect 30382 63758 30434 63810
rect 32398 63758 32450 63810
rect 34526 63758 34578 63810
rect 36654 63758 36706 63810
rect 37886 63758 37938 63810
rect 14814 63646 14866 63698
rect 21982 63646 22034 63698
rect 22206 63646 22258 63698
rect 23326 63646 23378 63698
rect 26574 63646 26626 63698
rect 38782 63758 38834 63810
rect 39902 63758 39954 63810
rect 45950 63758 46002 63810
rect 46398 63758 46450 63810
rect 47742 63758 47794 63810
rect 27806 63646 27858 63698
rect 28030 63646 28082 63698
rect 28366 63646 28418 63698
rect 41918 63646 41970 63698
rect 47182 63646 47234 63698
rect 48862 63646 48914 63698
rect 4478 63478 4530 63530
rect 4582 63478 4634 63530
rect 4686 63478 4738 63530
rect 35198 63478 35250 63530
rect 35302 63478 35354 63530
rect 35406 63478 35458 63530
rect 12574 63310 12626 63362
rect 24558 63310 24610 63362
rect 44382 63310 44434 63362
rect 12686 63198 12738 63250
rect 19854 63198 19906 63250
rect 24222 63198 24274 63250
rect 25118 63198 25170 63250
rect 31166 63198 31218 63250
rect 35982 63198 36034 63250
rect 38334 63198 38386 63250
rect 38894 63198 38946 63250
rect 39454 63198 39506 63250
rect 40238 63198 40290 63250
rect 18734 63086 18786 63138
rect 19182 63086 19234 63138
rect 19742 63086 19794 63138
rect 21982 63086 22034 63138
rect 22094 63086 22146 63138
rect 22766 63086 22818 63138
rect 22990 63086 23042 63138
rect 23550 63086 23602 63138
rect 24334 63086 24386 63138
rect 25006 63086 25058 63138
rect 25230 63086 25282 63138
rect 25566 63086 25618 63138
rect 34750 63086 34802 63138
rect 35870 63086 35922 63138
rect 36094 63086 36146 63138
rect 37214 63086 37266 63138
rect 37886 63086 37938 63138
rect 38110 63086 38162 63138
rect 40014 63086 40066 63138
rect 43150 63086 43202 63138
rect 48750 63086 48802 63138
rect 11790 62974 11842 63026
rect 14254 62974 14306 63026
rect 21646 62974 21698 63026
rect 22430 62974 22482 63026
rect 23102 62974 23154 63026
rect 37102 62974 37154 63026
rect 38446 62974 38498 63026
rect 42366 62974 42418 63026
rect 43822 62974 43874 63026
rect 45390 62974 45442 63026
rect 11454 62862 11506 62914
rect 11678 62862 11730 62914
rect 19966 62862 20018 62914
rect 20190 62862 20242 62914
rect 22318 62862 22370 62914
rect 26014 62862 26066 62914
rect 28478 62862 28530 62914
rect 35198 62862 35250 62914
rect 35646 62862 35698 62914
rect 36878 62862 36930 62914
rect 39342 62862 39394 62914
rect 39566 62862 39618 62914
rect 44046 62862 44098 62914
rect 44270 62862 44322 62914
rect 19838 62694 19890 62746
rect 19942 62694 19994 62746
rect 20046 62694 20098 62746
rect 50558 62694 50610 62746
rect 50662 62694 50714 62746
rect 50766 62694 50818 62746
rect 12686 62526 12738 62578
rect 12910 62526 12962 62578
rect 15822 62526 15874 62578
rect 16046 62526 16098 62578
rect 17950 62526 18002 62578
rect 24222 62526 24274 62578
rect 24558 62526 24610 62578
rect 24670 62526 24722 62578
rect 33070 62526 33122 62578
rect 33294 62526 33346 62578
rect 34078 62526 34130 62578
rect 36542 62526 36594 62578
rect 37662 62526 37714 62578
rect 38110 62526 38162 62578
rect 39118 62526 39170 62578
rect 41022 62526 41074 62578
rect 41134 62526 41186 62578
rect 41694 62526 41746 62578
rect 42030 62526 42082 62578
rect 42590 62526 42642 62578
rect 43262 62526 43314 62578
rect 43822 62526 43874 62578
rect 44606 62526 44658 62578
rect 16718 62414 16770 62466
rect 16830 62414 16882 62466
rect 18622 62414 18674 62466
rect 28142 62414 28194 62466
rect 28254 62414 28306 62466
rect 33518 62414 33570 62466
rect 34302 62414 34354 62466
rect 39454 62414 39506 62466
rect 40350 62414 40402 62466
rect 41358 62414 41410 62466
rect 41806 62414 41858 62466
rect 43598 62414 43650 62466
rect 44046 62414 44098 62466
rect 44158 62414 44210 62466
rect 9662 62302 9714 62354
rect 13022 62302 13074 62354
rect 15710 62302 15762 62354
rect 16270 62302 16322 62354
rect 16494 62302 16546 62354
rect 18398 62302 18450 62354
rect 24222 62302 24274 62354
rect 28478 62302 28530 62354
rect 28814 62302 28866 62354
rect 29486 62302 29538 62354
rect 33854 62302 33906 62354
rect 35198 62302 35250 62354
rect 39678 62302 39730 62354
rect 40014 62302 40066 62354
rect 40910 62302 40962 62354
rect 42366 62302 42418 62354
rect 42814 62302 42866 62354
rect 45390 62302 45442 62354
rect 48750 62302 48802 62354
rect 10334 62190 10386 62242
rect 12462 62190 12514 62242
rect 15934 62190 15986 62242
rect 21310 62190 21362 62242
rect 25342 62190 25394 62242
rect 26014 62190 26066 62242
rect 27470 62190 27522 62242
rect 27918 62190 27970 62242
rect 31614 62190 31666 62242
rect 32286 62190 32338 62242
rect 34750 62190 34802 62242
rect 35646 62190 35698 62242
rect 36094 62190 36146 62242
rect 37326 62190 37378 62242
rect 39902 62190 39954 62242
rect 46062 62190 46114 62242
rect 48190 62190 48242 62242
rect 50766 62190 50818 62242
rect 27134 62078 27186 62130
rect 27806 62078 27858 62130
rect 32958 62078 33010 62130
rect 33966 62078 34018 62130
rect 4478 61910 4530 61962
rect 4582 61910 4634 61962
rect 4686 61910 4738 61962
rect 35198 61910 35250 61962
rect 35302 61910 35354 61962
rect 35406 61910 35458 61962
rect 30494 61742 30546 61794
rect 40798 61742 40850 61794
rect 41134 61742 41186 61794
rect 41470 61742 41522 61794
rect 41806 61742 41858 61794
rect 42142 61742 42194 61794
rect 45726 61742 45778 61794
rect 9998 61630 10050 61682
rect 10558 61630 10610 61682
rect 15038 61630 15090 61682
rect 17166 61630 17218 61682
rect 20414 61630 20466 61682
rect 22094 61630 22146 61682
rect 24222 61630 24274 61682
rect 25118 61630 25170 61682
rect 31838 61630 31890 61682
rect 32398 61630 32450 61682
rect 33630 61630 33682 61682
rect 38110 61630 38162 61682
rect 40574 61630 40626 61682
rect 43598 61630 43650 61682
rect 45278 61630 45330 61682
rect 46286 61630 46338 61682
rect 48078 61630 48130 61682
rect 50206 61630 50258 61682
rect 10110 61518 10162 61570
rect 10446 61518 10498 61570
rect 10670 61518 10722 61570
rect 11118 61518 11170 61570
rect 11902 61518 11954 61570
rect 12126 61518 12178 61570
rect 14254 61518 14306 61570
rect 17614 61518 17666 61570
rect 21310 61518 21362 61570
rect 24558 61518 24610 61570
rect 25342 61518 25394 61570
rect 27470 61518 27522 61570
rect 27694 61518 27746 61570
rect 27918 61518 27970 61570
rect 28366 61518 28418 61570
rect 29038 61518 29090 61570
rect 29934 61518 29986 61570
rect 30830 61518 30882 61570
rect 31390 61518 31442 61570
rect 32174 61518 32226 61570
rect 32510 61518 32562 61570
rect 32734 61518 32786 61570
rect 33966 61518 34018 61570
rect 34638 61518 34690 61570
rect 35086 61518 35138 61570
rect 37550 61518 37602 61570
rect 38670 61518 38722 61570
rect 39902 61518 39954 61570
rect 40238 61518 40290 61570
rect 45950 61518 46002 61570
rect 46398 61518 46450 61570
rect 47294 61518 47346 61570
rect 50878 61518 50930 61570
rect 11454 61406 11506 61458
rect 12574 61406 12626 61458
rect 13918 61406 13970 61458
rect 18286 61406 18338 61458
rect 25678 61406 25730 61458
rect 26238 61406 26290 61458
rect 26350 61406 26402 61458
rect 29262 61406 29314 61458
rect 29374 61406 29426 61458
rect 29822 61406 29874 61458
rect 30046 61406 30098 61458
rect 31502 61406 31554 61458
rect 33742 61406 33794 61458
rect 37998 61406 38050 61458
rect 40126 61406 40178 61458
rect 42254 61406 42306 61458
rect 42702 61406 42754 61458
rect 44942 61406 44994 61458
rect 46174 61406 46226 61458
rect 10894 61294 10946 61346
rect 11678 61294 11730 61346
rect 11790 61294 11842 61346
rect 12910 61294 12962 61346
rect 13582 61294 13634 61346
rect 26574 61294 26626 61346
rect 26798 61294 26850 61346
rect 26910 61294 26962 61346
rect 27022 61294 27074 61346
rect 28142 61294 28194 61346
rect 35310 61294 35362 61346
rect 35758 61294 35810 61346
rect 36206 61294 36258 61346
rect 37326 61294 37378 61346
rect 39006 61294 39058 61346
rect 39342 61294 39394 61346
rect 41582 61294 41634 61346
rect 43150 61294 43202 61346
rect 44382 61294 44434 61346
rect 45166 61294 45218 61346
rect 45390 61294 45442 61346
rect 46958 61294 47010 61346
rect 50542 61294 50594 61346
rect 19838 61126 19890 61178
rect 19942 61126 19994 61178
rect 20046 61126 20098 61178
rect 50558 61126 50610 61178
rect 50662 61126 50714 61178
rect 50766 61126 50818 61178
rect 12798 60958 12850 61010
rect 14478 60958 14530 61010
rect 14814 60958 14866 61010
rect 18846 60958 18898 61010
rect 19630 60958 19682 61010
rect 20862 60958 20914 61010
rect 21758 60958 21810 61010
rect 22430 60958 22482 61010
rect 23102 60958 23154 61010
rect 24670 60958 24722 61010
rect 28926 60958 28978 61010
rect 30382 60958 30434 61010
rect 31502 60958 31554 61010
rect 41694 60958 41746 61010
rect 50318 60958 50370 61010
rect 10334 60846 10386 60898
rect 16046 60846 16098 60898
rect 16158 60846 16210 60898
rect 16830 60846 16882 60898
rect 18958 60846 19010 60898
rect 22206 60846 22258 60898
rect 22654 60846 22706 60898
rect 23214 60846 23266 60898
rect 28478 60846 28530 60898
rect 30270 60846 30322 60898
rect 30606 60846 30658 60898
rect 32062 60846 32114 60898
rect 48862 60846 48914 60898
rect 9550 60734 9602 60786
rect 13134 60734 13186 60786
rect 16606 60734 16658 60786
rect 17950 60734 18002 60786
rect 19518 60734 19570 60786
rect 19742 60734 19794 60786
rect 20190 60734 20242 60786
rect 20302 60734 20354 60786
rect 20638 60734 20690 60786
rect 21198 60734 21250 60786
rect 21534 60734 21586 60786
rect 22094 60734 22146 60786
rect 22990 60734 23042 60786
rect 24334 60734 24386 60786
rect 28142 60734 28194 60786
rect 28702 60734 28754 60786
rect 30158 60734 30210 60786
rect 32286 60734 32338 60786
rect 32510 60734 32562 60786
rect 32958 60734 33010 60786
rect 33742 60734 33794 60786
rect 34750 60734 34802 60786
rect 34974 60734 35026 60786
rect 35422 60734 35474 60786
rect 35758 60734 35810 60786
rect 38894 60734 38946 60786
rect 39118 60734 39170 60786
rect 39566 60734 39618 60786
rect 46174 60734 46226 60786
rect 46958 60734 47010 60786
rect 47518 60734 47570 60786
rect 49086 60734 49138 60786
rect 49870 60734 49922 60786
rect 12462 60622 12514 60674
rect 17502 60622 17554 60674
rect 21422 60622 21474 60674
rect 23998 60622 24050 60674
rect 25230 60622 25282 60674
rect 27358 60622 27410 60674
rect 28590 60622 28642 60674
rect 29710 60622 29762 60674
rect 31054 60622 31106 60674
rect 32398 60622 32450 60674
rect 33182 60622 33234 60674
rect 33630 60622 33682 60674
rect 34862 60622 34914 60674
rect 36430 60622 36482 60674
rect 38558 60622 38610 60674
rect 39006 60622 39058 60674
rect 40014 60622 40066 60674
rect 40350 60622 40402 60674
rect 41022 60622 41074 60674
rect 42366 60622 42418 60674
rect 43038 60622 43090 60674
rect 43262 60622 43314 60674
rect 45390 60622 45442 60674
rect 47406 60622 47458 60674
rect 48862 60622 48914 60674
rect 16046 60510 16098 60562
rect 17390 60510 17442 60562
rect 20526 60510 20578 60562
rect 47294 60510 47346 60562
rect 4478 60342 4530 60394
rect 4582 60342 4634 60394
rect 4686 60342 4738 60394
rect 35198 60342 35250 60394
rect 35302 60342 35354 60394
rect 35406 60342 35458 60394
rect 12126 60174 12178 60226
rect 26238 60174 26290 60226
rect 26574 60174 26626 60226
rect 28030 60174 28082 60226
rect 28366 60174 28418 60226
rect 36206 60174 36258 60226
rect 48078 60174 48130 60226
rect 48750 60174 48802 60226
rect 49086 60174 49138 60226
rect 49198 60174 49250 60226
rect 12238 60062 12290 60114
rect 23102 60062 23154 60114
rect 24334 60062 24386 60114
rect 29598 60062 29650 60114
rect 32846 60062 32898 60114
rect 34974 60062 35026 60114
rect 35982 60062 36034 60114
rect 38110 60062 38162 60114
rect 39566 60062 39618 60114
rect 46958 60062 47010 60114
rect 11454 59950 11506 60002
rect 15486 59950 15538 60002
rect 16046 59950 16098 60002
rect 19630 59950 19682 60002
rect 20526 59950 20578 60002
rect 22094 59950 22146 60002
rect 23662 59950 23714 60002
rect 23886 59950 23938 60002
rect 26014 59950 26066 60002
rect 26910 59950 26962 60002
rect 27134 59950 27186 60002
rect 28030 59950 28082 60002
rect 32174 59950 32226 60002
rect 37102 59950 37154 60002
rect 37326 59950 37378 60002
rect 37550 59950 37602 60002
rect 38222 59950 38274 60002
rect 39342 59950 39394 60002
rect 39790 59950 39842 60002
rect 40014 59950 40066 60002
rect 42030 59950 42082 60002
rect 42366 59950 42418 60002
rect 42590 59950 42642 60002
rect 42926 59950 42978 60002
rect 43710 59950 43762 60002
rect 46398 59950 46450 60002
rect 46734 59950 46786 60002
rect 47518 59950 47570 60002
rect 48862 59950 48914 60002
rect 11678 59838 11730 59890
rect 11790 59838 11842 59890
rect 16494 59838 16546 59890
rect 20750 59838 20802 59890
rect 21870 59838 21922 59890
rect 27246 59838 27298 59890
rect 30942 59838 30994 59890
rect 38558 59838 38610 59890
rect 40574 59838 40626 59890
rect 42254 59838 42306 59890
rect 43486 59838 43538 59890
rect 44830 59838 44882 59890
rect 45166 59838 45218 59890
rect 45502 59838 45554 59890
rect 45614 59838 45666 59890
rect 46958 59838 47010 59890
rect 47406 59838 47458 59890
rect 47630 59838 47682 59890
rect 15598 59726 15650 59778
rect 15710 59726 15762 59778
rect 15822 59726 15874 59778
rect 16382 59726 16434 59778
rect 20078 59726 20130 59778
rect 21534 59726 21586 59778
rect 22654 59726 22706 59778
rect 25230 59726 25282 59778
rect 25790 59726 25842 59778
rect 27694 59726 27746 59778
rect 31278 59726 31330 59778
rect 31838 59726 31890 59778
rect 35534 59726 35586 59778
rect 35646 59726 35698 59778
rect 35758 59726 35810 59778
rect 37438 59726 37490 59778
rect 39566 59726 39618 59778
rect 40238 59726 40290 59778
rect 40462 59726 40514 59778
rect 41022 59726 41074 59778
rect 41470 59726 41522 59778
rect 43150 59726 43202 59778
rect 43262 59726 43314 59778
rect 44046 59726 44098 59778
rect 46062 59726 46114 59778
rect 49758 59726 49810 59778
rect 50206 59726 50258 59778
rect 19838 59558 19890 59610
rect 19942 59558 19994 59610
rect 20046 59558 20098 59610
rect 50558 59558 50610 59610
rect 50662 59558 50714 59610
rect 50766 59558 50818 59610
rect 17502 59390 17554 59442
rect 18846 59390 18898 59442
rect 19070 59390 19122 59442
rect 19406 59390 19458 59442
rect 19966 59390 20018 59442
rect 24110 59390 24162 59442
rect 24558 59390 24610 59442
rect 27134 59390 27186 59442
rect 33070 59390 33122 59442
rect 14702 59278 14754 59330
rect 19742 59278 19794 59330
rect 21422 59278 21474 59330
rect 26238 59278 26290 59330
rect 20190 59222 20242 59274
rect 27470 59278 27522 59330
rect 33518 59278 33570 59330
rect 33630 59278 33682 59330
rect 34190 59334 34242 59386
rect 34526 59390 34578 59442
rect 37998 59390 38050 59442
rect 39342 59390 39394 59442
rect 39566 59390 39618 59442
rect 39678 59390 39730 59442
rect 39902 59390 39954 59442
rect 41134 59390 41186 59442
rect 42590 59390 42642 59442
rect 43710 59390 43762 59442
rect 47518 59390 47570 59442
rect 48638 59390 48690 59442
rect 48862 59390 48914 59442
rect 49422 59390 49474 59442
rect 49870 59390 49922 59442
rect 34302 59278 34354 59330
rect 35534 59278 35586 59330
rect 38446 59278 38498 59330
rect 38558 59278 38610 59330
rect 41582 59278 41634 59330
rect 47742 59278 47794 59330
rect 9550 59166 9602 59218
rect 14030 59166 14082 59218
rect 20750 59166 20802 59218
rect 21534 59166 21586 59218
rect 22766 59166 22818 59218
rect 24670 59166 24722 59218
rect 26126 59166 26178 59218
rect 26798 59166 26850 59218
rect 27134 59166 27186 59218
rect 29038 59166 29090 59218
rect 32286 59166 32338 59218
rect 33742 59166 33794 59218
rect 34862 59166 34914 59218
rect 38670 59166 38722 59218
rect 39230 59166 39282 59218
rect 40014 59166 40066 59218
rect 41134 59166 41186 59218
rect 41806 59166 41858 59218
rect 42478 59166 42530 59218
rect 42814 59166 42866 59218
rect 43486 59166 43538 59218
rect 43822 59166 43874 59218
rect 44046 59166 44098 59218
rect 44270 59166 44322 59218
rect 45166 59166 45218 59218
rect 46174 59166 46226 59218
rect 46510 59166 46562 59218
rect 46958 59166 47010 59218
rect 47294 59166 47346 59218
rect 48974 59166 49026 59218
rect 8990 59054 9042 59106
rect 10334 59054 10386 59106
rect 12462 59054 12514 59106
rect 16830 59054 16882 59106
rect 20078 59054 20130 59106
rect 21422 59054 21474 59106
rect 22430 59054 22482 59106
rect 23662 59054 23714 59106
rect 27918 59054 27970 59106
rect 28814 59054 28866 59106
rect 29822 59054 29874 59106
rect 31950 59054 32002 59106
rect 37662 59054 37714 59106
rect 43150 59054 43202 59106
rect 45502 59054 45554 59106
rect 47406 59054 47458 59106
rect 50318 59054 50370 59106
rect 8878 58942 8930 58994
rect 24558 58942 24610 58994
rect 25230 58942 25282 58994
rect 25342 58942 25394 58994
rect 25566 58942 25618 58994
rect 25678 58942 25730 58994
rect 26238 58942 26290 58994
rect 32398 58942 32450 58994
rect 45278 58942 45330 58994
rect 4478 58774 4530 58826
rect 4582 58774 4634 58826
rect 4686 58774 4738 58826
rect 35198 58774 35250 58826
rect 35302 58774 35354 58826
rect 35406 58774 35458 58826
rect 27694 58606 27746 58658
rect 29486 58606 29538 58658
rect 33182 58606 33234 58658
rect 33518 58606 33570 58658
rect 34302 58606 34354 58658
rect 40798 58606 40850 58658
rect 41806 58606 41858 58658
rect 9662 58494 9714 58546
rect 14926 58494 14978 58546
rect 15934 58494 15986 58546
rect 21534 58494 21586 58546
rect 24670 58494 24722 58546
rect 25790 58494 25842 58546
rect 30046 58494 30098 58546
rect 30942 58494 30994 58546
rect 32734 58494 32786 58546
rect 33406 58494 33458 58546
rect 39566 58494 39618 58546
rect 41470 58494 41522 58546
rect 45278 58494 45330 58546
rect 50094 58494 50146 58546
rect 12238 58382 12290 58434
rect 14814 58382 14866 58434
rect 15038 58382 15090 58434
rect 15486 58382 15538 58434
rect 16046 58382 16098 58434
rect 17166 58382 17218 58434
rect 17614 58382 17666 58434
rect 18846 58382 18898 58434
rect 19854 58382 19906 58434
rect 21870 58382 21922 58434
rect 24894 58382 24946 58434
rect 25678 58382 25730 58434
rect 26910 58382 26962 58434
rect 28030 58382 28082 58434
rect 29822 58382 29874 58434
rect 30158 58382 30210 58434
rect 32958 58382 33010 58434
rect 34190 58382 34242 58434
rect 37102 58382 37154 58434
rect 37550 58382 37602 58434
rect 38446 58382 38498 58434
rect 39230 58382 39282 58434
rect 39454 58382 39506 58434
rect 39790 58382 39842 58434
rect 40238 58382 40290 58434
rect 41358 58382 41410 58434
rect 45950 58382 46002 58434
rect 46846 58382 46898 58434
rect 47182 58382 47234 58434
rect 16494 58270 16546 58322
rect 17502 58270 17554 58322
rect 17950 58270 18002 58322
rect 20190 58270 20242 58322
rect 20526 58270 20578 58322
rect 20750 58270 20802 58322
rect 22542 58270 22594 58322
rect 26350 58270 26402 58322
rect 26686 58270 26738 58322
rect 28142 58270 28194 58322
rect 35198 58270 35250 58322
rect 36094 58270 36146 58322
rect 38110 58270 38162 58322
rect 38222 58270 38274 58322
rect 40126 58270 40178 58322
rect 40350 58270 40402 58322
rect 42926 58270 42978 58322
rect 12686 58158 12738 58210
rect 14030 58158 14082 58210
rect 14366 58158 14418 58210
rect 15262 58158 15314 58210
rect 15934 58158 15986 58210
rect 16270 58158 16322 58210
rect 17278 58158 17330 58210
rect 17838 58158 17890 58210
rect 18622 58158 18674 58210
rect 19518 58158 19570 58210
rect 19742 58158 19794 58210
rect 20302 58158 20354 58210
rect 28254 58158 28306 58210
rect 28366 58158 28418 58210
rect 29934 58158 29986 58210
rect 31502 58158 31554 58210
rect 31950 58158 32002 58210
rect 34302 58158 34354 58210
rect 34862 58158 34914 58210
rect 35646 58158 35698 58210
rect 37662 58158 37714 58210
rect 37774 58158 37826 58210
rect 38782 58158 38834 58210
rect 42590 58158 42642 58210
rect 43598 58214 43650 58266
rect 43710 58214 43762 58266
rect 44382 58270 44434 58322
rect 46734 58270 46786 58322
rect 47966 58270 48018 58322
rect 43934 58158 43986 58210
rect 44942 58158 44994 58210
rect 45166 58158 45218 58210
rect 45390 58158 45442 58210
rect 45838 58158 45890 58210
rect 19838 57990 19890 58042
rect 19942 57990 19994 58042
rect 20046 57990 20098 58042
rect 50558 57990 50610 58042
rect 50662 57990 50714 58042
rect 50766 57990 50818 58042
rect 10670 57822 10722 57874
rect 20750 57822 20802 57874
rect 20974 57822 21026 57874
rect 21422 57822 21474 57874
rect 21534 57822 21586 57874
rect 22766 57822 22818 57874
rect 22878 57822 22930 57874
rect 24558 57822 24610 57874
rect 30830 57822 30882 57874
rect 32622 57822 32674 57874
rect 41806 57822 41858 57874
rect 41918 57822 41970 57874
rect 42030 57822 42082 57874
rect 43486 57822 43538 57874
rect 43710 57822 43762 57874
rect 45166 57822 45218 57874
rect 46734 57822 46786 57874
rect 47182 57822 47234 57874
rect 9662 57710 9714 57762
rect 13470 57710 13522 57762
rect 18398 57710 18450 57762
rect 21086 57710 21138 57762
rect 23550 57710 23602 57762
rect 41134 57710 41186 57762
rect 42254 57710 42306 57762
rect 43822 57710 43874 57762
rect 48078 57710 48130 57762
rect 6190 57598 6242 57650
rect 9550 57598 9602 57650
rect 9886 57598 9938 57650
rect 10446 57598 10498 57650
rect 10558 57598 10610 57650
rect 10782 57598 10834 57650
rect 11006 57598 11058 57650
rect 12798 57598 12850 57650
rect 17614 57598 17666 57650
rect 21646 57598 21698 57650
rect 21982 57598 22034 57650
rect 22654 57598 22706 57650
rect 23326 57598 23378 57650
rect 23998 57598 24050 57650
rect 24670 57598 24722 57650
rect 25230 57598 25282 57650
rect 30942 57598 30994 57650
rect 33518 57598 33570 57650
rect 38558 57598 38610 57650
rect 41022 57598 41074 57650
rect 41358 57598 41410 57650
rect 41582 57598 41634 57650
rect 44942 57598 44994 57650
rect 45278 57598 45330 57650
rect 45614 57598 45666 57650
rect 46062 57598 46114 57650
rect 46174 57598 46226 57650
rect 46286 57598 46338 57650
rect 46958 57598 47010 57650
rect 47406 57598 47458 57650
rect 47630 57598 47682 57650
rect 47854 57598 47906 57650
rect 48190 57598 48242 57650
rect 6862 57486 6914 57538
rect 8990 57486 9042 57538
rect 20526 57486 20578 57538
rect 27246 57486 27298 57538
rect 31390 57486 31442 57538
rect 33182 57486 33234 57538
rect 34078 57486 34130 57538
rect 36878 57486 36930 57538
rect 40350 57486 40402 57538
rect 48862 57486 48914 57538
rect 49310 57486 49362 57538
rect 49758 57486 49810 57538
rect 4478 57206 4530 57258
rect 4582 57206 4634 57258
rect 4686 57206 4738 57258
rect 35198 57206 35250 57258
rect 35302 57206 35354 57258
rect 35406 57206 35458 57258
rect 11678 57038 11730 57090
rect 13806 57038 13858 57090
rect 18510 57038 18562 57090
rect 18846 57038 18898 57090
rect 19182 57038 19234 57090
rect 20302 57038 20354 57090
rect 21422 57038 21474 57090
rect 22990 57038 23042 57090
rect 24894 57038 24946 57090
rect 36318 57038 36370 57090
rect 8542 56926 8594 56978
rect 8990 56926 9042 56978
rect 11790 56926 11842 56978
rect 15710 56926 15762 56978
rect 17838 56926 17890 56978
rect 20414 56926 20466 56978
rect 23662 56926 23714 56978
rect 26462 56926 26514 56978
rect 28590 56926 28642 56978
rect 33966 56926 34018 56978
rect 39342 56926 39394 56978
rect 41470 56926 41522 56978
rect 45838 56926 45890 56978
rect 48750 56926 48802 56978
rect 5742 56814 5794 56866
rect 8878 56814 8930 56866
rect 9438 56814 9490 56866
rect 11006 56814 11058 56866
rect 14254 56814 14306 56866
rect 14926 56814 14978 56866
rect 18174 56814 18226 56866
rect 21310 56814 21362 56866
rect 22094 56814 22146 56866
rect 22318 56814 22370 56866
rect 23214 56814 23266 56866
rect 23550 56814 23602 56866
rect 23774 56814 23826 56866
rect 24222 56814 24274 56866
rect 25678 56814 25730 56866
rect 29150 56814 29202 56866
rect 31838 56814 31890 56866
rect 32846 56814 32898 56866
rect 34414 56814 34466 56866
rect 36430 56814 36482 56866
rect 42254 56814 42306 56866
rect 47294 56814 47346 56866
rect 6414 56702 6466 56754
rect 9102 56702 9154 56754
rect 10334 56702 10386 56754
rect 10782 56702 10834 56754
rect 11230 56702 11282 56754
rect 11342 56702 11394 56754
rect 13694 56702 13746 56754
rect 18398 56702 18450 56754
rect 19406 56702 19458 56754
rect 21422 56702 21474 56754
rect 22654 56702 22706 56754
rect 22878 56702 22930 56754
rect 24334 56702 24386 56754
rect 24446 56702 24498 56754
rect 30158 56702 30210 56754
rect 33518 56702 33570 56754
rect 35198 56702 35250 56754
rect 36990 56702 37042 56754
rect 37438 56702 37490 56754
rect 38670 56702 38722 56754
rect 44046 56702 44098 56754
rect 47406 56702 47458 56754
rect 47630 56702 47682 56754
rect 9326 56590 9378 56642
rect 9998 56590 10050 56642
rect 10222 56590 10274 56642
rect 10670 56590 10722 56642
rect 14478 56590 14530 56642
rect 25342 56590 25394 56642
rect 29486 56590 29538 56642
rect 30494 56590 30546 56642
rect 30942 56590 30994 56642
rect 31614 56590 31666 56642
rect 32286 56590 32338 56642
rect 33182 56590 33234 56642
rect 34862 56590 34914 56642
rect 37102 56590 37154 56642
rect 37550 56590 37602 56642
rect 37998 56590 38050 56642
rect 38334 56590 38386 56642
rect 39006 56590 39058 56642
rect 43710 56590 43762 56642
rect 43934 56590 43986 56642
rect 46734 56590 46786 56642
rect 47966 56646 48018 56698
rect 48302 56702 48354 56754
rect 19838 56422 19890 56474
rect 19942 56422 19994 56474
rect 20046 56422 20098 56474
rect 50558 56422 50610 56474
rect 50662 56422 50714 56474
rect 50766 56422 50818 56474
rect 9102 56254 9154 56306
rect 11566 56254 11618 56306
rect 15710 56254 15762 56306
rect 17390 56254 17442 56306
rect 17950 56254 18002 56306
rect 21646 56254 21698 56306
rect 22094 56254 22146 56306
rect 24446 56254 24498 56306
rect 25230 56254 25282 56306
rect 30382 56254 30434 56306
rect 32510 56254 32562 56306
rect 42366 56254 42418 56306
rect 44158 56254 44210 56306
rect 44494 56254 44546 56306
rect 45390 56254 45442 56306
rect 46398 56254 46450 56306
rect 46958 56254 47010 56306
rect 47294 56254 47346 56306
rect 7198 56142 7250 56194
rect 8430 56142 8482 56194
rect 8766 56142 8818 56194
rect 8878 56142 8930 56194
rect 9886 56142 9938 56194
rect 13022 56142 13074 56194
rect 16606 56142 16658 56194
rect 16718 56142 16770 56194
rect 17502 56142 17554 56194
rect 22318 56142 22370 56194
rect 23550 56142 23602 56194
rect 34302 56142 34354 56194
rect 38558 56142 38610 56194
rect 42702 56142 42754 56194
rect 43710 56142 43762 56194
rect 45166 56142 45218 56194
rect 45502 56142 45554 56194
rect 47854 56142 47906 56194
rect 48078 56142 48130 56194
rect 48974 56142 49026 56194
rect 49086 56142 49138 56194
rect 6974 56030 7026 56082
rect 7086 56030 7138 56082
rect 7310 56030 7362 56082
rect 7422 56030 7474 56082
rect 8318 56030 8370 56082
rect 10110 56030 10162 56082
rect 10334 56030 10386 56082
rect 10558 56030 10610 56082
rect 11342 56030 11394 56082
rect 12238 56030 12290 56082
rect 15486 56030 15538 56082
rect 15934 56030 15986 56082
rect 16158 56030 16210 56082
rect 16382 56030 16434 56082
rect 22542 56030 22594 56082
rect 23998 56030 24050 56082
rect 24334 56030 24386 56082
rect 25454 56030 25506 56082
rect 25902 56030 25954 56082
rect 26574 56030 26626 56082
rect 33070 56030 33122 56082
rect 33518 56030 33570 56082
rect 33966 56030 34018 56082
rect 34974 56030 35026 56082
rect 42926 56030 42978 56082
rect 43262 56030 43314 56082
rect 43934 56030 43986 56082
rect 44718 56030 44770 56082
rect 45054 56030 45106 56082
rect 47630 56030 47682 56082
rect 48862 56030 48914 56082
rect 7982 55918 8034 55970
rect 10446 55918 10498 55970
rect 15150 55918 15202 55970
rect 15822 55918 15874 55970
rect 20414 55918 20466 55970
rect 23102 55918 23154 55970
rect 25342 55918 25394 55970
rect 26350 55918 26402 55970
rect 27358 55918 27410 55970
rect 29486 55918 29538 55970
rect 29934 55918 29986 55970
rect 31838 55918 31890 55970
rect 40350 55918 40402 55970
rect 41022 55918 41074 55970
rect 42702 55918 42754 55970
rect 45838 55918 45890 55970
rect 7870 55806 7922 55858
rect 20302 55806 20354 55858
rect 44270 55806 44322 55858
rect 44382 55806 44434 55858
rect 45950 55806 46002 55858
rect 47742 55806 47794 55858
rect 49534 55806 49586 55858
rect 4478 55638 4530 55690
rect 4582 55638 4634 55690
rect 4686 55638 4738 55690
rect 35198 55638 35250 55690
rect 35302 55638 35354 55690
rect 35406 55638 35458 55690
rect 8542 55358 8594 55410
rect 9326 55358 9378 55410
rect 13470 55358 13522 55410
rect 15598 55358 15650 55410
rect 17838 55358 17890 55410
rect 28030 55358 28082 55410
rect 31726 55358 31778 55410
rect 34414 55358 34466 55410
rect 34974 55358 35026 55410
rect 37774 55358 37826 55410
rect 39902 55358 39954 55410
rect 43822 55358 43874 55410
rect 45950 55358 46002 55410
rect 48078 55358 48130 55410
rect 48638 55358 48690 55410
rect 5742 55246 5794 55298
rect 12238 55246 12290 55298
rect 16382 55246 16434 55298
rect 19630 55246 19682 55298
rect 26350 55246 26402 55298
rect 27022 55246 27074 55298
rect 28142 55246 28194 55298
rect 28366 55246 28418 55298
rect 28590 55246 28642 55298
rect 29262 55246 29314 55298
rect 32062 55246 32114 55298
rect 33966 55246 34018 55298
rect 36206 55246 36258 55298
rect 36542 55246 36594 55298
rect 36990 55246 37042 55298
rect 41582 55246 41634 55298
rect 42702 55246 42754 55298
rect 43374 55246 43426 55298
rect 43710 55246 43762 55298
rect 44382 55246 44434 55298
rect 45166 55246 45218 55298
rect 48750 55246 48802 55298
rect 49310 55246 49362 55298
rect 50430 55246 50482 55298
rect 6414 55134 6466 55186
rect 11454 55134 11506 55186
rect 19966 55134 20018 55186
rect 20526 55134 20578 55186
rect 20638 55134 20690 55186
rect 23438 55134 23490 55186
rect 27246 55134 27298 55186
rect 30270 55134 30322 55186
rect 32398 55134 32450 55186
rect 35646 55134 35698 55186
rect 41022 55134 41074 55186
rect 42254 55134 42306 55186
rect 48526 55134 48578 55186
rect 17390 55022 17442 55074
rect 18398 55022 18450 55074
rect 19854 55022 19906 55074
rect 20302 55022 20354 55074
rect 27918 55022 27970 55074
rect 29150 55022 29202 55074
rect 29934 55022 29986 55074
rect 30718 55022 30770 55074
rect 31166 55022 31218 55074
rect 35310 55022 35362 55074
rect 35870 55022 35922 55074
rect 35982 55022 36034 55074
rect 41134 55022 41186 55074
rect 41806 55022 41858 55074
rect 42142 55022 42194 55074
rect 42366 55022 42418 55074
rect 43038 55022 43090 55074
rect 43934 55022 43986 55074
rect 49870 55022 49922 55074
rect 49982 55022 50034 55074
rect 50094 55022 50146 55074
rect 19838 54854 19890 54906
rect 19942 54854 19994 54906
rect 20046 54854 20098 54906
rect 50558 54854 50610 54906
rect 50662 54854 50714 54906
rect 50766 54854 50818 54906
rect 6638 54686 6690 54738
rect 6750 54686 6802 54738
rect 6974 54686 7026 54738
rect 7422 54686 7474 54738
rect 7646 54686 7698 54738
rect 8654 54686 8706 54738
rect 15598 54686 15650 54738
rect 24558 54686 24610 54738
rect 26462 54686 26514 54738
rect 31166 54686 31218 54738
rect 31838 54686 31890 54738
rect 34078 54686 34130 54738
rect 34414 54686 34466 54738
rect 36318 54686 36370 54738
rect 47966 54686 48018 54738
rect 2046 54574 2098 54626
rect 7758 54574 7810 54626
rect 15150 54574 15202 54626
rect 15262 54574 15314 54626
rect 16494 54574 16546 54626
rect 26126 54574 26178 54626
rect 26798 54574 26850 54626
rect 26910 54574 26962 54626
rect 29150 54574 29202 54626
rect 29486 54574 29538 54626
rect 29822 54574 29874 54626
rect 30158 54574 30210 54626
rect 30494 54574 30546 54626
rect 34750 54574 34802 54626
rect 35086 54574 35138 54626
rect 37550 54574 37602 54626
rect 41694 54574 41746 54626
rect 48190 54574 48242 54626
rect 50878 54574 50930 54626
rect 1710 54462 1762 54514
rect 7198 54462 7250 54514
rect 8878 54462 8930 54514
rect 9662 54462 9714 54514
rect 14926 54462 14978 54514
rect 15710 54462 15762 54514
rect 16270 54462 16322 54514
rect 23438 54462 23490 54514
rect 24446 54462 24498 54514
rect 24782 54462 24834 54514
rect 25678 54462 25730 54514
rect 30942 54462 30994 54514
rect 32174 54462 32226 54514
rect 35310 54462 35362 54514
rect 35646 54462 35698 54514
rect 35758 54462 35810 54514
rect 36206 54462 36258 54514
rect 36430 54462 36482 54514
rect 36766 54462 36818 54514
rect 41022 54462 41074 54514
rect 44158 54462 44210 54514
rect 47630 54462 47682 54514
rect 51662 54462 51714 54514
rect 2494 54350 2546 54402
rect 6638 54350 6690 54402
rect 10334 54350 10386 54402
rect 12462 54350 12514 54402
rect 17502 54350 17554 54402
rect 18062 54350 18114 54402
rect 21310 54350 21362 54402
rect 27470 54350 27522 54402
rect 27918 54350 27970 54402
rect 28366 54350 28418 54402
rect 33294 54350 33346 54402
rect 39678 54350 39730 54402
rect 43822 54350 43874 54402
rect 44942 54350 44994 54402
rect 47070 54350 47122 54402
rect 48078 54350 48130 54402
rect 48750 54350 48802 54402
rect 25342 54238 25394 54290
rect 25454 54238 25506 54290
rect 25790 54238 25842 54290
rect 26910 54238 26962 54290
rect 33406 54238 33458 54290
rect 35422 54238 35474 54290
rect 4478 54070 4530 54122
rect 4582 54070 4634 54122
rect 4686 54070 4738 54122
rect 35198 54070 35250 54122
rect 35302 54070 35354 54122
rect 35406 54070 35458 54122
rect 44942 53902 44994 53954
rect 49534 53902 49586 53954
rect 49758 53902 49810 53954
rect 49870 53902 49922 53954
rect 6638 53790 6690 53842
rect 10446 53790 10498 53842
rect 20750 53790 20802 53842
rect 22094 53790 22146 53842
rect 24222 53790 24274 53842
rect 25342 53790 25394 53842
rect 26686 53790 26738 53842
rect 27918 53790 27970 53842
rect 31614 53790 31666 53842
rect 34974 53790 35026 53842
rect 37438 53790 37490 53842
rect 47854 53790 47906 53842
rect 48638 53790 48690 53842
rect 49422 53790 49474 53842
rect 6750 53678 6802 53730
rect 6974 53678 7026 53730
rect 7422 53678 7474 53730
rect 7758 53678 7810 53730
rect 8206 53678 8258 53730
rect 9662 53678 9714 53730
rect 10222 53678 10274 53730
rect 10558 53678 10610 53730
rect 10782 53678 10834 53730
rect 11118 53678 11170 53730
rect 11230 53678 11282 53730
rect 17950 53678 18002 53730
rect 18622 53678 18674 53730
rect 21310 53678 21362 53730
rect 24446 53678 24498 53730
rect 25566 53678 25618 53730
rect 26126 53678 26178 53730
rect 26798 53678 26850 53730
rect 27470 53678 27522 53730
rect 27694 53678 27746 53730
rect 28030 53678 28082 53730
rect 33742 53678 33794 53730
rect 34414 53678 34466 53730
rect 35086 53678 35138 53730
rect 35534 53678 35586 53730
rect 35758 53678 35810 53730
rect 35982 53678 36034 53730
rect 36430 53678 36482 53730
rect 37886 53678 37938 53730
rect 38222 53678 38274 53730
rect 40126 53678 40178 53730
rect 40798 53678 40850 53730
rect 42478 53678 42530 53730
rect 43038 53678 43090 53730
rect 43934 53678 43986 53730
rect 44270 53678 44322 53730
rect 46734 53678 46786 53730
rect 47070 53678 47122 53730
rect 47742 53678 47794 53730
rect 48526 53678 48578 53730
rect 50542 53678 50594 53730
rect 1710 53566 1762 53618
rect 7198 53566 7250 53618
rect 9438 53566 9490 53618
rect 16270 53566 16322 53618
rect 25230 53566 25282 53618
rect 27134 53566 27186 53618
rect 27246 53566 27298 53618
rect 30046 53566 30098 53618
rect 30382 53566 30434 53618
rect 37102 53566 37154 53618
rect 41358 53566 41410 53618
rect 41694 53566 41746 53618
rect 42702 53566 42754 53618
rect 43262 53566 43314 53618
rect 43374 53566 43426 53618
rect 43822 53566 43874 53618
rect 44830 53566 44882 53618
rect 50206 53566 50258 53618
rect 50318 53566 50370 53618
rect 50878 53566 50930 53618
rect 2046 53454 2098 53506
rect 2494 53454 2546 53506
rect 6638 53454 6690 53506
rect 7646 53454 7698 53506
rect 8094 53454 8146 53506
rect 10334 53454 10386 53506
rect 16382 53454 16434 53506
rect 16606 53454 16658 53506
rect 16942 53454 16994 53506
rect 17614 53454 17666 53506
rect 26574 53454 26626 53506
rect 28254 53454 28306 53506
rect 29710 53454 29762 53506
rect 34862 53454 34914 53506
rect 35870 53454 35922 53506
rect 37326 53454 37378 53506
rect 37550 53454 37602 53506
rect 37998 53454 38050 53506
rect 40462 53454 40514 53506
rect 41022 53454 41074 53506
rect 41246 53454 41298 53506
rect 41806 53454 41858 53506
rect 42030 53454 42082 53506
rect 42254 53454 42306 53506
rect 42366 53454 42418 53506
rect 43710 53454 43762 53506
rect 46510 53454 46562 53506
rect 46622 53454 46674 53506
rect 19838 53286 19890 53338
rect 19942 53286 19994 53338
rect 20046 53286 20098 53338
rect 50558 53286 50610 53338
rect 50662 53286 50714 53338
rect 50766 53286 50818 53338
rect 8430 53118 8482 53170
rect 9998 53118 10050 53170
rect 11678 53118 11730 53170
rect 14478 53118 14530 53170
rect 15598 53118 15650 53170
rect 22990 53118 23042 53170
rect 23326 53118 23378 53170
rect 24670 53118 24722 53170
rect 26686 53118 26738 53170
rect 27246 53118 27298 53170
rect 28366 53118 28418 53170
rect 30046 53118 30098 53170
rect 30270 53118 30322 53170
rect 30830 53118 30882 53170
rect 31054 53118 31106 53170
rect 32286 53118 32338 53170
rect 33070 53118 33122 53170
rect 35198 53118 35250 53170
rect 35422 53118 35474 53170
rect 35534 53118 35586 53170
rect 36430 53118 36482 53170
rect 36766 53118 36818 53170
rect 37438 53118 37490 53170
rect 46958 53118 47010 53170
rect 48302 53118 48354 53170
rect 49086 53118 49138 53170
rect 2046 53006 2098 53058
rect 5294 53006 5346 53058
rect 7758 53006 7810 53058
rect 13582 53006 13634 53058
rect 13918 53006 13970 53058
rect 14926 53006 14978 53058
rect 15934 53006 15986 53058
rect 16494 53006 16546 53058
rect 20974 53006 21026 53058
rect 23214 53006 23266 53058
rect 24110 53006 24162 53058
rect 26014 53006 26066 53058
rect 29038 53006 29090 53058
rect 33406 53006 33458 53058
rect 34526 53006 34578 53058
rect 34638 53006 34690 53058
rect 36542 53006 36594 53058
rect 39454 53006 39506 53058
rect 42590 53006 42642 53058
rect 1710 52894 1762 52946
rect 4622 52894 4674 52946
rect 8094 52894 8146 52946
rect 8766 52894 8818 52946
rect 9774 52894 9826 52946
rect 12014 52894 12066 52946
rect 14366 52894 14418 52946
rect 14702 52894 14754 52946
rect 15374 52894 15426 52946
rect 15486 52894 15538 52946
rect 15710 52894 15762 52946
rect 16718 52894 16770 52946
rect 17502 52894 17554 52946
rect 20750 52894 20802 52946
rect 21198 52894 21250 52946
rect 21646 52894 21698 52946
rect 21870 52894 21922 52946
rect 22766 52894 22818 52946
rect 23998 52894 24050 52946
rect 24222 52894 24274 52946
rect 25678 52894 25730 52946
rect 26350 52894 26402 52946
rect 27470 52894 27522 52946
rect 27918 52894 27970 52946
rect 28478 52894 28530 52946
rect 28814 52894 28866 52946
rect 29486 52894 29538 52946
rect 30606 52894 30658 52946
rect 31390 52894 31442 52946
rect 34862 52894 34914 52946
rect 37102 52894 37154 52946
rect 37214 52894 37266 52946
rect 37550 52894 37602 52946
rect 39006 52894 39058 52946
rect 39678 52894 39730 52946
rect 42254 52894 42306 52946
rect 42814 52950 42866 53002
rect 43150 53006 43202 53058
rect 45390 53006 45442 53058
rect 45950 53006 46002 53058
rect 46062 53006 46114 53058
rect 47966 53006 48018 53058
rect 48078 53006 48130 53058
rect 45726 52894 45778 52946
rect 47182 52894 47234 52946
rect 49310 52894 49362 52946
rect 2494 52782 2546 52834
rect 7422 52782 7474 52834
rect 14590 52782 14642 52834
rect 18174 52782 18226 52834
rect 20302 52782 20354 52834
rect 21758 52782 21810 52834
rect 25342 52782 25394 52834
rect 27358 52782 27410 52834
rect 28926 52782 28978 52834
rect 29486 52782 29538 52834
rect 29822 52782 29874 52834
rect 31838 52782 31890 52834
rect 39230 52782 39282 52834
rect 42478 52782 42530 52834
rect 47294 52782 47346 52834
rect 28366 52670 28418 52722
rect 29934 52670 29986 52722
rect 30718 52670 30770 52722
rect 34526 52670 34578 52722
rect 43262 52670 43314 52722
rect 46510 52670 46562 52722
rect 4478 52502 4530 52554
rect 4582 52502 4634 52554
rect 4686 52502 4738 52554
rect 35198 52502 35250 52554
rect 35302 52502 35354 52554
rect 35406 52502 35458 52554
rect 8094 52334 8146 52386
rect 11902 52334 11954 52386
rect 19182 52334 19234 52386
rect 20526 52334 20578 52386
rect 21198 52334 21250 52386
rect 21758 52334 21810 52386
rect 25342 52334 25394 52386
rect 29262 52334 29314 52386
rect 6638 52222 6690 52274
rect 15262 52222 15314 52274
rect 17390 52222 17442 52274
rect 20078 52222 20130 52274
rect 20638 52222 20690 52274
rect 21422 52222 21474 52274
rect 22430 52222 22482 52274
rect 23550 52222 23602 52274
rect 25230 52222 25282 52274
rect 28590 52222 28642 52274
rect 33294 52222 33346 52274
rect 34862 52222 34914 52274
rect 38894 52222 38946 52274
rect 45502 52222 45554 52274
rect 1710 52110 1762 52162
rect 2494 52110 2546 52162
rect 6526 52110 6578 52162
rect 6750 52110 6802 52162
rect 6974 52110 7026 52162
rect 7086 52110 7138 52162
rect 7422 52110 7474 52162
rect 8206 52110 8258 52162
rect 11454 52110 11506 52162
rect 12574 52110 12626 52162
rect 13022 52110 13074 52162
rect 13918 52110 13970 52162
rect 14590 52110 14642 52162
rect 18286 52110 18338 52162
rect 19406 52110 19458 52162
rect 19630 52110 19682 52162
rect 20190 52110 20242 52162
rect 22206 52110 22258 52162
rect 22878 52110 22930 52162
rect 24222 52110 24274 52162
rect 25678 52110 25730 52162
rect 29038 52110 29090 52162
rect 30158 52110 30210 52162
rect 30718 52110 30770 52162
rect 32398 52110 32450 52162
rect 33518 52110 33570 52162
rect 38222 52110 38274 52162
rect 38446 52110 38498 52162
rect 39790 52110 39842 52162
rect 39902 52110 39954 52162
rect 40014 52110 40066 52162
rect 44270 52110 44322 52162
rect 49422 52110 49474 52162
rect 7646 51998 7698 52050
rect 7758 51998 7810 52050
rect 11118 51998 11170 52050
rect 12014 51998 12066 52050
rect 14142 51998 14194 52050
rect 19070 51998 19122 52050
rect 19966 51998 20018 52050
rect 23102 51998 23154 52050
rect 23998 51998 24050 52050
rect 26462 51998 26514 52050
rect 29374 51998 29426 52050
rect 29598 51998 29650 52050
rect 30382 51998 30434 52050
rect 30942 51998 30994 52050
rect 31054 51998 31106 52050
rect 32734 51998 32786 52050
rect 33854 51998 33906 52050
rect 38670 51998 38722 52050
rect 39006 51998 39058 52050
rect 2046 51886 2098 51938
rect 11902 51886 11954 51938
rect 17950 51886 18002 51938
rect 18398 51886 18450 51938
rect 18622 51886 18674 51938
rect 18846 51886 18898 51938
rect 29934 51886 29986 51938
rect 30046 51886 30098 51938
rect 32622 51886 32674 51938
rect 34750 51886 34802 51938
rect 39342 51886 39394 51938
rect 19838 51718 19890 51770
rect 19942 51718 19994 51770
rect 20046 51718 20098 51770
rect 50558 51718 50610 51770
rect 50662 51718 50714 51770
rect 50766 51718 50818 51770
rect 16270 51550 16322 51602
rect 16718 51550 16770 51602
rect 17838 51550 17890 51602
rect 19742 51550 19794 51602
rect 20526 51550 20578 51602
rect 28478 51550 28530 51602
rect 36430 51550 36482 51602
rect 38558 51550 38610 51602
rect 39006 51550 39058 51602
rect 45054 51550 45106 51602
rect 47742 51550 47794 51602
rect 48078 51550 48130 51602
rect 48862 51550 48914 51602
rect 49758 51550 49810 51602
rect 2046 51438 2098 51490
rect 5294 51438 5346 51490
rect 9886 51438 9938 51490
rect 16830 51438 16882 51490
rect 18062 51438 18114 51490
rect 19966 51438 20018 51490
rect 21198 51438 21250 51490
rect 22878 51438 22930 51490
rect 23214 51438 23266 51490
rect 26014 51438 26066 51490
rect 28590 51438 28642 51490
rect 33966 51438 34018 51490
rect 37998 51438 38050 51490
rect 43374 51438 43426 51490
rect 44830 51438 44882 51490
rect 45166 51438 45218 51490
rect 45390 51438 45442 51490
rect 46734 51438 46786 51490
rect 47518 51438 47570 51490
rect 48750 51438 48802 51490
rect 49310 51438 49362 51490
rect 1710 51326 1762 51378
rect 4622 51326 4674 51378
rect 10110 51326 10162 51378
rect 15822 51326 15874 51378
rect 16046 51326 16098 51378
rect 16382 51326 16434 51378
rect 18286 51326 18338 51378
rect 19406 51326 19458 51378
rect 20302 51326 20354 51378
rect 20638 51326 20690 51378
rect 20750 51326 20802 51378
rect 21422 51326 21474 51378
rect 21870 51326 21922 51378
rect 22094 51326 22146 51378
rect 22542 51326 22594 51378
rect 23326 51326 23378 51378
rect 23438 51326 23490 51378
rect 23774 51326 23826 51378
rect 24222 51326 24274 51378
rect 25230 51326 25282 51378
rect 29038 51326 29090 51378
rect 33182 51326 33234 51378
rect 36766 51326 36818 51378
rect 37886 51326 37938 51378
rect 38782 51326 38834 51378
rect 38894 51326 38946 51378
rect 39454 51326 39506 51378
rect 39902 51326 39954 51378
rect 44158 51326 44210 51378
rect 46174 51326 46226 51378
rect 46958 51326 47010 51378
rect 47406 51326 47458 51378
rect 47966 51326 48018 51378
rect 48974 51326 49026 51378
rect 2494 51214 2546 51266
rect 2942 51214 2994 51266
rect 7422 51214 7474 51266
rect 11790 51214 11842 51266
rect 19294 51214 19346 51266
rect 19630 51214 19682 51266
rect 21310 51214 21362 51266
rect 28142 51214 28194 51266
rect 29710 51214 29762 51266
rect 31838 51214 31890 51266
rect 36094 51214 36146 51266
rect 37214 51214 37266 51266
rect 41246 51214 41298 51266
rect 46398 51214 46450 51266
rect 37998 51102 38050 51154
rect 39454 51102 39506 51154
rect 48078 51102 48130 51154
rect 4478 50934 4530 50986
rect 4582 50934 4634 50986
rect 4686 50934 4738 50986
rect 35198 50934 35250 50986
rect 35302 50934 35354 50986
rect 35406 50934 35458 50986
rect 7086 50766 7138 50818
rect 14478 50766 14530 50818
rect 22766 50766 22818 50818
rect 29934 50766 29986 50818
rect 36542 50766 36594 50818
rect 41806 50766 41858 50818
rect 10894 50654 10946 50706
rect 14590 50654 14642 50706
rect 16606 50654 16658 50706
rect 23326 50654 23378 50706
rect 30046 50654 30098 50706
rect 33854 50654 33906 50706
rect 35646 50654 35698 50706
rect 39230 50654 39282 50706
rect 41358 50654 41410 50706
rect 42366 50654 42418 50706
rect 46734 50654 46786 50706
rect 47070 50654 47122 50706
rect 49198 50654 49250 50706
rect 1822 50542 1874 50594
rect 7198 50542 7250 50594
rect 12238 50542 12290 50594
rect 12910 50542 12962 50594
rect 13694 50542 13746 50594
rect 20078 50542 20130 50594
rect 20750 50542 20802 50594
rect 22206 50542 22258 50594
rect 22318 50542 22370 50594
rect 26350 50542 26402 50594
rect 27022 50542 27074 50594
rect 31278 50542 31330 50594
rect 33406 50542 33458 50594
rect 35870 50542 35922 50594
rect 36990 50542 37042 50594
rect 37998 50542 38050 50594
rect 38558 50542 38610 50594
rect 41694 50542 41746 50594
rect 43150 50542 43202 50594
rect 43486 50542 43538 50594
rect 43822 50542 43874 50594
rect 49982 50542 50034 50594
rect 2046 50430 2098 50482
rect 2382 50430 2434 50482
rect 2718 50430 2770 50482
rect 3166 50430 3218 50482
rect 7086 50430 7138 50482
rect 9438 50430 9490 50482
rect 9774 50430 9826 50482
rect 10110 50430 10162 50482
rect 10446 50430 10498 50482
rect 10894 50430 10946 50482
rect 11006 50430 11058 50482
rect 11230 50430 11282 50482
rect 11454 50430 11506 50482
rect 12462 50430 12514 50482
rect 12798 50430 12850 50482
rect 13470 50430 13522 50482
rect 20638 50430 20690 50482
rect 22094 50430 22146 50482
rect 23662 50430 23714 50482
rect 37102 50430 37154 50482
rect 41806 50430 41858 50482
rect 43934 50430 43986 50482
rect 20414 50318 20466 50370
rect 21310 50318 21362 50370
rect 21646 50318 21698 50370
rect 26462 50318 26514 50370
rect 26574 50318 26626 50370
rect 30942 50318 30994 50370
rect 36206 50318 36258 50370
rect 36430 50318 36482 50370
rect 37886 50318 37938 50370
rect 44046 50318 44098 50370
rect 19838 50150 19890 50202
rect 19942 50150 19994 50202
rect 20046 50150 20098 50202
rect 50558 50150 50610 50202
rect 50662 50150 50714 50202
rect 50766 50150 50818 50202
rect 7086 49982 7138 50034
rect 7870 49982 7922 50034
rect 8206 49982 8258 50034
rect 16270 49982 16322 50034
rect 17502 49982 17554 50034
rect 27470 49982 27522 50034
rect 28142 49982 28194 50034
rect 36542 49982 36594 50034
rect 40126 49982 40178 50034
rect 2046 49870 2098 49922
rect 7534 49870 7586 49922
rect 13582 49870 13634 49922
rect 16046 49870 16098 49922
rect 25342 49870 25394 49922
rect 27694 49870 27746 49922
rect 28254 49870 28306 49922
rect 30382 49870 30434 49922
rect 30606 49870 30658 49922
rect 31726 49870 31778 49922
rect 35198 49870 35250 49922
rect 36206 49870 36258 49922
rect 38222 49870 38274 49922
rect 39230 49870 39282 49922
rect 42254 49870 42306 49922
rect 45838 49870 45890 49922
rect 51662 49870 51714 49922
rect 1710 49758 1762 49810
rect 6862 49758 6914 49810
rect 7198 49758 7250 49810
rect 8542 49758 8594 49810
rect 9662 49758 9714 49810
rect 12798 49758 12850 49810
rect 16494 49758 16546 49810
rect 16718 49758 16770 49810
rect 18510 49758 18562 49810
rect 19294 49758 19346 49810
rect 26350 49758 26402 49810
rect 26574 49758 26626 49810
rect 27022 49758 27074 49810
rect 27246 49758 27298 49810
rect 30158 49758 30210 49810
rect 31390 49758 31442 49810
rect 35310 49758 35362 49810
rect 36766 49758 36818 49810
rect 37550 49758 37602 49810
rect 39454 49758 39506 49810
rect 40014 49758 40066 49810
rect 42142 49758 42194 49810
rect 42478 49758 42530 49810
rect 43150 49758 43202 49810
rect 43486 49758 43538 49810
rect 43710 49758 43762 49810
rect 43934 49758 43986 49810
rect 44270 49758 44322 49810
rect 44494 49758 44546 49810
rect 49310 49758 49362 49810
rect 49646 49758 49698 49810
rect 2494 49646 2546 49698
rect 10334 49646 10386 49698
rect 12462 49646 12514 49698
rect 15710 49646 15762 49698
rect 16382 49646 16434 49698
rect 18062 49646 18114 49698
rect 18846 49646 18898 49698
rect 20078 49646 20130 49698
rect 22206 49646 22258 49698
rect 26462 49646 26514 49698
rect 28702 49646 28754 49698
rect 29598 49646 29650 49698
rect 34750 49646 34802 49698
rect 35870 49646 35922 49698
rect 37438 49646 37490 49698
rect 43598 49646 43650 49698
rect 44158 49646 44210 49698
rect 45390 49646 45442 49698
rect 17838 49534 17890 49586
rect 25230 49534 25282 49586
rect 27358 49534 27410 49586
rect 28142 49534 28194 49586
rect 29374 49534 29426 49586
rect 29598 49534 29650 49586
rect 30270 49534 30322 49586
rect 35198 49534 35250 49586
rect 4478 49366 4530 49418
rect 4582 49366 4634 49418
rect 4686 49366 4738 49418
rect 35198 49366 35250 49418
rect 35302 49366 35354 49418
rect 35406 49366 35458 49418
rect 43822 49198 43874 49250
rect 45950 49198 46002 49250
rect 1934 49086 1986 49138
rect 8542 49086 8594 49138
rect 8990 49086 9042 49138
rect 10222 49086 10274 49138
rect 12350 49086 12402 49138
rect 13582 49086 13634 49138
rect 15374 49086 15426 49138
rect 17502 49086 17554 49138
rect 21422 49086 21474 49138
rect 24334 49086 24386 49138
rect 26462 49086 26514 49138
rect 27246 49086 27298 49138
rect 28142 49086 28194 49138
rect 32622 49086 32674 49138
rect 37102 49086 37154 49138
rect 38670 49086 38722 49138
rect 40238 49086 40290 49138
rect 41134 49086 41186 49138
rect 43150 49086 43202 49138
rect 44942 49086 44994 49138
rect 49982 49086 50034 49138
rect 4286 48974 4338 49026
rect 5630 48974 5682 49026
rect 9550 48974 9602 49026
rect 12574 48974 12626 49026
rect 13470 48974 13522 49026
rect 13918 48974 13970 49026
rect 14030 48974 14082 49026
rect 14702 48974 14754 49026
rect 18286 48974 18338 49026
rect 20414 48974 20466 49026
rect 20750 48974 20802 49026
rect 23662 48974 23714 49026
rect 27694 48974 27746 49026
rect 29822 48974 29874 49026
rect 33406 48974 33458 49026
rect 34638 48974 34690 49026
rect 35758 48974 35810 49026
rect 35870 48974 35922 49026
rect 37550 48974 37602 49026
rect 38110 48974 38162 49026
rect 39006 48974 39058 49026
rect 39454 48974 39506 49026
rect 41806 48974 41858 49026
rect 42030 48974 42082 49026
rect 42702 48974 42754 49026
rect 46174 48974 46226 49026
rect 47182 48974 47234 49026
rect 50430 48974 50482 49026
rect 4734 48862 4786 48914
rect 6414 48862 6466 48914
rect 12910 48862 12962 48914
rect 13694 48862 13746 48914
rect 17838 48862 17890 48914
rect 18062 48862 18114 48914
rect 20190 48862 20242 48914
rect 20638 48862 20690 48914
rect 29374 48862 29426 48914
rect 30494 48862 30546 48914
rect 33742 48862 33794 48914
rect 35982 48862 36034 48914
rect 39678 48862 39730 48914
rect 39790 48862 39842 48914
rect 41470 48862 41522 48914
rect 42254 48862 42306 48914
rect 42366 48862 42418 48914
rect 43598 48862 43650 48914
rect 45278 48862 45330 48914
rect 46510 48862 46562 48914
rect 47854 48862 47906 48914
rect 8878 48750 8930 48802
rect 12798 48750 12850 48802
rect 18174 48750 18226 48802
rect 18398 48750 18450 48802
rect 19070 48750 19122 48802
rect 19630 48750 19682 48802
rect 19854 48750 19906 48802
rect 29038 48750 29090 48802
rect 29262 48750 29314 48802
rect 34414 48750 34466 48802
rect 34974 48750 35026 48802
rect 36430 48750 36482 48802
rect 36990 48750 37042 48802
rect 37214 48750 37266 48802
rect 37774 48750 37826 48802
rect 37998 48750 38050 48802
rect 39118 48750 39170 48802
rect 39342 48750 39394 48802
rect 41582 48750 41634 48802
rect 42926 48750 42978 48802
rect 43150 48750 43202 48802
rect 44158 48750 44210 48802
rect 45614 48750 45666 48802
rect 46398 48750 46450 48802
rect 46622 48750 46674 48802
rect 50318 48750 50370 48802
rect 19838 48582 19890 48634
rect 19942 48582 19994 48634
rect 20046 48582 20098 48634
rect 50558 48582 50610 48634
rect 50662 48582 50714 48634
rect 50766 48582 50818 48634
rect 6974 48414 7026 48466
rect 7086 48414 7138 48466
rect 8094 48414 8146 48466
rect 11678 48414 11730 48466
rect 16718 48414 16770 48466
rect 17502 48414 17554 48466
rect 17726 48414 17778 48466
rect 21198 48414 21250 48466
rect 22094 48414 22146 48466
rect 23774 48414 23826 48466
rect 33742 48414 33794 48466
rect 38222 48414 38274 48466
rect 39118 48414 39170 48466
rect 40014 48414 40066 48466
rect 41022 48414 41074 48466
rect 43374 48414 43426 48466
rect 43598 48414 43650 48466
rect 43822 48414 43874 48466
rect 44830 48414 44882 48466
rect 7198 48302 7250 48354
rect 7758 48302 7810 48354
rect 8654 48302 8706 48354
rect 10110 48302 10162 48354
rect 16830 48302 16882 48354
rect 17390 48302 17442 48354
rect 22206 48302 22258 48354
rect 31278 48302 31330 48354
rect 33070 48302 33122 48354
rect 37998 48302 38050 48354
rect 38446 48302 38498 48354
rect 43262 48302 43314 48354
rect 46062 48302 46114 48354
rect 4286 48190 4338 48242
rect 6862 48190 6914 48242
rect 7422 48190 7474 48242
rect 8878 48190 8930 48242
rect 9886 48190 9938 48242
rect 10222 48190 10274 48242
rect 11454 48190 11506 48242
rect 11790 48190 11842 48242
rect 15262 48190 15314 48242
rect 16046 48190 16098 48242
rect 18062 48190 18114 48242
rect 20974 48190 21026 48242
rect 21310 48190 21362 48242
rect 21534 48190 21586 48242
rect 21758 48190 21810 48242
rect 22430 48190 22482 48242
rect 24222 48190 24274 48242
rect 25230 48190 25282 48242
rect 30942 48190 30994 48242
rect 32062 48190 32114 48242
rect 33294 48190 33346 48242
rect 34638 48178 34690 48230
rect 38670 48190 38722 48242
rect 39342 48190 39394 48242
rect 39678 48190 39730 48242
rect 40238 48190 40290 48242
rect 41470 48190 41522 48242
rect 45390 48190 45442 48242
rect 4846 48078 4898 48130
rect 6302 48078 6354 48130
rect 11118 48078 11170 48130
rect 12462 48078 12514 48130
rect 14590 48078 14642 48130
rect 15710 48078 15762 48130
rect 15822 48078 15874 48130
rect 17950 48078 18002 48130
rect 18510 48078 18562 48130
rect 22878 48078 22930 48130
rect 24670 48078 24722 48130
rect 27246 48078 27298 48130
rect 31614 48078 31666 48130
rect 32510 48078 32562 48130
rect 34302 48078 34354 48130
rect 35422 48078 35474 48130
rect 37550 48078 37602 48130
rect 38446 48078 38498 48130
rect 39230 48078 39282 48130
rect 40126 48078 40178 48130
rect 40910 48078 40962 48130
rect 42478 48078 42530 48130
rect 42926 48078 42978 48130
rect 43934 48078 43986 48130
rect 44382 48078 44434 48130
rect 48190 48078 48242 48130
rect 1934 47966 1986 48018
rect 6414 47966 6466 48018
rect 42478 47966 42530 48018
rect 42702 47966 42754 48018
rect 4478 47798 4530 47850
rect 4582 47798 4634 47850
rect 4686 47798 4738 47850
rect 35198 47798 35250 47850
rect 35302 47798 35354 47850
rect 35406 47798 35458 47850
rect 12798 47630 12850 47682
rect 14478 47630 14530 47682
rect 38110 47630 38162 47682
rect 41022 47630 41074 47682
rect 42030 47630 42082 47682
rect 42254 47630 42306 47682
rect 1934 47518 1986 47570
rect 5854 47518 5906 47570
rect 12686 47518 12738 47570
rect 14366 47518 14418 47570
rect 16270 47518 16322 47570
rect 18398 47518 18450 47570
rect 27694 47518 27746 47570
rect 32622 47518 32674 47570
rect 37438 47518 37490 47570
rect 38894 47518 38946 47570
rect 39566 47518 39618 47570
rect 40574 47518 40626 47570
rect 42254 47518 42306 47570
rect 48302 47518 48354 47570
rect 48750 47518 48802 47570
rect 57934 47518 57986 47570
rect 4286 47406 4338 47458
rect 10110 47406 10162 47458
rect 11342 47406 11394 47458
rect 19182 47406 19234 47458
rect 21534 47406 21586 47458
rect 21982 47406 22034 47458
rect 22654 47406 22706 47458
rect 23326 47406 23378 47458
rect 24782 47406 24834 47458
rect 28030 47406 28082 47458
rect 28702 47406 28754 47458
rect 29822 47406 29874 47458
rect 30158 47406 30210 47458
rect 30494 47406 30546 47458
rect 31054 47406 31106 47458
rect 31278 47406 31330 47458
rect 31614 47406 31666 47458
rect 31838 47406 31890 47458
rect 32062 47406 32114 47458
rect 32174 47406 32226 47458
rect 32734 47406 32786 47458
rect 33742 47406 33794 47458
rect 34302 47406 34354 47458
rect 35198 47406 35250 47458
rect 35758 47406 35810 47458
rect 36206 47406 36258 47458
rect 36990 47406 37042 47458
rect 37886 47406 37938 47458
rect 38334 47406 38386 47458
rect 40126 47406 40178 47458
rect 40350 47406 40402 47458
rect 40798 47406 40850 47458
rect 43598 47406 43650 47458
rect 44046 47406 44098 47458
rect 45166 47406 45218 47458
rect 45278 47406 45330 47458
rect 45726 47406 45778 47458
rect 46398 47406 46450 47458
rect 46622 47406 46674 47458
rect 55582 47406 55634 47458
rect 14254 47294 14306 47346
rect 16046 47294 16098 47346
rect 21758 47294 21810 47346
rect 23102 47294 23154 47346
rect 23662 47294 23714 47346
rect 25566 47294 25618 47346
rect 29598 47294 29650 47346
rect 30942 47294 30994 47346
rect 32958 47294 33010 47346
rect 34750 47294 34802 47346
rect 39790 47294 39842 47346
rect 41134 47294 41186 47346
rect 41246 47294 41298 47346
rect 42926 47294 42978 47346
rect 43374 47294 43426 47346
rect 44270 47294 44322 47346
rect 45054 47294 45106 47346
rect 46062 47294 46114 47346
rect 46958 47294 47010 47346
rect 47182 47294 47234 47346
rect 47630 47294 47682 47346
rect 47742 47294 47794 47346
rect 4734 47182 4786 47234
rect 11454 47182 11506 47234
rect 11566 47182 11618 47234
rect 11678 47182 11730 47234
rect 11790 47182 11842 47234
rect 20078 47182 20130 47234
rect 20526 47182 20578 47234
rect 21870 47182 21922 47234
rect 22094 47182 22146 47234
rect 22542 47182 22594 47234
rect 23214 47182 23266 47234
rect 24446 47182 24498 47234
rect 28142 47182 28194 47234
rect 28254 47182 28306 47234
rect 29262 47182 29314 47234
rect 29710 47182 29762 47234
rect 32510 47182 32562 47234
rect 34974 47182 35026 47234
rect 35086 47182 35138 47234
rect 35534 47182 35586 47234
rect 35646 47182 35698 47234
rect 37998 47182 38050 47234
rect 39230 47182 39282 47234
rect 41806 47182 41858 47234
rect 42702 47182 42754 47234
rect 42814 47182 42866 47234
rect 43262 47182 43314 47234
rect 43934 47182 43986 47234
rect 46286 47182 46338 47234
rect 47070 47182 47122 47234
rect 47966 47182 48018 47234
rect 19838 47014 19890 47066
rect 19942 47014 19994 47066
rect 20046 47014 20098 47066
rect 50558 47014 50610 47066
rect 50662 47014 50714 47066
rect 50766 47014 50818 47066
rect 8206 46846 8258 46898
rect 17838 46846 17890 46898
rect 27134 46846 27186 46898
rect 27470 46846 27522 46898
rect 27694 46846 27746 46898
rect 32286 46846 32338 46898
rect 35758 46846 35810 46898
rect 40798 46846 40850 46898
rect 41022 46846 41074 46898
rect 41582 46846 41634 46898
rect 44494 46846 44546 46898
rect 45950 46846 46002 46898
rect 2046 46734 2098 46786
rect 11678 46734 11730 46786
rect 28590 46734 28642 46786
rect 29934 46734 29986 46786
rect 33966 46734 34018 46786
rect 34078 46734 34130 46786
rect 34974 46734 35026 46786
rect 41134 46734 41186 46786
rect 44382 46734 44434 46786
rect 46174 46734 46226 46786
rect 47070 46734 47122 46786
rect 47630 46734 47682 46786
rect 1710 46622 1762 46674
rect 4622 46622 4674 46674
rect 7758 46622 7810 46674
rect 7982 46622 8034 46674
rect 8430 46622 8482 46674
rect 12350 46622 12402 46674
rect 17614 46622 17666 46674
rect 17838 46622 17890 46674
rect 18174 46622 18226 46674
rect 21310 46622 21362 46674
rect 24670 46622 24722 46674
rect 25342 46622 25394 46674
rect 25790 46622 25842 46674
rect 26574 46622 26626 46674
rect 26798 46622 26850 46674
rect 28142 46622 28194 46674
rect 28366 46622 28418 46674
rect 28702 46622 28754 46674
rect 29262 46622 29314 46674
rect 29710 46622 29762 46674
rect 30382 46622 30434 46674
rect 31278 46622 31330 46674
rect 31502 46622 31554 46674
rect 32062 46622 32114 46674
rect 34190 46622 34242 46674
rect 34638 46622 34690 46674
rect 35198 46622 35250 46674
rect 35982 46622 36034 46674
rect 36430 46622 36482 46674
rect 37438 46622 37490 46674
rect 41806 46622 41858 46674
rect 42030 46622 42082 46674
rect 42478 46622 42530 46674
rect 42926 46622 42978 46674
rect 43038 46622 43090 46674
rect 43486 46622 43538 46674
rect 44606 46622 44658 46674
rect 44942 46622 44994 46674
rect 45502 46622 45554 46674
rect 46062 46622 46114 46674
rect 46510 46622 46562 46674
rect 46734 46622 46786 46674
rect 47406 46622 47458 46674
rect 47966 46622 48018 46674
rect 53454 46622 53506 46674
rect 2494 46510 2546 46562
rect 2942 46510 2994 46562
rect 5294 46510 5346 46562
rect 7422 46510 7474 46562
rect 8094 46510 8146 46562
rect 9550 46510 9602 46562
rect 16942 46510 16994 46562
rect 18510 46510 18562 46562
rect 20638 46510 20690 46562
rect 21758 46510 21810 46562
rect 23886 46510 23938 46562
rect 27582 46510 27634 46562
rect 33182 46510 33234 46562
rect 34750 46510 34802 46562
rect 35870 46510 35922 46562
rect 36766 46510 36818 46562
rect 38222 46510 38274 46562
rect 40350 46510 40402 46562
rect 41694 46510 41746 46562
rect 42254 46510 42306 46562
rect 42702 46510 42754 46562
rect 47518 46510 47570 46562
rect 53230 46510 53282 46562
rect 25230 46398 25282 46450
rect 30382 46398 30434 46450
rect 33518 46398 33570 46450
rect 36542 46398 36594 46450
rect 36878 46398 36930 46450
rect 43710 46398 43762 46450
rect 44046 46398 44098 46450
rect 55358 46398 55410 46450
rect 4478 46230 4530 46282
rect 4582 46230 4634 46282
rect 4686 46230 4738 46282
rect 35198 46230 35250 46282
rect 35302 46230 35354 46282
rect 35406 46230 35458 46282
rect 8990 46062 9042 46114
rect 11678 46062 11730 46114
rect 21534 46062 21586 46114
rect 35870 46062 35922 46114
rect 43262 46062 43314 46114
rect 6414 45950 6466 46002
rect 10670 45950 10722 46002
rect 11566 45950 11618 46002
rect 16606 45950 16658 46002
rect 17166 45950 17218 46002
rect 22430 45950 22482 46002
rect 23662 45950 23714 46002
rect 28478 45950 28530 46002
rect 36430 45950 36482 46002
rect 46398 45950 46450 46002
rect 48526 45950 48578 46002
rect 55022 45950 55074 46002
rect 57822 45950 57874 46002
rect 1822 45838 1874 45890
rect 6750 45838 6802 45890
rect 6974 45838 7026 45890
rect 8206 45838 8258 45890
rect 10110 45838 10162 45890
rect 10334 45838 10386 45890
rect 10558 45838 10610 45890
rect 10782 45838 10834 45890
rect 11118 45838 11170 45890
rect 12910 45838 12962 45890
rect 13806 45838 13858 45890
rect 20078 45838 20130 45890
rect 21982 45838 22034 45890
rect 22318 45838 22370 45890
rect 22542 45838 22594 45890
rect 23214 45838 23266 45890
rect 23550 45838 23602 45890
rect 23774 45838 23826 45890
rect 27694 45838 27746 45890
rect 28030 45838 28082 45890
rect 34638 45838 34690 45890
rect 35310 45838 35362 45890
rect 36206 45838 36258 45890
rect 36878 45838 36930 45890
rect 42814 45838 42866 45890
rect 43822 45838 43874 45890
rect 44046 45838 44098 45890
rect 44830 45838 44882 45890
rect 45054 45838 45106 45890
rect 45390 45838 45442 45890
rect 45838 45838 45890 45890
rect 49198 45838 49250 45890
rect 52670 45838 52722 45890
rect 55582 45838 55634 45890
rect 2382 45726 2434 45778
rect 3166 45726 3218 45778
rect 6526 45726 6578 45778
rect 7534 45726 7586 45778
rect 7982 45726 8034 45778
rect 8430 45726 8482 45778
rect 8542 45726 8594 45778
rect 8878 45726 8930 45778
rect 8990 45726 9042 45778
rect 11230 45726 11282 45778
rect 12574 45726 12626 45778
rect 14478 45726 14530 45778
rect 19294 45726 19346 45778
rect 20750 45726 20802 45778
rect 21422 45726 21474 45778
rect 28478 45726 28530 45778
rect 30270 45726 30322 45778
rect 34974 45726 35026 45778
rect 35534 45726 35586 45778
rect 37214 45726 37266 45778
rect 37774 45726 37826 45778
rect 43710 45726 43762 45778
rect 2046 45614 2098 45666
rect 2718 45614 2770 45666
rect 6414 45614 6466 45666
rect 7422 45614 7474 45666
rect 7646 45614 7698 45666
rect 7758 45614 7810 45666
rect 12686 45614 12738 45666
rect 20526 45614 20578 45666
rect 20638 45614 20690 45666
rect 22094 45614 22146 45666
rect 23326 45614 23378 45666
rect 35310 45614 35362 45666
rect 37102 45614 37154 45666
rect 44942 45614 44994 45666
rect 19838 45446 19890 45498
rect 19942 45446 19994 45498
rect 20046 45446 20098 45498
rect 50558 45446 50610 45498
rect 50662 45446 50714 45498
rect 50766 45446 50818 45498
rect 8654 45278 8706 45330
rect 8878 45278 8930 45330
rect 18286 45278 18338 45330
rect 18734 45278 18786 45330
rect 18958 45278 19010 45330
rect 27358 45278 27410 45330
rect 27582 45278 27634 45330
rect 28030 45278 28082 45330
rect 31502 45278 31554 45330
rect 32622 45278 32674 45330
rect 33406 45278 33458 45330
rect 33518 45278 33570 45330
rect 34638 45278 34690 45330
rect 38558 45278 38610 45330
rect 44158 45278 44210 45330
rect 44382 45278 44434 45330
rect 45390 45278 45442 45330
rect 45838 45278 45890 45330
rect 46398 45278 46450 45330
rect 2046 45166 2098 45218
rect 5966 45166 6018 45218
rect 8990 45166 9042 45218
rect 11678 45166 11730 45218
rect 13470 45166 13522 45218
rect 18174 45166 18226 45218
rect 27134 45166 27186 45218
rect 28590 45166 28642 45218
rect 29374 45166 29426 45218
rect 31278 45166 31330 45218
rect 32398 45166 32450 45218
rect 33630 45166 33682 45218
rect 33966 45166 34018 45218
rect 35646 45166 35698 45218
rect 38894 45166 38946 45218
rect 41694 45166 41746 45218
rect 1710 45054 1762 45106
rect 5182 45054 5234 45106
rect 12350 45054 12402 45106
rect 14030 45054 14082 45106
rect 17726 45054 17778 45106
rect 18510 45054 18562 45106
rect 19070 45054 19122 45106
rect 23214 45054 23266 45106
rect 25342 45054 25394 45106
rect 28478 45054 28530 45106
rect 28702 45054 28754 45106
rect 29150 45054 29202 45106
rect 29822 45054 29874 45106
rect 31614 45054 31666 45106
rect 31950 45054 32002 45106
rect 32286 45054 32338 45106
rect 34078 45054 34130 45106
rect 34862 45054 34914 45106
rect 40910 45054 40962 45106
rect 44830 45054 44882 45106
rect 45054 45054 45106 45106
rect 45614 45054 45666 45106
rect 45950 45054 46002 45106
rect 2494 44942 2546 44994
rect 8094 44942 8146 44994
rect 9550 44942 9602 44994
rect 13582 44942 13634 44994
rect 14702 44942 14754 44994
rect 16830 44942 16882 44994
rect 18286 44942 18338 44994
rect 21758 44942 21810 44994
rect 27470 44942 27522 44994
rect 29598 44942 29650 44994
rect 30942 44942 30994 44994
rect 31390 44942 31442 44994
rect 37774 44942 37826 44994
rect 43822 44942 43874 44994
rect 44270 44942 44322 44994
rect 13246 44830 13298 44882
rect 4478 44662 4530 44714
rect 4582 44662 4634 44714
rect 4686 44662 4738 44714
rect 35198 44662 35250 44714
rect 35302 44662 35354 44714
rect 35406 44662 35458 44714
rect 12462 44494 12514 44546
rect 12910 44494 12962 44546
rect 19630 44494 19682 44546
rect 21310 44494 21362 44546
rect 42814 44494 42866 44546
rect 43374 44494 43426 44546
rect 6526 44382 6578 44434
rect 8654 44382 8706 44434
rect 9102 44382 9154 44434
rect 11118 44382 11170 44434
rect 11454 44382 11506 44434
rect 11902 44382 11954 44434
rect 21422 44382 21474 44434
rect 22094 44382 22146 44434
rect 27134 44382 27186 44434
rect 27582 44382 27634 44434
rect 31278 44382 31330 44434
rect 33406 44382 33458 44434
rect 34526 44382 34578 44434
rect 35870 44382 35922 44434
rect 42926 44382 42978 44434
rect 45502 44382 45554 44434
rect 57934 44382 57986 44434
rect 5742 44270 5794 44322
rect 12574 44270 12626 44322
rect 12798 44270 12850 44322
rect 17614 44270 17666 44322
rect 19406 44270 19458 44322
rect 19854 44270 19906 44322
rect 22654 44270 22706 44322
rect 25118 44270 25170 44322
rect 27022 44270 27074 44322
rect 27358 44270 27410 44322
rect 27918 44270 27970 44322
rect 28366 44270 28418 44322
rect 30494 44270 30546 44322
rect 35310 44270 35362 44322
rect 44942 44270 44994 44322
rect 48414 44270 48466 44322
rect 48526 44270 48578 44322
rect 49086 44270 49138 44322
rect 49422 44270 49474 44322
rect 49646 44270 49698 44322
rect 55582 44270 55634 44322
rect 1710 44158 1762 44210
rect 8990 44158 9042 44210
rect 14030 44158 14082 44210
rect 20190 44158 20242 44210
rect 20750 44158 20802 44210
rect 24222 44158 24274 44210
rect 24558 44158 24610 44210
rect 24894 44158 24946 44210
rect 26686 44158 26738 44210
rect 35086 44158 35138 44210
rect 38670 44158 38722 44210
rect 41582 44158 41634 44210
rect 48862 44158 48914 44210
rect 2046 44046 2098 44098
rect 2494 44046 2546 44098
rect 11566 44046 11618 44098
rect 12014 44046 12066 44098
rect 20078 44046 20130 44098
rect 21534 44046 21586 44098
rect 23998 44046 24050 44098
rect 26462 44046 26514 44098
rect 29262 44046 29314 44098
rect 34078 44046 34130 44098
rect 38334 44046 38386 44098
rect 43374 44046 43426 44098
rect 48750 44046 48802 44098
rect 49310 44046 49362 44098
rect 19838 43878 19890 43930
rect 19942 43878 19994 43930
rect 20046 43878 20098 43930
rect 50558 43878 50610 43930
rect 50662 43878 50714 43930
rect 50766 43878 50818 43930
rect 11454 43710 11506 43762
rect 12574 43710 12626 43762
rect 7646 43598 7698 43650
rect 7758 43598 7810 43650
rect 11790 43598 11842 43650
rect 12350 43598 12402 43650
rect 14478 43598 14530 43650
rect 21534 43598 21586 43650
rect 24110 43598 24162 43650
rect 24334 43598 24386 43650
rect 28926 43598 28978 43650
rect 29150 43598 29202 43650
rect 32286 43598 32338 43650
rect 33966 43598 34018 43650
rect 35982 43598 36034 43650
rect 37998 43598 38050 43650
rect 38782 43598 38834 43650
rect 39566 43598 39618 43650
rect 41358 43598 41410 43650
rect 42142 43598 42194 43650
rect 43822 43598 43874 43650
rect 47966 43598 48018 43650
rect 4286 43486 4338 43538
rect 11678 43486 11730 43538
rect 12238 43486 12290 43538
rect 12910 43486 12962 43538
rect 13246 43486 13298 43538
rect 13694 43486 13746 43538
rect 18174 43486 18226 43538
rect 18398 43486 18450 43538
rect 19182 43486 19234 43538
rect 22206 43486 22258 43538
rect 22654 43486 22706 43538
rect 22878 43486 22930 43538
rect 23102 43486 23154 43538
rect 23326 43486 23378 43538
rect 23774 43486 23826 43538
rect 23886 43486 23938 43538
rect 25566 43486 25618 43538
rect 29486 43486 29538 43538
rect 29934 43486 29986 43538
rect 33742 43486 33794 43538
rect 34750 43486 34802 43538
rect 35758 43486 35810 43538
rect 37774 43486 37826 43538
rect 39118 43486 39170 43538
rect 40910 43486 40962 43538
rect 41582 43486 41634 43538
rect 41918 43486 41970 43538
rect 42590 43486 42642 43538
rect 43038 43486 43090 43538
rect 46846 43486 46898 43538
rect 47070 43486 47122 43538
rect 47406 43486 47458 43538
rect 47518 43486 47570 43538
rect 48190 43486 48242 43538
rect 48862 43486 48914 43538
rect 4846 43374 4898 43426
rect 10446 43374 10498 43426
rect 16606 43374 16658 43426
rect 17502 43374 17554 43426
rect 18510 43374 18562 43426
rect 19406 43374 19458 43426
rect 22990 43374 23042 43426
rect 26350 43374 26402 43426
rect 28478 43374 28530 43426
rect 29374 43374 29426 43426
rect 30382 43374 30434 43426
rect 34414 43374 34466 43426
rect 35198 43374 35250 43426
rect 36430 43374 36482 43426
rect 41134 43374 41186 43426
rect 42366 43374 42418 43426
rect 45950 43374 46002 43426
rect 46398 43374 46450 43426
rect 47182 43374 47234 43426
rect 47742 43374 47794 43426
rect 49534 43374 49586 43426
rect 51662 43374 51714 43426
rect 1934 43262 1986 43314
rect 10334 43262 10386 43314
rect 11790 43262 11842 43314
rect 13022 43262 13074 43314
rect 13358 43262 13410 43314
rect 36206 43262 36258 43314
rect 36430 43262 36482 43314
rect 4478 43094 4530 43146
rect 4582 43094 4634 43146
rect 4686 43094 4738 43146
rect 35198 43094 35250 43146
rect 35302 43094 35354 43146
rect 35406 43094 35458 43146
rect 9662 42926 9714 42978
rect 9886 42926 9938 42978
rect 10110 42926 10162 42978
rect 11454 42926 11506 42978
rect 17950 42926 18002 42978
rect 18174 42926 18226 42978
rect 19406 42926 19458 42978
rect 19742 42926 19794 42978
rect 22094 42926 22146 42978
rect 57934 42926 57986 42978
rect 9326 42814 9378 42866
rect 10222 42814 10274 42866
rect 17726 42814 17778 42866
rect 19182 42814 19234 42866
rect 20750 42814 20802 42866
rect 21982 42814 22034 42866
rect 25790 42814 25842 42866
rect 27918 42814 27970 42866
rect 32510 42814 32562 42866
rect 49534 42814 49586 42866
rect 50206 42814 50258 42866
rect 50654 42814 50706 42866
rect 10670 42702 10722 42754
rect 13694 42702 13746 42754
rect 14030 42702 14082 42754
rect 19966 42702 20018 42754
rect 23774 42702 23826 42754
rect 23998 42702 24050 42754
rect 24334 42702 24386 42754
rect 24558 42702 24610 42754
rect 25006 42702 25058 42754
rect 26238 42702 26290 42754
rect 26686 42702 26738 42754
rect 26798 42702 26850 42754
rect 27134 42702 27186 42754
rect 27582 42702 27634 42754
rect 29598 42702 29650 42754
rect 30158 42702 30210 42754
rect 30718 42702 30770 42754
rect 31054 42702 31106 42754
rect 31390 42702 31442 42754
rect 32734 42702 32786 42754
rect 33182 42702 33234 42754
rect 33630 42702 33682 42754
rect 34078 42702 34130 42754
rect 34190 42702 34242 42754
rect 34638 42702 34690 42754
rect 34974 42702 35026 42754
rect 35086 42702 35138 42754
rect 36206 42702 36258 42754
rect 37662 42702 37714 42754
rect 38110 42702 38162 42754
rect 38334 42702 38386 42754
rect 38670 42702 38722 42754
rect 38894 42702 38946 42754
rect 39678 42702 39730 42754
rect 39902 42702 39954 42754
rect 40238 42702 40290 42754
rect 40574 42702 40626 42754
rect 40686 42702 40738 42754
rect 41358 42702 41410 42754
rect 41582 42702 41634 42754
rect 42478 42702 42530 42754
rect 42702 42702 42754 42754
rect 45390 42702 45442 42754
rect 45838 42702 45890 42754
rect 46062 42702 46114 42754
rect 46398 42702 46450 42754
rect 46622 42702 46674 42754
rect 46958 42702 47010 42754
rect 47294 42702 47346 42754
rect 47630 42702 47682 42754
rect 47854 42702 47906 42754
rect 48190 42702 48242 42754
rect 48414 42702 48466 42754
rect 48750 42702 48802 42754
rect 49086 42702 49138 42754
rect 49758 42702 49810 42754
rect 55582 42702 55634 42754
rect 1710 42590 1762 42642
rect 10894 42590 10946 42642
rect 11006 42590 11058 42642
rect 13918 42590 13970 42642
rect 22430 42590 22482 42642
rect 25230 42590 25282 42642
rect 26014 42590 26066 42642
rect 29710 42590 29762 42642
rect 31614 42590 31666 42642
rect 31950 42590 32002 42642
rect 33406 42590 33458 42642
rect 35870 42590 35922 42642
rect 36430 42590 36482 42642
rect 37326 42590 37378 42642
rect 39230 42590 39282 42642
rect 41022 42590 41074 42642
rect 41918 42590 41970 42642
rect 42254 42590 42306 42642
rect 44830 42590 44882 42642
rect 2046 42478 2098 42530
rect 2494 42478 2546 42530
rect 10222 42478 10274 42530
rect 18622 42478 18674 42530
rect 21646 42478 21698 42530
rect 22766 42478 22818 42530
rect 23102 42478 23154 42530
rect 23438 42478 23490 42530
rect 23886 42478 23938 42530
rect 24782 42478 24834 42530
rect 26350 42478 26402 42530
rect 27022 42478 27074 42530
rect 29934 42478 29986 42530
rect 31166 42478 31218 42530
rect 32958 42478 33010 42530
rect 33854 42478 33906 42530
rect 34750 42478 34802 42530
rect 36318 42478 36370 42530
rect 36990 42478 37042 42530
rect 37998 42478 38050 42530
rect 39118 42478 39170 42530
rect 40014 42478 40066 42530
rect 40910 42478 40962 42530
rect 41806 42478 41858 42530
rect 42366 42478 42418 42530
rect 45166 42478 45218 42530
rect 45726 42478 45778 42530
rect 46622 42478 46674 42530
rect 47406 42478 47458 42530
rect 48526 42478 48578 42530
rect 49310 42478 49362 42530
rect 49534 42478 49586 42530
rect 50542 42478 50594 42530
rect 19838 42310 19890 42362
rect 19942 42310 19994 42362
rect 20046 42310 20098 42362
rect 50558 42310 50610 42362
rect 50662 42310 50714 42362
rect 50766 42310 50818 42362
rect 10894 42142 10946 42194
rect 25230 42142 25282 42194
rect 26686 42142 26738 42194
rect 26910 42142 26962 42194
rect 35422 42142 35474 42194
rect 37886 42142 37938 42194
rect 39342 42142 39394 42194
rect 42254 42142 42306 42194
rect 45838 42142 45890 42194
rect 46510 42142 46562 42194
rect 48078 42142 48130 42194
rect 2046 42030 2098 42082
rect 9886 42030 9938 42082
rect 13246 42030 13298 42082
rect 18846 42030 18898 42082
rect 22318 42030 22370 42082
rect 24558 42030 24610 42082
rect 27134 42030 27186 42082
rect 27246 42030 27298 42082
rect 30830 42030 30882 42082
rect 41022 42030 41074 42082
rect 47518 42030 47570 42082
rect 49310 42030 49362 42082
rect 49534 42030 49586 42082
rect 1710 41918 1762 41970
rect 9774 41918 9826 41970
rect 10334 41918 10386 41970
rect 10782 41918 10834 41970
rect 11006 41918 11058 41970
rect 12574 41918 12626 41970
rect 19070 41918 19122 41970
rect 23102 41918 23154 41970
rect 23886 41918 23938 41970
rect 24334 41918 24386 41970
rect 25454 41918 25506 41970
rect 26126 41918 26178 41970
rect 26462 41918 26514 41970
rect 27694 41918 27746 41970
rect 29150 41918 29202 41970
rect 29262 41918 29314 41970
rect 29486 41918 29538 41970
rect 29598 41918 29650 41970
rect 30494 41918 30546 41970
rect 33406 41918 33458 41970
rect 34302 41918 34354 41970
rect 34862 41918 34914 41970
rect 35646 41918 35698 41970
rect 36766 41918 36818 41970
rect 37326 41918 37378 41970
rect 37550 41918 37602 41970
rect 38558 41918 38610 41970
rect 39006 41918 39058 41970
rect 39678 41918 39730 41970
rect 41246 41918 41298 41970
rect 41470 41918 41522 41970
rect 41582 41918 41634 41970
rect 46174 41918 46226 41970
rect 46734 41918 46786 41970
rect 47182 41918 47234 41970
rect 49086 41918 49138 41970
rect 49758 41918 49810 41970
rect 53454 41918 53506 41970
rect 2494 41806 2546 41858
rect 10558 41806 10610 41858
rect 15374 41806 15426 41858
rect 20190 41806 20242 41858
rect 23774 41806 23826 41858
rect 24110 41806 24162 41858
rect 29374 41806 29426 41858
rect 33966 41806 34018 41858
rect 36318 41806 36370 41858
rect 41358 41806 41410 41858
rect 49422 41806 49474 41858
rect 53230 41806 53282 41858
rect 9886 41694 9938 41746
rect 55358 41694 55410 41746
rect 4478 41526 4530 41578
rect 4582 41526 4634 41578
rect 4686 41526 4738 41578
rect 35198 41526 35250 41578
rect 35302 41526 35354 41578
rect 35406 41526 35458 41578
rect 10782 41358 10834 41410
rect 11006 41358 11058 41410
rect 11678 41358 11730 41410
rect 34414 41358 34466 41410
rect 34974 41358 35026 41410
rect 50990 41358 51042 41410
rect 57934 41358 57986 41410
rect 10110 41246 10162 41298
rect 15486 41246 15538 41298
rect 16046 41246 16098 41298
rect 21982 41246 22034 41298
rect 26574 41246 26626 41298
rect 27470 41246 27522 41298
rect 28030 41246 28082 41298
rect 28702 41246 28754 41298
rect 29150 41246 29202 41298
rect 32510 41246 32562 41298
rect 34414 41246 34466 41298
rect 38110 41246 38162 41298
rect 41806 41246 41858 41298
rect 43934 41246 43986 41298
rect 48638 41246 48690 41298
rect 51102 41246 51154 41298
rect 55022 41246 55074 41298
rect 10558 41134 10610 41186
rect 11230 41134 11282 41186
rect 15710 41134 15762 41186
rect 16606 41134 16658 41186
rect 19406 41134 19458 41186
rect 19966 41134 20018 41186
rect 24110 41134 24162 41186
rect 25566 41134 25618 41186
rect 29262 41134 29314 41186
rect 29710 41134 29762 41186
rect 35198 41134 35250 41186
rect 41134 41134 41186 41186
rect 45166 41134 45218 41186
rect 49198 41134 49250 41186
rect 51550 41134 51602 41186
rect 52670 41134 52722 41186
rect 55582 41134 55634 41186
rect 1710 41022 1762 41074
rect 2382 41022 2434 41074
rect 2718 41022 2770 41074
rect 11566 41022 11618 41074
rect 12238 41022 12290 41074
rect 18734 41022 18786 41074
rect 21870 41022 21922 41074
rect 22654 41022 22706 41074
rect 22990 41022 23042 41074
rect 24782 41022 24834 41074
rect 25790 41022 25842 41074
rect 27022 41022 27074 41074
rect 30382 41022 30434 41074
rect 2046 40910 2098 40962
rect 3166 40910 3218 40962
rect 10670 40910 10722 40962
rect 11790 40910 11842 40962
rect 12014 40910 12066 40962
rect 12686 40910 12738 40962
rect 16382 40910 16434 40962
rect 18622 40910 18674 40962
rect 19070 40910 19122 40962
rect 19630 40910 19682 40962
rect 19854 40910 19906 40962
rect 23550 40910 23602 40962
rect 25118 40910 25170 40962
rect 26126 40910 26178 40962
rect 34750 40910 34802 40962
rect 51438 40910 51490 40962
rect 19838 40742 19890 40794
rect 19942 40742 19994 40794
rect 20046 40742 20098 40794
rect 50558 40742 50610 40794
rect 50662 40742 50714 40794
rect 50766 40742 50818 40794
rect 2494 40574 2546 40626
rect 21086 40574 21138 40626
rect 21422 40574 21474 40626
rect 23102 40574 23154 40626
rect 23886 40574 23938 40626
rect 24446 40574 24498 40626
rect 24670 40574 24722 40626
rect 25342 40574 25394 40626
rect 26910 40574 26962 40626
rect 35310 40574 35362 40626
rect 37214 40574 37266 40626
rect 2046 40462 2098 40514
rect 16046 40462 16098 40514
rect 18622 40462 18674 40514
rect 22094 40462 22146 40514
rect 22766 40462 22818 40514
rect 23438 40462 23490 40514
rect 24334 40462 24386 40514
rect 25790 40462 25842 40514
rect 30606 40462 30658 40514
rect 34190 40462 34242 40514
rect 35758 40462 35810 40514
rect 36318 40462 36370 40514
rect 38446 40462 38498 40514
rect 49534 40462 49586 40514
rect 1710 40350 1762 40402
rect 2942 40350 2994 40402
rect 11230 40350 11282 40402
rect 16830 40350 16882 40402
rect 17838 40350 17890 40402
rect 21870 40350 21922 40402
rect 23998 40350 24050 40402
rect 26462 40350 26514 40402
rect 27246 40350 27298 40402
rect 33854 40350 33906 40402
rect 33966 40350 34018 40402
rect 34414 40350 34466 40402
rect 34862 40350 34914 40402
rect 34974 40350 35026 40402
rect 35198 40350 35250 40402
rect 36206 40350 36258 40402
rect 38670 40350 38722 40402
rect 38894 40350 38946 40402
rect 39006 40350 39058 40402
rect 39566 40350 39618 40402
rect 39678 40350 39730 40402
rect 39902 40350 39954 40402
rect 40014 40350 40066 40402
rect 41246 40350 41298 40402
rect 42030 40350 42082 40402
rect 44942 40350 44994 40402
rect 48750 40350 48802 40402
rect 53454 40350 53506 40402
rect 13918 40238 13970 40290
rect 17390 40238 17442 40290
rect 20750 40238 20802 40290
rect 34078 40238 34130 40290
rect 35086 40238 35138 40290
rect 35870 40238 35922 40290
rect 36878 40238 36930 40290
rect 38782 40238 38834 40290
rect 39790 40238 39842 40290
rect 44158 40238 44210 40290
rect 45614 40238 45666 40290
rect 47742 40238 47794 40290
rect 51662 40238 51714 40290
rect 17502 40126 17554 40178
rect 23886 40126 23938 40178
rect 55358 40126 55410 40178
rect 4478 39958 4530 40010
rect 4582 39958 4634 40010
rect 4686 39958 4738 40010
rect 35198 39958 35250 40010
rect 35302 39958 35354 40010
rect 35406 39958 35458 40010
rect 12910 39790 12962 39842
rect 42926 39790 42978 39842
rect 57934 39790 57986 39842
rect 11118 39678 11170 39730
rect 13582 39678 13634 39730
rect 16830 39678 16882 39730
rect 18958 39678 19010 39730
rect 19742 39678 19794 39730
rect 19966 39678 20018 39730
rect 20750 39678 20802 39730
rect 21422 39678 21474 39730
rect 23214 39678 23266 39730
rect 31278 39678 31330 39730
rect 32398 39678 32450 39730
rect 33966 39678 34018 39730
rect 36094 39678 36146 39730
rect 37886 39678 37938 39730
rect 40014 39678 40066 39730
rect 41582 39678 41634 39730
rect 43374 39678 43426 39730
rect 43486 39678 43538 39730
rect 47742 39678 47794 39730
rect 51438 39678 51490 39730
rect 10446 39566 10498 39618
rect 11006 39566 11058 39618
rect 11678 39566 11730 39618
rect 12686 39566 12738 39618
rect 16046 39566 16098 39618
rect 19294 39566 19346 39618
rect 19518 39566 19570 39618
rect 26798 39566 26850 39618
rect 30718 39566 30770 39618
rect 31390 39566 31442 39618
rect 33294 39566 33346 39618
rect 37214 39566 37266 39618
rect 40686 39566 40738 39618
rect 41470 39566 41522 39618
rect 41918 39566 41970 39618
rect 43038 39566 43090 39618
rect 45390 39566 45442 39618
rect 45950 39566 46002 39618
rect 46286 39566 46338 39618
rect 46958 39566 47010 39618
rect 48638 39566 48690 39618
rect 55582 39566 55634 39618
rect 1710 39454 1762 39506
rect 2046 39454 2098 39506
rect 12910 39454 12962 39506
rect 15710 39454 15762 39506
rect 19966 39454 20018 39506
rect 29822 39454 29874 39506
rect 31838 39454 31890 39506
rect 40910 39454 40962 39506
rect 47294 39454 47346 39506
rect 49310 39454 49362 39506
rect 55358 39454 55410 39506
rect 2494 39342 2546 39394
rect 13470 39342 13522 39394
rect 14030 39342 14082 39394
rect 15374 39342 15426 39394
rect 15598 39342 15650 39394
rect 20190 39342 20242 39394
rect 27470 39342 27522 39394
rect 30158 39342 30210 39394
rect 30942 39342 30994 39394
rect 31166 39342 31218 39394
rect 31726 39342 31778 39394
rect 41358 39342 41410 39394
rect 41694 39342 41746 39394
rect 45614 39342 45666 39394
rect 46174 39342 46226 39394
rect 46398 39342 46450 39394
rect 46510 39342 46562 39394
rect 47630 39342 47682 39394
rect 19838 39174 19890 39226
rect 19942 39174 19994 39226
rect 20046 39174 20098 39226
rect 50558 39174 50610 39226
rect 50662 39174 50714 39226
rect 50766 39174 50818 39226
rect 14590 39006 14642 39058
rect 15262 39006 15314 39058
rect 16046 39006 16098 39058
rect 17502 39006 17554 39058
rect 18062 39006 18114 39058
rect 18510 39006 18562 39058
rect 25454 39006 25506 39058
rect 31726 39006 31778 39058
rect 32174 39006 32226 39058
rect 32510 39006 32562 39058
rect 39342 39006 39394 39058
rect 49086 39006 49138 39058
rect 49198 39006 49250 39058
rect 49310 39006 49362 39058
rect 11902 38894 11954 38946
rect 22094 38894 22146 38946
rect 24670 38894 24722 38946
rect 29598 38894 29650 38946
rect 31166 38894 31218 38946
rect 39454 38894 39506 38946
rect 49646 38894 49698 38946
rect 4286 38782 4338 38834
rect 11230 38782 11282 38834
rect 15038 38782 15090 38834
rect 20414 38782 20466 38834
rect 20862 38782 20914 38834
rect 21310 38782 21362 38834
rect 30270 38782 30322 38834
rect 31390 38782 31442 38834
rect 31614 38782 31666 38834
rect 38334 38782 38386 38834
rect 41022 38782 41074 38834
rect 49422 38782 49474 38834
rect 53454 38782 53506 38834
rect 10670 38670 10722 38722
rect 10782 38670 10834 38722
rect 14030 38670 14082 38722
rect 15710 38670 15762 38722
rect 16606 38670 16658 38722
rect 24222 38670 24274 38722
rect 24558 38670 24610 38722
rect 27246 38670 27298 38722
rect 27470 38670 27522 38722
rect 30830 38670 30882 38722
rect 31502 38670 31554 38722
rect 33294 38670 33346 38722
rect 38894 38670 38946 38722
rect 53230 38670 53282 38722
rect 1934 38558 1986 38610
rect 15598 38558 15650 38610
rect 20862 38558 20914 38610
rect 40910 38558 40962 38610
rect 55358 38558 55410 38610
rect 4478 38390 4530 38442
rect 4582 38390 4634 38442
rect 4686 38390 4738 38442
rect 35198 38390 35250 38442
rect 35302 38390 35354 38442
rect 35406 38390 35458 38442
rect 13470 38222 13522 38274
rect 20750 38222 20802 38274
rect 22094 38222 22146 38274
rect 27582 38222 27634 38274
rect 33854 38222 33906 38274
rect 57934 38222 57986 38274
rect 9774 38110 9826 38162
rect 11902 38110 11954 38162
rect 18286 38110 18338 38162
rect 21758 38110 21810 38162
rect 23886 38110 23938 38162
rect 27134 38110 27186 38162
rect 27918 38110 27970 38162
rect 31390 38110 31442 38162
rect 33518 38110 33570 38162
rect 33966 38110 34018 38162
rect 38222 38110 38274 38162
rect 40350 38110 40402 38162
rect 43262 38110 43314 38162
rect 9102 37998 9154 38050
rect 13694 37998 13746 38050
rect 14478 37998 14530 38050
rect 14590 37998 14642 38050
rect 15710 37998 15762 38050
rect 16158 37998 16210 38050
rect 16718 37998 16770 38050
rect 17502 37998 17554 38050
rect 17950 37998 18002 38050
rect 18062 37998 18114 38050
rect 18398 37998 18450 38050
rect 18622 37998 18674 38050
rect 19854 37998 19906 38050
rect 20190 37998 20242 38050
rect 20414 37998 20466 38050
rect 22990 37998 23042 38050
rect 24334 37998 24386 38050
rect 28478 37998 28530 38050
rect 29374 37998 29426 38050
rect 30270 37998 30322 38050
rect 30606 37998 30658 38050
rect 37438 37998 37490 38050
rect 42254 37998 42306 38050
rect 47182 37998 47234 38050
rect 47518 37998 47570 38050
rect 55358 37998 55410 38050
rect 55582 37998 55634 38050
rect 1710 37886 1762 37938
rect 13470 37886 13522 37938
rect 17390 37886 17442 37938
rect 19518 37886 19570 37938
rect 22206 37886 22258 37938
rect 25006 37886 25058 37938
rect 30158 37886 30210 37938
rect 43822 37886 43874 37938
rect 46846 37886 46898 37938
rect 48526 37886 48578 37938
rect 2046 37774 2098 37826
rect 2494 37774 2546 37826
rect 16494 37774 16546 37826
rect 17278 37774 17330 37826
rect 19294 37774 19346 37826
rect 22094 37774 22146 37826
rect 22654 37774 22706 37826
rect 23326 37774 23378 37826
rect 27806 37774 27858 37826
rect 28142 37774 28194 37826
rect 28366 37774 28418 37826
rect 29150 37774 29202 37826
rect 29262 37774 29314 37826
rect 29598 37774 29650 37826
rect 29934 37774 29986 37826
rect 34526 37774 34578 37826
rect 34862 37774 34914 37826
rect 35422 37774 35474 37826
rect 42366 37774 42418 37826
rect 42478 37774 42530 37826
rect 42590 37774 42642 37826
rect 42702 37774 42754 37826
rect 43710 37774 43762 37826
rect 46734 37774 46786 37826
rect 47406 37774 47458 37826
rect 47630 37774 47682 37826
rect 47742 37774 47794 37826
rect 48414 37774 48466 37826
rect 19838 37606 19890 37658
rect 19942 37606 19994 37658
rect 20046 37606 20098 37658
rect 50558 37606 50610 37658
rect 50662 37606 50714 37658
rect 50766 37606 50818 37658
rect 17614 37438 17666 37490
rect 17838 37438 17890 37490
rect 18958 37438 19010 37490
rect 21870 37438 21922 37490
rect 22990 37438 23042 37490
rect 24334 37438 24386 37490
rect 26126 37438 26178 37490
rect 26238 37438 26290 37490
rect 33630 37438 33682 37490
rect 41470 37438 41522 37490
rect 49310 37438 49362 37490
rect 2046 37326 2098 37378
rect 11790 37326 11842 37378
rect 20974 37326 21026 37378
rect 21198 37326 21250 37378
rect 22094 37326 22146 37378
rect 22766 37326 22818 37378
rect 24558 37326 24610 37378
rect 25342 37326 25394 37378
rect 29150 37326 29202 37378
rect 30382 37326 30434 37378
rect 30494 37326 30546 37378
rect 30942 37326 30994 37378
rect 31390 37326 31442 37378
rect 31502 37326 31554 37378
rect 34974 37326 35026 37378
rect 42590 37326 42642 37378
rect 1710 37214 1762 37266
rect 16718 37214 16770 37266
rect 18062 37214 18114 37266
rect 18398 37214 18450 37266
rect 18622 37214 18674 37266
rect 18846 37214 18898 37266
rect 20078 37214 20130 37266
rect 20526 37214 20578 37266
rect 22206 37214 22258 37266
rect 22654 37214 22706 37266
rect 23662 37214 23714 37266
rect 24110 37214 24162 37266
rect 24670 37214 24722 37266
rect 25454 37214 25506 37266
rect 25678 37214 25730 37266
rect 26350 37214 26402 37266
rect 29822 37214 29874 37266
rect 30158 37214 30210 37266
rect 34302 37214 34354 37266
rect 37438 37214 37490 37266
rect 41918 37214 41970 37266
rect 45166 37214 45218 37266
rect 48862 37214 48914 37266
rect 48974 37214 49026 37266
rect 49198 37214 49250 37266
rect 53454 37214 53506 37266
rect 2494 37102 2546 37154
rect 10334 37102 10386 37154
rect 17950 37102 18002 37154
rect 18958 37102 19010 37154
rect 19406 37102 19458 37154
rect 20862 37102 20914 37154
rect 21646 37102 21698 37154
rect 27022 37102 27074 37154
rect 37102 37102 37154 37154
rect 38222 37102 38274 37154
rect 40350 37102 40402 37154
rect 41134 37102 41186 37154
rect 44718 37102 44770 37154
rect 45838 37102 45890 37154
rect 47966 37102 48018 37154
rect 49086 37102 49138 37154
rect 10222 36990 10274 37042
rect 19518 36990 19570 37042
rect 25342 36990 25394 37042
rect 30830 36990 30882 37042
rect 31502 36990 31554 37042
rect 55358 36990 55410 37042
rect 4478 36822 4530 36874
rect 4582 36822 4634 36874
rect 4686 36822 4738 36874
rect 35198 36822 35250 36874
rect 35302 36822 35354 36874
rect 35406 36822 35458 36874
rect 16830 36654 16882 36706
rect 50430 36654 50482 36706
rect 57934 36654 57986 36706
rect 1934 36542 1986 36594
rect 4846 36542 4898 36594
rect 9214 36542 9266 36594
rect 11342 36542 11394 36594
rect 14254 36542 14306 36594
rect 16382 36542 16434 36594
rect 17502 36542 17554 36594
rect 19630 36542 19682 36594
rect 23662 36542 23714 36594
rect 24446 36542 24498 36594
rect 27470 36542 27522 36594
rect 29262 36542 29314 36594
rect 35086 36542 35138 36594
rect 43486 36542 43538 36594
rect 55022 36542 55074 36594
rect 4174 36430 4226 36482
rect 8430 36430 8482 36482
rect 13470 36430 13522 36482
rect 20414 36430 20466 36482
rect 21310 36430 21362 36482
rect 25902 36430 25954 36482
rect 29374 36430 29426 36482
rect 29822 36430 29874 36482
rect 30158 36430 30210 36482
rect 30718 36430 30770 36482
rect 31054 36430 31106 36482
rect 32174 36430 32226 36482
rect 35646 36430 35698 36482
rect 36318 36430 36370 36482
rect 42254 36430 42306 36482
rect 42814 36430 42866 36482
rect 46174 36430 46226 36482
rect 52782 36430 52834 36482
rect 55582 36430 55634 36482
rect 16718 36318 16770 36370
rect 21870 36318 21922 36370
rect 22206 36318 22258 36370
rect 22654 36318 22706 36370
rect 22766 36318 22818 36370
rect 25678 36318 25730 36370
rect 27246 36318 27298 36370
rect 32958 36318 33010 36370
rect 37214 36318 37266 36370
rect 42590 36318 42642 36370
rect 44270 36318 44322 36370
rect 48750 36318 48802 36370
rect 50542 36318 50594 36370
rect 50990 36318 51042 36370
rect 12910 36206 12962 36258
rect 16830 36206 16882 36258
rect 21422 36206 21474 36258
rect 21646 36206 21698 36258
rect 22430 36206 22482 36258
rect 23214 36206 23266 36258
rect 24894 36206 24946 36258
rect 28590 36206 28642 36258
rect 29150 36206 29202 36258
rect 30382 36206 30434 36258
rect 30830 36206 30882 36258
rect 35870 36206 35922 36258
rect 35982 36206 36034 36258
rect 36094 36206 36146 36258
rect 43374 36206 43426 36258
rect 44158 36206 44210 36258
rect 50878 36206 50930 36258
rect 52110 36206 52162 36258
rect 19838 36038 19890 36090
rect 19942 36038 19994 36090
rect 20046 36038 20098 36090
rect 50558 36038 50610 36090
rect 50662 36038 50714 36090
rect 50766 36038 50818 36090
rect 2718 35870 2770 35922
rect 18062 35870 18114 35922
rect 20750 35870 20802 35922
rect 23550 35870 23602 35922
rect 23998 35870 24050 35922
rect 26014 35870 26066 35922
rect 26462 35870 26514 35922
rect 26910 35870 26962 35922
rect 27358 35870 27410 35922
rect 33518 35870 33570 35922
rect 33630 35870 33682 35922
rect 33742 35870 33794 35922
rect 34414 35870 34466 35922
rect 39790 35870 39842 35922
rect 45166 35870 45218 35922
rect 45502 35870 45554 35922
rect 45838 35870 45890 35922
rect 46286 35870 46338 35922
rect 46398 35870 46450 35922
rect 46510 35870 46562 35922
rect 47966 35870 48018 35922
rect 48078 35870 48130 35922
rect 2046 35758 2098 35810
rect 14366 35758 14418 35810
rect 17502 35758 17554 35810
rect 18958 35758 19010 35810
rect 19406 35758 19458 35810
rect 19742 35758 19794 35810
rect 20414 35758 20466 35810
rect 22990 35758 23042 35810
rect 30382 35758 30434 35810
rect 33182 35758 33234 35810
rect 34526 35758 34578 35810
rect 35982 35758 36034 35810
rect 38446 35758 38498 35810
rect 38782 35758 38834 35810
rect 39454 35758 39506 35810
rect 41022 35758 41074 35810
rect 46846 35758 46898 35810
rect 49534 35758 49586 35810
rect 1710 35646 1762 35698
rect 2382 35646 2434 35698
rect 10558 35646 10610 35698
rect 10782 35646 10834 35698
rect 11790 35646 11842 35698
rect 12238 35646 12290 35698
rect 12686 35646 12738 35698
rect 13582 35646 13634 35698
rect 17390 35646 17442 35698
rect 18398 35646 18450 35698
rect 21422 35646 21474 35698
rect 22318 35646 22370 35698
rect 22654 35646 22706 35698
rect 25790 35646 25842 35698
rect 29598 35646 29650 35698
rect 33406 35646 33458 35698
rect 35310 35646 35362 35698
rect 39678 35646 39730 35698
rect 39902 35646 39954 35698
rect 40126 35646 40178 35698
rect 40910 35646 40962 35698
rect 41358 35646 41410 35698
rect 46622 35646 46674 35698
rect 47630 35646 47682 35698
rect 47742 35646 47794 35698
rect 48750 35646 48802 35698
rect 53454 35646 53506 35698
rect 3166 35534 3218 35586
rect 10222 35534 10274 35586
rect 13134 35534 13186 35586
rect 16494 35534 16546 35586
rect 21646 35534 21698 35586
rect 22094 35534 22146 35586
rect 22542 35534 22594 35586
rect 32510 35534 32562 35586
rect 38110 35534 38162 35586
rect 42142 35534 42194 35586
rect 44270 35534 44322 35586
rect 44718 35534 44770 35586
rect 47966 35534 48018 35586
rect 51662 35534 51714 35586
rect 53230 35534 53282 35586
rect 10110 35422 10162 35474
rect 11118 35422 11170 35474
rect 55358 35422 55410 35474
rect 4478 35254 4530 35306
rect 4582 35254 4634 35306
rect 4686 35254 4738 35306
rect 35198 35254 35250 35306
rect 35302 35254 35354 35306
rect 35406 35254 35458 35306
rect 16830 35086 16882 35138
rect 16942 35086 16994 35138
rect 17278 35086 17330 35138
rect 32062 35086 32114 35138
rect 33294 35086 33346 35138
rect 37102 35086 37154 35138
rect 37438 35086 37490 35138
rect 38110 35086 38162 35138
rect 43262 35086 43314 35138
rect 44942 35086 44994 35138
rect 56590 35086 56642 35138
rect 2494 34974 2546 35026
rect 9102 34974 9154 35026
rect 11230 34974 11282 35026
rect 12462 34974 12514 35026
rect 16382 34974 16434 35026
rect 17726 34974 17778 35026
rect 18510 34974 18562 35026
rect 19070 34974 19122 35026
rect 22654 34974 22706 35026
rect 30606 34974 30658 35026
rect 36542 34974 36594 35026
rect 37214 34974 37266 35026
rect 41694 34974 41746 35026
rect 47070 34974 47122 35026
rect 49198 34974 49250 35026
rect 8430 34862 8482 34914
rect 13470 34862 13522 34914
rect 17166 34862 17218 34914
rect 18062 34862 18114 34914
rect 18734 34862 18786 34914
rect 21646 34862 21698 34914
rect 22318 34862 22370 34914
rect 25566 34862 25618 34914
rect 26238 34862 26290 34914
rect 26910 34862 26962 34914
rect 27022 34862 27074 34914
rect 27470 34862 27522 34914
rect 27694 34862 27746 34914
rect 27918 34862 27970 34914
rect 31278 34862 31330 34914
rect 32510 34862 32562 34914
rect 34302 34862 34354 34914
rect 34750 34862 34802 34914
rect 35086 34862 35138 34914
rect 36094 34862 36146 34914
rect 38446 34862 38498 34914
rect 41246 34862 41298 34914
rect 41582 34862 41634 34914
rect 42254 34862 42306 34914
rect 42590 34862 42642 34914
rect 42702 34862 42754 34914
rect 45726 34862 45778 34914
rect 46398 34862 46450 34914
rect 55582 34862 55634 34914
rect 1710 34750 1762 34802
rect 14254 34750 14306 34802
rect 18286 34750 18338 34802
rect 20638 34750 20690 34802
rect 20750 34750 20802 34802
rect 21758 34750 21810 34802
rect 24782 34750 24834 34802
rect 28030 34750 28082 34802
rect 31614 34750 31666 34802
rect 31950 34750 32002 34802
rect 33182 34750 33234 34802
rect 35422 34750 35474 34802
rect 35758 34750 35810 34802
rect 38782 34750 38834 34802
rect 39678 34750 39730 34802
rect 40462 34750 40514 34802
rect 43150 34750 43202 34802
rect 43934 34750 43986 34802
rect 44830 34750 44882 34802
rect 2046 34638 2098 34690
rect 2942 34638 2994 34690
rect 12126 34638 12178 34690
rect 12910 34638 12962 34690
rect 20414 34638 20466 34690
rect 21870 34638 21922 34690
rect 25902 34638 25954 34690
rect 27246 34638 27298 34690
rect 28478 34638 28530 34690
rect 29262 34638 29314 34690
rect 32062 34638 32114 34690
rect 32846 34638 32898 34690
rect 33294 34638 33346 34690
rect 33854 34638 33906 34690
rect 35310 34638 35362 34690
rect 35870 34638 35922 34690
rect 37662 34638 37714 34690
rect 38222 34638 38274 34690
rect 38670 34638 38722 34690
rect 39342 34638 39394 34690
rect 40126 34638 40178 34690
rect 41358 34638 41410 34690
rect 41694 34638 41746 34690
rect 42366 34638 42418 34690
rect 42478 34638 42530 34690
rect 43262 34638 43314 34690
rect 43598 34638 43650 34690
rect 43822 34638 43874 34690
rect 44942 34638 44994 34690
rect 45950 34638 46002 34690
rect 19838 34470 19890 34522
rect 19942 34470 19994 34522
rect 20046 34470 20098 34522
rect 50558 34470 50610 34522
rect 50662 34470 50714 34522
rect 50766 34470 50818 34522
rect 15150 34302 15202 34354
rect 16158 34302 16210 34354
rect 24334 34302 24386 34354
rect 26574 34302 26626 34354
rect 27694 34302 27746 34354
rect 30942 34302 30994 34354
rect 31726 34302 31778 34354
rect 33854 34302 33906 34354
rect 34302 34302 34354 34354
rect 38782 34302 38834 34354
rect 39678 34302 39730 34354
rect 39790 34302 39842 34354
rect 41246 34302 41298 34354
rect 45950 34302 46002 34354
rect 46510 34302 46562 34354
rect 47406 34302 47458 34354
rect 47630 34302 47682 34354
rect 15710 34190 15762 34242
rect 23998 34190 24050 34242
rect 25230 34190 25282 34242
rect 26238 34190 26290 34242
rect 28030 34190 28082 34242
rect 29486 34190 29538 34242
rect 31278 34190 31330 34242
rect 39342 34190 39394 34242
rect 39454 34190 39506 34242
rect 40014 34190 40066 34242
rect 40126 34190 40178 34242
rect 40910 34190 40962 34242
rect 41022 34190 41074 34242
rect 42254 34190 42306 34242
rect 45614 34190 45666 34242
rect 46286 34190 46338 34242
rect 46734 34190 46786 34242
rect 46846 34190 46898 34242
rect 49534 34190 49586 34242
rect 4286 34078 4338 34130
rect 10558 34078 10610 34130
rect 11006 34078 11058 34130
rect 11790 34078 11842 34130
rect 12238 34078 12290 34130
rect 13022 34078 13074 34130
rect 13582 34078 13634 34130
rect 14030 34078 14082 34130
rect 16270 34078 16322 34130
rect 23662 34078 23714 34130
rect 24222 34078 24274 34130
rect 24446 34078 24498 34130
rect 24670 34078 24722 34130
rect 25454 34078 25506 34130
rect 25678 34078 25730 34130
rect 25790 34078 25842 34130
rect 26910 34078 26962 34130
rect 28366 34078 28418 34130
rect 28926 34078 28978 34130
rect 29598 34078 29650 34130
rect 29822 34078 29874 34130
rect 34414 34078 34466 34130
rect 34750 34078 34802 34130
rect 35086 34078 35138 34130
rect 35534 34078 35586 34130
rect 41470 34078 41522 34130
rect 47742 34078 47794 34130
rect 48750 34078 48802 34130
rect 53454 34078 53506 34130
rect 4734 33966 4786 34018
rect 13246 33966 13298 34018
rect 23214 33966 23266 34018
rect 23550 33966 23602 34018
rect 25566 33966 25618 34018
rect 27022 33966 27074 34018
rect 28590 33966 28642 34018
rect 32398 33966 32450 34018
rect 33294 33966 33346 34018
rect 34638 33966 34690 34018
rect 36206 33966 36258 34018
rect 38334 33966 38386 34018
rect 44382 33966 44434 34018
rect 44830 33966 44882 34018
rect 48190 33966 48242 34018
rect 51662 33966 51714 34018
rect 1934 33854 1986 33906
rect 11118 33854 11170 33906
rect 15486 33854 15538 33906
rect 16158 33854 16210 33906
rect 55358 33854 55410 33906
rect 4478 33686 4530 33738
rect 4582 33686 4634 33738
rect 4686 33686 4738 33738
rect 35198 33686 35250 33738
rect 35302 33686 35354 33738
rect 35406 33686 35458 33738
rect 14590 33518 14642 33570
rect 27470 33518 27522 33570
rect 34414 33518 34466 33570
rect 48078 33518 48130 33570
rect 48862 33518 48914 33570
rect 49422 33518 49474 33570
rect 50542 33518 50594 33570
rect 57934 33518 57986 33570
rect 11118 33406 11170 33458
rect 18062 33406 18114 33458
rect 18510 33406 18562 33458
rect 21982 33406 22034 33458
rect 23102 33406 23154 33458
rect 25230 33406 25282 33458
rect 32622 33406 32674 33458
rect 35982 33406 36034 33458
rect 8206 33294 8258 33346
rect 14926 33294 14978 33346
rect 15150 33294 15202 33346
rect 18846 33294 18898 33346
rect 19630 33294 19682 33346
rect 25902 33294 25954 33346
rect 27694 33294 27746 33346
rect 27918 33294 27970 33346
rect 28590 33294 28642 33346
rect 30046 33294 30098 33346
rect 31502 33294 31554 33346
rect 34862 33294 34914 33346
rect 35086 33294 35138 33346
rect 36542 33294 36594 33346
rect 36878 33294 36930 33346
rect 37214 33294 37266 33346
rect 37662 33294 37714 33346
rect 40910 33294 40962 33346
rect 41246 33294 41298 33346
rect 46062 33294 46114 33346
rect 46398 33294 46450 33346
rect 47966 33294 48018 33346
rect 48750 33294 48802 33346
rect 49534 33294 49586 33346
rect 49758 33294 49810 33346
rect 50094 33294 50146 33346
rect 50654 33294 50706 33346
rect 55582 33294 55634 33346
rect 1710 33182 1762 33234
rect 8990 33182 9042 33234
rect 14702 33182 14754 33234
rect 16942 33182 16994 33234
rect 27134 33182 27186 33234
rect 29374 33182 29426 33234
rect 32174 33182 32226 33234
rect 34974 33182 35026 33234
rect 55358 33182 55410 33234
rect 2046 33070 2098 33122
rect 2494 33070 2546 33122
rect 19182 33070 19234 33122
rect 26574 33070 26626 33122
rect 28366 33070 28418 33122
rect 28478 33070 28530 33122
rect 29150 33070 29202 33122
rect 29262 33070 29314 33122
rect 29598 33070 29650 33122
rect 30158 33070 30210 33122
rect 30382 33070 30434 33122
rect 30830 33070 30882 33122
rect 31166 33070 31218 33122
rect 31838 33070 31890 33122
rect 34190 33070 34242 33122
rect 34302 33070 34354 33122
rect 35534 33070 35586 33122
rect 35870 33070 35922 33122
rect 36094 33070 36146 33122
rect 37102 33070 37154 33122
rect 38110 33070 38162 33122
rect 39566 33070 39618 33122
rect 40686 33070 40738 33122
rect 41022 33070 41074 33122
rect 43374 33070 43426 33122
rect 46286 33070 46338 33122
rect 47742 33070 47794 33122
rect 48078 33070 48130 33122
rect 48862 33070 48914 33122
rect 49422 33070 49474 33122
rect 49982 33070 50034 33122
rect 50542 33070 50594 33122
rect 19838 32902 19890 32954
rect 19942 32902 19994 32954
rect 20046 32902 20098 32954
rect 50558 32902 50610 32954
rect 50662 32902 50714 32954
rect 50766 32902 50818 32954
rect 9438 32734 9490 32786
rect 9662 32734 9714 32786
rect 9886 32734 9938 32786
rect 14926 32734 14978 32786
rect 16158 32734 16210 32786
rect 18734 32734 18786 32786
rect 22430 32734 22482 32786
rect 24782 32734 24834 32786
rect 25118 32734 25170 32786
rect 30942 32734 30994 32786
rect 34190 32734 34242 32786
rect 34414 32734 34466 32786
rect 35198 32734 35250 32786
rect 35534 32734 35586 32786
rect 43038 32734 43090 32786
rect 2046 32622 2098 32674
rect 15150 32622 15202 32674
rect 16718 32622 16770 32674
rect 17614 32622 17666 32674
rect 17726 32622 17778 32674
rect 17950 32622 18002 32674
rect 19854 32622 19906 32674
rect 22542 32622 22594 32674
rect 24558 32622 24610 32674
rect 25342 32622 25394 32674
rect 26238 32622 26290 32674
rect 26574 32622 26626 32674
rect 29038 32622 29090 32674
rect 31278 32622 31330 32674
rect 33630 32622 33682 32674
rect 34750 32622 34802 32674
rect 35982 32622 36034 32674
rect 1710 32510 1762 32562
rect 11790 32510 11842 32562
rect 12126 32510 12178 32562
rect 12686 32510 12738 32562
rect 13134 32510 13186 32562
rect 13470 32510 13522 32562
rect 13582 32510 13634 32562
rect 14590 32510 14642 32562
rect 16494 32510 16546 32562
rect 18062 32510 18114 32562
rect 18510 32510 18562 32562
rect 19182 32510 19234 32562
rect 22766 32510 22818 32562
rect 22990 32510 23042 32562
rect 24446 32510 24498 32562
rect 25454 32510 25506 32562
rect 29822 32510 29874 32562
rect 31614 32510 31666 32562
rect 32174 32510 32226 32562
rect 33182 32510 33234 32562
rect 35422 32510 35474 32562
rect 35646 32510 35698 32562
rect 36318 32510 36370 32562
rect 36542 32510 36594 32562
rect 37438 32510 37490 32562
rect 43710 32510 43762 32562
rect 47070 32510 47122 32562
rect 53454 32510 53506 32562
rect 2494 32398 2546 32450
rect 8990 32398 9042 32450
rect 9998 32398 10050 32450
rect 15598 32398 15650 32450
rect 18622 32398 18674 32450
rect 21982 32398 22034 32450
rect 22430 32398 22482 32450
rect 23438 32398 23490 32450
rect 24222 32398 24274 32450
rect 26014 32398 26066 32450
rect 26910 32398 26962 32450
rect 30718 32398 30770 32450
rect 36430 32398 36482 32450
rect 38222 32398 38274 32450
rect 40350 32398 40402 32450
rect 43262 32398 43314 32450
rect 44158 32398 44210 32450
rect 46286 32398 46338 32450
rect 49198 32398 49250 32450
rect 8878 32286 8930 32338
rect 12014 32286 12066 32338
rect 14814 32286 14866 32338
rect 55358 32286 55410 32338
rect 4478 32118 4530 32170
rect 4582 32118 4634 32170
rect 4686 32118 4738 32170
rect 35198 32118 35250 32170
rect 35302 32118 35354 32170
rect 35406 32118 35458 32170
rect 14030 31950 14082 32002
rect 16270 31950 16322 32002
rect 21646 31950 21698 32002
rect 21982 31950 22034 32002
rect 24446 31950 24498 32002
rect 24782 31950 24834 32002
rect 36990 31950 37042 32002
rect 1934 31838 1986 31890
rect 4846 31838 4898 31890
rect 8654 31838 8706 31890
rect 10782 31838 10834 31890
rect 11678 31838 11730 31890
rect 14702 31838 14754 31890
rect 16718 31838 16770 31890
rect 18846 31838 18898 31890
rect 23102 31838 23154 31890
rect 24894 31838 24946 31890
rect 25678 31838 25730 31890
rect 37326 31838 37378 31890
rect 39006 31838 39058 31890
rect 44046 31838 44098 31890
rect 45502 31838 45554 31890
rect 50542 31838 50594 31890
rect 55022 31838 55074 31890
rect 57934 31838 57986 31890
rect 4174 31726 4226 31778
rect 7982 31726 8034 31778
rect 11342 31726 11394 31778
rect 12126 31726 12178 31778
rect 14478 31726 14530 31778
rect 15374 31726 15426 31778
rect 15598 31726 15650 31778
rect 15822 31726 15874 31778
rect 19630 31726 19682 31778
rect 27134 31726 27186 31778
rect 29374 31726 29426 31778
rect 34974 31726 35026 31778
rect 35310 31726 35362 31778
rect 37550 31726 37602 31778
rect 39454 31726 39506 31778
rect 39678 31726 39730 31778
rect 40014 31726 40066 31778
rect 41134 31726 41186 31778
rect 45614 31726 45666 31778
rect 46510 31726 46562 31778
rect 47630 31726 47682 31778
rect 52670 31726 52722 31778
rect 55582 31726 55634 31778
rect 14142 31614 14194 31666
rect 22654 31614 22706 31666
rect 25230 31614 25282 31666
rect 26350 31614 26402 31666
rect 26910 31614 26962 31666
rect 28590 31614 28642 31666
rect 29934 31614 29986 31666
rect 39902 31614 39954 31666
rect 41918 31614 41970 31666
rect 48414 31614 48466 31666
rect 12686 31502 12738 31554
rect 13694 31502 13746 31554
rect 14030 31502 14082 31554
rect 15038 31502 15090 31554
rect 21758 31502 21810 31554
rect 22318 31502 22370 31554
rect 23550 31502 23602 31554
rect 23998 31502 24050 31554
rect 24558 31502 24610 31554
rect 25454 31502 25506 31554
rect 25678 31502 25730 31554
rect 25790 31502 25842 31554
rect 26238 31502 26290 31554
rect 26798 31502 26850 31554
rect 27470 31502 27522 31554
rect 27694 31502 27746 31554
rect 27806 31502 27858 31554
rect 28142 31502 28194 31554
rect 35422 31502 35474 31554
rect 35534 31502 35586 31554
rect 35758 31502 35810 31554
rect 36318 31502 36370 31554
rect 38894 31502 38946 31554
rect 39118 31502 39170 31554
rect 45166 31502 45218 31554
rect 45390 31502 45442 31554
rect 45838 31502 45890 31554
rect 46286 31502 46338 31554
rect 46958 31502 47010 31554
rect 47294 31502 47346 31554
rect 19838 31334 19890 31386
rect 19942 31334 19994 31386
rect 20046 31334 20098 31386
rect 50558 31334 50610 31386
rect 50662 31334 50714 31386
rect 50766 31334 50818 31386
rect 2046 31166 2098 31218
rect 16046 31166 16098 31218
rect 31502 31166 31554 31218
rect 32174 31166 32226 31218
rect 38222 31166 38274 31218
rect 39006 31166 39058 31218
rect 41246 31166 41298 31218
rect 42142 31166 42194 31218
rect 42254 31166 42306 31218
rect 42702 31166 42754 31218
rect 45726 31166 45778 31218
rect 46174 31166 46226 31218
rect 2718 31054 2770 31106
rect 14926 31054 14978 31106
rect 16606 31054 16658 31106
rect 17502 31054 17554 31106
rect 17614 31054 17666 31106
rect 20862 31054 20914 31106
rect 23550 31054 23602 31106
rect 24110 31054 24162 31106
rect 30830 31054 30882 31106
rect 30942 31054 30994 31106
rect 31838 31054 31890 31106
rect 32510 31054 32562 31106
rect 33854 31054 33906 31106
rect 36318 31054 36370 31106
rect 36430 31054 36482 31106
rect 50766 31054 50818 31106
rect 1710 30942 1762 30994
rect 2382 30942 2434 30994
rect 10110 30942 10162 30994
rect 10558 30942 10610 30994
rect 11230 30942 11282 30994
rect 11902 30942 11954 30994
rect 15598 30942 15650 30994
rect 16382 30942 16434 30994
rect 20078 30942 20130 30994
rect 24446 30942 24498 30994
rect 25230 30942 25282 30994
rect 31166 30942 31218 30994
rect 33070 30942 33122 30994
rect 38110 30942 38162 30994
rect 38334 30942 38386 30994
rect 38670 30942 38722 30994
rect 39342 30942 39394 30994
rect 41358 30942 41410 30994
rect 41582 30942 41634 30994
rect 42030 30942 42082 30994
rect 42590 30942 42642 30994
rect 42814 30942 42866 30994
rect 43150 30942 43202 30994
rect 45166 30942 45218 30994
rect 45614 30942 45666 30994
rect 45838 30942 45890 30994
rect 47406 30942 47458 30994
rect 47854 30942 47906 30994
rect 48078 30942 48130 30994
rect 49086 30942 49138 30994
rect 3166 30830 3218 30882
rect 10894 30830 10946 30882
rect 12462 30830 12514 30882
rect 12798 30830 12850 30882
rect 22990 30830 23042 30882
rect 23214 30830 23266 30882
rect 27246 30830 27298 30882
rect 35982 30830 36034 30882
rect 36990 30830 37042 30882
rect 39566 30830 39618 30882
rect 46510 30830 46562 30882
rect 46734 30830 46786 30882
rect 47182 30830 47234 30882
rect 47966 30830 48018 30882
rect 10334 30718 10386 30770
rect 17502 30718 17554 30770
rect 36430 30718 36482 30770
rect 41246 30718 41298 30770
rect 4478 30550 4530 30602
rect 4582 30550 4634 30602
rect 4686 30550 4738 30602
rect 35198 30550 35250 30602
rect 35302 30550 35354 30602
rect 35406 30550 35458 30602
rect 42702 30382 42754 30434
rect 46734 30382 46786 30434
rect 2494 30270 2546 30322
rect 10782 30270 10834 30322
rect 16382 30270 16434 30322
rect 19406 30270 19458 30322
rect 23774 30270 23826 30322
rect 25902 30270 25954 30322
rect 29486 30270 29538 30322
rect 29822 30270 29874 30322
rect 31166 30270 31218 30322
rect 35198 30270 35250 30322
rect 35758 30270 35810 30322
rect 38782 30270 38834 30322
rect 42142 30270 42194 30322
rect 47630 30270 47682 30322
rect 48862 30270 48914 30322
rect 49870 30270 49922 30322
rect 55358 30270 55410 30322
rect 7982 30158 8034 30210
rect 11342 30158 11394 30210
rect 13582 30158 13634 30210
rect 19742 30158 19794 30210
rect 20302 30158 20354 30210
rect 21534 30158 21586 30210
rect 21870 30158 21922 30210
rect 22318 30158 22370 30210
rect 22542 30158 22594 30210
rect 22766 30158 22818 30210
rect 26574 30158 26626 30210
rect 27470 30158 27522 30210
rect 27582 30158 27634 30210
rect 28030 30158 28082 30210
rect 28702 30158 28754 30210
rect 29150 30158 29202 30210
rect 30270 30158 30322 30210
rect 31278 30158 31330 30210
rect 32062 30158 32114 30210
rect 32510 30158 32562 30210
rect 32958 30158 33010 30210
rect 33406 30158 33458 30210
rect 34078 30158 34130 30210
rect 37326 30158 37378 30210
rect 37886 30158 37938 30210
rect 38334 30158 38386 30210
rect 39230 30158 39282 30210
rect 40574 30158 40626 30210
rect 41470 30158 41522 30210
rect 42254 30158 42306 30210
rect 43262 30158 43314 30210
rect 44942 30158 44994 30210
rect 45614 30158 45666 30210
rect 45950 30158 46002 30210
rect 46846 30158 46898 30210
rect 47854 30158 47906 30210
rect 48750 30158 48802 30210
rect 49422 30158 49474 30210
rect 49646 30158 49698 30210
rect 50430 30158 50482 30210
rect 53230 30158 53282 30210
rect 53454 30158 53506 30210
rect 1710 30046 1762 30098
rect 2046 30046 2098 30098
rect 8654 30046 8706 30098
rect 14254 30046 14306 30098
rect 18398 30046 18450 30098
rect 22206 30046 22258 30098
rect 23326 30046 23378 30098
rect 27246 30046 27298 30098
rect 31390 30046 31442 30098
rect 33630 30046 33682 30098
rect 36990 30046 37042 30098
rect 39118 30046 39170 30098
rect 39566 30046 39618 30098
rect 41358 30046 41410 30098
rect 43374 30046 43426 30098
rect 45054 30046 45106 30098
rect 45390 30046 45442 30098
rect 46286 30046 46338 30098
rect 46734 30046 46786 30098
rect 48414 30046 48466 30098
rect 50766 30046 50818 30098
rect 2942 29934 2994 29986
rect 11902 29934 11954 29986
rect 12350 29934 12402 29986
rect 18286 29934 18338 29986
rect 20862 29934 20914 29986
rect 21310 29934 21362 29986
rect 21422 29934 21474 29986
rect 27694 29934 27746 29986
rect 28142 29934 28194 29986
rect 28254 29934 28306 29986
rect 37102 29934 37154 29986
rect 39342 29934 39394 29986
rect 40462 29934 40514 29986
rect 44382 29934 44434 29986
rect 45278 29934 45330 29986
rect 45838 29934 45890 29986
rect 48974 29934 49026 29986
rect 50206 29934 50258 29986
rect 50654 29934 50706 29986
rect 19838 29766 19890 29818
rect 19942 29766 19994 29818
rect 20046 29766 20098 29818
rect 50558 29766 50610 29818
rect 50662 29766 50714 29818
rect 50766 29766 50818 29818
rect 8878 29598 8930 29650
rect 16046 29598 16098 29650
rect 16270 29598 16322 29650
rect 22654 29598 22706 29650
rect 23102 29598 23154 29650
rect 25454 29598 25506 29650
rect 25566 29598 25618 29650
rect 31278 29598 31330 29650
rect 32286 29598 32338 29650
rect 33182 29598 33234 29650
rect 33630 29598 33682 29650
rect 38782 29598 38834 29650
rect 39342 29598 39394 29650
rect 40462 29598 40514 29650
rect 46510 29598 46562 29650
rect 46622 29598 46674 29650
rect 46734 29598 46786 29650
rect 47854 29598 47906 29650
rect 2046 29486 2098 29538
rect 12462 29486 12514 29538
rect 15822 29486 15874 29538
rect 16718 29486 16770 29538
rect 24558 29486 24610 29538
rect 29822 29486 29874 29538
rect 31502 29486 31554 29538
rect 34414 29486 34466 29538
rect 37550 29486 37602 29538
rect 40238 29486 40290 29538
rect 41134 29486 41186 29538
rect 47406 29486 47458 29538
rect 1710 29374 1762 29426
rect 10110 29374 10162 29426
rect 10558 29374 10610 29426
rect 11230 29374 11282 29426
rect 11454 29374 11506 29426
rect 12238 29374 12290 29426
rect 12798 29374 12850 29426
rect 13022 29374 13074 29426
rect 14030 29374 14082 29426
rect 15150 29374 15202 29426
rect 22654 29374 22706 29426
rect 23550 29374 23602 29426
rect 24446 29374 24498 29426
rect 24782 29374 24834 29426
rect 25790 29374 25842 29426
rect 25902 29374 25954 29426
rect 26686 29374 26738 29426
rect 30046 29374 30098 29426
rect 30494 29374 30546 29426
rect 31838 29374 31890 29426
rect 32174 29374 32226 29426
rect 34974 29374 35026 29426
rect 35758 29374 35810 29426
rect 36094 29374 36146 29426
rect 37214 29374 37266 29426
rect 38334 29374 38386 29426
rect 38558 29374 38610 29426
rect 39118 29374 39170 29426
rect 39454 29374 39506 29426
rect 40126 29374 40178 29426
rect 46174 29374 46226 29426
rect 47182 29374 47234 29426
rect 47630 29374 47682 29426
rect 2494 29262 2546 29314
rect 8990 29262 9042 29314
rect 13694 29262 13746 29314
rect 15486 29262 15538 29314
rect 15934 29262 15986 29314
rect 17614 29262 17666 29314
rect 23326 29262 23378 29314
rect 24110 29262 24162 29314
rect 25678 29262 25730 29314
rect 27358 29262 27410 29314
rect 29486 29262 29538 29314
rect 31390 29262 31442 29314
rect 34638 29262 34690 29314
rect 36654 29262 36706 29314
rect 38110 29262 38162 29314
rect 38670 29262 38722 29314
rect 48862 29262 48914 29314
rect 10334 29150 10386 29202
rect 13470 29150 13522 29202
rect 16606 29150 16658 29202
rect 32286 29150 32338 29202
rect 47518 29150 47570 29202
rect 4478 28982 4530 29034
rect 4582 28982 4634 29034
rect 4686 28982 4738 29034
rect 35198 28982 35250 29034
rect 35302 28982 35354 29034
rect 35406 28982 35458 29034
rect 22542 28814 22594 28866
rect 22878 28814 22930 28866
rect 28030 28814 28082 28866
rect 28366 28814 28418 28866
rect 29262 28814 29314 28866
rect 31390 28814 31442 28866
rect 33742 28814 33794 28866
rect 39790 28814 39842 28866
rect 40126 28814 40178 28866
rect 41358 28814 41410 28866
rect 42366 28814 42418 28866
rect 42702 28814 42754 28866
rect 45950 28814 46002 28866
rect 57934 28814 57986 28866
rect 17166 28702 17218 28754
rect 18286 28702 18338 28754
rect 20414 28702 20466 28754
rect 21646 28702 21698 28754
rect 24670 28702 24722 28754
rect 26798 28702 26850 28754
rect 27134 28702 27186 28754
rect 28590 28702 28642 28754
rect 31166 28702 31218 28754
rect 35646 28702 35698 28754
rect 37550 28702 37602 28754
rect 38670 28702 38722 28754
rect 40350 28702 40402 28754
rect 42926 28702 42978 28754
rect 47854 28702 47906 28754
rect 55358 28702 55410 28754
rect 1710 28590 1762 28642
rect 2494 28590 2546 28642
rect 12798 28590 12850 28642
rect 13470 28590 13522 28642
rect 14254 28590 14306 28642
rect 17502 28590 17554 28642
rect 21422 28590 21474 28642
rect 21870 28590 21922 28642
rect 21982 28590 22034 28642
rect 22654 28590 22706 28642
rect 23998 28590 24050 28642
rect 30606 28590 30658 28642
rect 31054 28590 31106 28642
rect 34526 28590 34578 28642
rect 34974 28590 35026 28642
rect 35534 28590 35586 28642
rect 35870 28590 35922 28642
rect 36094 28590 36146 28642
rect 36430 28590 36482 28642
rect 36990 28590 37042 28642
rect 39790 28590 39842 28642
rect 40798 28590 40850 28642
rect 41358 28590 41410 28642
rect 41806 28590 41858 28642
rect 43486 28590 43538 28642
rect 43598 28590 43650 28642
rect 44942 28590 44994 28642
rect 45054 28590 45106 28642
rect 45614 28590 45666 28642
rect 46286 28590 46338 28642
rect 46958 28590 47010 28642
rect 47518 28590 47570 28642
rect 55582 28590 55634 28642
rect 8430 28478 8482 28530
rect 13582 28478 13634 28530
rect 15038 28478 15090 28530
rect 22990 28478 23042 28530
rect 23214 28478 23266 28530
rect 23438 28478 23490 28530
rect 29150 28478 29202 28530
rect 29934 28478 29986 28530
rect 32398 28478 32450 28530
rect 32734 28478 32786 28530
rect 32846 28478 32898 28530
rect 33854 28478 33906 28530
rect 35198 28478 35250 28530
rect 36318 28478 36370 28530
rect 37998 28478 38050 28530
rect 39118 28478 39170 28530
rect 44270 28478 44322 28530
rect 45166 28478 45218 28530
rect 47182 28478 47234 28530
rect 2046 28366 2098 28418
rect 22542 28366 22594 28418
rect 27694 28366 27746 28418
rect 29262 28366 29314 28418
rect 30046 28366 30098 28418
rect 30158 28366 30210 28418
rect 32286 28366 32338 28418
rect 33070 28366 33122 28418
rect 33742 28366 33794 28418
rect 38110 28366 38162 28418
rect 38334 28366 38386 28418
rect 44046 28366 44098 28418
rect 44158 28366 44210 28418
rect 46062 28366 46114 28418
rect 47294 28366 47346 28418
rect 19838 28198 19890 28250
rect 19942 28198 19994 28250
rect 20046 28198 20098 28250
rect 50558 28198 50610 28250
rect 50662 28198 50714 28250
rect 50766 28198 50818 28250
rect 14366 28030 14418 28082
rect 15710 28030 15762 28082
rect 15822 28030 15874 28082
rect 15934 28030 15986 28082
rect 16718 28030 16770 28082
rect 17502 28030 17554 28082
rect 22542 28030 22594 28082
rect 23326 28030 23378 28082
rect 24670 28030 24722 28082
rect 25342 28030 25394 28082
rect 26798 28030 26850 28082
rect 27918 28030 27970 28082
rect 30270 28030 30322 28082
rect 30606 28030 30658 28082
rect 31166 28030 31218 28082
rect 32062 28030 32114 28082
rect 40910 28030 40962 28082
rect 45726 28030 45778 28082
rect 46510 28030 46562 28082
rect 2046 27918 2098 27970
rect 9998 27918 10050 27970
rect 11790 27918 11842 27970
rect 16494 27918 16546 27970
rect 16830 27918 16882 27970
rect 24110 27918 24162 27970
rect 29374 27918 29426 27970
rect 29710 27918 29762 27970
rect 29822 27918 29874 27970
rect 32286 27918 32338 27970
rect 41694 27918 41746 27970
rect 44494 27918 44546 27970
rect 49534 27918 49586 27970
rect 50318 27918 50370 27970
rect 50430 27918 50482 27970
rect 1710 27806 1762 27858
rect 11118 27806 11170 27858
rect 16382 27806 16434 27858
rect 19070 27806 19122 27858
rect 22318 27806 22370 27858
rect 22990 27806 23042 27858
rect 23550 27806 23602 27858
rect 24222 27806 24274 27858
rect 25230 27806 25282 27858
rect 25566 27806 25618 27858
rect 25902 27806 25954 27858
rect 29038 27806 29090 27858
rect 31502 27806 31554 27858
rect 31726 27806 31778 27858
rect 32510 27806 32562 27858
rect 33070 27806 33122 27858
rect 37438 27806 37490 27858
rect 41246 27806 41298 27858
rect 45278 27806 45330 27858
rect 48078 27806 48130 27858
rect 48750 27806 48802 27858
rect 49310 27806 49362 27858
rect 50094 27806 50146 27858
rect 2494 27694 2546 27746
rect 13918 27694 13970 27746
rect 18286 27694 18338 27746
rect 18846 27694 18898 27746
rect 19854 27694 19906 27746
rect 21982 27694 22034 27746
rect 22430 27694 22482 27746
rect 26238 27694 26290 27746
rect 28478 27694 28530 27746
rect 32398 27694 32450 27746
rect 33854 27694 33906 27746
rect 35982 27694 36034 27746
rect 38222 27694 38274 27746
rect 40350 27694 40402 27746
rect 41582 27694 41634 27746
rect 42366 27694 42418 27746
rect 47966 27694 48018 27746
rect 49646 27694 49698 27746
rect 9886 27582 9938 27634
rect 18510 27582 18562 27634
rect 18846 27582 18898 27634
rect 23214 27582 23266 27634
rect 24110 27582 24162 27634
rect 29822 27582 29874 27634
rect 41918 27582 41970 27634
rect 4478 27414 4530 27466
rect 4582 27414 4634 27466
rect 4686 27414 4738 27466
rect 35198 27414 35250 27466
rect 35302 27414 35354 27466
rect 35406 27414 35458 27466
rect 14030 27246 14082 27298
rect 18398 27246 18450 27298
rect 22542 27246 22594 27298
rect 35198 27246 35250 27298
rect 43038 27246 43090 27298
rect 46846 27246 46898 27298
rect 9102 27134 9154 27186
rect 11230 27134 11282 27186
rect 14366 27134 14418 27186
rect 16606 27134 16658 27186
rect 18510 27134 18562 27186
rect 20862 27134 20914 27186
rect 22654 27134 22706 27186
rect 24670 27134 24722 27186
rect 25902 27134 25954 27186
rect 26350 27134 26402 27186
rect 27134 27134 27186 27186
rect 29934 27134 29986 27186
rect 32062 27134 32114 27186
rect 32510 27134 32562 27186
rect 33966 27134 34018 27186
rect 37998 27134 38050 27186
rect 41582 27134 41634 27186
rect 43934 27134 43986 27186
rect 47406 27134 47458 27186
rect 48526 27134 48578 27186
rect 8430 27022 8482 27074
rect 13694 27022 13746 27074
rect 14142 27022 14194 27074
rect 14702 27022 14754 27074
rect 15486 27022 15538 27074
rect 15822 27022 15874 27074
rect 17614 27022 17666 27074
rect 18846 27022 18898 27074
rect 19630 27022 19682 27074
rect 21646 27022 21698 27074
rect 22430 27022 22482 27074
rect 23326 27022 23378 27074
rect 23998 27022 24050 27074
rect 24222 27022 24274 27074
rect 25118 27022 25170 27074
rect 27470 27022 27522 27074
rect 28030 27022 28082 27074
rect 29262 27022 29314 27074
rect 33294 27022 33346 27074
rect 33406 27022 33458 27074
rect 34078 27022 34130 27074
rect 34414 27022 34466 27074
rect 34526 27022 34578 27074
rect 34862 27022 34914 27074
rect 35758 27022 35810 27074
rect 37774 27022 37826 27074
rect 38334 27022 38386 27074
rect 39006 27022 39058 27074
rect 40014 27022 40066 27074
rect 40350 27022 40402 27074
rect 41806 27022 41858 27074
rect 42142 27022 42194 27074
rect 42478 27022 42530 27074
rect 42702 27022 42754 27074
rect 43262 27022 43314 27074
rect 43598 27022 43650 27074
rect 45390 27022 45442 27074
rect 45726 27022 45778 27074
rect 46062 27022 46114 27074
rect 46174 27022 46226 27074
rect 46510 27022 46562 27074
rect 47742 27022 47794 27074
rect 51326 27022 51378 27074
rect 1710 26910 1762 26962
rect 2382 26910 2434 26962
rect 2718 26910 2770 26962
rect 3166 26910 3218 26962
rect 16942 26910 16994 26962
rect 17054 26910 17106 26962
rect 17390 26910 17442 26962
rect 20078 26910 20130 26962
rect 21310 26910 21362 26962
rect 21534 26910 21586 26962
rect 24558 26910 24610 26962
rect 25454 26910 25506 26962
rect 33854 26910 33906 26962
rect 34750 26910 34802 26962
rect 35310 26910 35362 26962
rect 35534 26910 35586 26962
rect 36318 26910 36370 26962
rect 37326 26910 37378 26962
rect 37550 26910 37602 26962
rect 38446 26910 38498 26962
rect 39454 26910 39506 26962
rect 42926 26910 42978 26962
rect 43374 26910 43426 26962
rect 44830 26910 44882 26962
rect 45838 26910 45890 26962
rect 46734 26910 46786 26962
rect 48190 26910 48242 26962
rect 50654 26910 50706 26962
rect 2046 26798 2098 26850
rect 23774 26798 23826 26850
rect 23886 26798 23938 26850
rect 24782 26798 24834 26850
rect 37998 26798 38050 26850
rect 38558 26798 38610 26850
rect 42030 26798 42082 26850
rect 44942 26798 44994 26850
rect 19838 26630 19890 26682
rect 19942 26630 19994 26682
rect 20046 26630 20098 26682
rect 50558 26630 50610 26682
rect 50662 26630 50714 26682
rect 50766 26630 50818 26682
rect 2046 26462 2098 26514
rect 2494 26462 2546 26514
rect 25118 26462 25170 26514
rect 25230 26462 25282 26514
rect 26014 26462 26066 26514
rect 28926 26462 28978 26514
rect 38334 26462 38386 26514
rect 38782 26462 38834 26514
rect 46174 26462 46226 26514
rect 46846 26462 46898 26514
rect 47182 26462 47234 26514
rect 47742 26462 47794 26514
rect 48078 26462 48130 26514
rect 48190 26462 48242 26514
rect 49646 26462 49698 26514
rect 49758 26462 49810 26514
rect 50094 26462 50146 26514
rect 15598 26350 15650 26402
rect 16830 26350 16882 26402
rect 20078 26350 20130 26402
rect 23662 26350 23714 26402
rect 23998 26350 24050 26402
rect 24446 26350 24498 26402
rect 24558 26350 24610 26402
rect 25454 26350 25506 26402
rect 26350 26350 26402 26402
rect 39006 26350 39058 26402
rect 47966 26350 48018 26402
rect 1710 26238 1762 26290
rect 11118 26238 11170 26290
rect 11678 26238 11730 26290
rect 12014 26238 12066 26290
rect 15374 26238 15426 26290
rect 16494 26238 16546 26290
rect 17614 26238 17666 26290
rect 18062 26238 18114 26290
rect 18846 26238 18898 26290
rect 19070 26238 19122 26290
rect 19518 26238 19570 26290
rect 20414 26238 20466 26290
rect 20638 26238 20690 26290
rect 21646 26238 21698 26290
rect 22542 26238 22594 26290
rect 23438 26238 23490 26290
rect 24222 26238 24274 26290
rect 25790 26238 25842 26290
rect 28590 26238 28642 26290
rect 34302 26238 34354 26290
rect 34750 26238 34802 26290
rect 35198 26238 35250 26290
rect 36094 26238 36146 26290
rect 36430 26238 36482 26290
rect 37886 26238 37938 26290
rect 38558 26238 38610 26290
rect 39118 26238 39170 26290
rect 43150 26238 43202 26290
rect 43934 26238 43986 26290
rect 44382 26238 44434 26290
rect 44942 26238 44994 26290
rect 45278 26238 45330 26290
rect 48974 26238 49026 26290
rect 49870 26238 49922 26290
rect 2942 26126 2994 26178
rect 8318 26126 8370 26178
rect 12798 26126 12850 26178
rect 14926 26126 14978 26178
rect 16158 26126 16210 26178
rect 21534 26126 21586 26178
rect 23102 26126 23154 26178
rect 23886 26126 23938 26178
rect 26798 26126 26850 26178
rect 27246 26126 27298 26178
rect 27694 26126 27746 26178
rect 28142 26126 28194 26178
rect 33742 26126 33794 26178
rect 36878 26126 36930 26178
rect 37326 26126 37378 26178
rect 42926 26126 42978 26178
rect 46622 26126 46674 26178
rect 48750 26126 48802 26178
rect 8206 26014 8258 26066
rect 17950 26014 18002 26066
rect 20974 26014 21026 26066
rect 35870 26014 35922 26066
rect 36766 26014 36818 26066
rect 37438 26014 37490 26066
rect 44830 26014 44882 26066
rect 49310 26014 49362 26066
rect 4478 25846 4530 25898
rect 4582 25846 4634 25898
rect 4686 25846 4738 25898
rect 35198 25846 35250 25898
rect 35302 25846 35354 25898
rect 35406 25846 35458 25898
rect 11118 25678 11170 25730
rect 13470 25678 13522 25730
rect 20638 25678 20690 25730
rect 33518 25678 33570 25730
rect 7198 25566 7250 25618
rect 9326 25566 9378 25618
rect 11342 25566 11394 25618
rect 13582 25566 13634 25618
rect 14702 25566 14754 25618
rect 16270 25566 16322 25618
rect 18398 25566 18450 25618
rect 19070 25566 19122 25618
rect 19742 25566 19794 25618
rect 35198 25566 35250 25618
rect 37774 25566 37826 25618
rect 39902 25566 39954 25618
rect 41246 25566 41298 25618
rect 45614 25566 45666 25618
rect 47742 25566 47794 25618
rect 6526 25454 6578 25506
rect 10446 25454 10498 25506
rect 11678 25454 11730 25506
rect 12350 25454 12402 25506
rect 14254 25454 14306 25506
rect 15150 25454 15202 25506
rect 15486 25454 15538 25506
rect 19406 25454 19458 25506
rect 26574 25454 26626 25506
rect 27134 25454 27186 25506
rect 28142 25454 28194 25506
rect 31278 25454 31330 25506
rect 32174 25454 32226 25506
rect 33294 25454 33346 25506
rect 33406 25454 33458 25506
rect 33742 25454 33794 25506
rect 33966 25454 34018 25506
rect 34862 25454 34914 25506
rect 37102 25454 37154 25506
rect 40574 25454 40626 25506
rect 44158 25454 44210 25506
rect 44830 25454 44882 25506
rect 1710 25342 1762 25394
rect 2046 25342 2098 25394
rect 10222 25342 10274 25394
rect 12910 25342 12962 25394
rect 20750 25342 20802 25394
rect 21870 25342 21922 25394
rect 27470 25342 27522 25394
rect 28366 25342 28418 25394
rect 31726 25342 31778 25394
rect 40238 25342 40290 25394
rect 43374 25342 43426 25394
rect 57598 25342 57650 25394
rect 58158 25342 58210 25394
rect 2494 25230 2546 25282
rect 13918 25230 13970 25282
rect 20638 25230 20690 25282
rect 31054 25230 31106 25282
rect 35870 25230 35922 25282
rect 40350 25230 40402 25282
rect 41022 25230 41074 25282
rect 57822 25230 57874 25282
rect 19838 25062 19890 25114
rect 19942 25062 19994 25114
rect 20046 25062 20098 25114
rect 50558 25062 50610 25114
rect 50662 25062 50714 25114
rect 50766 25062 50818 25114
rect 10222 24894 10274 24946
rect 14590 24894 14642 24946
rect 14926 24894 14978 24946
rect 15486 24894 15538 24946
rect 18734 24894 18786 24946
rect 19182 24894 19234 24946
rect 19966 24894 20018 24946
rect 23774 24894 23826 24946
rect 24334 24894 24386 24946
rect 24558 24894 24610 24946
rect 34190 24894 34242 24946
rect 48078 24894 48130 24946
rect 57822 24894 57874 24946
rect 2046 24782 2098 24834
rect 11118 24782 11170 24834
rect 14254 24782 14306 24834
rect 18062 24782 18114 24834
rect 22430 24782 22482 24834
rect 23886 24782 23938 24834
rect 24670 24782 24722 24834
rect 25342 24782 25394 24834
rect 25454 24782 25506 24834
rect 25790 24782 25842 24834
rect 26798 24782 26850 24834
rect 33406 24782 33458 24834
rect 33854 24782 33906 24834
rect 33966 24782 34018 24834
rect 43598 24782 43650 24834
rect 48190 24782 48242 24834
rect 48750 24782 48802 24834
rect 50654 24782 50706 24834
rect 1710 24670 1762 24722
rect 5630 24670 5682 24722
rect 11790 24670 11842 24722
rect 12238 24670 12290 24722
rect 13022 24670 13074 24722
rect 14030 24670 14082 24722
rect 23214 24670 23266 24722
rect 23550 24670 23602 24722
rect 23998 24670 24050 24722
rect 25118 24670 25170 24722
rect 26126 24670 26178 24722
rect 26574 24670 26626 24722
rect 30270 24670 30322 24722
rect 31166 24670 31218 24722
rect 32062 24670 32114 24722
rect 36206 24670 36258 24722
rect 41470 24670 41522 24722
rect 41582 24670 41634 24722
rect 42366 24670 42418 24722
rect 43374 24670 43426 24722
rect 44046 24670 44098 24722
rect 47854 24670 47906 24722
rect 49422 24670 49474 24722
rect 49982 24670 50034 24722
rect 50542 24670 50594 24722
rect 58158 24670 58210 24722
rect 2494 24558 2546 24610
rect 6302 24558 6354 24610
rect 8430 24558 8482 24610
rect 8766 24558 8818 24610
rect 8878 24558 8930 24610
rect 9662 24558 9714 24610
rect 12574 24558 12626 24610
rect 17726 24558 17778 24610
rect 19630 24558 19682 24610
rect 20302 24558 20354 24610
rect 27246 24558 27298 24610
rect 29486 24558 29538 24610
rect 31502 24558 31554 24610
rect 32398 24558 32450 24610
rect 33294 24558 33346 24610
rect 34638 24558 34690 24610
rect 37102 24558 37154 24610
rect 42702 24558 42754 24610
rect 44718 24558 44770 24610
rect 46846 24558 46898 24610
rect 47294 24558 47346 24610
rect 48974 24558 49026 24610
rect 57598 24558 57650 24610
rect 11230 24446 11282 24498
rect 13358 24446 13410 24498
rect 18174 24446 18226 24498
rect 18510 24446 18562 24498
rect 19294 24446 19346 24498
rect 19854 24446 19906 24498
rect 43038 24446 43090 24498
rect 50430 24446 50482 24498
rect 4478 24278 4530 24330
rect 4582 24278 4634 24330
rect 4686 24278 4738 24330
rect 35198 24278 35250 24330
rect 35302 24278 35354 24330
rect 35406 24278 35458 24330
rect 8318 24110 8370 24162
rect 23550 24110 23602 24162
rect 29262 24110 29314 24162
rect 43486 24110 43538 24162
rect 9998 23998 10050 24050
rect 12126 23998 12178 24050
rect 19854 23998 19906 24050
rect 21534 23998 21586 24050
rect 23214 23998 23266 24050
rect 23662 23998 23714 24050
rect 27694 23998 27746 24050
rect 28254 23998 28306 24050
rect 28590 23998 28642 24050
rect 32734 23998 32786 24050
rect 34862 23998 34914 24050
rect 36206 23998 36258 24050
rect 38782 23998 38834 24050
rect 39118 23998 39170 24050
rect 43598 23998 43650 24050
rect 7198 23886 7250 23938
rect 7646 23886 7698 23938
rect 7758 23886 7810 23938
rect 8094 23886 8146 23938
rect 12910 23886 12962 23938
rect 17278 23886 17330 23938
rect 19294 23886 19346 23938
rect 22654 23886 22706 23938
rect 22990 23886 23042 23938
rect 24894 23886 24946 23938
rect 31950 23886 32002 23938
rect 35758 23886 35810 23938
rect 37438 23886 37490 23938
rect 37998 23886 38050 23938
rect 42030 23886 42082 23938
rect 43150 23886 43202 23938
rect 50094 23886 50146 23938
rect 50654 23886 50706 23938
rect 1710 23774 1762 23826
rect 2046 23774 2098 23826
rect 6974 23774 7026 23826
rect 8318 23774 8370 23826
rect 13694 23774 13746 23826
rect 19070 23774 19122 23826
rect 20750 23774 20802 23826
rect 24334 23774 24386 23826
rect 24446 23774 24498 23826
rect 25566 23774 25618 23826
rect 29150 23774 29202 23826
rect 29598 23774 29650 23826
rect 36990 23774 37042 23826
rect 41246 23774 41298 23826
rect 43934 23774 43986 23826
rect 44046 23774 44098 23826
rect 46958 23774 47010 23826
rect 50430 23774 50482 23826
rect 58158 23774 58210 23826
rect 2494 23662 2546 23714
rect 20302 23662 20354 23714
rect 21870 23662 21922 23714
rect 29934 23662 29986 23714
rect 35198 23662 35250 23714
rect 42590 23662 42642 23714
rect 57598 23662 57650 23714
rect 57822 23662 57874 23714
rect 19838 23494 19890 23546
rect 19942 23494 19994 23546
rect 20046 23494 20098 23546
rect 50558 23494 50610 23546
rect 50662 23494 50714 23546
rect 50766 23494 50818 23546
rect 14366 23326 14418 23378
rect 15150 23326 15202 23378
rect 22206 23326 22258 23378
rect 39230 23326 39282 23378
rect 40238 23326 40290 23378
rect 49982 23326 50034 23378
rect 50206 23326 50258 23378
rect 2046 23214 2098 23266
rect 13470 23214 13522 23266
rect 13806 23214 13858 23266
rect 18174 23214 18226 23266
rect 20974 23214 21026 23266
rect 22654 23214 22706 23266
rect 27470 23214 27522 23266
rect 27806 23214 27858 23266
rect 28366 23214 28418 23266
rect 35646 23214 35698 23266
rect 47854 23214 47906 23266
rect 47966 23214 48018 23266
rect 50318 23214 50370 23266
rect 1710 23102 1762 23154
rect 5406 23102 5458 23154
rect 9774 23102 9826 23154
rect 10334 23102 10386 23154
rect 11118 23102 11170 23154
rect 11230 23102 11282 23154
rect 11790 23102 11842 23154
rect 13022 23102 13074 23154
rect 17502 23102 17554 23154
rect 20638 23102 20690 23154
rect 23550 23102 23602 23154
rect 24558 23102 24610 23154
rect 25342 23102 25394 23154
rect 25678 23102 25730 23154
rect 26014 23102 26066 23154
rect 26350 23102 26402 23154
rect 27134 23102 27186 23154
rect 31838 23102 31890 23154
rect 34638 23102 34690 23154
rect 39790 23102 39842 23154
rect 40910 23102 40962 23154
rect 41358 23102 41410 23154
rect 42142 23102 42194 23154
rect 42590 23102 42642 23154
rect 42926 23102 42978 23154
rect 43038 23102 43090 23154
rect 44382 23102 44434 23154
rect 44606 23102 44658 23154
rect 44942 23102 44994 23154
rect 45166 23102 45218 23154
rect 45950 23102 46002 23154
rect 46398 23102 46450 23154
rect 46846 23102 46898 23154
rect 47294 23102 47346 23154
rect 47518 23102 47570 23154
rect 49422 23102 49474 23154
rect 49646 23102 49698 23154
rect 2494 22990 2546 23042
rect 6078 22990 6130 23042
rect 8206 22990 8258 23042
rect 12126 22990 12178 23042
rect 12686 22990 12738 23042
rect 14702 22990 14754 23042
rect 16718 22990 16770 23042
rect 20302 22990 20354 23042
rect 21422 22990 21474 23042
rect 23102 22990 23154 23042
rect 24110 22990 24162 23042
rect 26126 22990 26178 23042
rect 26574 22990 26626 23042
rect 28926 22990 28978 23042
rect 31054 22990 31106 23042
rect 33182 22990 33234 23042
rect 47406 22990 47458 23042
rect 48750 22990 48802 23042
rect 10110 22878 10162 22930
rect 14590 22878 14642 22930
rect 16830 22878 16882 22930
rect 22094 22878 22146 22930
rect 23102 22878 23154 22930
rect 42814 22878 42866 22930
rect 43934 22878 43986 22930
rect 47966 22878 48018 22930
rect 4478 22710 4530 22762
rect 4582 22710 4634 22762
rect 4686 22710 4738 22762
rect 35198 22710 35250 22762
rect 35302 22710 35354 22762
rect 35406 22710 35458 22762
rect 6974 22542 7026 22594
rect 7758 22542 7810 22594
rect 20526 22542 20578 22594
rect 26910 22542 26962 22594
rect 30942 22542 30994 22594
rect 7086 22430 7138 22482
rect 10782 22430 10834 22482
rect 11790 22430 11842 22482
rect 14366 22430 14418 22482
rect 14814 22430 14866 22482
rect 16942 22430 16994 22482
rect 23326 22430 23378 22482
rect 28142 22430 28194 22482
rect 31166 22430 31218 22482
rect 33518 22430 33570 22482
rect 35646 22430 35698 22482
rect 40462 22430 40514 22482
rect 41246 22430 41298 22482
rect 42142 22430 42194 22482
rect 43150 22430 43202 22482
rect 43486 22430 43538 22482
rect 45278 22430 45330 22482
rect 47854 22430 47906 22482
rect 49982 22430 50034 22482
rect 7982 22318 8034 22370
rect 8430 22318 8482 22370
rect 8766 22318 8818 22370
rect 9214 22318 9266 22370
rect 10110 22318 10162 22370
rect 10446 22318 10498 22370
rect 11230 22318 11282 22370
rect 17726 22318 17778 22370
rect 18398 22318 18450 22370
rect 18846 22318 18898 22370
rect 19518 22318 19570 22370
rect 19742 22318 19794 22370
rect 20414 22318 20466 22370
rect 25230 22318 25282 22370
rect 27694 22318 27746 22370
rect 30270 22318 30322 22370
rect 30718 22318 30770 22370
rect 31726 22318 31778 22370
rect 32286 22318 32338 22370
rect 32398 22318 32450 22370
rect 36318 22318 36370 22370
rect 37550 22318 37602 22370
rect 40798 22318 40850 22370
rect 41694 22318 41746 22370
rect 43598 22318 43650 22370
rect 44830 22318 44882 22370
rect 45502 22318 45554 22370
rect 46174 22318 46226 22370
rect 47070 22318 47122 22370
rect 1710 22206 1762 22258
rect 2382 22206 2434 22258
rect 13582 22206 13634 22258
rect 20750 22206 20802 22258
rect 27134 22206 27186 22258
rect 38334 22206 38386 22258
rect 44158 22206 44210 22258
rect 45950 22206 46002 22258
rect 57598 22206 57650 22258
rect 58158 22206 58210 22258
rect 2046 22094 2098 22146
rect 2718 22094 2770 22146
rect 3166 22094 3218 22146
rect 12238 22094 12290 22146
rect 13470 22094 13522 22146
rect 13918 22094 13970 22146
rect 27022 22094 27074 22146
rect 28590 22094 28642 22146
rect 42590 22094 42642 22146
rect 44046 22094 44098 22146
rect 45054 22094 45106 22146
rect 45278 22094 45330 22146
rect 45838 22094 45890 22146
rect 46622 22094 46674 22146
rect 57822 22094 57874 22146
rect 19838 21926 19890 21978
rect 19942 21926 19994 21978
rect 20046 21926 20098 21978
rect 50558 21926 50610 21978
rect 50662 21926 50714 21978
rect 50766 21926 50818 21978
rect 2494 21758 2546 21810
rect 18174 21758 18226 21810
rect 22878 21758 22930 21810
rect 23102 21758 23154 21810
rect 25342 21758 25394 21810
rect 31054 21758 31106 21810
rect 32510 21758 32562 21810
rect 33070 21758 33122 21810
rect 34526 21758 34578 21810
rect 40126 21758 40178 21810
rect 41022 21758 41074 21810
rect 41470 21758 41522 21810
rect 41918 21758 41970 21810
rect 46510 21758 46562 21810
rect 47518 21758 47570 21810
rect 47854 21758 47906 21810
rect 2046 21646 2098 21698
rect 8990 21646 9042 21698
rect 11006 21646 11058 21698
rect 14254 21646 14306 21698
rect 23774 21646 23826 21698
rect 24558 21646 24610 21698
rect 25454 21646 25506 21698
rect 26350 21646 26402 21698
rect 30494 21646 30546 21698
rect 30942 21646 30994 21698
rect 35534 21646 35586 21698
rect 35870 21646 35922 21698
rect 36430 21646 36482 21698
rect 37102 21646 37154 21698
rect 39790 21646 39842 21698
rect 42254 21646 42306 21698
rect 44046 21646 44098 21698
rect 47294 21646 47346 21698
rect 1710 21534 1762 21586
rect 6302 21534 6354 21586
rect 6526 21534 6578 21586
rect 7870 21534 7922 21586
rect 7982 21534 8034 21586
rect 8766 21534 8818 21586
rect 10222 21534 10274 21586
rect 13470 21534 13522 21586
rect 18510 21534 18562 21586
rect 19518 21534 19570 21586
rect 23550 21534 23602 21586
rect 24110 21534 24162 21586
rect 24334 21534 24386 21586
rect 24670 21534 24722 21586
rect 25118 21534 25170 21586
rect 26014 21534 26066 21586
rect 26238 21534 26290 21586
rect 27246 21534 27298 21586
rect 30606 21534 30658 21586
rect 33966 21534 34018 21586
rect 35198 21534 35250 21586
rect 37550 21534 37602 21586
rect 38558 21534 38610 21586
rect 39566 21534 39618 21586
rect 43374 21534 43426 21586
rect 46846 21534 46898 21586
rect 47182 21534 47234 21586
rect 2942 21422 2994 21474
rect 9662 21422 9714 21474
rect 13134 21422 13186 21474
rect 16382 21422 16434 21474
rect 16718 21422 16770 21474
rect 17614 21422 17666 21474
rect 18958 21422 19010 21474
rect 20190 21422 20242 21474
rect 22318 21422 22370 21474
rect 22990 21422 23042 21474
rect 27918 21422 27970 21474
rect 30046 21422 30098 21474
rect 31502 21422 31554 21474
rect 31950 21422 32002 21474
rect 33518 21422 33570 21474
rect 37998 21422 38050 21474
rect 40238 21422 40290 21474
rect 42702 21422 42754 21474
rect 46174 21422 46226 21474
rect 8990 21310 9042 21362
rect 9550 21310 9602 21362
rect 16830 21310 16882 21362
rect 26798 21310 26850 21362
rect 30494 21310 30546 21362
rect 38670 21310 38722 21362
rect 4478 21142 4530 21194
rect 4582 21142 4634 21194
rect 4686 21142 4738 21194
rect 35198 21142 35250 21194
rect 35302 21142 35354 21194
rect 35406 21142 35458 21194
rect 10110 20974 10162 21026
rect 16606 20974 16658 21026
rect 20302 20974 20354 21026
rect 23438 20974 23490 21026
rect 30270 20974 30322 21026
rect 40238 20974 40290 21026
rect 6862 20862 6914 20914
rect 8990 20862 9042 20914
rect 10334 20862 10386 20914
rect 11902 20862 11954 20914
rect 19966 20862 20018 20914
rect 20414 20862 20466 20914
rect 21310 20862 21362 20914
rect 23102 20862 23154 20914
rect 24334 20862 24386 20914
rect 28142 20862 28194 20914
rect 32062 20862 32114 20914
rect 38446 20862 38498 20914
rect 44046 20862 44098 20914
rect 45278 20862 45330 20914
rect 48302 20862 48354 20914
rect 6078 20750 6130 20802
rect 9550 20750 9602 20802
rect 10558 20750 10610 20802
rect 11454 20750 11506 20802
rect 12910 20750 12962 20802
rect 14254 20750 14306 20802
rect 15374 20750 15426 20802
rect 15710 20750 15762 20802
rect 16046 20750 16098 20802
rect 16158 20750 16210 20802
rect 17166 20750 17218 20802
rect 17838 20750 17890 20802
rect 21534 20750 21586 20802
rect 22430 20750 22482 20802
rect 23774 20750 23826 20802
rect 23998 20750 24050 20802
rect 27246 20750 27298 20802
rect 28254 20750 28306 20802
rect 28702 20750 28754 20802
rect 29598 20750 29650 20802
rect 30158 20750 30210 20802
rect 30830 20750 30882 20802
rect 31054 20750 31106 20802
rect 31502 20750 31554 20802
rect 36206 20750 36258 20802
rect 37550 20750 37602 20802
rect 37998 20750 38050 20802
rect 39006 20750 39058 20802
rect 39566 20750 39618 20802
rect 40014 20750 40066 20802
rect 41582 20750 41634 20802
rect 42926 20750 42978 20802
rect 47854 20750 47906 20802
rect 1710 20638 1762 20690
rect 9326 20638 9378 20690
rect 14030 20638 14082 20690
rect 26462 20638 26514 20690
rect 34302 20638 34354 20690
rect 34974 20638 35026 20690
rect 41470 20638 41522 20690
rect 41694 20638 41746 20690
rect 42366 20638 42418 20690
rect 42590 20638 42642 20690
rect 47742 20638 47794 20690
rect 2046 20526 2098 20578
rect 2494 20526 2546 20578
rect 12350 20526 12402 20578
rect 13694 20526 13746 20578
rect 27806 20526 27858 20578
rect 28030 20526 28082 20578
rect 34750 20526 34802 20578
rect 34862 20526 34914 20578
rect 35534 20526 35586 20578
rect 35646 20526 35698 20578
rect 35758 20526 35810 20578
rect 37102 20526 37154 20578
rect 40686 20526 40738 20578
rect 42814 20526 42866 20578
rect 43598 20526 43650 20578
rect 45838 20526 45890 20578
rect 46286 20526 46338 20578
rect 46846 20526 46898 20578
rect 47294 20526 47346 20578
rect 47518 20526 47570 20578
rect 19838 20358 19890 20410
rect 19942 20358 19994 20410
rect 20046 20358 20098 20410
rect 50558 20358 50610 20410
rect 50662 20358 50714 20410
rect 50766 20358 50818 20410
rect 15150 20190 15202 20242
rect 17950 20190 18002 20242
rect 18510 20190 18562 20242
rect 38670 20190 38722 20242
rect 41246 20190 41298 20242
rect 42478 20190 42530 20242
rect 47406 20190 47458 20242
rect 2046 20078 2098 20130
rect 16046 20078 16098 20130
rect 22542 20078 22594 20130
rect 25342 20078 25394 20130
rect 31390 20078 31442 20130
rect 33070 20078 33122 20130
rect 33406 20078 33458 20130
rect 33966 20078 34018 20130
rect 34190 20078 34242 20130
rect 36094 20078 36146 20130
rect 39454 20078 39506 20130
rect 39678 20078 39730 20130
rect 40014 20078 40066 20130
rect 42926 20078 42978 20130
rect 45614 20078 45666 20130
rect 46846 20078 46898 20130
rect 47742 20078 47794 20130
rect 1710 19966 1762 20018
rect 6078 19966 6130 20018
rect 14814 19966 14866 20018
rect 18734 19966 18786 20018
rect 19182 19966 19234 20018
rect 19966 19966 20018 20018
rect 20862 19966 20914 20018
rect 21870 19966 21922 20018
rect 25678 19966 25730 20018
rect 31166 19966 31218 20018
rect 31502 19966 31554 20018
rect 34414 19966 34466 20018
rect 34862 19966 34914 20018
rect 35422 19966 35474 20018
rect 41694 19966 41746 20018
rect 41806 19966 41858 20018
rect 42030 19966 42082 20018
rect 43374 19966 43426 20018
rect 44494 19966 44546 20018
rect 45166 19966 45218 20018
rect 47630 19966 47682 20018
rect 47854 19966 47906 20018
rect 2494 19854 2546 19906
rect 6862 19854 6914 19906
rect 8990 19854 9042 19906
rect 10222 19854 10274 19906
rect 15710 19854 15762 19906
rect 16606 19854 16658 19906
rect 17502 19854 17554 19906
rect 19630 19854 19682 19906
rect 21310 19854 21362 19906
rect 24670 19854 24722 19906
rect 27694 19854 27746 19906
rect 31950 19854 32002 19906
rect 34302 19854 34354 19906
rect 38222 19854 38274 19906
rect 43822 19854 43874 19906
rect 46062 19854 46114 19906
rect 48862 19854 48914 19906
rect 17390 19742 17442 19794
rect 19294 19742 19346 19794
rect 44046 19742 44098 19794
rect 45838 19742 45890 19794
rect 46398 19742 46450 19794
rect 46622 19742 46674 19794
rect 46958 19742 47010 19794
rect 4478 19574 4530 19626
rect 4582 19574 4634 19626
rect 4686 19574 4738 19626
rect 35198 19574 35250 19626
rect 35302 19574 35354 19626
rect 35406 19574 35458 19626
rect 6862 19406 6914 19458
rect 9774 19406 9826 19458
rect 12798 19406 12850 19458
rect 14702 19406 14754 19458
rect 16830 19406 16882 19458
rect 22318 19406 22370 19458
rect 27246 19406 27298 19458
rect 35310 19406 35362 19458
rect 37102 19406 37154 19458
rect 37438 19406 37490 19458
rect 37886 19406 37938 19458
rect 38222 19406 38274 19458
rect 6750 19294 6802 19346
rect 14590 19294 14642 19346
rect 19854 19294 19906 19346
rect 20414 19294 20466 19346
rect 21310 19294 21362 19346
rect 24782 19294 24834 19346
rect 34974 19294 35026 19346
rect 37662 19294 37714 19346
rect 38110 19294 38162 19346
rect 42254 19294 42306 19346
rect 42702 19294 42754 19346
rect 47966 19294 48018 19346
rect 50094 19294 50146 19346
rect 7198 19182 7250 19234
rect 7422 19182 7474 19234
rect 8766 19182 8818 19234
rect 8878 19182 8930 19234
rect 9662 19182 9714 19234
rect 10446 19182 10498 19234
rect 11006 19182 11058 19234
rect 11454 19182 11506 19234
rect 11902 19182 11954 19234
rect 12350 19182 12402 19234
rect 13918 19182 13970 19234
rect 14366 19182 14418 19234
rect 14926 19182 14978 19234
rect 15822 19182 15874 19234
rect 16942 19182 16994 19234
rect 17726 19182 17778 19234
rect 17838 19182 17890 19234
rect 18622 19182 18674 19234
rect 19070 19182 19122 19234
rect 21758 19182 21810 19234
rect 22766 19182 22818 19234
rect 23326 19182 23378 19234
rect 25118 19182 25170 19234
rect 25566 19182 25618 19234
rect 26014 19182 26066 19234
rect 27470 19182 27522 19234
rect 27694 19182 27746 19234
rect 28142 19182 28194 19234
rect 28254 19182 28306 19234
rect 29262 19182 29314 19234
rect 30270 19182 30322 19234
rect 30942 19182 30994 19234
rect 31166 19182 31218 19234
rect 31502 19182 31554 19234
rect 32174 19182 32226 19234
rect 35758 19182 35810 19234
rect 36094 19182 36146 19234
rect 37214 19182 37266 19234
rect 39342 19182 39394 19234
rect 42590 19182 42642 19234
rect 43710 19182 43762 19234
rect 45502 19182 45554 19234
rect 46398 19182 46450 19234
rect 47182 19182 47234 19234
rect 9886 19070 9938 19122
rect 12910 19070 12962 19122
rect 16382 19070 16434 19122
rect 16718 19070 16770 19122
rect 20750 19070 20802 19122
rect 22430 19070 22482 19122
rect 23550 19070 23602 19122
rect 24110 19070 24162 19122
rect 25454 19070 25506 19122
rect 26910 19070 26962 19122
rect 29710 19070 29762 19122
rect 29934 19070 29986 19122
rect 32846 19070 32898 19122
rect 35870 19070 35922 19122
rect 37102 19070 37154 19122
rect 38558 19070 38610 19122
rect 40126 19070 40178 19122
rect 42926 19070 42978 19122
rect 43150 19070 43202 19122
rect 44942 19070 44994 19122
rect 45054 19070 45106 19122
rect 46174 19070 46226 19122
rect 46286 19070 46338 19122
rect 22318 18958 22370 19010
rect 22878 18958 22930 19010
rect 22990 18958 23042 19010
rect 23662 18958 23714 19010
rect 23886 18958 23938 19010
rect 25678 18958 25730 19010
rect 26126 18958 26178 19010
rect 26238 18958 26290 19010
rect 26462 18958 26514 19010
rect 28030 18958 28082 19010
rect 29598 18958 29650 19010
rect 30382 18958 30434 19010
rect 30494 18958 30546 19010
rect 31390 18958 31442 19010
rect 39006 18958 39058 19010
rect 43486 18958 43538 19010
rect 43598 18958 43650 19010
rect 43934 18958 43986 19010
rect 44718 18958 44770 19010
rect 46846 18958 46898 19010
rect 19838 18790 19890 18842
rect 19942 18790 19994 18842
rect 20046 18790 20098 18842
rect 50558 18790 50610 18842
rect 50662 18790 50714 18842
rect 50766 18790 50818 18842
rect 11790 18622 11842 18674
rect 22430 18622 22482 18674
rect 24558 18622 24610 18674
rect 33630 18622 33682 18674
rect 40126 18622 40178 18674
rect 40350 18622 40402 18674
rect 47854 18622 47906 18674
rect 2046 18510 2098 18562
rect 24670 18510 24722 18562
rect 34078 18510 34130 18562
rect 36318 18510 36370 18562
rect 37326 18510 37378 18562
rect 39454 18510 39506 18562
rect 39902 18510 39954 18562
rect 40910 18510 40962 18562
rect 45950 18510 46002 18562
rect 46846 18510 46898 18562
rect 1710 18398 1762 18450
rect 6526 18398 6578 18450
rect 6974 18398 7026 18450
rect 7870 18398 7922 18450
rect 7982 18398 8034 18450
rect 8766 18398 8818 18450
rect 10110 18398 10162 18450
rect 12238 18398 12290 18450
rect 16046 18398 16098 18450
rect 16270 18398 16322 18450
rect 16494 18398 16546 18450
rect 16718 18398 16770 18450
rect 17726 18398 17778 18450
rect 18958 18398 19010 18450
rect 19182 18398 19234 18450
rect 20190 18398 20242 18450
rect 20638 18398 20690 18450
rect 20974 18398 21026 18450
rect 21086 18398 21138 18450
rect 22206 18398 22258 18450
rect 22542 18398 22594 18450
rect 22766 18398 22818 18450
rect 23662 18398 23714 18450
rect 23998 18398 24050 18450
rect 24334 18398 24386 18450
rect 25790 18398 25842 18450
rect 29038 18398 29090 18450
rect 29710 18398 29762 18450
rect 32286 18398 32338 18450
rect 33742 18398 33794 18450
rect 33854 18398 33906 18450
rect 34526 18398 34578 18450
rect 34862 18398 34914 18450
rect 35310 18398 35362 18450
rect 35534 18398 35586 18450
rect 35758 18398 35810 18450
rect 35870 18398 35922 18450
rect 36542 18398 36594 18450
rect 36766 18398 36818 18450
rect 37102 18398 37154 18450
rect 37774 18398 37826 18450
rect 38670 18398 38722 18450
rect 39118 18398 39170 18450
rect 40238 18398 40290 18450
rect 41134 18398 41186 18450
rect 41470 18398 41522 18450
rect 42142 18398 42194 18450
rect 42926 18398 42978 18450
rect 45726 18398 45778 18450
rect 46286 18398 46338 18450
rect 46622 18398 46674 18450
rect 47406 18398 47458 18450
rect 47742 18398 47794 18450
rect 48078 18398 48130 18450
rect 51662 18398 51714 18450
rect 2494 18286 2546 18338
rect 8878 18286 8930 18338
rect 9550 18286 9602 18338
rect 10558 18286 10610 18338
rect 11342 18286 11394 18338
rect 12910 18286 12962 18338
rect 15038 18286 15090 18338
rect 15374 18286 15426 18338
rect 18062 18286 18114 18338
rect 18622 18286 18674 18338
rect 24110 18286 24162 18338
rect 25342 18286 25394 18338
rect 28590 18286 28642 18338
rect 31838 18286 31890 18338
rect 33406 18286 33458 18338
rect 35086 18286 35138 18338
rect 36318 18286 36370 18338
rect 37214 18286 37266 18338
rect 38334 18286 38386 18338
rect 41022 18286 41074 18338
rect 45054 18286 45106 18338
rect 46734 18286 46786 18338
rect 48750 18286 48802 18338
rect 50878 18286 50930 18338
rect 8206 18174 8258 18226
rect 10446 18174 10498 18226
rect 15598 18174 15650 18226
rect 16718 18174 16770 18226
rect 18510 18174 18562 18226
rect 19630 18174 19682 18226
rect 4478 18006 4530 18058
rect 4582 18006 4634 18058
rect 4686 18006 4738 18058
rect 35198 18006 35250 18058
rect 35302 18006 35354 18058
rect 35406 18006 35458 18058
rect 14030 17838 14082 17890
rect 17054 17838 17106 17890
rect 28254 17838 28306 17890
rect 28590 17838 28642 17890
rect 34078 17838 34130 17890
rect 40910 17838 40962 17890
rect 41246 17838 41298 17890
rect 48974 17838 49026 17890
rect 7870 17726 7922 17778
rect 9998 17726 10050 17778
rect 11118 17726 11170 17778
rect 12126 17726 12178 17778
rect 16158 17726 16210 17778
rect 17390 17726 17442 17778
rect 19630 17726 19682 17778
rect 20078 17726 20130 17778
rect 22094 17726 22146 17778
rect 24222 17726 24274 17778
rect 25342 17726 25394 17778
rect 28254 17726 28306 17778
rect 30046 17726 30098 17778
rect 30830 17726 30882 17778
rect 31614 17726 31666 17778
rect 32398 17726 32450 17778
rect 33630 17726 33682 17778
rect 34862 17726 34914 17778
rect 35982 17726 36034 17778
rect 37774 17726 37826 17778
rect 39902 17726 39954 17778
rect 40686 17726 40738 17778
rect 43038 17726 43090 17778
rect 43598 17726 43650 17778
rect 43934 17726 43986 17778
rect 46398 17726 46450 17778
rect 49758 17726 49810 17778
rect 50206 17726 50258 17778
rect 7086 17614 7138 17666
rect 12350 17614 12402 17666
rect 12910 17614 12962 17666
rect 13694 17614 13746 17666
rect 14254 17614 14306 17666
rect 14814 17614 14866 17666
rect 15150 17614 15202 17666
rect 15598 17614 15650 17666
rect 16494 17614 16546 17666
rect 16942 17614 16994 17666
rect 18062 17614 18114 17666
rect 18510 17614 18562 17666
rect 18958 17614 19010 17666
rect 21422 17614 21474 17666
rect 24782 17614 24834 17666
rect 30270 17614 30322 17666
rect 31054 17614 31106 17666
rect 33182 17614 33234 17666
rect 33966 17614 34018 17666
rect 34974 17614 35026 17666
rect 35310 17614 35362 17666
rect 35870 17614 35922 17666
rect 36206 17614 36258 17666
rect 37102 17614 37154 17666
rect 41470 17614 41522 17666
rect 41806 17614 41858 17666
rect 44718 17614 44770 17666
rect 47294 17614 47346 17666
rect 48190 17614 48242 17666
rect 48414 17614 48466 17666
rect 48750 17614 48802 17666
rect 1710 17502 1762 17554
rect 2382 17502 2434 17554
rect 2718 17502 2770 17554
rect 19518 17502 19570 17554
rect 31614 17502 31666 17554
rect 32846 17502 32898 17554
rect 34078 17502 34130 17554
rect 34750 17502 34802 17554
rect 36430 17502 36482 17554
rect 45726 17502 45778 17554
rect 45838 17502 45890 17554
rect 47406 17502 47458 17554
rect 2046 17390 2098 17442
rect 3166 17390 3218 17442
rect 11006 17390 11058 17442
rect 24558 17390 24610 17442
rect 31390 17390 31442 17442
rect 31950 17390 32002 17442
rect 40350 17390 40402 17442
rect 41694 17390 41746 17442
rect 42590 17390 42642 17442
rect 45054 17390 45106 17442
rect 45278 17390 45330 17442
rect 45390 17390 45442 17442
rect 45502 17390 45554 17442
rect 46734 17390 46786 17442
rect 47630 17390 47682 17442
rect 47966 17390 48018 17442
rect 48302 17390 48354 17442
rect 49310 17390 49362 17442
rect 19838 17222 19890 17274
rect 19942 17222 19994 17274
rect 20046 17222 20098 17274
rect 50558 17222 50610 17274
rect 50662 17222 50714 17274
rect 50766 17222 50818 17274
rect 2494 17054 2546 17106
rect 13358 17054 13410 17106
rect 23214 17054 23266 17106
rect 24334 17054 24386 17106
rect 25342 17054 25394 17106
rect 26910 17054 26962 17106
rect 28142 17054 28194 17106
rect 28590 17054 28642 17106
rect 28926 17054 28978 17106
rect 30270 17054 30322 17106
rect 30830 17054 30882 17106
rect 31502 17054 31554 17106
rect 32062 17054 32114 17106
rect 33182 17054 33234 17106
rect 33966 17054 34018 17106
rect 34190 17054 34242 17106
rect 35198 17054 35250 17106
rect 35758 17054 35810 17106
rect 36542 17054 36594 17106
rect 38894 17054 38946 17106
rect 39678 17054 39730 17106
rect 40126 17054 40178 17106
rect 41358 17054 41410 17106
rect 42814 17054 42866 17106
rect 46398 17054 46450 17106
rect 46958 17054 47010 17106
rect 47406 17054 47458 17106
rect 48862 17054 48914 17106
rect 49086 17054 49138 17106
rect 49310 17054 49362 17106
rect 49758 17054 49810 17106
rect 2046 16942 2098 16994
rect 10558 16942 10610 16994
rect 13470 16942 13522 16994
rect 14702 16942 14754 16994
rect 23550 16942 23602 16994
rect 24446 16942 24498 16994
rect 25454 16942 25506 16994
rect 36430 16942 36482 16994
rect 36990 16942 37042 16994
rect 39118 16942 39170 16994
rect 39230 16942 39282 16994
rect 43374 16942 43426 16994
rect 43710 16942 43762 16994
rect 43934 16942 43986 16994
rect 44270 16942 44322 16994
rect 45838 16942 45890 16994
rect 46286 16942 46338 16994
rect 49198 16942 49250 16994
rect 1822 16830 1874 16882
rect 9886 16830 9938 16882
rect 14030 16830 14082 16882
rect 21870 16830 21922 16882
rect 23886 16830 23938 16882
rect 26798 16830 26850 16882
rect 27022 16830 27074 16882
rect 27470 16830 27522 16882
rect 27694 16830 27746 16882
rect 27918 16830 27970 16882
rect 31950 16830 32002 16882
rect 34750 16830 34802 16882
rect 34974 16830 35026 16882
rect 35310 16830 35362 16882
rect 37662 16830 37714 16882
rect 38670 16830 38722 16882
rect 40798 16830 40850 16882
rect 41134 16830 41186 16882
rect 41806 16830 41858 16882
rect 42030 16830 42082 16882
rect 42366 16830 42418 16882
rect 44942 16830 44994 16882
rect 46622 16830 46674 16882
rect 8878 16718 8930 16770
rect 12686 16718 12738 16770
rect 16830 16718 16882 16770
rect 17614 16718 17666 16770
rect 26462 16718 26514 16770
rect 27806 16718 27858 16770
rect 30606 16718 30658 16770
rect 37886 16718 37938 16770
rect 38334 16718 38386 16770
rect 41918 16718 41970 16770
rect 43486 16718 43538 16770
rect 45166 16718 45218 16770
rect 47854 16718 47906 16770
rect 8990 16606 9042 16658
rect 23886 16606 23938 16658
rect 24334 16606 24386 16658
rect 25342 16606 25394 16658
rect 25902 16606 25954 16658
rect 26238 16606 26290 16658
rect 30942 16606 30994 16658
rect 32062 16606 32114 16658
rect 36542 16606 36594 16658
rect 38670 16606 38722 16658
rect 41022 16606 41074 16658
rect 45614 16606 45666 16658
rect 45950 16606 46002 16658
rect 4478 16438 4530 16490
rect 4582 16438 4634 16490
rect 4686 16438 4738 16490
rect 35198 16438 35250 16490
rect 35302 16438 35354 16490
rect 35406 16438 35458 16490
rect 38334 16270 38386 16322
rect 38670 16270 38722 16322
rect 49086 16270 49138 16322
rect 1822 16158 1874 16210
rect 9102 16158 9154 16210
rect 11230 16158 11282 16210
rect 12686 16158 12738 16210
rect 17278 16158 17330 16210
rect 18622 16158 18674 16210
rect 20750 16158 20802 16210
rect 22878 16158 22930 16210
rect 25342 16158 25394 16210
rect 28590 16158 28642 16210
rect 30046 16158 30098 16210
rect 30606 16158 30658 16210
rect 37102 16158 37154 16210
rect 46286 16158 46338 16210
rect 47294 16158 47346 16210
rect 49982 16158 50034 16210
rect 8430 16046 8482 16098
rect 14478 16046 14530 16098
rect 17838 16046 17890 16098
rect 23662 16046 23714 16098
rect 23886 16046 23938 16098
rect 24558 16046 24610 16098
rect 25790 16046 25842 16098
rect 35646 16046 35698 16098
rect 37998 16046 38050 16098
rect 42814 16046 42866 16098
rect 44830 16046 44882 16098
rect 45054 16046 45106 16098
rect 45502 16046 45554 16098
rect 45838 16046 45890 16098
rect 46622 16046 46674 16098
rect 47630 16046 47682 16098
rect 47854 16046 47906 16098
rect 48414 16046 48466 16098
rect 49534 16046 49586 16098
rect 50430 16046 50482 16098
rect 15150 15934 15202 15986
rect 23774 15934 23826 15986
rect 26462 15934 26514 15986
rect 29374 15934 29426 15986
rect 37886 15934 37938 15986
rect 39230 15934 39282 15986
rect 46734 15934 46786 15986
rect 49422 15934 49474 15986
rect 12798 15822 12850 15874
rect 29038 15822 29090 15874
rect 29262 15822 29314 15874
rect 36206 15822 36258 15874
rect 37662 15822 37714 15874
rect 38446 15822 38498 15874
rect 44942 15822 44994 15874
rect 46958 15822 47010 15874
rect 48190 15822 48242 15874
rect 48750 15822 48802 15874
rect 48974 15822 49026 15874
rect 49198 15822 49250 15874
rect 19838 15654 19890 15706
rect 19942 15654 19994 15706
rect 20046 15654 20098 15706
rect 50558 15654 50610 15706
rect 50662 15654 50714 15706
rect 50766 15654 50818 15706
rect 16382 15486 16434 15538
rect 16718 15486 16770 15538
rect 22990 15486 23042 15538
rect 25342 15486 25394 15538
rect 26238 15486 26290 15538
rect 26350 15486 26402 15538
rect 26462 15486 26514 15538
rect 28030 15486 28082 15538
rect 29598 15486 29650 15538
rect 32286 15486 32338 15538
rect 33294 15486 33346 15538
rect 35198 15486 35250 15538
rect 35870 15486 35922 15538
rect 35982 15486 36034 15538
rect 36878 15486 36930 15538
rect 39118 15486 39170 15538
rect 40350 15486 40402 15538
rect 42702 15486 42754 15538
rect 48750 15486 48802 15538
rect 48862 15486 48914 15538
rect 49758 15486 49810 15538
rect 50430 15486 50482 15538
rect 13694 15374 13746 15426
rect 16830 15374 16882 15426
rect 22318 15374 22370 15426
rect 22654 15374 22706 15426
rect 22766 15374 22818 15426
rect 26798 15374 26850 15426
rect 28142 15374 28194 15426
rect 29822 15374 29874 15426
rect 29934 15374 29986 15426
rect 32174 15374 32226 15426
rect 33518 15374 33570 15426
rect 39006 15374 39058 15426
rect 42030 15374 42082 15426
rect 48078 15374 48130 15426
rect 14478 15262 14530 15314
rect 17726 15262 17778 15314
rect 21870 15262 21922 15314
rect 23774 15262 23826 15314
rect 24110 15262 24162 15314
rect 24334 15262 24386 15314
rect 24670 15262 24722 15314
rect 25230 15262 25282 15314
rect 25566 15262 25618 15314
rect 25790 15262 25842 15314
rect 27246 15262 27298 15314
rect 27694 15262 27746 15314
rect 28366 15262 28418 15314
rect 28702 15262 28754 15314
rect 29150 15262 29202 15314
rect 30158 15262 30210 15314
rect 30494 15262 30546 15314
rect 30942 15262 30994 15314
rect 31838 15262 31890 15314
rect 32510 15262 32562 15314
rect 33070 15262 33122 15314
rect 33966 15262 34018 15314
rect 34190 15262 34242 15314
rect 34638 15262 34690 15314
rect 34750 15262 34802 15314
rect 35310 15262 35362 15314
rect 35422 15262 35474 15314
rect 35758 15262 35810 15314
rect 36430 15262 36482 15314
rect 37662 15262 37714 15314
rect 38334 15262 38386 15314
rect 39790 15262 39842 15314
rect 40014 15262 40066 15314
rect 41022 15262 41074 15314
rect 41582 15262 41634 15314
rect 43038 15262 43090 15314
rect 43822 15262 43874 15314
rect 46622 15262 46674 15314
rect 47294 15262 47346 15314
rect 48974 15262 49026 15314
rect 49310 15262 49362 15314
rect 50990 15262 51042 15314
rect 11566 15150 11618 15202
rect 18398 15150 18450 15202
rect 20526 15150 20578 15202
rect 23550 15150 23602 15202
rect 24222 15150 24274 15202
rect 33182 15150 33234 15202
rect 34078 15150 34130 15202
rect 37886 15150 37938 15202
rect 41918 15150 41970 15202
rect 45950 15150 46002 15202
rect 46510 15150 46562 15202
rect 52782 15150 52834 15202
rect 21870 15038 21922 15090
rect 22318 15038 22370 15090
rect 23214 15038 23266 15090
rect 31278 15038 31330 15090
rect 38110 15038 38162 15090
rect 39118 15038 39170 15090
rect 46734 15038 46786 15090
rect 4478 14870 4530 14922
rect 4582 14870 4634 14922
rect 4686 14870 4738 14922
rect 35198 14870 35250 14922
rect 35302 14870 35354 14922
rect 35406 14870 35458 14922
rect 10110 14702 10162 14754
rect 18734 14702 18786 14754
rect 27918 14702 27970 14754
rect 28478 14702 28530 14754
rect 29374 14702 29426 14754
rect 36318 14702 36370 14754
rect 36878 14702 36930 14754
rect 10446 14590 10498 14642
rect 12126 14590 12178 14642
rect 21870 14590 21922 14642
rect 23102 14590 23154 14642
rect 23886 14590 23938 14642
rect 25454 14590 25506 14642
rect 27134 14590 27186 14642
rect 27806 14590 27858 14642
rect 28142 14590 28194 14642
rect 28590 14590 28642 14642
rect 30718 14590 30770 14642
rect 31838 14590 31890 14642
rect 33406 14590 33458 14642
rect 35534 14590 35586 14642
rect 40910 14590 40962 14642
rect 43038 14590 43090 14642
rect 44046 14590 44098 14642
rect 45502 14590 45554 14642
rect 47518 14590 47570 14642
rect 50766 14590 50818 14642
rect 9550 14478 9602 14530
rect 9774 14478 9826 14530
rect 11118 14478 11170 14530
rect 11902 14478 11954 14530
rect 17950 14478 18002 14530
rect 18174 14478 18226 14530
rect 19294 14478 19346 14530
rect 19630 14478 19682 14530
rect 19966 14478 20018 14530
rect 20414 14478 20466 14530
rect 24110 14478 24162 14530
rect 24334 14478 24386 14530
rect 24782 14478 24834 14530
rect 25230 14478 25282 14530
rect 26126 14478 26178 14530
rect 26462 14478 26514 14530
rect 29710 14478 29762 14530
rect 29934 14478 29986 14530
rect 30270 14478 30322 14530
rect 30606 14478 30658 14530
rect 31166 14478 31218 14530
rect 32174 14478 32226 14530
rect 32622 14478 32674 14530
rect 36206 14478 36258 14530
rect 38110 14478 38162 14530
rect 38334 14478 38386 14530
rect 38670 14478 38722 14530
rect 39790 14478 39842 14530
rect 40238 14478 40290 14530
rect 44830 14478 44882 14530
rect 45166 14478 45218 14530
rect 46286 14478 46338 14530
rect 46622 14478 46674 14530
rect 47070 14478 47122 14530
rect 47966 14478 48018 14530
rect 21422 14366 21474 14418
rect 25118 14366 25170 14418
rect 26574 14366 26626 14418
rect 30830 14366 30882 14418
rect 31278 14366 31330 14418
rect 36990 14366 37042 14418
rect 37438 14366 37490 14418
rect 37886 14366 37938 14418
rect 38782 14366 38834 14418
rect 45950 14366 46002 14418
rect 46062 14366 46114 14418
rect 48638 14366 48690 14418
rect 21310 14254 21362 14306
rect 22318 14254 22370 14306
rect 22654 14254 22706 14306
rect 24222 14254 24274 14306
rect 36318 14254 36370 14306
rect 37214 14254 37266 14306
rect 38222 14254 38274 14306
rect 39678 14254 39730 14306
rect 43486 14254 43538 14306
rect 44942 14254 44994 14306
rect 19838 14086 19890 14138
rect 19942 14086 19994 14138
rect 20046 14086 20098 14138
rect 50558 14086 50610 14138
rect 50662 14086 50714 14138
rect 50766 14086 50818 14138
rect 27582 13918 27634 13970
rect 28254 13918 28306 13970
rect 35086 13918 35138 13970
rect 36318 13918 36370 13970
rect 38782 13918 38834 13970
rect 39230 13918 39282 13970
rect 40126 13918 40178 13970
rect 40238 13918 40290 13970
rect 40350 13918 40402 13970
rect 42142 13918 42194 13970
rect 42366 13918 42418 13970
rect 43038 13918 43090 13970
rect 43486 13918 43538 13970
rect 44494 13918 44546 13970
rect 47854 13918 47906 13970
rect 48750 13918 48802 13970
rect 49198 13918 49250 13970
rect 49870 13918 49922 13970
rect 19294 13806 19346 13858
rect 22542 13806 22594 13858
rect 25230 13806 25282 13858
rect 26910 13806 26962 13858
rect 27246 13806 27298 13858
rect 27918 13806 27970 13858
rect 28590 13806 28642 13858
rect 31166 13806 31218 13858
rect 33406 13806 33458 13858
rect 35198 13806 35250 13858
rect 36766 13806 36818 13858
rect 37438 13806 37490 13858
rect 41918 13806 41970 13858
rect 42478 13806 42530 13858
rect 46734 13806 46786 13858
rect 47630 13806 47682 13858
rect 18510 13694 18562 13746
rect 21870 13694 21922 13746
rect 25902 13694 25954 13746
rect 31950 13694 32002 13746
rect 34302 13694 34354 13746
rect 34526 13694 34578 13746
rect 34862 13694 34914 13746
rect 37326 13694 37378 13746
rect 37886 13694 37938 13746
rect 38446 13694 38498 13746
rect 39006 13694 39058 13746
rect 39678 13694 39730 13746
rect 41470 13694 41522 13746
rect 45614 13694 45666 13746
rect 46174 13694 46226 13746
rect 47070 13694 47122 13746
rect 47406 13694 47458 13746
rect 48974 13694 49026 13746
rect 21422 13582 21474 13634
rect 24670 13582 24722 13634
rect 26014 13582 26066 13634
rect 29038 13582 29090 13634
rect 32398 13582 32450 13634
rect 33630 13582 33682 13634
rect 35870 13582 35922 13634
rect 38894 13582 38946 13634
rect 41134 13582 41186 13634
rect 43934 13582 43986 13634
rect 46734 13582 46786 13634
rect 47518 13582 47570 13634
rect 48862 13582 48914 13634
rect 32286 13470 32338 13522
rect 37438 13470 37490 13522
rect 38110 13470 38162 13522
rect 4478 13302 4530 13354
rect 4582 13302 4634 13354
rect 4686 13302 4738 13354
rect 35198 13302 35250 13354
rect 35302 13302 35354 13354
rect 35406 13302 35458 13354
rect 24446 13134 24498 13186
rect 30830 13134 30882 13186
rect 33406 13134 33458 13186
rect 33742 13134 33794 13186
rect 40350 13134 40402 13186
rect 46846 13134 46898 13186
rect 20750 13022 20802 13074
rect 27582 13022 27634 13074
rect 28254 13022 28306 13074
rect 29374 13022 29426 13074
rect 30270 13022 30322 13074
rect 31054 13022 31106 13074
rect 32398 13022 32450 13074
rect 33182 13022 33234 13074
rect 35310 13022 35362 13074
rect 35870 13022 35922 13074
rect 37886 13022 37938 13074
rect 40014 13022 40066 13074
rect 44270 13022 44322 13074
rect 45502 13022 45554 13074
rect 48526 13022 48578 13074
rect 49422 13022 49474 13074
rect 22990 12910 23042 12962
rect 23662 12910 23714 12962
rect 24110 12910 24162 12962
rect 24670 12910 24722 12962
rect 25006 12910 25058 12962
rect 25342 12910 25394 12962
rect 25454 12910 25506 12962
rect 26238 12910 26290 12962
rect 26574 12910 26626 12962
rect 31502 12910 31554 12962
rect 31950 12910 32002 12962
rect 36430 12910 36482 12962
rect 37102 12910 37154 12962
rect 40798 12910 40850 12962
rect 41134 12910 41186 12962
rect 41470 12910 41522 12962
rect 45838 12910 45890 12962
rect 46286 12910 46338 12962
rect 46622 12910 46674 12962
rect 47518 12910 47570 12962
rect 48190 12910 48242 12962
rect 48414 12910 48466 12962
rect 49086 12910 49138 12962
rect 32510 12798 32562 12850
rect 34190 12798 34242 12850
rect 34750 12798 34802 12850
rect 40462 12798 40514 12850
rect 42142 12798 42194 12850
rect 47182 12798 47234 12850
rect 47742 12798 47794 12850
rect 26462 12686 26514 12738
rect 27022 12686 27074 12738
rect 32286 12686 32338 12738
rect 34638 12686 34690 12738
rect 40910 12686 40962 12738
rect 47630 12686 47682 12738
rect 48638 12686 48690 12738
rect 19838 12518 19890 12570
rect 19942 12518 19994 12570
rect 20046 12518 20098 12570
rect 50558 12518 50610 12570
rect 50662 12518 50714 12570
rect 50766 12518 50818 12570
rect 19966 12350 20018 12402
rect 24782 12350 24834 12402
rect 25230 12350 25282 12402
rect 30270 12350 30322 12402
rect 31054 12350 31106 12402
rect 32398 12350 32450 12402
rect 33294 12350 33346 12402
rect 40238 12350 40290 12402
rect 41134 12350 41186 12402
rect 42590 12350 42642 12402
rect 43934 12350 43986 12402
rect 44606 12350 44658 12402
rect 47966 12350 48018 12402
rect 48190 12350 48242 12402
rect 48862 12350 48914 12402
rect 20974 12238 21026 12290
rect 23998 12238 24050 12290
rect 31278 12238 31330 12290
rect 31390 12238 31442 12290
rect 38670 12238 38722 12290
rect 44270 12238 44322 12290
rect 44382 12238 44434 12290
rect 47854 12238 47906 12290
rect 20302 12126 20354 12178
rect 20750 12126 20802 12178
rect 21534 12126 21586 12178
rect 21982 12126 22034 12178
rect 22542 12126 22594 12178
rect 23774 12126 23826 12178
rect 25454 12126 25506 12178
rect 25790 12126 25842 12178
rect 27694 12126 27746 12178
rect 28030 12126 28082 12178
rect 28702 12126 28754 12178
rect 29262 12126 29314 12178
rect 29710 12126 29762 12178
rect 30830 12126 30882 12178
rect 33966 12126 34018 12178
rect 34750 12126 34802 12178
rect 36206 12126 36258 12178
rect 36766 12126 36818 12178
rect 37886 12126 37938 12178
rect 38334 12126 38386 12178
rect 38894 12126 38946 12178
rect 39566 12126 39618 12178
rect 41470 12126 41522 12178
rect 42814 12126 42866 12178
rect 45054 12126 45106 12178
rect 45502 12126 45554 12178
rect 46062 12126 46114 12178
rect 47294 12126 47346 12178
rect 22206 12014 22258 12066
rect 25566 12014 25618 12066
rect 26126 12014 26178 12066
rect 26574 12014 26626 12066
rect 28142 12014 28194 12066
rect 31838 12014 31890 12066
rect 33630 12014 33682 12066
rect 35310 12014 35362 12066
rect 35758 12014 35810 12066
rect 37326 12014 37378 12066
rect 43262 12014 43314 12066
rect 45726 12014 45778 12066
rect 47406 12014 47458 12066
rect 22094 11902 22146 11954
rect 28814 11902 28866 11954
rect 36542 11902 36594 11954
rect 45390 11902 45442 11954
rect 4478 11734 4530 11786
rect 4582 11734 4634 11786
rect 4686 11734 4738 11786
rect 35198 11734 35250 11786
rect 35302 11734 35354 11786
rect 35406 11734 35458 11786
rect 19742 11566 19794 11618
rect 21198 11566 21250 11618
rect 21422 11566 21474 11618
rect 32062 11566 32114 11618
rect 38670 11566 38722 11618
rect 41470 11566 41522 11618
rect 19854 11454 19906 11506
rect 21534 11454 21586 11506
rect 22654 11454 22706 11506
rect 31950 11454 32002 11506
rect 32510 11454 32562 11506
rect 34302 11454 34354 11506
rect 36430 11454 36482 11506
rect 40462 11454 40514 11506
rect 46174 11454 46226 11506
rect 46510 11454 46562 11506
rect 48638 11454 48690 11506
rect 18398 11342 18450 11394
rect 18734 11342 18786 11394
rect 19518 11342 19570 11394
rect 20526 11342 20578 11394
rect 23326 11342 23378 11394
rect 29374 11342 29426 11394
rect 29822 11342 29874 11394
rect 30830 11342 30882 11394
rect 31054 11342 31106 11394
rect 31502 11342 31554 11394
rect 32958 11342 33010 11394
rect 33630 11342 33682 11394
rect 37214 11342 37266 11394
rect 37998 11342 38050 11394
rect 38110 11342 38162 11394
rect 39230 11342 39282 11394
rect 39902 11342 39954 11394
rect 41358 11342 41410 11394
rect 42142 11342 42194 11394
rect 42590 11342 42642 11394
rect 42926 11342 42978 11394
rect 43038 11342 43090 11394
rect 44830 11342 44882 11394
rect 45166 11342 45218 11394
rect 49310 11342 49362 11394
rect 20750 11230 20802 11282
rect 25342 11230 25394 11282
rect 33182 11230 33234 11282
rect 36990 11230 37042 11282
rect 39678 11230 39730 11282
rect 40462 11230 40514 11282
rect 40910 11230 40962 11282
rect 45502 11230 45554 11282
rect 46062 11230 46114 11282
rect 23102 11118 23154 11170
rect 32398 11118 32450 11170
rect 40238 11118 40290 11170
rect 44382 11118 44434 11170
rect 45390 11118 45442 11170
rect 19838 10950 19890 11002
rect 19942 10950 19994 11002
rect 20046 10950 20098 11002
rect 50558 10950 50610 11002
rect 50662 10950 50714 11002
rect 50766 10950 50818 11002
rect 32510 10782 32562 10834
rect 39678 10782 39730 10834
rect 41134 10782 41186 10834
rect 42254 10782 42306 10834
rect 31950 10670 32002 10722
rect 33070 10670 33122 10722
rect 35758 10670 35810 10722
rect 38782 10670 38834 10722
rect 21422 10558 21474 10610
rect 21870 10558 21922 10610
rect 27022 10558 27074 10610
rect 30382 10558 30434 10610
rect 33406 10558 33458 10610
rect 34302 10558 34354 10610
rect 34750 10558 34802 10610
rect 35534 10558 35586 10610
rect 36654 10558 36706 10610
rect 36766 10558 36818 10610
rect 37214 10558 37266 10610
rect 38334 10558 38386 10610
rect 46510 10558 46562 10610
rect 20974 10446 21026 10498
rect 22542 10446 22594 10498
rect 24670 10446 24722 10498
rect 27806 10446 27858 10498
rect 29934 10446 29986 10498
rect 30718 10446 30770 10498
rect 31614 10446 31666 10498
rect 37662 10446 37714 10498
rect 41918 10446 41970 10498
rect 42366 10446 42418 10498
rect 44830 10446 44882 10498
rect 31502 10334 31554 10386
rect 34078 10334 34130 10386
rect 36206 10334 36258 10386
rect 4478 10166 4530 10218
rect 4582 10166 4634 10218
rect 4686 10166 4738 10218
rect 35198 10166 35250 10218
rect 35302 10166 35354 10218
rect 35406 10166 35458 10218
rect 31614 9998 31666 10050
rect 25118 9886 25170 9938
rect 28366 9886 28418 9938
rect 31054 9886 31106 9938
rect 35982 9886 36034 9938
rect 36430 9886 36482 9938
rect 37438 9886 37490 9938
rect 38558 9886 38610 9938
rect 42254 9886 42306 9938
rect 43038 9886 43090 9938
rect 44382 9886 44434 9938
rect 47742 9886 47794 9938
rect 22206 9774 22258 9826
rect 25454 9774 25506 9826
rect 30494 9774 30546 9826
rect 30718 9774 30770 9826
rect 31278 9774 31330 9826
rect 32062 9774 32114 9826
rect 32510 9774 32562 9826
rect 33182 9774 33234 9826
rect 36990 9774 37042 9826
rect 38894 9774 38946 9826
rect 39342 9774 39394 9826
rect 42590 9774 42642 9826
rect 44830 9774 44882 9826
rect 22990 9662 23042 9714
rect 26238 9662 26290 9714
rect 33854 9662 33906 9714
rect 40126 9662 40178 9714
rect 45614 9662 45666 9714
rect 21646 9550 21698 9602
rect 29710 9550 29762 9602
rect 38110 9550 38162 9602
rect 19838 9382 19890 9434
rect 19942 9382 19994 9434
rect 20046 9382 20098 9434
rect 50558 9382 50610 9434
rect 50662 9382 50714 9434
rect 50766 9382 50818 9434
rect 22878 9214 22930 9266
rect 24446 9214 24498 9266
rect 32622 9214 32674 9266
rect 38782 9214 38834 9266
rect 39230 9214 39282 9266
rect 40238 9214 40290 9266
rect 40910 9214 40962 9266
rect 45614 9214 45666 9266
rect 46622 9214 46674 9266
rect 22990 9102 23042 9154
rect 24558 9102 24610 9154
rect 25342 9102 25394 9154
rect 30830 9102 30882 9154
rect 39678 9102 39730 9154
rect 40350 9102 40402 9154
rect 45502 9102 45554 9154
rect 23438 8990 23490 9042
rect 23886 8990 23938 9042
rect 25790 8990 25842 9042
rect 26574 8990 26626 9042
rect 27806 8990 27858 9042
rect 31614 8990 31666 9042
rect 38334 8990 38386 9042
rect 42366 8990 42418 9042
rect 26238 8878 26290 8930
rect 27918 8878 27970 8930
rect 28702 8878 28754 8930
rect 36318 8878 36370 8930
rect 41470 8878 41522 8930
rect 43038 8878 43090 8930
rect 45166 8878 45218 8930
rect 46062 8878 46114 8930
rect 26574 8766 26626 8818
rect 39566 8766 39618 8818
rect 45950 8766 46002 8818
rect 4478 8598 4530 8650
rect 4582 8598 4634 8650
rect 4686 8598 4738 8650
rect 35198 8598 35250 8650
rect 35302 8598 35354 8650
rect 35406 8598 35458 8650
rect 26462 8430 26514 8482
rect 33966 8430 34018 8482
rect 42478 8430 42530 8482
rect 24222 8318 24274 8370
rect 26574 8318 26626 8370
rect 28030 8318 28082 8370
rect 28142 8318 28194 8370
rect 31502 8318 31554 8370
rect 33630 8318 33682 8370
rect 34078 8318 34130 8370
rect 36318 8318 36370 8370
rect 39902 8318 39954 8370
rect 40686 8318 40738 8370
rect 42702 8318 42754 8370
rect 45726 8318 45778 8370
rect 47854 8318 47906 8370
rect 30830 8206 30882 8258
rect 36990 8206 37042 8258
rect 41806 8206 41858 8258
rect 42366 8206 42418 8258
rect 42926 8206 42978 8258
rect 43822 8206 43874 8258
rect 44942 8206 44994 8258
rect 36430 8094 36482 8146
rect 37774 8094 37826 8146
rect 44270 8094 44322 8146
rect 19838 7814 19890 7866
rect 19942 7814 19994 7866
rect 20046 7814 20098 7866
rect 50558 7814 50610 7866
rect 50662 7814 50714 7866
rect 50766 7814 50818 7866
rect 42254 7646 42306 7698
rect 45726 7646 45778 7698
rect 39566 7534 39618 7586
rect 40350 7422 40402 7474
rect 42926 7422 42978 7474
rect 43374 7422 43426 7474
rect 43822 7422 43874 7474
rect 44718 7422 44770 7474
rect 37438 7310 37490 7362
rect 42142 7310 42194 7362
rect 43710 7310 43762 7362
rect 45166 7310 45218 7362
rect 43150 7198 43202 7250
rect 4478 7030 4530 7082
rect 4582 7030 4634 7082
rect 4686 7030 4738 7082
rect 35198 7030 35250 7082
rect 35302 7030 35354 7082
rect 35406 7030 35458 7082
rect 19838 6246 19890 6298
rect 19942 6246 19994 6298
rect 20046 6246 20098 6298
rect 50558 6246 50610 6298
rect 50662 6246 50714 6298
rect 50766 6246 50818 6298
rect 42590 6078 42642 6130
rect 45614 5966 45666 6018
rect 43374 5854 43426 5906
rect 43598 5854 43650 5906
rect 44494 5854 44546 5906
rect 45278 5854 45330 5906
rect 29598 5742 29650 5794
rect 43822 5742 43874 5794
rect 45054 5630 45106 5682
rect 4478 5462 4530 5514
rect 4582 5462 4634 5514
rect 4686 5462 4738 5514
rect 35198 5462 35250 5514
rect 35302 5462 35354 5514
rect 35406 5462 35458 5514
rect 28702 5070 28754 5122
rect 29150 5070 29202 5122
rect 30046 5070 30098 5122
rect 29486 4958 29538 5010
rect 29822 4958 29874 5010
rect 19838 4678 19890 4730
rect 19942 4678 19994 4730
rect 20046 4678 20098 4730
rect 50558 4678 50610 4730
rect 50662 4678 50714 4730
rect 50766 4678 50818 4730
rect 26910 4510 26962 4562
rect 30830 4510 30882 4562
rect 27358 4286 27410 4338
rect 30494 4286 30546 4338
rect 16830 4174 16882 4226
rect 18398 4174 18450 4226
rect 19070 4174 19122 4226
rect 19742 4174 19794 4226
rect 20862 4174 20914 4226
rect 23550 4174 23602 4226
rect 24334 4174 24386 4226
rect 24670 4174 24722 4226
rect 30270 4174 30322 4226
rect 31390 4174 31442 4226
rect 33630 4174 33682 4226
rect 34302 4174 34354 4226
rect 36430 4174 36482 4226
rect 37102 4174 37154 4226
rect 37774 4174 37826 4226
rect 38446 4174 38498 4226
rect 39678 4174 39730 4226
rect 40350 4174 40402 4226
rect 41134 4174 41186 4226
rect 43374 4174 43426 4226
rect 44046 4174 44098 4226
rect 24222 4062 24274 4114
rect 24670 4062 24722 4114
rect 28142 4062 28194 4114
rect 4478 3894 4530 3946
rect 4582 3894 4634 3946
rect 4686 3894 4738 3946
rect 35198 3894 35250 3946
rect 35302 3894 35354 3946
rect 35406 3894 35458 3946
rect 29374 3614 29426 3666
rect 16270 3502 16322 3554
rect 17278 3502 17330 3554
rect 17950 3502 18002 3554
rect 18622 3502 18674 3554
rect 23214 3502 23266 3554
rect 23886 3502 23938 3554
rect 26014 3502 26066 3554
rect 27246 3502 27298 3554
rect 27582 3502 27634 3554
rect 28366 3502 28418 3554
rect 31502 3502 31554 3554
rect 33854 3502 33906 3554
rect 34526 3502 34578 3554
rect 36654 3502 36706 3554
rect 37326 3502 37378 3554
rect 38222 3502 38274 3554
rect 12686 3390 12738 3442
rect 13134 3390 13186 3442
rect 13470 3390 13522 3442
rect 15822 3390 15874 3442
rect 16046 3390 16098 3442
rect 17054 3390 17106 3442
rect 18174 3390 18226 3442
rect 18846 3390 18898 3442
rect 19182 3390 19234 3442
rect 19518 3390 19570 3442
rect 19854 3390 19906 3442
rect 20190 3390 20242 3442
rect 21086 3390 21138 3442
rect 21422 3390 21474 3442
rect 21870 3390 21922 3442
rect 22990 3390 23042 3442
rect 23662 3390 23714 3442
rect 24558 3390 24610 3442
rect 24894 3390 24946 3442
rect 25566 3390 25618 3442
rect 25790 3390 25842 3442
rect 26798 3390 26850 3442
rect 27806 3390 27858 3442
rect 31278 3390 31330 3442
rect 32958 3390 33010 3442
rect 33182 3390 33234 3442
rect 33518 3390 33570 3442
rect 34190 3390 34242 3442
rect 34862 3390 34914 3442
rect 35534 3390 35586 3442
rect 35982 3390 36034 3442
rect 36318 3390 36370 3442
rect 36990 3390 37042 3442
rect 37662 3390 37714 3442
rect 37998 3390 38050 3442
rect 38670 3390 38722 3442
rect 39006 3390 39058 3442
rect 39902 3390 39954 3442
rect 40238 3390 40290 3442
rect 40574 3390 40626 3442
rect 40910 3390 40962 3442
rect 41246 3390 41298 3442
rect 41582 3390 41634 3442
rect 42366 3390 42418 3442
rect 42590 3390 42642 3442
rect 42926 3390 42978 3442
rect 43598 3390 43650 3442
rect 43934 3390 43986 3442
rect 44270 3390 44322 3442
rect 44606 3390 44658 3442
rect 19838 3110 19890 3162
rect 19942 3110 19994 3162
rect 20046 3110 20098 3162
rect 50558 3110 50610 3162
rect 50662 3110 50714 3162
rect 50766 3110 50818 3162
<< metal2 >>
rect 19836 76860 20100 76870
rect 19892 76804 19940 76860
rect 19996 76804 20044 76860
rect 19836 76794 20100 76804
rect 50556 76860 50820 76870
rect 50612 76804 50660 76860
rect 50716 76804 50764 76860
rect 50556 76794 50820 76804
rect 4476 76076 4740 76086
rect 4532 76020 4580 76076
rect 4636 76020 4684 76076
rect 4476 76010 4740 76020
rect 35196 76076 35460 76086
rect 35252 76020 35300 76076
rect 35356 76020 35404 76076
rect 35196 76010 35460 76020
rect 19836 75292 20100 75302
rect 19892 75236 19940 75292
rect 19996 75236 20044 75292
rect 19836 75226 20100 75236
rect 50556 75292 50820 75302
rect 50612 75236 50660 75292
rect 50716 75236 50764 75292
rect 50556 75226 50820 75236
rect 4476 74508 4740 74518
rect 4532 74452 4580 74508
rect 4636 74452 4684 74508
rect 4476 74442 4740 74452
rect 35196 74508 35460 74518
rect 35252 74452 35300 74508
rect 35356 74452 35404 74508
rect 35196 74442 35460 74452
rect 19836 73724 20100 73734
rect 19892 73668 19940 73724
rect 19996 73668 20044 73724
rect 19836 73658 20100 73668
rect 50556 73724 50820 73734
rect 50612 73668 50660 73724
rect 50716 73668 50764 73724
rect 50556 73658 50820 73668
rect 4476 72940 4740 72950
rect 4532 72884 4580 72940
rect 4636 72884 4684 72940
rect 4476 72874 4740 72884
rect 35196 72940 35460 72950
rect 35252 72884 35300 72940
rect 35356 72884 35404 72940
rect 35196 72874 35460 72884
rect 19836 72156 20100 72166
rect 19892 72100 19940 72156
rect 19996 72100 20044 72156
rect 19836 72090 20100 72100
rect 50556 72156 50820 72166
rect 50612 72100 50660 72156
rect 50716 72100 50764 72156
rect 50556 72090 50820 72100
rect 40236 71988 40292 71998
rect 39116 71986 40292 71988
rect 39116 71934 40238 71986
rect 40290 71934 40292 71986
rect 39116 71932 40292 71934
rect 39116 71874 39172 71932
rect 40236 71922 40292 71932
rect 39116 71822 39118 71874
rect 39170 71822 39172 71874
rect 39116 71810 39172 71822
rect 39900 71762 39956 71774
rect 39900 71710 39902 71762
rect 39954 71710 39956 71762
rect 36988 71650 37044 71662
rect 36988 71598 36990 71650
rect 37042 71598 37044 71650
rect 4476 71372 4740 71382
rect 4532 71316 4580 71372
rect 4636 71316 4684 71372
rect 4476 71306 4740 71316
rect 35196 71372 35460 71382
rect 35252 71316 35300 71372
rect 35356 71316 35404 71372
rect 35196 71306 35460 71316
rect 34412 71092 34468 71102
rect 34412 71090 35028 71092
rect 34412 71038 34414 71090
rect 34466 71038 35028 71090
rect 34412 71036 35028 71038
rect 34412 71026 34468 71036
rect 31612 70978 31668 70990
rect 31612 70926 31614 70978
rect 31666 70926 31668 70978
rect 4172 70644 4228 70654
rect 2044 54628 2100 54638
rect 2044 54626 3332 54628
rect 2044 54574 2046 54626
rect 2098 54574 3332 54626
rect 2044 54572 3332 54574
rect 2044 54562 2100 54572
rect 1708 54514 1764 54526
rect 1708 54462 1710 54514
rect 1762 54462 1764 54514
rect 1708 54404 1764 54462
rect 1708 53844 1764 54348
rect 2492 54404 2548 54414
rect 2492 54310 2548 54348
rect 1708 53778 1764 53788
rect 1708 53618 1764 53630
rect 1708 53566 1710 53618
rect 1762 53566 1764 53618
rect 1708 53172 1764 53566
rect 2044 53508 2100 53518
rect 2044 53506 2324 53508
rect 2044 53454 2046 53506
rect 2098 53454 2324 53506
rect 2044 53452 2324 53454
rect 2044 53442 2100 53452
rect 1708 53106 1764 53116
rect 1596 53060 1652 53070
rect 1484 50596 1540 50606
rect 1484 43652 1540 50540
rect 1484 43586 1540 43596
rect 1596 41412 1652 53004
rect 2044 53060 2100 53070
rect 2044 52966 2100 53004
rect 1708 52946 1764 52958
rect 1708 52894 1710 52946
rect 1762 52894 1764 52946
rect 1708 52500 1764 52894
rect 1708 52434 1764 52444
rect 1708 52162 1764 52174
rect 1708 52110 1710 52162
rect 1762 52110 1764 52162
rect 1708 51828 1764 52110
rect 2044 51940 2100 51950
rect 2044 51938 2212 51940
rect 2044 51886 2046 51938
rect 2098 51886 2212 51938
rect 2044 51884 2212 51886
rect 2044 51874 2100 51884
rect 1708 51762 1764 51772
rect 2044 51492 2100 51502
rect 1932 51490 2100 51492
rect 1932 51438 2046 51490
rect 2098 51438 2100 51490
rect 1932 51436 2100 51438
rect 1708 51378 1764 51390
rect 1708 51326 1710 51378
rect 1762 51326 1764 51378
rect 1708 51156 1764 51326
rect 1708 51090 1764 51100
rect 1820 50594 1876 50606
rect 1820 50542 1822 50594
rect 1874 50542 1876 50594
rect 1820 50372 1876 50542
rect 1708 49810 1764 49822
rect 1708 49758 1710 49810
rect 1762 49758 1764 49810
rect 1708 49700 1764 49758
rect 1820 49812 1876 50316
rect 1820 49746 1876 49756
rect 1708 49140 1764 49644
rect 1932 49364 1988 51436
rect 2044 51426 2100 51436
rect 2044 50708 2100 50718
rect 2044 50482 2100 50652
rect 2044 50430 2046 50482
rect 2098 50430 2100 50482
rect 2044 50418 2100 50430
rect 1708 49074 1764 49084
rect 1820 49308 1988 49364
rect 2044 49922 2100 49934
rect 2044 49870 2046 49922
rect 2098 49870 2100 49922
rect 1708 46674 1764 46686
rect 1708 46622 1710 46674
rect 1762 46622 1764 46674
rect 1708 46452 1764 46622
rect 1708 46386 1764 46396
rect 1820 46116 1876 49308
rect 2044 49252 2100 49870
rect 2044 49186 2100 49196
rect 1932 49138 1988 49150
rect 1932 49086 1934 49138
rect 1986 49086 1988 49138
rect 1932 48468 1988 49086
rect 1932 48402 1988 48412
rect 1932 48020 1988 48030
rect 1932 47926 1988 47964
rect 1932 47570 1988 47582
rect 1932 47518 1934 47570
rect 1986 47518 1988 47570
rect 1932 47124 1988 47518
rect 1932 47058 1988 47068
rect 2044 46788 2100 46798
rect 2044 46694 2100 46732
rect 1820 46060 1988 46116
rect 1820 45890 1876 45902
rect 1820 45838 1822 45890
rect 1874 45838 1876 45890
rect 1708 45106 1764 45118
rect 1708 45054 1710 45106
rect 1762 45054 1764 45106
rect 1708 44996 1764 45054
rect 1820 45108 1876 45838
rect 1820 45042 1876 45052
rect 1708 44436 1764 44940
rect 1932 44884 1988 46060
rect 2044 45668 2100 45678
rect 2044 45574 2100 45612
rect 2044 45220 2100 45230
rect 2044 45126 2100 45164
rect 1932 44818 1988 44828
rect 1708 44370 1764 44380
rect 1708 44210 1764 44222
rect 1708 44158 1710 44210
rect 1762 44158 1764 44210
rect 1708 43764 1764 44158
rect 2044 44100 2100 44110
rect 2044 44006 2100 44044
rect 1708 43698 1764 43708
rect 2156 43428 2212 51884
rect 2268 48580 2324 53452
rect 2492 53506 2548 53518
rect 2492 53454 2494 53506
rect 2546 53454 2548 53506
rect 2492 53172 2548 53454
rect 2492 53106 2548 53116
rect 2492 52834 2548 52846
rect 2492 52782 2494 52834
rect 2546 52782 2548 52834
rect 2492 52500 2548 52782
rect 2492 52434 2548 52444
rect 2492 52162 2548 52174
rect 2492 52110 2494 52162
rect 2546 52110 2548 52162
rect 2492 51828 2548 52110
rect 2492 51762 2548 51772
rect 2492 51266 2548 51278
rect 2492 51214 2494 51266
rect 2546 51214 2548 51266
rect 2380 50484 2436 50494
rect 2380 50390 2436 50428
rect 2492 50372 2548 51214
rect 2940 51266 2996 51278
rect 2940 51214 2942 51266
rect 2994 51214 2996 51266
rect 2940 51156 2996 51214
rect 2940 51090 2996 51100
rect 2716 50596 2772 50606
rect 2716 50482 2772 50540
rect 2716 50430 2718 50482
rect 2770 50430 2772 50482
rect 2716 50418 2772 50430
rect 3164 50484 3220 50494
rect 3164 50390 3220 50428
rect 2492 50306 2548 50316
rect 2492 49700 2548 49710
rect 2492 49606 2548 49644
rect 2268 48524 2884 48580
rect 2492 46562 2548 46574
rect 2492 46510 2494 46562
rect 2546 46510 2548 46562
rect 2492 46004 2548 46510
rect 2268 45948 2548 46004
rect 2268 45108 2324 45948
rect 2380 45780 2436 45790
rect 2380 45686 2436 45724
rect 2268 45042 2324 45052
rect 2716 45666 2772 45678
rect 2716 45614 2718 45666
rect 2770 45614 2772 45666
rect 2492 44996 2548 45006
rect 2492 44902 2548 44940
rect 2716 44436 2772 45614
rect 2716 44370 2772 44380
rect 2492 44098 2548 44110
rect 2492 44046 2494 44098
rect 2546 44046 2548 44098
rect 2492 43764 2548 44046
rect 2492 43698 2548 43708
rect 2156 43362 2212 43372
rect 1932 43316 1988 43326
rect 1932 43222 1988 43260
rect 2828 42868 2884 48524
rect 3276 47124 3332 54572
rect 3276 47068 3444 47124
rect 2940 46562 2996 46574
rect 2940 46510 2942 46562
rect 2994 46510 2996 46562
rect 2940 46452 2996 46510
rect 2940 46386 2996 46396
rect 3164 45780 3220 45790
rect 3164 45686 3220 45724
rect 3388 44548 3444 47068
rect 3388 44482 3444 44492
rect 2828 42802 2884 42812
rect 1708 42642 1764 42654
rect 1708 42590 1710 42642
rect 1762 42590 1764 42642
rect 1708 42420 1764 42590
rect 1708 42354 1764 42364
rect 2044 42530 2100 42542
rect 2044 42478 2046 42530
rect 2098 42478 2100 42530
rect 2044 42308 2100 42478
rect 2492 42530 2548 42542
rect 2492 42478 2494 42530
rect 2546 42478 2548 42530
rect 2492 42420 2548 42478
rect 2492 42354 2548 42364
rect 2044 42242 2100 42252
rect 2044 42082 2100 42094
rect 2044 42030 2046 42082
rect 2098 42030 2100 42082
rect 1708 41970 1764 41982
rect 1708 41918 1710 41970
rect 1762 41918 1764 41970
rect 1708 41748 1764 41918
rect 2044 41972 2100 42030
rect 2044 41906 2100 41916
rect 1708 41682 1764 41692
rect 2492 41858 2548 41870
rect 2492 41806 2494 41858
rect 2546 41806 2548 41858
rect 2492 41748 2548 41806
rect 2492 41682 2548 41692
rect 1596 41346 1652 41356
rect 1708 41076 1764 41086
rect 1708 40982 1764 41020
rect 2380 41074 2436 41086
rect 2380 41022 2382 41074
rect 2434 41022 2436 41074
rect 2044 40964 2100 40974
rect 2044 40870 2100 40908
rect 2044 40514 2100 40526
rect 2044 40462 2046 40514
rect 2098 40462 2100 40514
rect 1708 40402 1764 40414
rect 1708 40350 1710 40402
rect 1762 40350 1764 40402
rect 1708 39732 1764 40350
rect 2044 40292 2100 40462
rect 2380 40404 2436 41022
rect 2492 41076 2548 41086
rect 2492 40626 2548 41020
rect 2716 41076 2772 41086
rect 2716 40982 2772 41020
rect 2492 40574 2494 40626
rect 2546 40574 2548 40626
rect 2492 40562 2548 40574
rect 3164 40962 3220 40974
rect 3164 40910 3166 40962
rect 3218 40910 3220 40962
rect 2380 40338 2436 40348
rect 2940 40402 2996 40414
rect 2940 40350 2942 40402
rect 2994 40350 2996 40402
rect 2044 40226 2100 40236
rect 1708 39666 1764 39676
rect 2940 39732 2996 40350
rect 3164 40404 3220 40910
rect 4172 40628 4228 70588
rect 19836 70588 20100 70598
rect 19892 70532 19940 70588
rect 19996 70532 20044 70588
rect 19836 70522 20100 70532
rect 31612 70532 31668 70926
rect 31612 70466 31668 70476
rect 32284 70866 32340 70878
rect 32284 70814 32286 70866
rect 32338 70814 32340 70866
rect 31052 70420 31108 70430
rect 30268 70418 31108 70420
rect 30268 70366 31054 70418
rect 31106 70366 31108 70418
rect 30268 70364 31108 70366
rect 32284 70420 32340 70814
rect 34860 70866 34916 70878
rect 34860 70814 34862 70866
rect 34914 70814 34916 70866
rect 34748 70756 34804 70766
rect 33964 70754 34804 70756
rect 33964 70702 34750 70754
rect 34802 70702 34804 70754
rect 33964 70700 34804 70702
rect 33180 70532 33236 70542
rect 32396 70420 32452 70430
rect 32284 70418 32452 70420
rect 32284 70366 32398 70418
rect 32450 70366 32452 70418
rect 32284 70364 32452 70366
rect 27804 70194 27860 70206
rect 27804 70142 27806 70194
rect 27858 70142 27860 70194
rect 23996 70084 24052 70094
rect 23996 70082 24612 70084
rect 23996 70030 23998 70082
rect 24050 70030 24612 70082
rect 23996 70028 24612 70030
rect 23996 70018 24052 70028
rect 22876 69972 22932 69982
rect 4476 69804 4740 69814
rect 4532 69748 4580 69804
rect 4636 69748 4684 69804
rect 4476 69738 4740 69748
rect 22876 69522 22932 69916
rect 23884 69972 23940 69982
rect 23884 69878 23940 69916
rect 22876 69470 22878 69522
rect 22930 69470 22932 69522
rect 22876 69458 22932 69470
rect 22204 69410 22260 69422
rect 22204 69358 22206 69410
rect 22258 69358 22260 69410
rect 19836 69020 20100 69030
rect 19892 68964 19940 69020
rect 19996 68964 20044 69020
rect 19836 68954 20100 68964
rect 22204 68964 22260 69358
rect 22204 68898 22260 68908
rect 22988 68964 23044 68974
rect 22764 68628 22820 68638
rect 22988 68628 23044 68908
rect 24556 68850 24612 70028
rect 25452 70082 25508 70094
rect 25452 70030 25454 70082
rect 25506 70030 25508 70082
rect 25004 69524 25060 69534
rect 24556 68798 24558 68850
rect 24610 68798 24612 68850
rect 24556 68786 24612 68798
rect 24668 69522 25060 69524
rect 24668 69470 25006 69522
rect 25058 69470 25060 69522
rect 24668 69468 25060 69470
rect 24668 68850 24724 69468
rect 25004 69458 25060 69468
rect 25340 69412 25396 69422
rect 25340 68964 25396 69356
rect 25340 68898 25396 68908
rect 24668 68798 24670 68850
rect 24722 68798 24724 68850
rect 23772 68738 23828 68750
rect 23772 68686 23774 68738
rect 23826 68686 23828 68738
rect 22764 68626 23044 68628
rect 22764 68574 22766 68626
rect 22818 68574 23044 68626
rect 22764 68572 23044 68574
rect 22764 68562 22820 68572
rect 19852 68514 19908 68526
rect 21980 68516 22036 68526
rect 19852 68462 19854 68514
rect 19906 68462 19908 68514
rect 4476 68236 4740 68246
rect 4532 68180 4580 68236
rect 4636 68180 4684 68236
rect 4476 68170 4740 68180
rect 19852 67844 19908 68462
rect 21420 68514 22036 68516
rect 21420 68462 21982 68514
rect 22034 68462 22036 68514
rect 21420 68460 22036 68462
rect 20748 68180 20804 68190
rect 21308 68180 21364 68190
rect 20748 67954 20804 68124
rect 20748 67902 20750 67954
rect 20802 67902 20804 67954
rect 20748 67890 20804 67902
rect 21196 68124 21308 68180
rect 19852 67778 19908 67788
rect 19836 67452 20100 67462
rect 19892 67396 19940 67452
rect 19996 67396 20044 67452
rect 19836 67386 20100 67396
rect 20524 67284 20580 67294
rect 20524 67190 20580 67228
rect 20300 67058 20356 67070
rect 20300 67006 20302 67058
rect 20354 67006 20356 67058
rect 15372 66946 15428 66958
rect 15372 66894 15374 66946
rect 15426 66894 15428 66946
rect 14252 66836 14308 66846
rect 4476 66668 4740 66678
rect 4532 66612 4580 66668
rect 4636 66612 4684 66668
rect 4476 66602 4740 66612
rect 14028 66500 14084 66510
rect 13692 66498 14084 66500
rect 13692 66446 14030 66498
rect 14082 66446 14084 66498
rect 13692 66444 14084 66446
rect 9884 65490 9940 65502
rect 9884 65438 9886 65490
rect 9938 65438 9940 65490
rect 4476 65100 4740 65110
rect 4532 65044 4580 65100
rect 4636 65044 4684 65100
rect 4476 65034 4740 65044
rect 9884 64820 9940 65438
rect 13132 65490 13188 65502
rect 13132 65438 13134 65490
rect 13186 65438 13188 65490
rect 10556 65378 10612 65390
rect 10556 65326 10558 65378
rect 10610 65326 10612 65378
rect 10108 64820 10164 64830
rect 9884 64764 10108 64820
rect 10108 64706 10164 64764
rect 10108 64654 10110 64706
rect 10162 64654 10164 64706
rect 10108 64642 10164 64654
rect 10556 63812 10612 65326
rect 12684 65380 12740 65390
rect 12684 65286 12740 65324
rect 12908 64818 12964 64830
rect 12908 64766 12910 64818
rect 12962 64766 12964 64818
rect 10780 64596 10836 64606
rect 10780 64594 11732 64596
rect 10780 64542 10782 64594
rect 10834 64542 11732 64594
rect 10780 64540 11732 64542
rect 10780 64530 10836 64540
rect 11676 64146 11732 64540
rect 11676 64094 11678 64146
rect 11730 64094 11732 64146
rect 11676 64082 11732 64094
rect 11788 64204 12852 64260
rect 11788 64146 11844 64204
rect 11788 64094 11790 64146
rect 11842 64094 11844 64146
rect 10556 63746 10612 63756
rect 11452 63922 11508 63934
rect 11452 63870 11454 63922
rect 11506 63870 11508 63922
rect 4476 63532 4740 63542
rect 4532 63476 4580 63532
rect 4636 63476 4684 63532
rect 4476 63466 4740 63476
rect 11452 63364 11508 63870
rect 11564 63924 11620 63934
rect 11564 63830 11620 63868
rect 11452 63298 11508 63308
rect 11788 63252 11844 64094
rect 12796 64146 12852 64204
rect 12796 64094 12798 64146
rect 12850 64094 12852 64146
rect 12796 64082 12852 64094
rect 12460 64036 12516 64046
rect 12460 63942 12516 63980
rect 11564 63196 11844 63252
rect 11900 63924 11956 63934
rect 11452 62916 11508 62926
rect 11116 62914 11508 62916
rect 11116 62862 11454 62914
rect 11506 62862 11508 62914
rect 11116 62860 11508 62862
rect 9660 62354 9716 62366
rect 9660 62302 9662 62354
rect 9714 62302 9716 62354
rect 4476 61964 4740 61974
rect 4532 61908 4580 61964
rect 4636 61908 4684 61964
rect 4476 61898 4740 61908
rect 9548 60786 9604 60798
rect 9548 60734 9550 60786
rect 9602 60734 9604 60786
rect 4476 60396 4740 60406
rect 4532 60340 4580 60396
rect 4636 60340 4684 60396
rect 4476 60330 4740 60340
rect 9548 59218 9604 60734
rect 9548 59166 9550 59218
rect 9602 59166 9604 59218
rect 8988 59106 9044 59118
rect 8988 59054 8990 59106
rect 9042 59054 9044 59106
rect 8876 58994 8932 59006
rect 8876 58942 8878 58994
rect 8930 58942 8932 58994
rect 4476 58828 4740 58838
rect 4532 58772 4580 58828
rect 4636 58772 4684 58828
rect 4476 58762 4740 58772
rect 6188 58548 6244 58558
rect 6188 57652 6244 58492
rect 5740 57650 6244 57652
rect 5740 57598 6190 57650
rect 6242 57598 6244 57650
rect 5740 57596 6244 57598
rect 4476 57260 4740 57270
rect 4532 57204 4580 57260
rect 4636 57204 4684 57260
rect 4476 57194 4740 57204
rect 5740 56866 5796 57596
rect 6188 57586 6244 57596
rect 6860 57538 6916 57550
rect 6860 57486 6862 57538
rect 6914 57486 6916 57538
rect 6860 56980 6916 57486
rect 6860 56914 6916 56924
rect 8540 56978 8596 56990
rect 8540 56926 8542 56978
rect 8594 56926 8596 56978
rect 5740 56814 5742 56866
rect 5794 56814 5796 56866
rect 4476 55692 4740 55702
rect 4532 55636 4580 55692
rect 4636 55636 4684 55692
rect 4476 55626 4740 55636
rect 5740 55298 5796 56814
rect 6412 56754 6468 56766
rect 6412 56702 6414 56754
rect 6466 56702 6468 56754
rect 6412 56308 6468 56702
rect 6412 56242 6468 56252
rect 7084 56308 7140 56318
rect 7140 56252 7252 56308
rect 7084 56242 7140 56252
rect 7196 56194 7252 56252
rect 7196 56142 7198 56194
rect 7250 56142 7252 56194
rect 7196 56130 7252 56142
rect 8428 56196 8484 56206
rect 8540 56196 8596 56926
rect 8876 56866 8932 58942
rect 8988 57652 9044 59054
rect 9548 57876 9604 59166
rect 9660 58548 9716 62302
rect 9996 62244 10052 62254
rect 9996 61682 10052 62188
rect 10332 62244 10388 62254
rect 10332 62242 10612 62244
rect 10332 62190 10334 62242
rect 10386 62190 10612 62242
rect 10332 62188 10612 62190
rect 10332 62178 10388 62188
rect 9996 61630 9998 61682
rect 10050 61630 10052 61682
rect 9996 61618 10052 61630
rect 10556 61682 10612 62188
rect 10556 61630 10558 61682
rect 10610 61630 10612 61682
rect 10556 61618 10612 61630
rect 10108 61572 10164 61582
rect 10444 61572 10500 61582
rect 10108 61570 10500 61572
rect 10108 61518 10110 61570
rect 10162 61518 10446 61570
rect 10498 61518 10500 61570
rect 10108 61516 10500 61518
rect 10108 61506 10164 61516
rect 10444 61506 10500 61516
rect 10668 61572 10724 61582
rect 10668 61478 10724 61516
rect 11116 61570 11172 62860
rect 11452 62850 11508 62860
rect 11452 62580 11508 62590
rect 11340 62524 11452 62580
rect 11340 62188 11396 62524
rect 11452 62514 11508 62524
rect 11564 62188 11620 63196
rect 11788 63026 11844 63038
rect 11788 62974 11790 63026
rect 11842 62974 11844 63026
rect 11676 62914 11732 62926
rect 11676 62862 11678 62914
rect 11730 62862 11732 62914
rect 11676 62580 11732 62862
rect 11676 62514 11732 62524
rect 11340 62132 11508 62188
rect 11564 62132 11732 62188
rect 11452 61684 11508 62132
rect 11452 61628 11620 61684
rect 11116 61518 11118 61570
rect 11170 61518 11172 61570
rect 11116 61506 11172 61518
rect 11452 61458 11508 61470
rect 11452 61406 11454 61458
rect 11506 61406 11508 61458
rect 10332 61348 10388 61358
rect 10332 60898 10388 61292
rect 10892 61346 10948 61358
rect 10892 61294 10894 61346
rect 10946 61294 10948 61346
rect 10892 61012 10948 61294
rect 10892 60946 10948 60956
rect 10332 60846 10334 60898
rect 10386 60846 10388 60898
rect 10332 60834 10388 60846
rect 11452 60002 11508 61406
rect 11452 59950 11454 60002
rect 11506 59950 11508 60002
rect 11452 59938 11508 59950
rect 11564 59892 11620 61628
rect 11676 61346 11732 62132
rect 11788 61796 11844 62974
rect 11900 62132 11956 63868
rect 12012 63924 12068 63934
rect 12572 63924 12628 63934
rect 12012 63922 12404 63924
rect 12012 63870 12014 63922
rect 12066 63870 12404 63922
rect 12012 63868 12404 63870
rect 12012 63858 12068 63868
rect 12348 63140 12404 63868
rect 12572 63830 12628 63868
rect 12460 63812 12516 63822
rect 12460 63718 12516 63756
rect 12908 63588 12964 64766
rect 13132 64820 13188 65438
rect 13132 64754 13188 64764
rect 13692 64706 13748 66444
rect 14028 66434 14084 66444
rect 13916 66162 13972 66174
rect 13916 66110 13918 66162
rect 13970 66110 13972 66162
rect 13804 65378 13860 65390
rect 13804 65326 13806 65378
rect 13858 65326 13860 65378
rect 13804 64820 13860 65326
rect 13916 65380 13972 66110
rect 14028 66050 14084 66062
rect 14028 65998 14030 66050
rect 14082 65998 14084 66050
rect 14028 65716 14084 65998
rect 14028 65650 14084 65660
rect 13916 65044 13972 65324
rect 13916 64988 14196 65044
rect 13916 64820 13972 64830
rect 13804 64818 13972 64820
rect 13804 64766 13918 64818
rect 13970 64766 13972 64818
rect 13804 64764 13972 64766
rect 13916 64754 13972 64764
rect 13692 64654 13694 64706
rect 13746 64654 13748 64706
rect 13692 64642 13748 64654
rect 13804 64482 13860 64494
rect 13804 64430 13806 64482
rect 13858 64430 13860 64482
rect 13804 64260 13860 64430
rect 14028 64484 14084 64494
rect 14028 64390 14084 64428
rect 13468 64034 13524 64046
rect 13468 63982 13470 64034
rect 13522 63982 13524 64034
rect 13020 63924 13076 63934
rect 13020 63830 13076 63868
rect 13356 63922 13412 63934
rect 13356 63870 13358 63922
rect 13410 63870 13412 63922
rect 13356 63588 13412 63870
rect 13468 63812 13524 63982
rect 13692 63924 13748 63934
rect 13692 63830 13748 63868
rect 13468 63746 13524 63756
rect 12684 63532 13412 63588
rect 12572 63364 12628 63374
rect 12572 63270 12628 63308
rect 12684 63250 12740 63532
rect 12684 63198 12686 63250
rect 12738 63198 12740 63250
rect 12684 63186 12740 63198
rect 12348 63084 12516 63140
rect 12460 62580 12516 63084
rect 12684 62580 12740 62590
rect 12460 62578 12740 62580
rect 12460 62526 12686 62578
rect 12738 62526 12740 62578
rect 12460 62524 12740 62526
rect 12684 62514 12740 62524
rect 12908 62580 12964 62590
rect 12908 62486 12964 62524
rect 13020 62354 13076 62366
rect 13020 62302 13022 62354
rect 13074 62302 13076 62354
rect 12460 62244 12516 62254
rect 12460 62150 12516 62188
rect 13020 62244 13076 62302
rect 13020 62178 13076 62188
rect 11900 62066 11956 62076
rect 11788 61740 12516 61796
rect 11900 61572 11956 61582
rect 11900 61478 11956 61516
rect 12124 61570 12180 61582
rect 12124 61518 12126 61570
rect 12178 61518 12180 61570
rect 11676 61294 11678 61346
rect 11730 61294 11732 61346
rect 11676 61012 11732 61294
rect 11788 61348 11844 61358
rect 11788 61254 11844 61292
rect 11676 60946 11732 60956
rect 12124 60226 12180 61518
rect 12460 60676 12516 61740
rect 12572 61572 12628 61582
rect 12572 61458 12628 61516
rect 12572 61406 12574 61458
rect 12626 61406 12628 61458
rect 12572 61394 12628 61406
rect 13804 61460 13860 64204
rect 13916 64036 13972 64046
rect 13916 63942 13972 63980
rect 14028 64036 14084 64046
rect 14140 64036 14196 64988
rect 14252 64706 14308 66780
rect 15260 66836 15316 66846
rect 15260 66742 15316 66780
rect 14476 66274 14532 66286
rect 14476 66222 14478 66274
rect 14530 66222 14532 66274
rect 14252 64654 14254 64706
rect 14306 64654 14308 64706
rect 14252 64642 14308 64654
rect 14364 64820 14420 64830
rect 14476 64820 14532 66222
rect 15260 66162 15316 66174
rect 15260 66110 15262 66162
rect 15314 66110 15316 66162
rect 14924 65716 14980 65726
rect 14812 65660 14924 65716
rect 14420 64764 14644 64820
rect 14028 64034 14196 64036
rect 14028 63982 14030 64034
rect 14082 63982 14196 64034
rect 14028 63980 14196 63982
rect 14028 63970 14084 63980
rect 14252 63028 14308 63038
rect 14364 63028 14420 64764
rect 14588 64706 14644 64764
rect 14588 64654 14590 64706
rect 14642 64654 14644 64706
rect 14588 64642 14644 64654
rect 14476 64596 14532 64606
rect 14476 63140 14532 64540
rect 14812 64148 14868 65660
rect 14924 65650 14980 65660
rect 15260 65492 15316 66110
rect 15260 65426 15316 65436
rect 15372 65380 15428 66894
rect 19852 66948 19908 66958
rect 19852 66946 20020 66948
rect 19852 66894 19854 66946
rect 19906 66894 20020 66946
rect 19852 66892 20020 66894
rect 19852 66882 19908 66892
rect 17388 66388 17444 66398
rect 17388 66386 17556 66388
rect 17388 66334 17390 66386
rect 17442 66334 17556 66386
rect 17388 66332 17556 66334
rect 17388 66322 17444 66332
rect 16380 65716 16436 65726
rect 16380 65622 16436 65660
rect 16492 65604 16548 65614
rect 16492 65510 16548 65548
rect 17500 65604 17556 66332
rect 19964 66276 20020 66892
rect 20300 66276 20356 67006
rect 21084 67060 21140 67070
rect 21084 66966 21140 67004
rect 19964 66274 20356 66276
rect 19964 66222 19966 66274
rect 20018 66222 20356 66274
rect 19964 66220 20356 66222
rect 19964 66210 20020 66220
rect 20188 66052 20244 66062
rect 19836 65884 20100 65894
rect 19892 65828 19940 65884
rect 19996 65828 20044 65884
rect 19836 65818 20100 65828
rect 17500 65538 17556 65548
rect 18508 65604 18564 65614
rect 18508 65510 18564 65548
rect 16156 65492 16212 65502
rect 16044 65490 16212 65492
rect 16044 65438 16158 65490
rect 16210 65438 16212 65490
rect 16044 65436 16212 65438
rect 15932 65380 15988 65390
rect 15372 65378 15988 65380
rect 15372 65326 15934 65378
rect 15986 65326 15988 65378
rect 15372 65324 15988 65326
rect 14700 64146 14868 64148
rect 14700 64094 14814 64146
rect 14866 64094 14868 64146
rect 14700 64092 14868 64094
rect 14700 63812 14756 64092
rect 14812 64082 14868 64092
rect 15036 64596 15092 64606
rect 14924 64036 14980 64046
rect 14924 63942 14980 63980
rect 15036 63812 15092 64540
rect 15372 64594 15428 64606
rect 15372 64542 15374 64594
rect 15426 64542 15428 64594
rect 14700 63746 14756 63756
rect 14812 63756 15092 63812
rect 15148 64484 15204 64494
rect 14812 63698 14868 63756
rect 14812 63646 14814 63698
rect 14866 63646 14868 63698
rect 14812 63634 14868 63646
rect 14476 63084 14756 63140
rect 14252 63026 14420 63028
rect 14252 62974 14254 63026
rect 14306 62974 14420 63026
rect 14252 62972 14420 62974
rect 14252 61570 14308 62972
rect 14700 62188 14756 63084
rect 15148 62580 15204 64428
rect 15372 64148 15428 64542
rect 15372 64082 15428 64092
rect 15596 64260 15652 64270
rect 15596 64146 15652 64204
rect 15596 64094 15598 64146
rect 15650 64094 15652 64146
rect 15596 64082 15652 64094
rect 15260 64034 15316 64046
rect 15260 63982 15262 64034
rect 15314 63982 15316 64034
rect 15260 63812 15316 63982
rect 15932 64036 15988 65324
rect 15932 63970 15988 63980
rect 16044 63922 16100 65436
rect 16156 65426 16212 65436
rect 17388 65490 17444 65502
rect 17388 65438 17390 65490
rect 17442 65438 17444 65490
rect 16380 64932 16436 64942
rect 16380 64484 16436 64876
rect 17388 64596 17444 65438
rect 17612 65490 17668 65502
rect 17612 65438 17614 65490
rect 17666 65438 17668 65490
rect 17388 64530 17444 64540
rect 17500 64818 17556 64830
rect 17500 64766 17502 64818
rect 17554 64766 17556 64818
rect 16044 63870 16046 63922
rect 16098 63870 16100 63922
rect 16044 63858 16100 63870
rect 16156 64372 16212 64382
rect 16156 64146 16212 64316
rect 16156 64094 16158 64146
rect 16210 64094 16212 64146
rect 15260 63746 15316 63756
rect 15820 62580 15876 62590
rect 14252 61518 14254 61570
rect 14306 61518 14308 61570
rect 13916 61460 13972 61470
rect 13804 61458 13972 61460
rect 13804 61406 13918 61458
rect 13970 61406 13972 61458
rect 13804 61404 13972 61406
rect 13916 61394 13972 61404
rect 12908 61348 12964 61358
rect 12908 61254 12964 61292
rect 13580 61346 13636 61358
rect 13580 61294 13582 61346
rect 13634 61294 13636 61346
rect 12796 61012 12852 61022
rect 12796 60918 12852 60956
rect 13132 60788 13188 60798
rect 13132 60694 13188 60732
rect 13580 60788 13636 61294
rect 13580 60722 13636 60732
rect 13916 60788 13972 60798
rect 12124 60174 12126 60226
rect 12178 60174 12180 60226
rect 12124 60162 12180 60174
rect 12236 60674 12516 60676
rect 12236 60622 12462 60674
rect 12514 60622 12516 60674
rect 12236 60620 12516 60622
rect 12236 60114 12292 60620
rect 12460 60610 12516 60620
rect 12236 60062 12238 60114
rect 12290 60062 12292 60114
rect 12236 60050 12292 60062
rect 11676 59892 11732 59902
rect 11564 59890 11732 59892
rect 11564 59838 11678 59890
rect 11730 59838 11732 59890
rect 11564 59836 11732 59838
rect 10332 59108 10388 59118
rect 10332 59106 10724 59108
rect 10332 59054 10334 59106
rect 10386 59054 10724 59106
rect 10332 59052 10724 59054
rect 10332 59042 10388 59052
rect 9660 58454 9716 58492
rect 9548 57810 9604 57820
rect 10668 57874 10724 59052
rect 11564 58660 11620 59836
rect 11676 59826 11732 59836
rect 11788 59890 11844 59902
rect 11788 59838 11790 59890
rect 11842 59838 11844 59890
rect 10668 57822 10670 57874
rect 10722 57822 10724 57874
rect 10668 57810 10724 57822
rect 11228 58604 11620 58660
rect 11788 58660 11844 59838
rect 12460 59106 12516 59118
rect 12460 59054 12462 59106
rect 12514 59054 12516 59106
rect 12460 58660 12516 59054
rect 11788 58604 12516 58660
rect 9660 57762 9716 57774
rect 9660 57710 9662 57762
rect 9714 57710 9716 57762
rect 9548 57652 9604 57662
rect 8988 57650 9604 57652
rect 8988 57598 9550 57650
rect 9602 57598 9604 57650
rect 8988 57596 9604 57598
rect 8988 57538 9044 57596
rect 9548 57586 9604 57596
rect 8988 57486 8990 57538
rect 9042 57486 9044 57538
rect 8988 57474 9044 57486
rect 8988 56980 9044 56990
rect 8988 56886 9044 56924
rect 9436 56868 9492 56878
rect 8876 56814 8878 56866
rect 8930 56814 8932 56866
rect 8876 56802 8932 56814
rect 9212 56866 9492 56868
rect 9212 56814 9438 56866
rect 9490 56814 9492 56866
rect 9212 56812 9492 56814
rect 9100 56756 9156 56766
rect 9100 56662 9156 56700
rect 8876 56644 8932 56654
rect 8764 56196 8820 56206
rect 8428 56194 8820 56196
rect 8428 56142 8430 56194
rect 8482 56142 8766 56194
rect 8818 56142 8820 56194
rect 8428 56140 8820 56142
rect 8428 56130 8484 56140
rect 8764 56130 8820 56140
rect 8876 56194 8932 56588
rect 9100 56308 9156 56318
rect 9212 56308 9268 56812
rect 9436 56802 9492 56812
rect 9324 56644 9380 56654
rect 9660 56644 9716 57710
rect 9324 56642 9492 56644
rect 9324 56590 9326 56642
rect 9378 56590 9492 56642
rect 9324 56588 9492 56590
rect 9324 56578 9380 56588
rect 9100 56306 9268 56308
rect 9100 56254 9102 56306
rect 9154 56254 9268 56306
rect 9100 56252 9268 56254
rect 9324 56420 9380 56430
rect 9100 56242 9156 56252
rect 8876 56142 8878 56194
rect 8930 56142 8932 56194
rect 6972 56084 7028 56094
rect 6972 55990 7028 56028
rect 7084 56082 7140 56094
rect 7084 56030 7086 56082
rect 7138 56030 7140 56082
rect 5740 55246 5742 55298
rect 5794 55246 5796 55298
rect 5740 55234 5796 55246
rect 6636 55860 6692 55870
rect 6412 55188 6468 55198
rect 6412 55186 6580 55188
rect 6412 55134 6414 55186
rect 6466 55134 6580 55186
rect 6412 55132 6580 55134
rect 6412 55122 6468 55132
rect 6524 54404 6580 55132
rect 6636 54738 6692 55804
rect 7084 54964 7140 56030
rect 6636 54686 6638 54738
rect 6690 54686 6692 54738
rect 6636 54674 6692 54686
rect 6748 54908 7140 54964
rect 7308 56082 7364 56094
rect 7308 56030 7310 56082
rect 7362 56030 7364 56082
rect 6748 54738 6804 54908
rect 6748 54686 6750 54738
rect 6802 54686 6804 54738
rect 6636 54404 6692 54414
rect 6524 54402 6692 54404
rect 6524 54350 6638 54402
rect 6690 54350 6692 54402
rect 6524 54348 6692 54350
rect 6636 54338 6692 54348
rect 4476 54124 4740 54134
rect 4532 54068 4580 54124
rect 4636 54068 4684 54124
rect 4476 54058 4740 54068
rect 5292 53844 5348 53854
rect 5292 53058 5348 53788
rect 6636 53844 6692 53854
rect 6636 53750 6692 53788
rect 6748 53730 6804 54686
rect 6748 53678 6750 53730
rect 6802 53678 6804 53730
rect 6636 53508 6692 53518
rect 6636 53414 6692 53452
rect 5292 53006 5294 53058
rect 5346 53006 5348 53058
rect 5292 52994 5348 53006
rect 6748 53060 6804 53678
rect 4620 52948 4676 52958
rect 4620 52946 4900 52948
rect 4620 52894 4622 52946
rect 4674 52894 4900 52946
rect 4620 52892 4900 52894
rect 4620 52882 4676 52892
rect 4476 52556 4740 52566
rect 4532 52500 4580 52556
rect 4636 52500 4684 52556
rect 4476 52490 4740 52500
rect 4620 51380 4676 51390
rect 4844 51380 4900 52892
rect 6524 52388 6580 52398
rect 5292 52276 5348 52286
rect 5292 51490 5348 52220
rect 6524 52162 6580 52332
rect 6636 52276 6692 52286
rect 6636 52182 6692 52220
rect 6524 52110 6526 52162
rect 6578 52110 6580 52162
rect 6524 52098 6580 52110
rect 6748 52162 6804 53004
rect 6748 52110 6750 52162
rect 6802 52110 6804 52162
rect 6748 52098 6804 52110
rect 6972 54740 7028 54750
rect 7308 54740 7364 56030
rect 6972 54738 7364 54740
rect 6972 54686 6974 54738
rect 7026 54686 7364 54738
rect 6972 54684 7364 54686
rect 7420 56082 7476 56094
rect 7420 56030 7422 56082
rect 7474 56030 7476 56082
rect 7420 54738 7476 56030
rect 8092 56084 8148 56094
rect 8316 56084 8372 56094
rect 8148 56082 8372 56084
rect 8148 56030 8318 56082
rect 8370 56030 8372 56082
rect 8148 56028 8372 56030
rect 8092 56018 8148 56028
rect 8316 56018 8372 56028
rect 7980 55970 8036 55982
rect 7980 55918 7982 55970
rect 8034 55918 8036 55970
rect 7868 55860 7924 55870
rect 7868 55766 7924 55804
rect 7980 55412 8036 55918
rect 8540 55412 8596 55422
rect 7980 55410 8596 55412
rect 7980 55358 8542 55410
rect 8594 55358 8596 55410
rect 7980 55356 8596 55358
rect 7420 54686 7422 54738
rect 7474 54686 7476 54738
rect 6972 53730 7028 54684
rect 7420 54674 7476 54686
rect 7644 54740 7700 54750
rect 7644 54646 7700 54684
rect 7756 54628 7812 54638
rect 7980 54628 8036 55356
rect 8540 55346 8596 55356
rect 8652 54740 8708 54750
rect 8876 54740 8932 56142
rect 9324 55410 9380 56364
rect 9436 56084 9492 56588
rect 9660 56578 9716 56588
rect 9884 57650 9940 57662
rect 9884 57598 9886 57650
rect 9938 57598 9940 57650
rect 9884 56194 9940 57598
rect 10444 57652 10500 57662
rect 10444 57558 10500 57596
rect 10556 57650 10612 57662
rect 10556 57598 10558 57650
rect 10610 57598 10612 57650
rect 10332 56754 10388 56766
rect 10332 56702 10334 56754
rect 10386 56702 10388 56754
rect 9996 56644 10052 56654
rect 10220 56644 10276 56654
rect 9996 56642 10164 56644
rect 9996 56590 9998 56642
rect 10050 56590 10164 56642
rect 9996 56588 10164 56590
rect 9996 56578 10052 56588
rect 10108 56308 10164 56588
rect 10220 56550 10276 56588
rect 10332 56420 10388 56702
rect 10332 56354 10388 56364
rect 10444 56756 10500 56766
rect 10556 56756 10612 57598
rect 10780 57652 10836 57662
rect 10780 57650 10948 57652
rect 10780 57598 10782 57650
rect 10834 57598 10948 57650
rect 10780 57596 10948 57598
rect 10780 57586 10836 57596
rect 10500 56700 10612 56756
rect 10780 56754 10836 56766
rect 10780 56702 10782 56754
rect 10834 56702 10836 56754
rect 10108 56252 10276 56308
rect 9884 56142 9886 56194
rect 9938 56142 9940 56194
rect 9884 56130 9940 56142
rect 9548 56084 9604 56094
rect 10108 56084 10164 56094
rect 9436 56028 9548 56084
rect 9548 56018 9604 56028
rect 9996 56028 10108 56084
rect 9324 55358 9326 55410
rect 9378 55358 9380 55410
rect 9324 55346 9380 55358
rect 8708 54684 8932 54740
rect 8652 54646 8708 54684
rect 7756 54626 8036 54628
rect 7756 54574 7758 54626
rect 7810 54574 8036 54626
rect 7756 54572 8036 54574
rect 7756 54562 7812 54572
rect 7196 54516 7252 54526
rect 8876 54516 8932 54526
rect 9660 54516 9716 54526
rect 7196 54514 7476 54516
rect 7196 54462 7198 54514
rect 7250 54462 7476 54514
rect 7196 54460 7476 54462
rect 7196 54450 7252 54460
rect 6972 53678 6974 53730
rect 7026 53678 7028 53730
rect 6972 53172 7028 53678
rect 7420 53730 7476 54460
rect 8652 54514 8932 54516
rect 8652 54462 8878 54514
rect 8930 54462 8932 54514
rect 8652 54460 8932 54462
rect 7756 53732 7812 53742
rect 8204 53732 8260 53742
rect 7420 53678 7422 53730
rect 7474 53678 7476 53730
rect 7420 53666 7476 53678
rect 7532 53730 8260 53732
rect 7532 53678 7758 53730
rect 7810 53678 8206 53730
rect 8258 53678 8260 53730
rect 7532 53676 8260 53678
rect 7196 53620 7252 53630
rect 7196 53618 7364 53620
rect 7196 53566 7198 53618
rect 7250 53566 7364 53618
rect 7196 53564 7364 53566
rect 7196 53554 7252 53564
rect 6972 52162 7028 53116
rect 6972 52110 6974 52162
rect 7026 52110 7028 52162
rect 6972 52098 7028 52110
rect 7084 52162 7140 52174
rect 7084 52110 7086 52162
rect 7138 52110 7140 52162
rect 5292 51438 5294 51490
rect 5346 51438 5348 51490
rect 5292 51426 5348 51438
rect 4620 51378 4900 51380
rect 4620 51326 4622 51378
rect 4674 51326 4900 51378
rect 4620 51324 4900 51326
rect 4620 51314 4676 51324
rect 4476 50988 4740 50998
rect 4532 50932 4580 50988
rect 4636 50932 4684 50988
rect 4476 50922 4740 50932
rect 4476 49420 4740 49430
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4476 49354 4740 49364
rect 4844 49140 4900 51324
rect 7084 50818 7140 52110
rect 7308 52164 7364 53564
rect 7420 52836 7476 52846
rect 7532 52836 7588 53676
rect 7756 53666 7812 53676
rect 8204 53666 8260 53676
rect 7420 52834 7588 52836
rect 7420 52782 7422 52834
rect 7474 52782 7588 52834
rect 7420 52780 7588 52782
rect 7644 53506 7700 53518
rect 7644 53454 7646 53506
rect 7698 53454 7700 53506
rect 7420 52770 7476 52780
rect 7420 52164 7476 52174
rect 7308 52162 7476 52164
rect 7308 52110 7422 52162
rect 7474 52110 7476 52162
rect 7308 52108 7476 52110
rect 7420 52098 7476 52108
rect 7644 52052 7700 53454
rect 8092 53508 8148 53518
rect 8092 53414 8148 53452
rect 8428 53172 8484 53182
rect 8428 53078 8484 53116
rect 8652 53172 8708 54460
rect 8876 54450 8932 54460
rect 9548 54514 9716 54516
rect 9548 54462 9662 54514
rect 9714 54462 9716 54514
rect 9548 54460 9716 54462
rect 9436 53732 9492 53742
rect 9436 53618 9492 53676
rect 9436 53566 9438 53618
rect 9490 53566 9492 53618
rect 9436 53554 9492 53566
rect 7756 53060 7812 53070
rect 7756 52966 7812 53004
rect 8092 52948 8148 52958
rect 8316 52948 8372 52958
rect 8092 52946 8316 52948
rect 8092 52894 8094 52946
rect 8146 52894 8316 52946
rect 8092 52892 8316 52894
rect 8092 52882 8148 52892
rect 8092 52388 8148 52398
rect 8092 52294 8148 52332
rect 8204 52164 8260 52174
rect 7980 52162 8260 52164
rect 7980 52110 8206 52162
rect 8258 52110 8260 52162
rect 7980 52108 8260 52110
rect 7532 52050 7700 52052
rect 7532 51998 7646 52050
rect 7698 51998 7700 52050
rect 7532 51996 7700 51998
rect 7532 51492 7588 51996
rect 7644 51986 7700 51996
rect 7756 52052 7812 52062
rect 7980 52052 8036 52108
rect 8204 52098 8260 52108
rect 7756 52050 8036 52052
rect 7756 51998 7758 52050
rect 7810 51998 8036 52050
rect 7756 51996 8036 51998
rect 7084 50766 7086 50818
rect 7138 50766 7140 50818
rect 7084 50754 7140 50766
rect 7308 51436 7588 51492
rect 4844 49074 4900 49084
rect 5404 50708 5460 50718
rect 4284 49026 4340 49038
rect 4284 48974 4286 49026
rect 4338 48974 4340 49026
rect 4284 48916 4340 48974
rect 4284 48850 4340 48860
rect 4732 48916 4788 48926
rect 4732 48822 4788 48860
rect 4284 48242 4340 48254
rect 4284 48190 4286 48242
rect 4338 48190 4340 48242
rect 4284 48132 4340 48190
rect 4844 48132 4900 48142
rect 4284 48130 4900 48132
rect 4284 48078 4846 48130
rect 4898 48078 4900 48130
rect 4284 48076 4900 48078
rect 4476 47852 4740 47862
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4476 47786 4740 47796
rect 4284 47458 4340 47470
rect 4284 47406 4286 47458
rect 4338 47406 4340 47458
rect 4284 47236 4340 47406
rect 4844 47460 4900 48076
rect 4844 47394 4900 47404
rect 4732 47236 4788 47246
rect 4284 47234 4788 47236
rect 4284 47182 4734 47234
rect 4786 47182 4788 47234
rect 4284 47180 4788 47182
rect 4732 47124 4788 47180
rect 4732 47068 5124 47124
rect 4620 47012 4676 47022
rect 4620 46674 4676 46956
rect 4620 46622 4622 46674
rect 4674 46622 4676 46674
rect 4620 46610 4676 46622
rect 4476 46284 4740 46294
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4476 46218 4740 46228
rect 4476 44716 4740 44726
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4476 44650 4740 44660
rect 5068 44660 5124 47068
rect 5292 47012 5348 47022
rect 5180 46956 5292 47012
rect 5180 45108 5236 46956
rect 5292 46946 5348 46956
rect 5292 46564 5348 46574
rect 5292 46470 5348 46508
rect 5404 46340 5460 50652
rect 7308 50708 7364 51436
rect 7420 51268 7476 51278
rect 7756 51268 7812 51996
rect 7420 51266 7812 51268
rect 7420 51214 7422 51266
rect 7474 51214 7812 51266
rect 7420 51212 7812 51214
rect 7420 51202 7476 51212
rect 7308 50652 8260 50708
rect 7196 50594 7252 50606
rect 7196 50542 7198 50594
rect 7250 50542 7252 50594
rect 7084 50484 7140 50522
rect 6748 49980 7028 50036
rect 5628 49140 5684 49150
rect 5628 49028 5684 49084
rect 5628 49026 5908 49028
rect 5628 48974 5630 49026
rect 5682 48974 5908 49026
rect 5628 48972 5908 48974
rect 5628 48962 5684 48972
rect 5852 47570 5908 48972
rect 6412 48914 6468 48926
rect 6412 48862 6414 48914
rect 6466 48862 6468 48914
rect 6412 48468 6468 48862
rect 6412 48402 6468 48412
rect 6300 48130 6356 48142
rect 6300 48078 6302 48130
rect 6354 48078 6356 48130
rect 6300 48020 6356 48078
rect 6300 47954 6356 47964
rect 6412 48018 6468 48030
rect 6412 47966 6414 48018
rect 6466 47966 6468 48018
rect 5852 47518 5854 47570
rect 5906 47518 5908 47570
rect 5852 47012 5908 47518
rect 5852 46946 5908 46956
rect 6412 46900 6468 47966
rect 6748 48020 6804 49980
rect 6860 49810 6916 49822
rect 6860 49758 6862 49810
rect 6914 49758 6916 49810
rect 6860 48242 6916 49758
rect 6972 49812 7028 49980
rect 7084 50034 7140 50428
rect 7084 49982 7086 50034
rect 7138 49982 7140 50034
rect 7084 49970 7140 49982
rect 7196 50036 7252 50542
rect 7308 50484 7364 50652
rect 7308 50418 7364 50428
rect 7868 50484 7924 50494
rect 7196 49970 7252 49980
rect 7756 50372 7812 50382
rect 7532 49924 7588 49934
rect 7308 49922 7700 49924
rect 7308 49870 7534 49922
rect 7586 49870 7700 49922
rect 7308 49868 7700 49870
rect 7196 49812 7252 49822
rect 6972 49810 7252 49812
rect 6972 49758 7198 49810
rect 7250 49758 7252 49810
rect 6972 49756 7252 49758
rect 7196 49746 7252 49756
rect 7308 49252 7364 49868
rect 7532 49858 7588 49868
rect 6860 48190 6862 48242
rect 6914 48190 6916 48242
rect 6860 48178 6916 48190
rect 6972 49196 7364 49252
rect 6972 48466 7028 49196
rect 7420 48804 7476 48814
rect 6972 48414 6974 48466
rect 7026 48414 7028 48466
rect 6860 48020 6916 48030
rect 6748 47964 6860 48020
rect 6860 47954 6916 47964
rect 6412 46834 6468 46844
rect 5404 46274 5460 46284
rect 6972 46116 7028 48414
rect 7084 48468 7140 48478
rect 7084 48374 7140 48412
rect 7196 48356 7252 48366
rect 7196 48262 7252 48300
rect 7420 48242 7476 48748
rect 7644 48580 7700 49868
rect 7756 49812 7812 50316
rect 7868 50034 7924 50428
rect 8204 50372 8260 50652
rect 7868 49982 7870 50034
rect 7922 49982 7924 50034
rect 7868 49970 7924 49982
rect 7980 50316 8260 50372
rect 8316 50372 8372 52892
rect 8652 50428 8708 53116
rect 7980 50036 8036 50316
rect 8316 50306 8372 50316
rect 8540 50372 8708 50428
rect 8764 52946 8820 52958
rect 8764 52894 8766 52946
rect 8818 52894 8820 52946
rect 8764 50484 8820 52894
rect 8764 50418 8820 50428
rect 9436 50484 9492 50522
rect 9436 50418 9492 50428
rect 9548 50428 9604 54460
rect 9660 54450 9716 54460
rect 9660 53730 9716 53742
rect 9660 53678 9662 53730
rect 9714 53678 9716 53730
rect 9660 52948 9716 53678
rect 9996 53508 10052 56028
rect 10108 55990 10164 56028
rect 10220 53730 10276 56252
rect 10444 56196 10500 56700
rect 10668 56644 10724 56654
rect 10332 56140 10500 56196
rect 10556 56642 10724 56644
rect 10556 56590 10670 56642
rect 10722 56590 10724 56642
rect 10556 56588 10724 56590
rect 10332 56082 10388 56140
rect 10332 56030 10334 56082
rect 10386 56030 10388 56082
rect 10332 55524 10388 56030
rect 10556 56082 10612 56588
rect 10668 56578 10724 56588
rect 10780 56420 10836 56702
rect 10780 56354 10836 56364
rect 10556 56030 10558 56082
rect 10610 56030 10612 56082
rect 10556 56018 10612 56030
rect 10892 56084 10948 57596
rect 11004 57650 11060 57662
rect 11004 57598 11006 57650
rect 11058 57598 11060 57650
rect 11004 56866 11060 57598
rect 11004 56814 11006 56866
rect 11058 56814 11060 56866
rect 11004 56802 11060 56814
rect 11228 56980 11284 58604
rect 11340 57652 11396 57662
rect 11396 57596 11732 57652
rect 11340 57586 11396 57596
rect 11676 57090 11732 57596
rect 11676 57038 11678 57090
rect 11730 57038 11732 57090
rect 11676 57026 11732 57038
rect 11788 56980 11844 56990
rect 12124 56980 12180 58604
rect 13020 58548 13076 58558
rect 12236 58434 12292 58446
rect 12236 58382 12238 58434
rect 12290 58382 12292 58434
rect 12236 58212 12292 58382
rect 12684 58212 12740 58222
rect 12236 58210 12852 58212
rect 12236 58158 12686 58210
rect 12738 58158 12852 58210
rect 12236 58156 12852 58158
rect 12684 58146 12740 58156
rect 11228 56924 11620 56980
rect 11228 56754 11284 56924
rect 11228 56702 11230 56754
rect 11282 56702 11284 56754
rect 11228 56690 11284 56702
rect 11340 56754 11396 56766
rect 11340 56702 11342 56754
rect 11394 56702 11396 56754
rect 11340 56308 11396 56702
rect 10892 56018 10948 56028
rect 11004 56252 11396 56308
rect 11564 56306 11620 56924
rect 11788 56978 12180 56980
rect 11788 56926 11790 56978
rect 11842 56926 12180 56978
rect 11788 56924 12180 56926
rect 12236 57876 12292 57886
rect 11788 56914 11844 56924
rect 11564 56254 11566 56306
rect 11618 56254 11620 56306
rect 10444 55970 10500 55982
rect 10444 55918 10446 55970
rect 10498 55918 10500 55970
rect 10444 55636 10500 55918
rect 10444 55580 10724 55636
rect 10332 55468 10612 55524
rect 10332 54402 10388 54414
rect 10332 54350 10334 54402
rect 10386 54350 10388 54402
rect 10332 53844 10388 54350
rect 10444 53844 10500 53854
rect 10332 53842 10500 53844
rect 10332 53790 10446 53842
rect 10498 53790 10500 53842
rect 10332 53788 10500 53790
rect 10444 53778 10500 53788
rect 10220 53678 10222 53730
rect 10274 53678 10276 53730
rect 10220 53666 10276 53678
rect 10556 53732 10612 55468
rect 10668 55188 10724 55580
rect 10668 55122 10724 55132
rect 11004 54292 11060 56252
rect 11564 56242 11620 56254
rect 11340 56082 11396 56094
rect 11340 56030 11342 56082
rect 11394 56030 11396 56082
rect 11340 55748 11396 56030
rect 12236 56082 12292 57820
rect 12796 57652 12852 58156
rect 12796 57558 12852 57596
rect 13020 56194 13076 58492
rect 13804 58436 13860 58446
rect 13468 57876 13524 57886
rect 13468 57762 13524 57820
rect 13468 57710 13470 57762
rect 13522 57710 13524 57762
rect 13468 57698 13524 57710
rect 13804 57090 13860 58380
rect 13804 57038 13806 57090
rect 13858 57038 13860 57090
rect 13804 57026 13860 57038
rect 13916 58212 13972 60732
rect 14028 59220 14084 59230
rect 14252 59220 14308 61518
rect 14588 62132 14756 62188
rect 14812 62578 15876 62580
rect 14812 62526 15822 62578
rect 15874 62526 15876 62578
rect 14812 62524 15876 62526
rect 14028 59218 14308 59220
rect 14028 59166 14030 59218
rect 14082 59166 14308 59218
rect 14028 59164 14308 59166
rect 14476 61348 14532 61358
rect 14476 61010 14532 61292
rect 14476 60958 14478 61010
rect 14530 60958 14532 61010
rect 14028 59154 14084 59164
rect 14028 58212 14084 58222
rect 13916 58210 14084 58212
rect 13916 58158 14030 58210
rect 14082 58158 14084 58210
rect 13916 58156 14084 58158
rect 13916 56868 13972 58156
rect 14028 58146 14084 58156
rect 14364 58212 14420 58222
rect 14364 58118 14420 58156
rect 14476 56980 14532 60958
rect 14252 56924 14532 56980
rect 14252 56868 14308 56924
rect 13804 56812 13972 56868
rect 14028 56866 14308 56868
rect 14028 56814 14254 56866
rect 14306 56814 14308 56866
rect 14028 56812 14308 56814
rect 13692 56756 13748 56766
rect 13692 56662 13748 56700
rect 13020 56142 13022 56194
rect 13074 56142 13076 56194
rect 13020 56130 13076 56142
rect 12236 56030 12238 56082
rect 12290 56030 12292 56082
rect 11340 55692 11620 55748
rect 11452 55188 11508 55198
rect 11452 55094 11508 55132
rect 11228 54292 11284 54302
rect 11004 54236 11228 54292
rect 10556 53638 10612 53676
rect 10780 53732 10836 53742
rect 11116 53732 11172 53742
rect 10780 53730 11172 53732
rect 10780 53678 10782 53730
rect 10834 53678 11118 53730
rect 11170 53678 11172 53730
rect 10780 53676 11172 53678
rect 10780 53666 10836 53676
rect 11116 53666 11172 53676
rect 11228 53730 11284 54236
rect 11228 53678 11230 53730
rect 11282 53678 11284 53730
rect 11228 53666 11284 53678
rect 10332 53508 10388 53518
rect 9996 53506 10388 53508
rect 9996 53454 10334 53506
rect 10386 53454 10388 53506
rect 9996 53452 10388 53454
rect 9996 53170 10052 53452
rect 10332 53442 10388 53452
rect 9996 53118 9998 53170
rect 10050 53118 10052 53170
rect 9996 53106 10052 53118
rect 11564 53172 11620 55692
rect 12236 55298 12292 56030
rect 13468 55412 13524 55422
rect 13468 55318 13524 55356
rect 12236 55246 12238 55298
rect 12290 55246 12292 55298
rect 12236 55234 12292 55246
rect 12460 54402 12516 54414
rect 12460 54350 12462 54402
rect 12514 54350 12516 54402
rect 12460 54292 12516 54350
rect 12460 54226 12516 54236
rect 11676 53172 11732 53182
rect 11564 53116 11676 53172
rect 11676 53078 11732 53116
rect 12684 53060 12740 53070
rect 9660 52882 9716 52892
rect 9772 52948 9828 52958
rect 11116 52948 11172 52958
rect 9772 52946 9940 52948
rect 9772 52894 9774 52946
rect 9826 52894 9940 52946
rect 9772 52892 9940 52894
rect 9772 52882 9828 52892
rect 9884 51490 9940 52892
rect 11116 52050 11172 52892
rect 12012 52948 12068 52958
rect 12012 52854 12068 52892
rect 11900 52388 11956 52398
rect 11788 52386 11956 52388
rect 11788 52334 11902 52386
rect 11954 52334 11956 52386
rect 11788 52332 11956 52334
rect 11452 52164 11508 52174
rect 11452 52070 11508 52108
rect 11116 51998 11118 52050
rect 11170 51998 11172 52050
rect 11116 51986 11172 51998
rect 9884 51438 9886 51490
rect 9938 51438 9940 51490
rect 9772 50596 9828 50606
rect 9772 50482 9828 50540
rect 9772 50430 9774 50482
rect 9826 50430 9828 50482
rect 9548 50372 9716 50428
rect 9772 50418 9828 50430
rect 9884 50484 9940 51438
rect 11788 51492 11844 52332
rect 11900 52322 11956 52332
rect 12572 52164 12628 52174
rect 12572 52070 12628 52108
rect 12012 52052 12068 52062
rect 12012 52050 12180 52052
rect 12012 51998 12014 52050
rect 12066 51998 12180 52050
rect 12012 51996 12180 51998
rect 12012 51986 12068 51996
rect 11788 51426 11844 51436
rect 11900 51938 11956 51950
rect 11900 51886 11902 51938
rect 11954 51886 11956 51938
rect 10108 51378 10164 51390
rect 10108 51326 10110 51378
rect 10162 51326 10164 51378
rect 10108 50820 10164 51326
rect 10108 50754 10164 50764
rect 11788 51266 11844 51278
rect 11788 51214 11790 51266
rect 11842 51214 11844 51266
rect 10892 50708 10948 50718
rect 10220 50706 10948 50708
rect 10220 50654 10894 50706
rect 10946 50654 10948 50706
rect 10220 50652 10948 50654
rect 10108 50482 10164 50494
rect 10108 50430 10110 50482
rect 10162 50430 10164 50482
rect 10108 50428 10164 50430
rect 9884 50418 9940 50428
rect 8204 50036 8260 50046
rect 7980 50034 8260 50036
rect 7980 49982 8206 50034
rect 8258 49982 8260 50034
rect 7980 49980 8260 49982
rect 8204 49970 8260 49980
rect 8316 50036 8372 50046
rect 8372 49980 8484 50036
rect 8316 49970 8372 49980
rect 7756 49756 8148 49812
rect 7644 48524 8036 48580
rect 7756 48356 7812 48366
rect 7812 48300 7924 48356
rect 7756 48262 7812 48300
rect 7420 48190 7422 48242
rect 7474 48190 7476 48242
rect 7420 48178 7476 48190
rect 7420 48020 7476 48030
rect 7420 46562 7476 47964
rect 7756 46900 7812 46910
rect 7756 46674 7812 46844
rect 7756 46622 7758 46674
rect 7810 46622 7812 46674
rect 7756 46610 7812 46622
rect 7868 46676 7924 48300
rect 7980 47236 8036 48524
rect 8092 48466 8148 49756
rect 8428 49140 8484 49980
rect 8540 49812 8596 50372
rect 9660 49812 9716 50372
rect 9996 50372 10164 50428
rect 9996 50306 10052 50316
rect 8540 49810 8820 49812
rect 8540 49758 8542 49810
rect 8594 49758 8820 49810
rect 8540 49756 8820 49758
rect 8540 49746 8596 49756
rect 8540 49140 8596 49150
rect 8428 49084 8540 49140
rect 8540 49046 8596 49084
rect 8092 48414 8094 48466
rect 8146 48414 8148 48466
rect 8092 48402 8148 48414
rect 8428 48916 8484 48926
rect 7980 47180 8260 47236
rect 8204 46898 8260 47180
rect 8204 46846 8206 46898
rect 8258 46846 8260 46898
rect 8204 46834 8260 46846
rect 8428 46900 8484 48860
rect 8652 48356 8708 48366
rect 8652 48262 8708 48300
rect 8764 48244 8820 49756
rect 9548 49756 9660 49812
rect 8988 49140 9044 49150
rect 8988 49046 9044 49084
rect 9548 49026 9604 49756
rect 9660 49718 9716 49756
rect 10220 49138 10276 50652
rect 10892 50642 10948 50652
rect 11228 50596 11284 50606
rect 10444 50484 10500 50494
rect 10892 50484 10948 50522
rect 10444 50482 10612 50484
rect 10444 50430 10446 50482
rect 10498 50430 10612 50482
rect 10444 50428 10612 50430
rect 10444 50418 10500 50428
rect 10556 50260 10612 50428
rect 10892 50418 10948 50428
rect 11004 50482 11060 50494
rect 11004 50430 11006 50482
rect 11058 50430 11060 50482
rect 11004 50260 11060 50430
rect 10556 50204 11060 50260
rect 11228 50482 11284 50540
rect 11228 50430 11230 50482
rect 11282 50430 11284 50482
rect 10332 49700 10388 49710
rect 10332 49606 10388 49644
rect 10220 49086 10222 49138
rect 10274 49086 10276 49138
rect 10220 49074 10276 49086
rect 9548 48974 9550 49026
rect 9602 48974 9604 49026
rect 9548 48962 9604 48974
rect 10556 48916 10612 50204
rect 8876 48804 8932 48814
rect 8876 48710 8932 48748
rect 8988 48356 9044 48366
rect 10108 48356 10164 48366
rect 9044 48300 9156 48356
rect 8988 48290 9044 48300
rect 8876 48244 8932 48254
rect 8764 48242 8932 48244
rect 8764 48190 8878 48242
rect 8930 48190 8932 48242
rect 8764 48188 8932 48190
rect 8876 48178 8932 48188
rect 8428 46834 8484 46844
rect 7980 46676 8036 46686
rect 7868 46674 8036 46676
rect 7868 46622 7982 46674
rect 8034 46622 8036 46674
rect 7868 46620 8036 46622
rect 7420 46510 7422 46562
rect 7474 46510 7476 46562
rect 7420 46498 7476 46510
rect 7980 46228 8036 46620
rect 8428 46676 8484 46686
rect 8428 46674 9044 46676
rect 8428 46622 8430 46674
rect 8482 46622 9044 46674
rect 8428 46620 9044 46622
rect 8428 46610 8484 46620
rect 8092 46564 8148 46574
rect 8092 46470 8148 46508
rect 7980 46162 8036 46172
rect 6748 46060 7028 46116
rect 8988 46114 9044 46620
rect 8988 46062 8990 46114
rect 9042 46062 9044 46114
rect 6412 46004 6468 46014
rect 5964 46002 6468 46004
rect 5964 45950 6414 46002
rect 6466 45950 6468 46002
rect 5964 45948 6468 45950
rect 5964 45218 6020 45948
rect 6412 45938 6468 45948
rect 6748 45890 6804 46060
rect 6748 45838 6750 45890
rect 6802 45838 6804 45890
rect 6748 45826 6804 45838
rect 6524 45780 6580 45790
rect 6524 45686 6580 45724
rect 5964 45166 5966 45218
rect 6018 45166 6020 45218
rect 5964 45154 6020 45166
rect 6412 45666 6468 45678
rect 6412 45614 6414 45666
rect 6466 45614 6468 45666
rect 5180 45106 5796 45108
rect 5180 45054 5182 45106
rect 5234 45054 5796 45106
rect 5180 45052 5796 45054
rect 5180 45042 5236 45052
rect 5180 44660 5236 44670
rect 5068 44604 5180 44660
rect 5180 44594 5236 44604
rect 5740 44322 5796 45052
rect 5740 44270 5742 44322
rect 5794 44270 5796 44322
rect 5740 44258 5796 44270
rect 6412 43764 6468 45614
rect 6636 45668 6692 45678
rect 6524 44436 6580 44446
rect 6636 44436 6692 45612
rect 6860 45556 6916 46060
rect 8988 46050 9044 46062
rect 6972 45948 8148 46004
rect 6972 45890 7028 45948
rect 6972 45838 6974 45890
rect 7026 45838 7028 45890
rect 6972 45826 7028 45838
rect 8092 45892 8148 45948
rect 8204 45892 8260 45902
rect 8092 45890 8260 45892
rect 8092 45838 8206 45890
rect 8258 45838 8260 45890
rect 8092 45836 8260 45838
rect 8204 45826 8260 45836
rect 7532 45780 7588 45790
rect 7532 45686 7588 45724
rect 7980 45778 8036 45790
rect 7980 45726 7982 45778
rect 8034 45726 8036 45778
rect 6860 45490 6916 45500
rect 7420 45666 7476 45678
rect 7420 45614 7422 45666
rect 7474 45614 7476 45666
rect 6524 44434 6692 44436
rect 6524 44382 6526 44434
rect 6578 44382 6692 44434
rect 6524 44380 6692 44382
rect 6524 44370 6580 44380
rect 7420 44212 7476 45614
rect 7644 45668 7700 45678
rect 7644 45574 7700 45612
rect 7756 45666 7812 45678
rect 7756 45614 7758 45666
rect 7810 45614 7812 45666
rect 7756 45556 7812 45614
rect 7756 45490 7812 45500
rect 7980 45332 8036 45726
rect 8428 45780 8484 45790
rect 8428 45686 8484 45724
rect 8540 45778 8596 45790
rect 8540 45726 8542 45778
rect 8594 45726 8596 45778
rect 7980 45266 8036 45276
rect 8092 45556 8148 45566
rect 8092 44996 8148 45500
rect 7420 44146 7476 44156
rect 7756 44994 8148 44996
rect 7756 44942 8094 44994
rect 8146 44942 8148 44994
rect 7756 44940 8148 44942
rect 6412 43698 6468 43708
rect 6636 44100 6692 44110
rect 4284 43538 4340 43550
rect 4284 43486 4286 43538
rect 4338 43486 4340 43538
rect 4284 43428 4340 43486
rect 4844 43428 4900 43438
rect 4284 43426 4900 43428
rect 4284 43374 4846 43426
rect 4898 43374 4900 43426
rect 4284 43372 4900 43374
rect 4476 43148 4740 43158
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4476 43082 4740 43092
rect 4844 42980 4900 43372
rect 4844 42914 4900 42924
rect 6636 41860 6692 44044
rect 7644 43764 7700 43774
rect 7644 43650 7700 43708
rect 7644 43598 7646 43650
rect 7698 43598 7700 43650
rect 7644 43586 7700 43598
rect 7756 43650 7812 44940
rect 8092 44930 8148 44940
rect 8540 44436 8596 45726
rect 8764 45780 8820 45790
rect 8652 45332 8708 45342
rect 8764 45332 8820 45724
rect 8876 45778 8932 45790
rect 8876 45726 8878 45778
rect 8930 45726 8932 45778
rect 8876 45556 8932 45726
rect 8988 45780 9044 45790
rect 9100 45780 9156 48300
rect 10108 48262 10164 48300
rect 9884 48244 9940 48254
rect 9884 48242 10052 48244
rect 9884 48190 9886 48242
rect 9938 48190 10052 48242
rect 9884 48188 10052 48190
rect 9884 48178 9940 48188
rect 9548 46562 9604 46574
rect 9548 46510 9550 46562
rect 9602 46510 9604 46562
rect 9548 46452 9604 46510
rect 9548 46386 9604 46396
rect 9996 45892 10052 48188
rect 10220 48242 10276 48254
rect 10220 48190 10222 48242
rect 10274 48190 10276 48242
rect 10108 48132 10164 48142
rect 10108 47458 10164 48076
rect 10108 47406 10110 47458
rect 10162 47406 10164 47458
rect 10108 46228 10164 47406
rect 10220 46452 10276 48190
rect 10556 47236 10612 48860
rect 10220 46386 10276 46396
rect 10332 47012 10388 47022
rect 10108 46172 10276 46228
rect 10108 45892 10164 45902
rect 9996 45890 10164 45892
rect 9996 45838 10110 45890
rect 10162 45838 10164 45890
rect 9996 45836 10164 45838
rect 10108 45826 10164 45836
rect 9044 45724 9156 45780
rect 9548 45780 9604 45790
rect 8988 45686 9044 45724
rect 8876 45490 8932 45500
rect 8876 45332 8932 45342
rect 8764 45330 8932 45332
rect 8764 45278 8878 45330
rect 8930 45278 8932 45330
rect 8764 45276 8932 45278
rect 8652 45238 8708 45276
rect 8876 45266 8932 45276
rect 8988 45220 9044 45230
rect 9548 45220 9604 45724
rect 8988 45218 9604 45220
rect 8988 45166 8990 45218
rect 9042 45166 9604 45218
rect 8988 45164 9604 45166
rect 8988 45154 9044 45164
rect 9548 44994 9604 45164
rect 9548 44942 9550 44994
rect 9602 44942 9604 44994
rect 9548 44930 9604 44942
rect 9772 45220 9828 45230
rect 9660 44884 9716 44894
rect 8652 44436 8708 44446
rect 9100 44436 9156 44446
rect 8540 44434 9156 44436
rect 8540 44382 8654 44434
rect 8706 44382 9102 44434
rect 9154 44382 9156 44434
rect 8540 44380 9156 44382
rect 8652 44370 8708 44380
rect 9100 44370 9156 44380
rect 8988 44212 9044 44222
rect 8988 44118 9044 44156
rect 7756 43598 7758 43650
rect 7810 43598 7812 43650
rect 7756 43586 7812 43598
rect 9548 43876 9604 43886
rect 9324 42868 9380 42878
rect 9324 42774 9380 42812
rect 6636 41794 6692 41804
rect 4476 41580 4740 41590
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4476 41514 4740 41524
rect 4172 40562 4228 40572
rect 9436 40628 9492 40638
rect 3164 40338 3220 40348
rect 9436 40404 9492 40572
rect 9436 40338 9492 40348
rect 4476 40012 4740 40022
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4476 39946 4740 39956
rect 5852 39956 5908 39966
rect 2940 39666 2996 39676
rect 4284 39844 4340 39854
rect 1708 39506 1764 39518
rect 1708 39454 1710 39506
rect 1762 39454 1764 39506
rect 1708 39060 1764 39454
rect 2044 39508 2100 39518
rect 2044 39414 2100 39452
rect 1708 38994 1764 39004
rect 2492 39394 2548 39406
rect 2492 39342 2494 39394
rect 2546 39342 2548 39394
rect 2492 39060 2548 39342
rect 2492 38994 2548 39004
rect 4284 38834 4340 39788
rect 4284 38782 4286 38834
rect 4338 38782 4340 38834
rect 4284 38770 4340 38782
rect 1932 38612 1988 38622
rect 1932 38518 1988 38556
rect 4476 38444 4740 38454
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4476 38378 4740 38388
rect 1708 37938 1764 37950
rect 1708 37886 1710 37938
rect 1762 37886 1764 37938
rect 1708 37716 1764 37886
rect 2044 37828 2100 37838
rect 2044 37734 2100 37772
rect 2492 37826 2548 37838
rect 2492 37774 2494 37826
rect 2546 37774 2548 37826
rect 1708 37650 1764 37660
rect 2492 37716 2548 37774
rect 2492 37650 2548 37660
rect 2716 37716 2772 37726
rect 2044 37380 2100 37390
rect 2044 37378 2212 37380
rect 2044 37326 2046 37378
rect 2098 37326 2212 37378
rect 2044 37324 2212 37326
rect 2044 37314 2100 37324
rect 1708 37266 1764 37278
rect 1708 37214 1710 37266
rect 1762 37214 1764 37266
rect 1708 37044 1764 37214
rect 1708 36978 1764 36988
rect 1932 36596 1988 36606
rect 1932 36502 1988 36540
rect 2044 35812 2100 35822
rect 2044 35718 2100 35756
rect 1708 35700 1764 35710
rect 1708 35606 1764 35644
rect 2156 35588 2212 37324
rect 2492 37154 2548 37166
rect 2492 37102 2494 37154
rect 2546 37102 2548 37154
rect 2492 37044 2548 37102
rect 2492 36978 2548 36988
rect 2716 35922 2772 37660
rect 4844 36932 4900 36942
rect 4476 36876 4740 36886
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4476 36810 4740 36820
rect 4844 36594 4900 36876
rect 4844 36542 4846 36594
rect 4898 36542 4900 36594
rect 4172 36484 4228 36494
rect 4172 36390 4228 36428
rect 4844 36484 4900 36542
rect 4844 36418 4900 36428
rect 2716 35870 2718 35922
rect 2770 35870 2772 35922
rect 2716 35858 2772 35870
rect 2156 35522 2212 35532
rect 2380 35698 2436 35710
rect 2380 35646 2382 35698
rect 2434 35646 2436 35698
rect 2380 35028 2436 35646
rect 2380 34962 2436 34972
rect 2492 35700 2548 35710
rect 2492 35026 2548 35644
rect 2492 34974 2494 35026
rect 2546 34974 2548 35026
rect 2492 34962 2548 34974
rect 3164 35586 3220 35598
rect 3164 35534 3166 35586
rect 3218 35534 3220 35586
rect 3164 35028 3220 35534
rect 4476 35308 4740 35318
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4476 35242 4740 35252
rect 3164 34962 3220 34972
rect 1708 34802 1764 34814
rect 1708 34750 1710 34802
rect 1762 34750 1764 34802
rect 1708 34356 1764 34750
rect 2044 34692 2100 34702
rect 2044 34598 2100 34636
rect 2940 34690 2996 34702
rect 2940 34638 2942 34690
rect 2994 34638 2996 34690
rect 1708 34290 1764 34300
rect 2940 34356 2996 34638
rect 2940 34290 2996 34300
rect 4284 34130 4340 34142
rect 4284 34078 4286 34130
rect 4338 34078 4340 34130
rect 4284 34020 4340 34078
rect 4284 33954 4340 33964
rect 4732 34020 4788 34030
rect 4732 33926 4788 33964
rect 1932 33908 1988 33918
rect 1932 33814 1988 33852
rect 4476 33740 4740 33750
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4476 33674 4740 33684
rect 1708 33234 1764 33246
rect 1708 33182 1710 33234
rect 1762 33182 1764 33234
rect 1708 33012 1764 33182
rect 2044 33124 2100 33134
rect 2044 33030 2100 33068
rect 2492 33122 2548 33134
rect 2492 33070 2494 33122
rect 2546 33070 2548 33122
rect 1708 32946 1764 32956
rect 2492 33012 2548 33070
rect 2492 32946 2548 32956
rect 5068 33012 5124 33022
rect 2044 32674 2100 32686
rect 2044 32622 2046 32674
rect 2098 32622 2100 32674
rect 1708 32562 1764 32574
rect 1708 32510 1710 32562
rect 1762 32510 1764 32562
rect 1708 32340 1764 32510
rect 1708 32274 1764 32284
rect 1932 31892 1988 31902
rect 1932 31798 1988 31836
rect 2044 31556 2100 32622
rect 2492 32450 2548 32462
rect 2492 32398 2494 32450
rect 2546 32398 2548 32450
rect 2492 32340 2548 32398
rect 2492 32274 2548 32284
rect 4476 32172 4740 32182
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4476 32106 4740 32116
rect 4844 31892 4900 31902
rect 5068 31892 5124 32956
rect 4844 31890 5124 31892
rect 4844 31838 4846 31890
rect 4898 31838 5124 31890
rect 4844 31836 5124 31838
rect 4172 31780 4228 31790
rect 4172 31686 4228 31724
rect 4844 31780 4900 31836
rect 4844 31714 4900 31724
rect 2044 31490 2100 31500
rect 2044 31220 2100 31230
rect 2044 31126 2100 31164
rect 5852 31220 5908 39900
rect 6748 39620 6804 39630
rect 6748 37716 6804 39564
rect 6748 37650 6804 37660
rect 8428 38052 8484 38062
rect 8428 36482 8484 37996
rect 9100 38052 9156 38062
rect 9100 37958 9156 37996
rect 9212 37044 9268 37054
rect 9212 36594 9268 36988
rect 9212 36542 9214 36594
rect 9266 36542 9268 36594
rect 9212 36530 9268 36542
rect 8428 36430 8430 36482
rect 8482 36430 8484 36482
rect 8428 34914 8484 36430
rect 9100 35476 9156 35486
rect 9100 35026 9156 35420
rect 9100 34974 9102 35026
rect 9154 34974 9156 35026
rect 9100 34962 9156 34974
rect 8428 34862 8430 34914
rect 8482 34862 8484 34914
rect 8428 34850 8484 34862
rect 8204 33346 8260 33358
rect 8204 33294 8206 33346
rect 8258 33294 8260 33346
rect 5852 31154 5908 31164
rect 7980 31780 8036 31790
rect 8204 31780 8260 33294
rect 8988 33236 9044 33246
rect 8988 33234 9492 33236
rect 8988 33182 8990 33234
rect 9042 33182 9492 33234
rect 8988 33180 9492 33182
rect 8988 33170 9044 33180
rect 9436 32786 9492 33180
rect 9436 32734 9438 32786
rect 9490 32734 9492 32786
rect 9436 32722 9492 32734
rect 8988 32450 9044 32462
rect 8988 32398 8990 32450
rect 9042 32398 9044 32450
rect 8876 32340 8932 32350
rect 8652 32338 8932 32340
rect 8652 32286 8878 32338
rect 8930 32286 8932 32338
rect 8652 32284 8932 32286
rect 8652 31890 8708 32284
rect 8876 32274 8932 32284
rect 8652 31838 8654 31890
rect 8706 31838 8708 31890
rect 8652 31826 8708 31838
rect 7980 31778 8260 31780
rect 7980 31726 7982 31778
rect 8034 31726 8260 31778
rect 7980 31724 8260 31726
rect 2716 31106 2772 31118
rect 2716 31054 2718 31106
rect 2770 31054 2772 31106
rect 1708 30996 1764 31006
rect 1708 30902 1764 30940
rect 2380 30994 2436 31006
rect 2380 30942 2382 30994
rect 2434 30942 2436 30994
rect 2380 30884 2436 30942
rect 2044 30548 2100 30558
rect 1708 30098 1764 30110
rect 1708 30046 1710 30098
rect 1762 30046 1764 30098
rect 1708 29652 1764 30046
rect 2044 30098 2100 30492
rect 2380 30324 2436 30828
rect 2380 30258 2436 30268
rect 2492 30996 2548 31006
rect 2492 30322 2548 30940
rect 2716 30436 2772 31054
rect 3164 30884 3220 30894
rect 3164 30790 3220 30828
rect 4476 30604 4740 30614
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4476 30538 4740 30548
rect 2716 30370 2772 30380
rect 2492 30270 2494 30322
rect 2546 30270 2548 30322
rect 2492 30258 2548 30270
rect 7980 30212 8036 31724
rect 8988 30772 9044 32398
rect 9548 31220 9604 43820
rect 9660 42978 9716 44828
rect 9772 43204 9828 45164
rect 10220 44324 10276 46172
rect 10332 45890 10388 46956
rect 10332 45838 10334 45890
rect 10386 45838 10388 45890
rect 10332 45826 10388 45838
rect 10444 46340 10500 46350
rect 10444 45668 10500 46284
rect 10556 45890 10612 47180
rect 10892 49252 10948 49262
rect 10668 46004 10724 46014
rect 10668 45910 10724 45948
rect 10556 45838 10558 45890
rect 10610 45838 10612 45890
rect 10556 45826 10612 45838
rect 10780 45892 10836 45902
rect 10780 45798 10836 45836
rect 10444 45612 10836 45668
rect 10220 44258 10276 44268
rect 9772 43138 9828 43148
rect 9884 43652 9940 43662
rect 9660 42926 9662 42978
rect 9714 42926 9716 42978
rect 9660 42914 9716 42926
rect 9884 42978 9940 43596
rect 10444 43428 10500 43438
rect 10444 43334 10500 43372
rect 10332 43316 10388 43326
rect 9884 42926 9886 42978
rect 9938 42926 9940 42978
rect 9884 42914 9940 42926
rect 10108 43314 10388 43316
rect 10108 43262 10334 43314
rect 10386 43262 10388 43314
rect 10108 43260 10388 43262
rect 10108 42978 10164 43260
rect 10332 43250 10388 43260
rect 10108 42926 10110 42978
rect 10162 42926 10164 42978
rect 10108 42914 10164 42926
rect 10220 42868 10276 42878
rect 10220 42774 10276 42812
rect 10668 42754 10724 42766
rect 10668 42702 10670 42754
rect 10722 42702 10724 42754
rect 10220 42532 10276 42542
rect 10220 42438 10276 42476
rect 9996 42196 10052 42206
rect 9884 42082 9940 42094
rect 9884 42030 9886 42082
rect 9938 42030 9940 42082
rect 9772 41970 9828 41982
rect 9772 41918 9774 41970
rect 9826 41918 9828 41970
rect 9772 41076 9828 41918
rect 9884 41972 9940 42030
rect 9884 41906 9940 41916
rect 9884 41748 9940 41758
rect 9884 41654 9940 41692
rect 9772 41010 9828 41020
rect 9772 38724 9828 38734
rect 9772 38162 9828 38668
rect 9772 38110 9774 38162
rect 9826 38110 9828 38162
rect 9772 38098 9828 38110
rect 9660 32788 9716 32798
rect 9884 32788 9940 32798
rect 9660 32786 9940 32788
rect 9660 32734 9662 32786
rect 9714 32734 9886 32786
rect 9938 32734 9940 32786
rect 9660 32732 9940 32734
rect 9660 32722 9716 32732
rect 9884 32722 9940 32732
rect 9996 32676 10052 42140
rect 10444 42084 10500 42094
rect 10332 41970 10388 41982
rect 10332 41918 10334 41970
rect 10386 41918 10388 41970
rect 10108 41412 10164 41422
rect 10332 41412 10388 41918
rect 10164 41356 10388 41412
rect 10444 41412 10500 42028
rect 10556 41860 10612 41870
rect 10556 41766 10612 41804
rect 10108 41298 10164 41356
rect 10444 41346 10500 41356
rect 10108 41246 10110 41298
rect 10162 41246 10164 41298
rect 10108 41234 10164 41246
rect 10556 41186 10612 41198
rect 10556 41134 10558 41186
rect 10610 41134 10612 41186
rect 10444 39620 10500 39630
rect 10444 39526 10500 39564
rect 10556 39508 10612 41134
rect 10668 40962 10724 42702
rect 10780 41970 10836 45612
rect 10892 45444 10948 49196
rect 11228 49028 11284 50430
rect 11452 50482 11508 50494
rect 11452 50430 11454 50482
rect 11506 50430 11508 50482
rect 11452 49252 11508 50430
rect 11788 49812 11844 51214
rect 11900 50428 11956 51886
rect 12124 50428 12180 51996
rect 12684 51940 12740 53004
rect 13580 53060 13636 53070
rect 13804 53060 13860 56812
rect 13636 53004 13860 53060
rect 13916 53058 13972 53070
rect 13916 53006 13918 53058
rect 13970 53006 13972 53058
rect 13580 52966 13636 53004
rect 13916 52836 13972 53006
rect 13916 52770 13972 52780
rect 13804 52724 13860 52734
rect 13580 52668 13804 52724
rect 13020 52164 13076 52174
rect 13020 52070 13076 52108
rect 12572 51884 12740 51940
rect 12236 50820 12292 50830
rect 12236 50594 12292 50764
rect 12572 50708 12628 51884
rect 12460 50652 12628 50708
rect 12236 50542 12238 50594
rect 12290 50542 12292 50594
rect 12236 50530 12292 50542
rect 12348 50596 12404 50606
rect 12348 50428 12404 50540
rect 11900 50372 12068 50428
rect 12124 50372 12404 50428
rect 12460 50482 12516 50652
rect 12908 50596 12964 50606
rect 12460 50430 12462 50482
rect 12514 50430 12516 50482
rect 12460 50418 12516 50430
rect 12796 50484 12852 50522
rect 12908 50502 12964 50540
rect 13132 50596 13188 50606
rect 12796 50418 12852 50428
rect 11788 49746 11844 49756
rect 11452 49186 11508 49196
rect 11116 48132 11172 48142
rect 11116 48038 11172 48076
rect 11228 47012 11284 48972
rect 11676 48804 11732 48814
rect 11676 48466 11732 48748
rect 12012 48804 12068 50316
rect 12348 49138 12404 50372
rect 13132 50372 13188 50540
rect 13468 50484 13524 50522
rect 13468 50418 13524 50428
rect 13132 50306 13188 50316
rect 13580 49922 13636 52668
rect 13804 52658 13860 52668
rect 13692 52164 13748 52174
rect 13692 50594 13748 52108
rect 13692 50542 13694 50594
rect 13746 50542 13748 50594
rect 13692 50428 13748 50542
rect 13916 52164 13972 52174
rect 14028 52164 14084 56812
rect 14252 56802 14308 56812
rect 14476 56644 14532 56654
rect 14476 56550 14532 56588
rect 14588 56308 14644 62132
rect 14812 61010 14868 62524
rect 15820 62514 15876 62524
rect 16044 62580 16100 62590
rect 16156 62580 16212 64094
rect 16268 64148 16324 64158
rect 16268 64054 16324 64092
rect 16380 64146 16436 64428
rect 16604 64260 16660 64270
rect 16660 64204 16772 64260
rect 16604 64194 16660 64204
rect 16380 64094 16382 64146
rect 16434 64094 16436 64146
rect 16380 64082 16436 64094
rect 16604 63924 16660 63934
rect 16604 63830 16660 63868
rect 16716 63252 16772 64204
rect 17388 63924 17444 63934
rect 17388 63830 17444 63868
rect 17500 63810 17556 64766
rect 17612 64372 17668 65438
rect 17724 65492 17780 65502
rect 17724 65398 17780 65436
rect 17836 65490 17892 65502
rect 17836 65438 17838 65490
rect 17890 65438 17892 65490
rect 17836 64932 17892 65438
rect 18060 65492 18116 65502
rect 18396 65492 18452 65502
rect 18060 65490 18452 65492
rect 18060 65438 18062 65490
rect 18114 65438 18398 65490
rect 18450 65438 18452 65490
rect 18060 65436 18452 65438
rect 18060 65426 18116 65436
rect 18396 65426 18452 65436
rect 19964 65490 20020 65502
rect 19964 65438 19966 65490
rect 20018 65438 20020 65490
rect 17836 64866 17892 64876
rect 17948 64820 18004 64830
rect 17948 64708 18004 64764
rect 19964 64820 20020 65438
rect 19964 64754 20020 64764
rect 17612 64306 17668 64316
rect 17724 64706 18004 64708
rect 17724 64654 17950 64706
rect 18002 64654 18004 64706
rect 17724 64652 18004 64654
rect 17500 63758 17502 63810
rect 17554 63758 17556 63810
rect 17500 63700 17556 63758
rect 16044 62578 16212 62580
rect 16044 62526 16046 62578
rect 16098 62526 16212 62578
rect 16044 62524 16212 62526
rect 16604 63196 16772 63252
rect 17276 63644 17556 63700
rect 16044 62514 16100 62524
rect 15708 62354 15764 62366
rect 15708 62302 15710 62354
rect 15762 62302 15764 62354
rect 15036 62244 15092 62254
rect 15036 61682 15092 62188
rect 15036 61630 15038 61682
rect 15090 61630 15092 61682
rect 15036 61618 15092 61630
rect 14812 60958 14814 61010
rect 14866 60958 14868 61010
rect 14812 60946 14868 60958
rect 15708 60564 15764 62302
rect 16268 62356 16324 62366
rect 16492 62356 16548 62366
rect 16268 62354 16548 62356
rect 16268 62302 16270 62354
rect 16322 62302 16494 62354
rect 16546 62302 16548 62354
rect 16268 62300 16548 62302
rect 16268 62290 16324 62300
rect 16492 62290 16548 62300
rect 15932 62244 15988 62282
rect 15932 62178 15988 62188
rect 16044 60898 16100 60910
rect 16044 60846 16046 60898
rect 16098 60846 16100 60898
rect 16044 60788 16100 60846
rect 16156 60900 16212 60910
rect 16156 60806 16212 60844
rect 16044 60722 16100 60732
rect 16604 60788 16660 63196
rect 16716 62466 16772 62478
rect 16716 62414 16718 62466
rect 16770 62414 16772 62466
rect 16716 60900 16772 62414
rect 16828 62468 16884 62478
rect 17276 62468 17332 63644
rect 16828 62466 17332 62468
rect 16828 62414 16830 62466
rect 16882 62414 17332 62466
rect 16828 62412 17332 62414
rect 17500 63140 17556 63150
rect 16828 62402 16884 62412
rect 17164 61682 17220 61694
rect 17164 61630 17166 61682
rect 17218 61630 17220 61682
rect 16828 60900 16884 60910
rect 16716 60898 16884 60900
rect 16716 60846 16830 60898
rect 16882 60846 16884 60898
rect 16716 60844 16884 60846
rect 17164 60900 17220 61630
rect 17388 60900 17444 60910
rect 17164 60844 17388 60900
rect 17500 60900 17556 63084
rect 17612 61572 17668 61582
rect 17724 61572 17780 64652
rect 17948 64642 18004 64652
rect 18620 64596 18676 64606
rect 18620 64594 19348 64596
rect 18620 64542 18622 64594
rect 18674 64542 19348 64594
rect 18620 64540 19348 64542
rect 18620 64530 18676 64540
rect 17948 64260 18004 64270
rect 17948 64146 18004 64204
rect 17948 64094 17950 64146
rect 18002 64094 18004 64146
rect 17948 64082 18004 64094
rect 19292 64146 19348 64540
rect 19836 64316 20100 64326
rect 19892 64260 19940 64316
rect 19996 64260 20044 64316
rect 19836 64250 20100 64260
rect 19292 64094 19294 64146
rect 19346 64094 19348 64146
rect 19292 64082 19348 64094
rect 20188 64148 20244 65996
rect 20300 65716 20356 66220
rect 20524 66948 20580 66958
rect 20524 66052 20580 66892
rect 21196 66724 21252 68124
rect 21308 68114 21364 68124
rect 21420 68066 21476 68460
rect 21980 68450 22036 68460
rect 21420 68014 21422 68066
rect 21474 68014 21476 68066
rect 21420 68002 21476 68014
rect 22876 68180 22932 68190
rect 21868 67844 21924 67854
rect 21868 67750 21924 67788
rect 22428 67844 22484 67854
rect 21308 67732 21364 67742
rect 21308 67638 21364 67676
rect 21980 67732 22036 67742
rect 21980 67638 22036 67676
rect 22092 67620 22148 67630
rect 21980 67284 22036 67294
rect 22092 67284 22148 67564
rect 21980 67282 22148 67284
rect 21980 67230 21982 67282
rect 22034 67230 22148 67282
rect 21980 67228 22148 67230
rect 22204 67396 22260 67406
rect 21980 67218 22036 67228
rect 21308 67170 21364 67182
rect 21308 67118 21310 67170
rect 21362 67118 21364 67170
rect 21308 66948 21364 67118
rect 21420 67058 21476 67070
rect 21420 67006 21422 67058
rect 21474 67006 21476 67058
rect 21420 66948 21476 67006
rect 21756 67058 21812 67070
rect 21756 67006 21758 67058
rect 21810 67006 21812 67058
rect 21756 66948 21812 67006
rect 21420 66892 21812 66948
rect 21308 66882 21364 66892
rect 21196 66668 21588 66724
rect 21420 66388 21476 66398
rect 21420 66294 21476 66332
rect 20524 65986 20580 65996
rect 20636 66050 20692 66062
rect 21308 66052 21364 66062
rect 20636 65998 20638 66050
rect 20690 65998 20692 66050
rect 20636 65716 20692 65998
rect 20300 65660 20692 65716
rect 20748 66050 21364 66052
rect 20748 65998 21310 66050
rect 21362 65998 21364 66050
rect 20748 65996 21364 65998
rect 20300 64148 20356 64158
rect 20188 64146 20356 64148
rect 20188 64094 20302 64146
rect 20354 64094 20356 64146
rect 20188 64092 20356 64094
rect 20300 64082 20356 64092
rect 20188 63922 20244 63934
rect 20188 63870 20190 63922
rect 20242 63870 20244 63922
rect 19404 63812 19460 63822
rect 19404 63810 19908 63812
rect 19404 63758 19406 63810
rect 19458 63758 19908 63810
rect 19404 63756 19908 63758
rect 19404 63746 19460 63756
rect 19852 63250 19908 63756
rect 19852 63198 19854 63250
rect 19906 63198 19908 63250
rect 19852 63186 19908 63198
rect 18732 63140 18788 63150
rect 19180 63140 19236 63150
rect 18788 63138 19236 63140
rect 18788 63086 19182 63138
rect 19234 63086 19236 63138
rect 18788 63084 19236 63086
rect 18732 63046 18788 63084
rect 19180 63074 19236 63084
rect 19740 63140 19796 63178
rect 20188 63140 20244 63870
rect 20412 63700 20468 65660
rect 20748 65602 20804 65996
rect 21308 65986 21364 65996
rect 21420 66052 21476 66062
rect 20748 65550 20750 65602
rect 20802 65550 20804 65602
rect 20748 65538 20804 65550
rect 20748 64818 20804 64830
rect 20748 64766 20750 64818
rect 20802 64766 20804 64818
rect 20748 64596 20804 64766
rect 21308 64596 21364 64606
rect 20748 64594 21364 64596
rect 20748 64542 21310 64594
rect 21362 64542 21364 64594
rect 20748 64540 21364 64542
rect 20524 63924 20580 63934
rect 20524 63922 21252 63924
rect 20524 63870 20526 63922
rect 20578 63870 21252 63922
rect 20524 63868 21252 63870
rect 20524 63858 20580 63868
rect 20412 63644 20692 63700
rect 20188 63084 20468 63140
rect 19740 63074 19796 63084
rect 19964 62916 20020 62926
rect 19628 62914 20020 62916
rect 19628 62862 19966 62914
rect 20018 62862 20020 62914
rect 19628 62860 20020 62862
rect 17948 62580 18004 62590
rect 17948 62486 18004 62524
rect 18508 62580 18564 62590
rect 18396 62356 18452 62366
rect 18508 62356 18564 62524
rect 18396 62354 18564 62356
rect 18396 62302 18398 62354
rect 18450 62302 18564 62354
rect 18396 62300 18564 62302
rect 18396 62290 18452 62300
rect 17612 61570 17724 61572
rect 17612 61518 17614 61570
rect 17666 61518 17724 61570
rect 17612 61516 17724 61518
rect 17612 61506 17668 61516
rect 17500 60844 17668 60900
rect 15708 60498 15764 60508
rect 16044 60562 16100 60574
rect 16044 60510 16046 60562
rect 16098 60510 16100 60562
rect 15484 60004 15540 60014
rect 15484 60002 15988 60004
rect 15484 59950 15486 60002
rect 15538 59950 15988 60002
rect 15484 59948 15988 59950
rect 15484 59938 15540 59948
rect 14700 59780 14756 59790
rect 14700 59330 14756 59724
rect 14700 59278 14702 59330
rect 14754 59278 14756 59330
rect 14700 59266 14756 59278
rect 15596 59778 15652 59790
rect 15596 59726 15598 59778
rect 15650 59726 15652 59778
rect 15596 58772 15652 59726
rect 15708 59780 15764 59790
rect 15708 59686 15764 59724
rect 15820 59778 15876 59790
rect 15820 59726 15822 59778
rect 15874 59726 15876 59778
rect 15820 58884 15876 59726
rect 15932 59780 15988 59948
rect 16044 60002 16100 60510
rect 16044 59950 16046 60002
rect 16098 59950 16100 60002
rect 16044 59938 16100 59950
rect 16492 59892 16548 59902
rect 16492 59798 16548 59836
rect 16380 59780 16436 59790
rect 15932 59778 16436 59780
rect 15932 59726 16382 59778
rect 16434 59726 16436 59778
rect 15932 59724 16436 59726
rect 16380 59714 16436 59724
rect 15820 58828 16212 58884
rect 15036 58716 16100 58772
rect 14924 58548 14980 58558
rect 14924 58454 14980 58492
rect 14812 58436 14868 58446
rect 14812 58342 14868 58380
rect 15036 58434 15092 58716
rect 15036 58382 15038 58434
rect 15090 58382 15092 58434
rect 15036 58370 15092 58382
rect 15484 58436 15540 58446
rect 15484 58342 15540 58380
rect 15260 58210 15316 58222
rect 15260 58158 15262 58210
rect 15314 58158 15316 58210
rect 15260 58100 15316 58158
rect 15260 58034 15316 58044
rect 14924 57876 14980 57886
rect 14924 56866 14980 57820
rect 14924 56814 14926 56866
rect 14978 56814 14980 56866
rect 14924 56802 14980 56814
rect 15148 56756 15204 56766
rect 14588 56252 14868 56308
rect 14476 53172 14532 53182
rect 14252 53170 14532 53172
rect 14252 53118 14478 53170
rect 14530 53118 14532 53170
rect 14252 53116 14532 53118
rect 14252 53060 14308 53116
rect 14476 53106 14532 53116
rect 13916 52162 14084 52164
rect 13916 52110 13918 52162
rect 13970 52110 14084 52162
rect 13916 52108 14084 52110
rect 14140 53004 14308 53060
rect 14140 52612 14196 53004
rect 13916 50484 13972 52108
rect 14140 52050 14196 52556
rect 14140 51998 14142 52050
rect 14194 51998 14196 52050
rect 14140 51986 14196 51998
rect 14364 52946 14420 52958
rect 14364 52894 14366 52946
rect 14418 52894 14420 52946
rect 13692 50372 13860 50428
rect 13916 50418 13972 50428
rect 14028 51492 14084 51502
rect 13580 49870 13582 49922
rect 13634 49870 13636 49922
rect 13580 49858 13636 49870
rect 12796 49812 12852 49822
rect 12796 49718 12852 49756
rect 12348 49086 12350 49138
rect 12402 49086 12404 49138
rect 12348 49074 12404 49086
rect 12460 49698 12516 49710
rect 12460 49646 12462 49698
rect 12514 49646 12516 49698
rect 12012 48738 12068 48748
rect 11676 48414 11678 48466
rect 11730 48414 11732 48466
rect 11676 48402 11732 48414
rect 12460 48468 12516 49646
rect 13580 49700 13636 49710
rect 12572 49252 12628 49262
rect 12572 49026 12628 49196
rect 13580 49138 13636 49644
rect 13580 49086 13582 49138
rect 13634 49086 13636 49138
rect 13580 49074 13636 49086
rect 13468 49028 13524 49038
rect 12572 48974 12574 49026
rect 12626 48974 12628 49026
rect 12572 48962 12628 48974
rect 13020 49026 13524 49028
rect 13020 48974 13470 49026
rect 13522 48974 13524 49026
rect 13020 48972 13524 48974
rect 12908 48914 12964 48926
rect 12908 48862 12910 48914
rect 12962 48862 12964 48914
rect 12796 48804 12852 48814
rect 12796 48710 12852 48748
rect 12460 48412 12628 48468
rect 11452 48244 11508 48254
rect 11340 48242 11508 48244
rect 11340 48190 11454 48242
rect 11506 48190 11508 48242
rect 11340 48188 11508 48190
rect 11340 47458 11396 48188
rect 11452 48178 11508 48188
rect 11788 48242 11844 48254
rect 11788 48190 11790 48242
rect 11842 48190 11844 48242
rect 11788 47572 11844 48190
rect 12460 48132 12516 48142
rect 12460 48038 12516 48076
rect 12572 47572 12628 48412
rect 12908 48244 12964 48862
rect 12908 48178 12964 48188
rect 13020 48020 13076 48972
rect 13468 48962 13524 48972
rect 13692 48916 13748 48926
rect 13692 48822 13748 48860
rect 12796 47964 13076 48020
rect 12796 47682 12852 47964
rect 12796 47630 12798 47682
rect 12850 47630 12852 47682
rect 12796 47618 12852 47630
rect 12684 47572 12740 47582
rect 11788 47570 12740 47572
rect 11788 47518 12686 47570
rect 12738 47518 12740 47570
rect 11788 47516 12740 47518
rect 12684 47506 12740 47516
rect 11340 47406 11342 47458
rect 11394 47406 11396 47458
rect 11340 47394 11396 47406
rect 11452 47234 11508 47246
rect 11452 47182 11454 47234
rect 11506 47182 11508 47234
rect 11452 47012 11508 47182
rect 11284 46956 11508 47012
rect 11564 47234 11620 47246
rect 11564 47182 11566 47234
rect 11618 47182 11620 47234
rect 11228 46946 11284 46956
rect 11564 46788 11620 47182
rect 11676 47236 11732 47246
rect 11676 47142 11732 47180
rect 11788 47234 11844 47246
rect 11788 47182 11790 47234
rect 11842 47182 11844 47234
rect 11676 46788 11732 46798
rect 11564 46786 11732 46788
rect 11564 46734 11678 46786
rect 11730 46734 11732 46786
rect 11564 46732 11732 46734
rect 11676 46722 11732 46732
rect 11788 46564 11844 47182
rect 12236 47236 12292 47246
rect 11676 46508 11844 46564
rect 12124 46788 12180 46798
rect 11564 46452 11620 46462
rect 11340 46004 11396 46014
rect 11396 45948 11508 46004
rect 11340 45938 11396 45948
rect 11116 45892 11172 45902
rect 11116 45798 11172 45836
rect 11228 45780 11284 45790
rect 11228 45686 11284 45724
rect 10892 45388 11060 45444
rect 11004 42868 11060 45388
rect 11452 45332 11508 45948
rect 11564 46002 11620 46396
rect 11676 46114 11732 46508
rect 11676 46062 11678 46114
rect 11730 46062 11732 46114
rect 11676 46050 11732 46062
rect 11564 45950 11566 46002
rect 11618 45950 11620 46002
rect 11564 45938 11620 45950
rect 11452 45276 11732 45332
rect 11676 45218 11732 45276
rect 11676 45166 11678 45218
rect 11730 45166 11732 45218
rect 11676 45154 11732 45166
rect 11116 44548 11172 44558
rect 11116 44436 11172 44492
rect 11452 44436 11508 44446
rect 11116 44434 11508 44436
rect 11116 44382 11118 44434
rect 11170 44382 11454 44434
rect 11506 44382 11508 44434
rect 11116 44380 11508 44382
rect 11116 44370 11172 44380
rect 11340 43764 11396 43774
rect 11004 42812 11172 42868
rect 10892 42642 10948 42654
rect 10892 42590 10894 42642
rect 10946 42590 10948 42642
rect 10892 42194 10948 42590
rect 11004 42642 11060 42654
rect 11004 42590 11006 42642
rect 11058 42590 11060 42642
rect 11004 42532 11060 42590
rect 11004 42466 11060 42476
rect 11116 42308 11172 42812
rect 10892 42142 10894 42194
rect 10946 42142 10948 42194
rect 10892 42130 10948 42142
rect 11004 42252 11172 42308
rect 10780 41918 10782 41970
rect 10834 41918 10836 41970
rect 10780 41906 10836 41918
rect 11004 41970 11060 42252
rect 11004 41918 11006 41970
rect 11058 41918 11060 41970
rect 11004 41906 11060 41918
rect 11340 41860 11396 43708
rect 11452 43762 11508 44380
rect 11900 44436 11956 44446
rect 11900 44212 11956 44380
rect 11900 44146 11956 44156
rect 11564 44100 11620 44110
rect 11564 44098 11732 44100
rect 11564 44046 11566 44098
rect 11618 44046 11732 44098
rect 11564 44044 11732 44046
rect 11564 44034 11620 44044
rect 11452 43710 11454 43762
rect 11506 43710 11508 43762
rect 11452 43652 11508 43710
rect 11676 43764 11732 44044
rect 12012 44098 12068 44110
rect 12012 44046 12014 44098
rect 12066 44046 12068 44098
rect 11676 43708 11844 43764
rect 11452 43586 11508 43596
rect 11788 43650 11844 43708
rect 11788 43598 11790 43650
rect 11842 43598 11844 43650
rect 11788 43586 11844 43598
rect 11676 43540 11732 43550
rect 11452 42980 11508 42990
rect 11676 42980 11732 43484
rect 11900 43428 11956 43438
rect 11788 43316 11844 43326
rect 11900 43316 11956 43372
rect 11788 43314 11956 43316
rect 11788 43262 11790 43314
rect 11842 43262 11956 43314
rect 11788 43260 11956 43262
rect 11788 43250 11844 43260
rect 11452 42978 11732 42980
rect 11452 42926 11454 42978
rect 11506 42926 11732 42978
rect 11452 42924 11732 42926
rect 11452 42914 11508 42924
rect 12012 42644 12068 44046
rect 12124 44100 12180 46732
rect 12124 43316 12180 44044
rect 12236 43764 12292 47180
rect 12348 46674 12404 46686
rect 12348 46622 12350 46674
rect 12402 46622 12404 46674
rect 12348 45106 12404 46622
rect 13804 46116 13860 50372
rect 13916 49028 13972 49038
rect 13916 48934 13972 48972
rect 14028 49026 14084 51436
rect 14364 50820 14420 52894
rect 14700 52946 14756 52958
rect 14700 52894 14702 52946
rect 14754 52894 14756 52946
rect 14588 52834 14644 52846
rect 14588 52782 14590 52834
rect 14642 52782 14644 52834
rect 14588 52724 14644 52782
rect 14700 52836 14756 52894
rect 14700 52770 14756 52780
rect 14588 52658 14644 52668
rect 14588 52164 14644 52174
rect 14588 52070 14644 52108
rect 14476 50820 14532 50830
rect 14364 50818 14532 50820
rect 14364 50766 14478 50818
rect 14530 50766 14532 50818
rect 14364 50764 14532 50766
rect 14476 50754 14532 50764
rect 14588 50708 14644 50718
rect 14588 50614 14644 50652
rect 14812 50428 14868 56252
rect 15148 56196 15204 56700
rect 15596 56644 15652 58716
rect 15932 58548 15988 58558
rect 15708 58546 15988 58548
rect 15708 58494 15934 58546
rect 15986 58494 15988 58546
rect 15708 58492 15988 58494
rect 15708 56978 15764 58492
rect 15932 58482 15988 58492
rect 16044 58434 16100 58716
rect 16044 58382 16046 58434
rect 16098 58382 16100 58434
rect 16044 58370 16100 58382
rect 15708 56926 15710 56978
rect 15762 56926 15764 56978
rect 15708 56914 15764 56926
rect 15932 58210 15988 58222
rect 15932 58158 15934 58210
rect 15986 58158 15988 58210
rect 15596 56308 15652 56588
rect 15708 56308 15764 56318
rect 15596 56306 15764 56308
rect 15596 56254 15710 56306
rect 15762 56254 15764 56306
rect 15596 56252 15764 56254
rect 15708 56242 15764 56252
rect 15932 56308 15988 58158
rect 15932 56242 15988 56252
rect 16044 58100 16100 58110
rect 16156 58100 16212 58828
rect 16492 58324 16548 58334
rect 16492 58230 16548 58268
rect 16268 58210 16324 58222
rect 16268 58158 16270 58210
rect 16322 58158 16324 58210
rect 16268 58100 16324 58158
rect 16604 58100 16660 60732
rect 16828 60676 16884 60844
rect 17388 60788 17444 60844
rect 17388 60732 17556 60788
rect 16828 60610 16884 60620
rect 17500 60674 17556 60732
rect 17500 60622 17502 60674
rect 17554 60622 17556 60674
rect 17500 60610 17556 60622
rect 17388 60564 17444 60574
rect 17388 60470 17444 60508
rect 16828 59892 16884 59902
rect 16828 59108 16884 59836
rect 17500 59444 17556 59454
rect 17612 59444 17668 60844
rect 16828 59014 16884 59052
rect 16940 59442 17668 59444
rect 16940 59390 17502 59442
rect 17554 59390 17668 59442
rect 16940 59388 17668 59390
rect 16100 58044 16324 58100
rect 16492 58044 16660 58100
rect 15148 55970 15204 56140
rect 15148 55918 15150 55970
rect 15202 55918 15204 55970
rect 15148 55906 15204 55918
rect 15484 56082 15540 56094
rect 15484 56030 15486 56082
rect 15538 56030 15540 56082
rect 15260 55412 15316 55422
rect 15148 54628 15204 54638
rect 15148 54534 15204 54572
rect 15260 54628 15316 55356
rect 15484 54740 15540 56030
rect 15932 56084 15988 56094
rect 16044 56084 16100 58044
rect 15932 56082 16100 56084
rect 15932 56030 15934 56082
rect 15986 56030 16100 56082
rect 15932 56028 16100 56030
rect 16156 56084 16212 56094
rect 16380 56084 16436 56094
rect 16156 56082 16436 56084
rect 16156 56030 16158 56082
rect 16210 56030 16382 56082
rect 16434 56030 16436 56082
rect 16156 56028 16436 56030
rect 15932 56018 15988 56028
rect 16156 56018 16212 56028
rect 16380 56018 16436 56028
rect 15820 55970 15876 55982
rect 15820 55918 15822 55970
rect 15874 55918 15876 55970
rect 15820 55468 15876 55918
rect 16492 55468 16548 58044
rect 16940 57652 16996 59388
rect 17500 59378 17556 59388
rect 17724 59276 17780 61516
rect 18284 61458 18340 61470
rect 18284 61406 18286 61458
rect 18338 61406 18340 61458
rect 18284 61348 18340 61406
rect 18284 61282 18340 61292
rect 17948 60788 18004 60798
rect 17948 60694 18004 60732
rect 17388 59220 17780 59276
rect 17836 60676 17892 60686
rect 17164 59108 17220 59118
rect 17164 58434 17220 59052
rect 17164 58382 17166 58434
rect 17218 58382 17220 58434
rect 17164 58370 17220 58382
rect 17276 58212 17332 58250
rect 17276 58146 17332 58156
rect 17388 57988 17444 59220
rect 17612 58436 17668 58446
rect 17612 58342 17668 58380
rect 17500 58324 17556 58334
rect 17500 58230 17556 58268
rect 17836 58212 17892 60620
rect 18508 59220 18564 62300
rect 18620 62466 18676 62478
rect 18620 62414 18622 62466
rect 18674 62414 18676 62466
rect 18620 61572 18676 62414
rect 19628 61572 19684 62860
rect 19964 62850 20020 62860
rect 20188 62916 20244 62926
rect 20188 62822 20244 62860
rect 19836 62748 20100 62758
rect 19892 62692 19940 62748
rect 19996 62692 20044 62748
rect 19836 62682 20100 62692
rect 20412 61684 20468 63084
rect 20636 62188 20692 63644
rect 20636 62132 20804 62188
rect 18620 61516 19684 61572
rect 20188 61682 20468 61684
rect 20188 61630 20414 61682
rect 20466 61630 20468 61682
rect 20188 61628 20468 61630
rect 18844 61348 18900 61358
rect 18844 61010 18900 61292
rect 18956 61236 19012 61516
rect 18956 61170 19012 61180
rect 19836 61180 20100 61190
rect 19892 61124 19940 61180
rect 19996 61124 20044 61180
rect 19836 61114 20100 61124
rect 19628 61012 19684 61022
rect 18844 60958 18846 61010
rect 18898 60958 18900 61010
rect 18844 60946 18900 60958
rect 18956 61010 19684 61012
rect 18956 60958 19630 61010
rect 19682 60958 19684 61010
rect 18956 60956 19684 60958
rect 18956 60898 19012 60956
rect 19628 60946 19684 60956
rect 19740 61012 19796 61022
rect 20188 61012 20244 61628
rect 20412 61618 20468 61628
rect 18956 60846 18958 60898
rect 19010 60846 19012 60898
rect 18956 60834 19012 60846
rect 19516 60788 19572 60798
rect 19516 60694 19572 60732
rect 19740 60786 19796 60956
rect 19740 60734 19742 60786
rect 19794 60734 19796 60786
rect 19404 60676 19460 60686
rect 19292 60620 19404 60676
rect 19180 59892 19236 59902
rect 18844 59444 18900 59454
rect 19068 59444 19124 59454
rect 18844 59442 19124 59444
rect 18844 59390 18846 59442
rect 18898 59390 19070 59442
rect 19122 59390 19124 59442
rect 18844 59388 19124 59390
rect 18844 59378 18900 59388
rect 18508 59164 18900 59220
rect 18844 58996 18900 59164
rect 18844 58940 19012 58996
rect 18732 58884 18788 58894
rect 17836 58146 17892 58156
rect 17948 58322 18004 58334
rect 17948 58270 17950 58322
rect 18002 58270 18004 58322
rect 17388 57932 17668 57988
rect 15596 55412 15876 55468
rect 16268 55412 16548 55468
rect 16604 56194 16660 56206
rect 16604 56142 16606 56194
rect 16658 56142 16660 56194
rect 15596 55410 15652 55412
rect 15596 55358 15598 55410
rect 15650 55358 15652 55410
rect 15596 55346 15652 55358
rect 15596 54740 15652 54750
rect 15484 54738 15652 54740
rect 15484 54686 15598 54738
rect 15650 54686 15652 54738
rect 15484 54684 15652 54686
rect 15596 54674 15652 54684
rect 15260 54626 15540 54628
rect 15260 54574 15262 54626
rect 15314 54574 15540 54626
rect 15260 54572 15540 54574
rect 15260 54562 15316 54572
rect 14924 54514 14980 54526
rect 14924 54462 14926 54514
rect 14978 54462 14980 54514
rect 14924 53058 14980 54462
rect 15484 54516 15540 54572
rect 15708 54516 15764 54526
rect 15484 54514 15764 54516
rect 15484 54462 15710 54514
rect 15762 54462 15764 54514
rect 15484 54460 15764 54462
rect 15708 54450 15764 54460
rect 16268 54514 16324 55412
rect 16268 54462 16270 54514
rect 16322 54462 16324 54514
rect 16268 54180 16324 54462
rect 16268 54114 16324 54124
rect 16380 55298 16436 55310
rect 16380 55246 16382 55298
rect 16434 55246 16436 55298
rect 16380 53844 16436 55246
rect 16380 53778 16436 53788
rect 16492 54628 16548 54638
rect 16604 54628 16660 56142
rect 16716 56196 16772 56206
rect 16716 56102 16772 56140
rect 16548 54572 16660 54628
rect 16268 53618 16324 53630
rect 16268 53566 16270 53618
rect 16322 53566 16324 53618
rect 16156 53508 16212 53518
rect 15932 53452 16156 53508
rect 15596 53172 15652 53182
rect 14924 53006 14926 53058
rect 14978 53006 14980 53058
rect 14924 52994 14980 53006
rect 15260 53170 15652 53172
rect 15260 53118 15598 53170
rect 15650 53118 15652 53170
rect 15260 53116 15652 53118
rect 15260 52274 15316 53116
rect 15596 53106 15652 53116
rect 15932 53058 15988 53452
rect 16156 53442 16212 53452
rect 15932 53006 15934 53058
rect 15986 53006 15988 53058
rect 15932 52994 15988 53006
rect 15372 52946 15428 52958
rect 15372 52894 15374 52946
rect 15426 52894 15428 52946
rect 15372 52612 15428 52894
rect 15372 52546 15428 52556
rect 15484 52946 15540 52958
rect 15708 52948 15764 52958
rect 15484 52894 15486 52946
rect 15538 52894 15540 52946
rect 15484 52724 15540 52894
rect 15260 52222 15262 52274
rect 15314 52222 15316 52274
rect 15260 52210 15316 52222
rect 14700 50372 14756 50382
rect 14812 50372 14980 50428
rect 14028 48974 14030 49026
rect 14082 48974 14084 49026
rect 14028 48962 14084 48974
rect 14252 50036 14308 50046
rect 14252 47346 14308 49980
rect 14700 49028 14756 50316
rect 14700 48934 14756 48972
rect 14588 48132 14644 48142
rect 14364 48130 14644 48132
rect 14364 48078 14590 48130
rect 14642 48078 14644 48130
rect 14364 48076 14644 48078
rect 14364 47570 14420 48076
rect 14588 48066 14644 48076
rect 14476 47684 14532 47694
rect 14476 47590 14532 47628
rect 14364 47518 14366 47570
rect 14418 47518 14420 47570
rect 14364 47506 14420 47518
rect 14252 47294 14254 47346
rect 14306 47294 14308 47346
rect 14252 47282 14308 47294
rect 14924 46228 14980 50372
rect 15484 49812 15540 52668
rect 15596 52946 15764 52948
rect 15596 52894 15710 52946
rect 15762 52894 15764 52946
rect 15596 52892 15764 52894
rect 15596 52836 15652 52892
rect 15708 52882 15764 52892
rect 15596 50036 15652 52780
rect 16268 51828 16324 53566
rect 15596 49970 15652 49980
rect 15708 51772 16324 51828
rect 16380 53508 16436 53518
rect 16492 53508 16548 54572
rect 16604 54180 16660 54190
rect 16660 54124 16772 54180
rect 16604 54114 16660 54124
rect 16380 53506 16548 53508
rect 16380 53454 16382 53506
rect 16434 53454 16548 53506
rect 16380 53452 16548 53454
rect 16604 53508 16660 53518
rect 15708 50708 15764 51772
rect 16268 51604 16324 51614
rect 16380 51604 16436 53452
rect 16604 53414 16660 53452
rect 16716 53284 16772 54124
rect 16604 53228 16772 53284
rect 16940 53506 16996 57596
rect 17612 57650 17668 57932
rect 17612 57598 17614 57650
rect 17666 57598 17668 57650
rect 17612 57586 17668 57598
rect 17836 56980 17892 56990
rect 17948 56980 18004 58270
rect 18620 58212 18676 58222
rect 18396 58210 18676 58212
rect 18396 58158 18622 58210
rect 18674 58158 18676 58210
rect 18396 58156 18676 58158
rect 18396 57762 18452 58156
rect 18620 58146 18676 58156
rect 18396 57710 18398 57762
rect 18450 57710 18452 57762
rect 18396 57698 18452 57710
rect 18620 57988 18676 57998
rect 18508 57092 18564 57102
rect 18508 56998 18564 57036
rect 17500 56978 18004 56980
rect 17500 56926 17838 56978
rect 17890 56926 18004 56978
rect 17500 56924 18004 56926
rect 17388 56308 17444 56318
rect 17388 56214 17444 56252
rect 17500 56194 17556 56924
rect 17836 56914 17892 56924
rect 18172 56868 18228 56878
rect 17500 56142 17502 56194
rect 17554 56142 17556 56194
rect 17500 56130 17556 56142
rect 17948 56866 18228 56868
rect 17948 56814 18174 56866
rect 18226 56814 18228 56866
rect 17948 56812 18228 56814
rect 17948 56306 18004 56812
rect 18172 56802 18228 56812
rect 18396 56756 18452 56766
rect 18396 56662 18452 56700
rect 17948 56254 17950 56306
rect 18002 56254 18004 56306
rect 17948 55468 18004 56254
rect 16940 53454 16942 53506
rect 16994 53454 16996 53506
rect 16492 53060 16548 53070
rect 16604 53060 16660 53228
rect 16492 53058 16660 53060
rect 16492 53006 16494 53058
rect 16546 53006 16660 53058
rect 16492 53004 16660 53006
rect 16492 52994 16548 53004
rect 16716 52948 16772 52958
rect 16716 52854 16772 52892
rect 16604 52612 16660 52622
rect 16660 52556 16772 52612
rect 16604 52546 16660 52556
rect 16268 51602 16436 51604
rect 16268 51550 16270 51602
rect 16322 51550 16436 51602
rect 16268 51548 16436 51550
rect 16604 52164 16660 52174
rect 16268 51538 16324 51548
rect 16492 51492 16548 51502
rect 16380 51436 16492 51492
rect 15484 49746 15540 49756
rect 15708 49698 15764 50652
rect 15820 51378 15876 51390
rect 15820 51326 15822 51378
rect 15874 51326 15876 51378
rect 15820 50484 15876 51326
rect 15820 50418 15876 50428
rect 16044 51378 16100 51390
rect 16044 51326 16046 51378
rect 16098 51326 16100 51378
rect 16044 49922 16100 51326
rect 16380 51378 16436 51436
rect 16492 51426 16548 51436
rect 16380 51326 16382 51378
rect 16434 51326 16436 51378
rect 16380 51314 16436 51326
rect 16604 50706 16660 52108
rect 16716 51602 16772 52556
rect 16716 51550 16718 51602
rect 16770 51550 16772 51602
rect 16716 51538 16772 51550
rect 16828 51492 16884 51502
rect 16828 51398 16884 51436
rect 16604 50654 16606 50706
rect 16658 50654 16660 50706
rect 16604 50372 16660 50654
rect 16940 50484 16996 53454
rect 17276 55412 18004 55468
rect 18396 55524 18452 55534
rect 16940 50418 16996 50428
rect 17052 52052 17108 52062
rect 16604 50306 16660 50316
rect 16268 50036 16324 50046
rect 16268 49942 16324 49980
rect 17052 49924 17108 51996
rect 16044 49870 16046 49922
rect 16098 49870 16100 49922
rect 16044 49858 16100 49870
rect 16828 49868 17108 49924
rect 17164 50596 17220 50606
rect 17164 49924 17220 50540
rect 17276 50148 17332 55412
rect 17836 55410 17892 55412
rect 17836 55358 17838 55410
rect 17890 55358 17892 55410
rect 17836 55336 17892 55358
rect 17388 55076 17444 55086
rect 17388 54982 17444 55020
rect 18396 55076 18452 55468
rect 18620 55468 18676 57932
rect 18732 56196 18788 58828
rect 18844 58434 18900 58446
rect 18844 58382 18846 58434
rect 18898 58382 18900 58434
rect 18844 57090 18900 58382
rect 18844 57038 18846 57090
rect 18898 57038 18900 57090
rect 18844 57026 18900 57038
rect 18956 56420 19012 58940
rect 19068 56980 19124 59388
rect 19180 58884 19236 59836
rect 19180 58818 19236 58828
rect 19180 58212 19236 58222
rect 19180 57090 19236 58156
rect 19180 57038 19182 57090
rect 19234 57038 19236 57090
rect 19180 57026 19236 57038
rect 19068 56420 19124 56924
rect 19292 56532 19348 60620
rect 19404 60610 19460 60620
rect 19628 60004 19684 60014
rect 19404 59948 19628 60004
rect 19404 59442 19460 59948
rect 19628 59910 19684 59948
rect 19740 59780 19796 60734
rect 19964 60956 20244 61012
rect 19964 60788 20020 60956
rect 19964 60722 20020 60732
rect 20076 60116 20132 60956
rect 20188 60786 20244 60798
rect 20188 60734 20190 60786
rect 20242 60734 20244 60786
rect 20188 60564 20244 60734
rect 20300 60788 20356 60798
rect 20300 60694 20356 60732
rect 20636 60786 20692 60798
rect 20636 60734 20638 60786
rect 20690 60734 20692 60786
rect 20524 60564 20580 60574
rect 20188 60562 20580 60564
rect 20188 60510 20526 60562
rect 20578 60510 20580 60562
rect 20188 60508 20580 60510
rect 20524 60498 20580 60508
rect 20636 60452 20692 60734
rect 20748 60564 20804 62132
rect 20860 61012 20916 61022
rect 20860 60918 20916 60956
rect 21196 60786 21252 63868
rect 21308 63140 21364 64540
rect 21420 64594 21476 65996
rect 21420 64542 21422 64594
rect 21474 64542 21476 64594
rect 21420 64530 21476 64542
rect 21308 63074 21364 63084
rect 21308 62916 21364 62926
rect 21364 62860 21476 62916
rect 21308 62850 21364 62860
rect 21308 62242 21364 62254
rect 21308 62190 21310 62242
rect 21362 62190 21364 62242
rect 21308 61572 21364 62190
rect 21308 61478 21364 61516
rect 21196 60734 21198 60786
rect 21250 60734 21252 60786
rect 21196 60722 21252 60734
rect 21420 60674 21476 62860
rect 21532 61348 21588 66668
rect 21644 66274 21700 66286
rect 21644 66222 21646 66274
rect 21698 66222 21700 66274
rect 21644 64706 21700 66222
rect 21756 65380 21812 66892
rect 21868 66946 21924 66958
rect 21868 66894 21870 66946
rect 21922 66894 21924 66946
rect 21868 66388 21924 66894
rect 21868 66322 21924 66332
rect 21980 66276 22036 66286
rect 22204 66276 22260 67340
rect 22316 67058 22372 67070
rect 22316 67006 22318 67058
rect 22370 67006 22372 67058
rect 22316 66498 22372 67006
rect 22428 66836 22484 67788
rect 22540 67842 22596 67854
rect 22540 67790 22542 67842
rect 22594 67790 22596 67842
rect 22540 67282 22596 67790
rect 22876 67842 22932 68124
rect 22876 67790 22878 67842
rect 22930 67790 22932 67842
rect 22876 67778 22932 67790
rect 22540 67230 22542 67282
rect 22594 67230 22596 67282
rect 22540 67218 22596 67230
rect 22876 67396 22932 67406
rect 22876 67282 22932 67340
rect 22876 67230 22878 67282
rect 22930 67230 22932 67282
rect 22876 67218 22932 67230
rect 22428 66770 22484 66780
rect 22652 67170 22708 67182
rect 22652 67118 22654 67170
rect 22706 67118 22708 67170
rect 22316 66446 22318 66498
rect 22370 66446 22372 66498
rect 22316 66434 22372 66446
rect 21980 66274 22260 66276
rect 21980 66222 21982 66274
rect 22034 66222 22260 66274
rect 21980 66220 22260 66222
rect 21980 66210 22036 66220
rect 21756 65314 21812 65324
rect 22204 66052 22260 66062
rect 22652 66052 22708 67118
rect 22876 66836 22932 66846
rect 22204 66050 22708 66052
rect 22204 65998 22206 66050
rect 22258 65998 22708 66050
rect 22204 65996 22708 65998
rect 22764 66780 22876 66836
rect 22204 65044 22260 65996
rect 21644 64654 21646 64706
rect 21698 64654 21700 64706
rect 21644 64642 21700 64654
rect 21868 64988 22260 65044
rect 21644 63028 21700 63038
rect 21644 62934 21700 62972
rect 21868 62188 21924 64988
rect 22764 64708 22820 66780
rect 22876 66770 22932 66780
rect 22988 65492 23044 68572
rect 23324 68626 23380 68638
rect 23324 68574 23326 68626
rect 23378 68574 23380 68626
rect 23100 67618 23156 67630
rect 23100 67566 23102 67618
rect 23154 67566 23156 67618
rect 23100 67396 23156 67566
rect 23100 67330 23156 67340
rect 23324 67172 23380 68574
rect 23548 68626 23604 68638
rect 23548 68574 23550 68626
rect 23602 68574 23604 68626
rect 23436 68068 23492 68078
rect 23436 67842 23492 68012
rect 23436 67790 23438 67842
rect 23490 67790 23492 67842
rect 23436 67172 23492 67790
rect 23548 67396 23604 68574
rect 23772 67956 23828 68686
rect 23996 68628 24052 68638
rect 24444 68628 24500 68638
rect 23884 68626 24052 68628
rect 23884 68574 23998 68626
rect 24050 68574 24052 68626
rect 23884 68572 24052 68574
rect 23884 68514 23940 68572
rect 23996 68562 24052 68572
rect 24332 68626 24500 68628
rect 24332 68574 24446 68626
rect 24498 68574 24500 68626
rect 24332 68572 24500 68574
rect 23884 68462 23886 68514
rect 23938 68462 23940 68514
rect 23884 68450 23940 68462
rect 23772 67900 23940 67956
rect 23772 67620 23828 67630
rect 23772 67526 23828 67564
rect 23884 67508 23940 67900
rect 24332 67620 24388 68572
rect 24444 68562 24500 68572
rect 24668 67844 24724 68798
rect 25452 68626 25508 70030
rect 25452 68574 25454 68626
rect 25506 68574 25508 68626
rect 24780 67956 24836 67966
rect 24780 67954 25172 67956
rect 24780 67902 24782 67954
rect 24834 67902 25172 67954
rect 24780 67900 25172 67902
rect 24780 67890 24836 67900
rect 24668 67778 24724 67788
rect 25116 67842 25172 67900
rect 25116 67790 25118 67842
rect 25170 67790 25172 67842
rect 25116 67778 25172 67790
rect 24892 67732 24948 67742
rect 24892 67638 24948 67676
rect 24332 67554 24388 67564
rect 24444 67618 24500 67630
rect 24444 67566 24446 67618
rect 24498 67566 24500 67618
rect 23996 67508 24052 67518
rect 23884 67452 23996 67508
rect 23996 67442 24052 67452
rect 24444 67508 24500 67566
rect 24444 67442 24500 67452
rect 24668 67618 24724 67630
rect 24668 67566 24670 67618
rect 24722 67566 24724 67618
rect 23548 67330 23604 67340
rect 24668 67396 24724 67566
rect 24668 67330 24724 67340
rect 23548 67172 23604 67182
rect 23996 67172 24052 67182
rect 23436 67170 23716 67172
rect 23436 67118 23550 67170
rect 23602 67118 23716 67170
rect 23436 67116 23716 67118
rect 23324 67106 23380 67116
rect 23548 67106 23604 67116
rect 23100 67060 23156 67070
rect 23100 66966 23156 67004
rect 23212 65602 23268 65614
rect 23212 65550 23214 65602
rect 23266 65550 23268 65602
rect 23100 65492 23156 65502
rect 22988 65436 23100 65492
rect 22876 65378 22932 65390
rect 22876 65326 22878 65378
rect 22930 65326 22932 65378
rect 22876 65268 22932 65326
rect 22876 65202 22932 65212
rect 22764 64652 22932 64708
rect 22764 64482 22820 64494
rect 22764 64430 22766 64482
rect 22818 64430 22820 64482
rect 22540 64146 22596 64158
rect 22540 64094 22542 64146
rect 22594 64094 22596 64146
rect 22316 63922 22372 63934
rect 22316 63870 22318 63922
rect 22370 63870 22372 63922
rect 22204 63810 22260 63822
rect 22204 63758 22206 63810
rect 22258 63758 22260 63810
rect 21980 63698 22036 63710
rect 21980 63646 21982 63698
rect 22034 63646 22036 63698
rect 21980 63138 22036 63646
rect 22204 63698 22260 63758
rect 22204 63646 22206 63698
rect 22258 63646 22260 63698
rect 22204 63634 22260 63646
rect 22204 63364 22260 63374
rect 21980 63086 21982 63138
rect 22034 63086 22036 63138
rect 21980 62804 22036 63086
rect 22092 63308 22204 63364
rect 22092 63138 22148 63308
rect 22204 63298 22260 63308
rect 22316 63140 22372 63870
rect 22092 63086 22094 63138
rect 22146 63086 22148 63138
rect 22092 63074 22148 63086
rect 22204 63084 22372 63140
rect 22428 63476 22484 63486
rect 22092 62804 22148 62814
rect 21980 62748 22092 62804
rect 22092 62738 22148 62748
rect 21868 62132 22036 62188
rect 21756 62076 22036 62132
rect 21532 61292 21700 61348
rect 21420 60622 21422 60674
rect 21474 60622 21476 60674
rect 21420 60610 21476 60622
rect 21532 60786 21588 60798
rect 21532 60734 21534 60786
rect 21586 60734 21588 60786
rect 20748 60508 21252 60564
rect 20076 60060 20244 60116
rect 19404 59390 19406 59442
rect 19458 59390 19460 59442
rect 19404 59378 19460 59390
rect 19628 59724 19796 59780
rect 19852 59780 19908 59790
rect 20076 59780 20132 59790
rect 19908 59778 20132 59780
rect 19908 59726 20078 59778
rect 20130 59726 20132 59778
rect 19908 59724 20132 59726
rect 19628 59276 19684 59724
rect 19852 59714 19908 59724
rect 20076 59714 20132 59724
rect 19836 59612 20100 59622
rect 19892 59556 19940 59612
rect 19996 59556 20044 59612
rect 19836 59546 20100 59556
rect 19964 59444 20020 59454
rect 20188 59444 20244 60060
rect 20524 60004 20580 60014
rect 20524 59910 20580 59948
rect 20636 59892 20692 60396
rect 20748 59892 20804 59902
rect 20636 59836 20748 59892
rect 20748 59798 20804 59836
rect 19964 59442 20356 59444
rect 19964 59390 19966 59442
rect 20018 59390 20356 59442
rect 19964 59388 20356 59390
rect 19964 59378 20020 59388
rect 19404 59220 19684 59276
rect 19740 59332 19796 59342
rect 19740 59238 19796 59276
rect 20188 59274 20244 59286
rect 20076 59220 20132 59230
rect 19404 57988 19460 59220
rect 20076 59106 20132 59164
rect 20076 59054 20078 59106
rect 20130 59054 20132 59106
rect 20076 59042 20132 59054
rect 20188 59222 20190 59274
rect 20242 59222 20244 59274
rect 20188 58548 20244 59222
rect 20300 58996 20356 59388
rect 20748 59220 20804 59230
rect 20748 59126 20804 59164
rect 20300 58940 20916 58996
rect 20188 58492 20468 58548
rect 19852 58436 19908 58446
rect 19852 58342 19908 58380
rect 20188 58322 20244 58334
rect 20188 58270 20190 58322
rect 20242 58270 20244 58322
rect 19404 57922 19460 57932
rect 19516 58210 19572 58222
rect 19740 58212 19796 58222
rect 19516 58158 19518 58210
rect 19570 58158 19572 58210
rect 19516 56868 19572 58158
rect 19628 58210 19796 58212
rect 19628 58158 19742 58210
rect 19794 58158 19796 58210
rect 19628 58156 19796 58158
rect 19628 57092 19684 58156
rect 19740 58146 19796 58156
rect 20188 58100 20244 58270
rect 20300 58212 20356 58222
rect 20300 58118 20356 58156
rect 19836 58044 20100 58054
rect 19892 57988 19940 58044
rect 19996 57988 20044 58044
rect 20188 58034 20244 58044
rect 19836 57978 20100 57988
rect 20412 57540 20468 58492
rect 20636 58436 20692 58446
rect 20524 58322 20580 58334
rect 20524 58270 20526 58322
rect 20578 58270 20580 58322
rect 20524 57764 20580 58270
rect 20636 57876 20692 58380
rect 20748 58324 20804 58334
rect 20748 58230 20804 58268
rect 20748 57876 20804 57886
rect 20636 57874 20804 57876
rect 20636 57822 20750 57874
rect 20802 57822 20804 57874
rect 20636 57820 20804 57822
rect 20860 57876 20916 58940
rect 20972 57876 21028 57886
rect 20860 57874 21028 57876
rect 20860 57822 20974 57874
rect 21026 57822 21028 57874
rect 20860 57820 21028 57822
rect 20748 57810 20804 57820
rect 20972 57810 21028 57820
rect 21084 57764 21140 57774
rect 20524 57708 20692 57764
rect 20524 57540 20580 57550
rect 20412 57538 20580 57540
rect 20412 57486 20526 57538
rect 20578 57486 20580 57538
rect 20412 57484 20580 57486
rect 19628 57026 19684 57036
rect 20300 57092 20356 57102
rect 20300 56998 20356 57036
rect 20412 56980 20468 57484
rect 20524 57474 20580 57484
rect 20636 57092 20692 57708
rect 21084 57670 21140 57708
rect 21196 57540 21252 60508
rect 21532 60452 21588 60734
rect 21532 60386 21588 60396
rect 21532 60116 21588 60126
rect 21420 59892 21476 59902
rect 21420 59330 21476 59836
rect 21532 59778 21588 60060
rect 21644 60004 21700 61292
rect 21756 61012 21812 62076
rect 22092 61684 22148 61694
rect 22204 61684 22260 63084
rect 22428 63026 22484 63420
rect 22428 62974 22430 63026
rect 22482 62974 22484 63026
rect 22316 62916 22372 62926
rect 22316 62822 22372 62860
rect 22092 61682 22260 61684
rect 22092 61630 22094 61682
rect 22146 61630 22260 61682
rect 22092 61628 22260 61630
rect 22092 61618 22148 61628
rect 22428 61572 22484 62974
rect 22428 61506 22484 61516
rect 22204 61460 22260 61470
rect 21812 60956 21924 61012
rect 21756 60918 21812 60956
rect 21644 59938 21700 59948
rect 21868 59890 21924 60956
rect 22204 60898 22260 61404
rect 22428 61012 22484 61022
rect 22540 61012 22596 64094
rect 22652 63922 22708 63934
rect 22652 63870 22654 63922
rect 22706 63870 22708 63922
rect 22652 63812 22708 63870
rect 22652 63746 22708 63756
rect 22764 63476 22820 64430
rect 22764 63410 22820 63420
rect 22876 63364 22932 64652
rect 22988 64706 23044 65436
rect 23100 65426 23156 65436
rect 22988 64654 22990 64706
rect 23042 64654 23044 64706
rect 22988 64642 23044 64654
rect 23212 65380 23268 65550
rect 22988 64148 23044 64158
rect 22988 64054 23044 64092
rect 22428 61010 22596 61012
rect 22428 60958 22430 61010
rect 22482 60958 22596 61010
rect 22428 60956 22596 60958
rect 22764 63138 22820 63150
rect 22764 63086 22766 63138
rect 22818 63086 22820 63138
rect 22764 62804 22820 63086
rect 22876 63140 22932 63308
rect 22988 63140 23044 63150
rect 22876 63138 23044 63140
rect 22876 63086 22990 63138
rect 23042 63086 23044 63138
rect 22876 63084 23044 63086
rect 22988 63074 23044 63084
rect 22428 60946 22484 60956
rect 22204 60846 22206 60898
rect 22258 60846 22260 60898
rect 22092 60788 22148 60798
rect 22092 60694 22148 60732
rect 22204 60116 22260 60846
rect 22652 60900 22708 60910
rect 22652 60806 22708 60844
rect 22204 60050 22260 60060
rect 22764 60788 22820 62748
rect 23100 63028 23156 63038
rect 23100 62356 23156 62972
rect 23100 62290 23156 62300
rect 23212 62188 23268 65324
rect 23436 65490 23492 65502
rect 23436 65438 23438 65490
rect 23490 65438 23492 65490
rect 23436 65268 23492 65438
rect 23324 63700 23380 63710
rect 23324 63606 23380 63644
rect 23436 62188 23492 65212
rect 23548 64484 23604 64494
rect 23548 64034 23604 64428
rect 23548 63982 23550 64034
rect 23602 63982 23604 64034
rect 23548 63970 23604 63982
rect 23548 63140 23604 63150
rect 23548 63046 23604 63084
rect 23660 62580 23716 67116
rect 23996 67078 24052 67116
rect 24220 67170 24276 67182
rect 24220 67118 24222 67170
rect 24274 67118 24276 67170
rect 24220 66948 24276 67118
rect 24220 66882 24276 66892
rect 24332 67058 24388 67070
rect 24332 67006 24334 67058
rect 24386 67006 24388 67058
rect 24332 66836 24388 67006
rect 24332 66770 24388 66780
rect 25452 66388 25508 68574
rect 25788 70082 25844 70094
rect 25788 70030 25790 70082
rect 25842 70030 25844 70082
rect 25676 67956 25732 67966
rect 25788 67956 25844 70030
rect 25900 69972 25956 69982
rect 25900 69970 26180 69972
rect 25900 69918 25902 69970
rect 25954 69918 26180 69970
rect 25900 69916 26180 69918
rect 25900 69906 25956 69916
rect 26124 69522 26180 69916
rect 26124 69470 26126 69522
rect 26178 69470 26180 69522
rect 26124 69458 26180 69470
rect 27804 69412 27860 70142
rect 28588 70084 28644 70094
rect 29708 70084 29764 70094
rect 28588 70082 28868 70084
rect 28588 70030 28590 70082
rect 28642 70030 28868 70082
rect 28588 70028 28868 70030
rect 28588 70018 28644 70028
rect 28252 69524 28308 69534
rect 28252 69522 28420 69524
rect 28252 69470 28254 69522
rect 28306 69470 28420 69522
rect 28252 69468 28420 69470
rect 28252 69458 28308 69468
rect 27804 68738 27860 69356
rect 27804 68686 27806 68738
rect 27858 68686 27860 68738
rect 27804 68674 27860 68686
rect 25676 67954 25844 67956
rect 25676 67902 25678 67954
rect 25730 67902 25844 67954
rect 25676 67900 25844 67902
rect 25676 67890 25732 67900
rect 26124 67844 26180 67854
rect 26124 67750 26180 67788
rect 28028 67844 28084 67854
rect 28252 67844 28308 67854
rect 28084 67842 28308 67844
rect 28084 67790 28254 67842
rect 28306 67790 28308 67842
rect 28084 67788 28308 67790
rect 28028 67750 28084 67788
rect 28252 67778 28308 67788
rect 26348 67732 26404 67742
rect 25564 67620 25620 67630
rect 25564 67526 25620 67564
rect 25788 67620 25844 67630
rect 25788 67526 25844 67564
rect 26236 67618 26292 67630
rect 26236 67566 26238 67618
rect 26290 67566 26292 67618
rect 26236 67284 26292 67566
rect 26348 67620 26404 67676
rect 26460 67620 26516 67630
rect 26348 67618 26516 67620
rect 26348 67566 26462 67618
rect 26514 67566 26516 67618
rect 26348 67564 26516 67566
rect 26460 67554 26516 67564
rect 28364 67620 28420 69468
rect 28812 67956 28868 70028
rect 29036 69300 29092 69310
rect 29036 69206 29092 69244
rect 29372 69298 29428 69310
rect 29372 69246 29374 69298
rect 29426 69246 29428 69298
rect 29260 69188 29316 69198
rect 29260 69094 29316 69132
rect 29372 68852 29428 69246
rect 29708 69186 29764 70028
rect 29708 69134 29710 69186
rect 29762 69134 29764 69186
rect 29708 68964 29764 69134
rect 29708 68898 29764 68908
rect 29820 69186 29876 69198
rect 29820 69134 29822 69186
rect 29874 69134 29876 69186
rect 29372 68786 29428 68796
rect 29820 68516 29876 69134
rect 29932 69186 29988 69198
rect 29932 69134 29934 69186
rect 29986 69134 29988 69186
rect 29932 69076 29988 69134
rect 29988 69020 30212 69076
rect 29932 69010 29988 69020
rect 29596 68460 29876 68516
rect 30044 68852 30100 68862
rect 29148 67956 29204 67966
rect 28812 67954 29204 67956
rect 28812 67902 29150 67954
rect 29202 67902 29204 67954
rect 28812 67900 29204 67902
rect 29148 67890 29204 67900
rect 29260 67956 29316 67966
rect 29596 67956 29652 68460
rect 29260 67954 29652 67956
rect 29260 67902 29262 67954
rect 29314 67902 29652 67954
rect 29260 67900 29652 67902
rect 29260 67890 29316 67900
rect 29708 67844 29764 67854
rect 29708 67842 29988 67844
rect 29708 67790 29710 67842
rect 29762 67790 29988 67842
rect 29708 67788 29988 67790
rect 29708 67778 29764 67788
rect 26236 67218 26292 67228
rect 28364 67172 28420 67564
rect 28140 67116 28364 67172
rect 25676 66946 25732 66958
rect 26124 66948 26180 66958
rect 25676 66894 25678 66946
rect 25730 66894 25732 66946
rect 25676 66834 25732 66894
rect 25676 66782 25678 66834
rect 25730 66782 25732 66834
rect 24892 66332 25508 66388
rect 25564 66386 25620 66398
rect 25564 66334 25566 66386
rect 25618 66334 25620 66386
rect 24668 66164 24724 66174
rect 24556 66162 24724 66164
rect 24556 66110 24670 66162
rect 24722 66110 24724 66162
rect 24556 66108 24724 66110
rect 24444 66050 24500 66062
rect 24444 65998 24446 66050
rect 24498 65998 24500 66050
rect 24444 65716 24500 65998
rect 24444 65650 24500 65660
rect 24220 65602 24276 65614
rect 24220 65550 24222 65602
rect 24274 65550 24276 65602
rect 23772 64820 23828 64830
rect 24220 64820 24276 65550
rect 23772 64818 24276 64820
rect 23772 64766 23774 64818
rect 23826 64766 24276 64818
rect 23772 64764 24276 64766
rect 24444 65490 24500 65502
rect 24444 65438 24446 65490
rect 24498 65438 24500 65490
rect 23772 64754 23828 64764
rect 24444 64148 24500 65438
rect 24556 64260 24612 66108
rect 24668 66098 24724 66108
rect 24780 66052 24836 66062
rect 24780 65958 24836 65996
rect 24892 65044 24948 66332
rect 25452 66164 25508 66174
rect 25452 66070 25508 66108
rect 24556 64194 24612 64204
rect 24668 64988 24948 65044
rect 25004 66050 25060 66062
rect 25004 65998 25006 66050
rect 25058 65998 25060 66050
rect 25004 65716 25060 65998
rect 25228 66050 25284 66062
rect 25228 65998 25230 66050
rect 25282 65998 25284 66050
rect 25228 65828 25284 65998
rect 25228 65762 25284 65772
rect 25564 66052 25620 66334
rect 25564 65716 25620 65996
rect 25676 65828 25732 66782
rect 26012 66946 26180 66948
rect 26012 66894 26126 66946
rect 26178 66894 26180 66946
rect 26012 66892 26180 66894
rect 25788 66276 25844 66286
rect 25788 66274 25956 66276
rect 25788 66222 25790 66274
rect 25842 66222 25956 66274
rect 25788 66220 25956 66222
rect 25788 66210 25844 66220
rect 25676 65762 25732 65772
rect 24444 64082 24500 64092
rect 23660 62514 23716 62524
rect 23772 63922 23828 63934
rect 24220 63924 24276 63934
rect 23772 63870 23774 63922
rect 23826 63870 23828 63922
rect 23212 62132 23380 62188
rect 23436 62132 23604 62188
rect 21868 59838 21870 59890
rect 21922 59838 21924 59890
rect 21868 59826 21924 59838
rect 22092 60002 22148 60014
rect 22092 59950 22094 60002
rect 22146 59950 22148 60002
rect 21532 59726 21534 59778
rect 21586 59726 21588 59778
rect 21532 59556 21588 59726
rect 21532 59490 21588 59500
rect 22092 59780 22148 59950
rect 22652 59780 22708 59790
rect 22092 59724 22652 59780
rect 21420 59278 21422 59330
rect 21474 59278 21476 59330
rect 21420 59266 21476 59278
rect 21532 59220 21588 59230
rect 21756 59220 21812 59230
rect 21532 59218 21700 59220
rect 21532 59166 21534 59218
rect 21586 59166 21700 59218
rect 21532 59164 21700 59166
rect 21532 59154 21588 59164
rect 20636 57026 20692 57036
rect 20972 57484 21252 57540
rect 21420 59106 21476 59118
rect 21420 59054 21422 59106
rect 21474 59054 21476 59106
rect 21420 58100 21476 59054
rect 21532 58548 21588 58558
rect 21532 58454 21588 58492
rect 21420 57874 21476 58044
rect 21420 57822 21422 57874
rect 21474 57822 21476 57874
rect 20412 56978 20580 56980
rect 20412 56926 20414 56978
rect 20466 56926 20580 56978
rect 20412 56924 20580 56926
rect 20412 56914 20468 56924
rect 19516 56802 19572 56812
rect 19404 56756 19460 56766
rect 19404 56662 19460 56700
rect 19292 56476 19684 56532
rect 19068 56364 19348 56420
rect 18956 56354 19012 56364
rect 18732 56140 19012 56196
rect 18956 56084 19012 56140
rect 18956 56028 19236 56084
rect 18956 55860 19012 55870
rect 18620 55412 18788 55468
rect 18396 54982 18452 55020
rect 18620 55300 18676 55310
rect 17500 54402 17556 54414
rect 17500 54350 17502 54402
rect 17554 54350 17556 54402
rect 17500 54180 17556 54350
rect 17500 54114 17556 54124
rect 18060 54402 18116 54414
rect 18060 54350 18062 54402
rect 18114 54350 18116 54402
rect 17948 53732 18004 53742
rect 17948 53638 18004 53676
rect 18060 53620 18116 54350
rect 18620 53730 18676 55244
rect 18620 53678 18622 53730
rect 18674 53678 18676 53730
rect 18620 53666 18676 53678
rect 18060 53564 18340 53620
rect 17612 53508 17668 53518
rect 17612 53506 18116 53508
rect 17612 53454 17614 53506
rect 17666 53454 18116 53506
rect 17612 53452 18116 53454
rect 17612 53442 17668 53452
rect 18060 53172 18116 53452
rect 17500 52946 17556 52958
rect 17500 52894 17502 52946
rect 17554 52894 17556 52946
rect 17388 52274 17444 52286
rect 17388 52222 17390 52274
rect 17442 52222 17444 52274
rect 17388 51492 17444 52222
rect 17500 52164 17556 52894
rect 17500 52098 17556 52108
rect 17948 51938 18004 51950
rect 17948 51886 17950 51938
rect 18002 51886 18004 51938
rect 17948 51828 18004 51886
rect 18060 51828 18116 53116
rect 18172 52836 18228 52846
rect 18172 52742 18228 52780
rect 18284 52162 18340 53564
rect 18284 52110 18286 52162
rect 18338 52110 18340 52162
rect 18172 52052 18228 52062
rect 18284 52052 18340 52110
rect 18732 52164 18788 55412
rect 18732 52098 18788 52108
rect 18228 51996 18340 52052
rect 18172 51986 18228 51996
rect 18396 51938 18452 51950
rect 18396 51886 18398 51938
rect 18450 51886 18452 51938
rect 18060 51772 18340 51828
rect 17836 51604 17892 51614
rect 17948 51604 18004 51772
rect 17836 51602 18004 51604
rect 17836 51550 17838 51602
rect 17890 51550 18004 51602
rect 17836 51548 18004 51550
rect 17836 51538 17892 51548
rect 17388 51426 17444 51436
rect 18060 51490 18116 51502
rect 18060 51438 18062 51490
rect 18114 51438 18116 51490
rect 17276 50082 17332 50092
rect 17500 50820 17556 50830
rect 17500 50034 17556 50764
rect 18060 50596 18116 51438
rect 18284 51378 18340 51772
rect 18284 51326 18286 51378
rect 18338 51326 18340 51378
rect 18284 51314 18340 51326
rect 18396 50820 18452 51886
rect 18620 51940 18676 51950
rect 18620 51846 18676 51884
rect 18844 51938 18900 51950
rect 18844 51886 18846 51938
rect 18898 51886 18900 51938
rect 18844 51828 18900 51886
rect 18844 51492 18900 51772
rect 18844 51426 18900 51436
rect 18396 50754 18452 50764
rect 18060 50530 18116 50540
rect 18956 50428 19012 55804
rect 19180 55468 19236 56028
rect 19068 55412 19236 55468
rect 19068 52050 19124 55412
rect 19180 52948 19236 52958
rect 19180 52386 19236 52892
rect 19180 52334 19182 52386
rect 19234 52334 19236 52386
rect 19180 52322 19236 52334
rect 19068 51998 19070 52050
rect 19122 51998 19124 52050
rect 19068 51604 19124 51998
rect 19068 51538 19124 51548
rect 19292 51492 19348 56364
rect 19628 55298 19684 56476
rect 19836 56476 20100 56486
rect 19892 56420 19940 56476
rect 19996 56420 20044 56476
rect 19836 56410 20100 56420
rect 20412 55970 20468 55982
rect 20412 55918 20414 55970
rect 20466 55918 20468 55970
rect 19628 55246 19630 55298
rect 19682 55246 19684 55298
rect 19628 55234 19684 55246
rect 20300 55858 20356 55870
rect 20300 55806 20302 55858
rect 20354 55806 20356 55858
rect 20300 55300 20356 55806
rect 20300 55234 20356 55244
rect 19852 55188 19908 55198
rect 19404 55076 19460 55086
rect 19852 55076 19908 55132
rect 19404 52162 19460 55020
rect 19628 55074 19908 55076
rect 19628 55022 19854 55074
rect 19906 55022 19908 55074
rect 19628 55020 19908 55022
rect 19964 55186 20020 55198
rect 19964 55134 19966 55186
rect 20018 55134 20020 55186
rect 19964 55076 20020 55134
rect 20300 55076 20356 55086
rect 19964 55020 20244 55076
rect 19628 54964 19684 55020
rect 19852 55010 19908 55020
rect 19404 52110 19406 52162
rect 19458 52110 19460 52162
rect 19404 52098 19460 52110
rect 19516 54908 19684 54964
rect 19836 54908 20100 54918
rect 17500 49982 17502 50034
rect 17554 49982 17556 50034
rect 17500 49970 17556 49982
rect 18844 50372 19012 50428
rect 19180 51436 19348 51492
rect 19404 51940 19460 51950
rect 17164 49868 17444 49924
rect 16492 49812 16548 49822
rect 15708 49646 15710 49698
rect 15762 49646 15764 49698
rect 15708 49634 15764 49646
rect 16380 49698 16436 49710
rect 16380 49646 16382 49698
rect 16434 49646 16436 49698
rect 16380 49252 16436 49646
rect 15372 49196 16436 49252
rect 15372 49138 15428 49196
rect 15372 49086 15374 49138
rect 15426 49086 15428 49138
rect 15372 49074 15428 49086
rect 15260 49028 15316 49038
rect 14924 46162 14980 46172
rect 15036 48804 15092 48814
rect 13804 46060 14196 46116
rect 12908 45890 12964 45902
rect 12908 45838 12910 45890
rect 12962 45838 12964 45890
rect 12348 45054 12350 45106
rect 12402 45054 12404 45106
rect 12348 43988 12404 45054
rect 12572 45778 12628 45790
rect 12572 45726 12574 45778
rect 12626 45726 12628 45778
rect 12572 44996 12628 45726
rect 12796 45780 12852 45790
rect 12684 45666 12740 45678
rect 12684 45614 12686 45666
rect 12738 45614 12740 45666
rect 12684 45108 12740 45614
rect 12684 45042 12740 45052
rect 12796 44996 12852 45724
rect 12908 45220 12964 45838
rect 13804 45890 13860 45902
rect 13804 45838 13806 45890
rect 13858 45838 13860 45890
rect 13468 45220 13524 45230
rect 12908 45218 13524 45220
rect 12908 45166 13470 45218
rect 13522 45166 13524 45218
rect 12908 45164 13524 45166
rect 13020 44996 13076 45006
rect 12796 44940 12964 44996
rect 12572 44930 12628 44940
rect 12460 44884 12516 44894
rect 12460 44546 12516 44828
rect 12460 44494 12462 44546
rect 12514 44494 12516 44546
rect 12460 44482 12516 44494
rect 12684 44884 12740 44894
rect 12572 44322 12628 44334
rect 12572 44270 12574 44322
rect 12626 44270 12628 44322
rect 12460 44100 12516 44110
rect 12572 44100 12628 44270
rect 12516 44044 12628 44100
rect 12460 44034 12516 44044
rect 12348 43922 12404 43932
rect 12236 43698 12292 43708
rect 12572 43764 12628 43774
rect 12684 43764 12740 44828
rect 12908 44546 12964 44940
rect 12908 44494 12910 44546
rect 12962 44494 12964 44546
rect 12908 44482 12964 44494
rect 12796 44322 12852 44334
rect 12796 44270 12798 44322
rect 12850 44270 12852 44322
rect 12796 44212 12852 44270
rect 12796 44146 12852 44156
rect 12572 43762 12740 43764
rect 12572 43710 12574 43762
rect 12626 43710 12740 43762
rect 12572 43708 12740 43710
rect 12796 43988 12852 43998
rect 12796 43764 12852 43932
rect 12572 43698 12628 43708
rect 12348 43652 12404 43662
rect 12348 43558 12404 43596
rect 12236 43540 12292 43550
rect 12236 43446 12292 43484
rect 12124 43250 12180 43260
rect 12012 42578 12068 42588
rect 12572 41972 12628 41982
rect 12796 41972 12852 43708
rect 12908 43540 12964 43550
rect 13020 43540 13076 44940
rect 13244 44884 13300 44894
rect 13244 44790 13300 44828
rect 12908 43538 13076 43540
rect 12908 43486 12910 43538
rect 12962 43486 13076 43538
rect 12908 43484 13076 43486
rect 13244 44212 13300 44222
rect 13244 43538 13300 44156
rect 13244 43486 13246 43538
rect 13298 43486 13300 43538
rect 12908 43428 12964 43484
rect 13244 43474 13300 43486
rect 12908 43362 12964 43372
rect 13020 43316 13076 43326
rect 13020 43222 13076 43260
rect 13356 43314 13412 43326
rect 13356 43262 13358 43314
rect 13410 43262 13412 43314
rect 13244 42084 13300 42094
rect 13356 42084 13412 43262
rect 13468 42756 13524 45164
rect 13804 45108 13860 45838
rect 14028 45108 14084 45118
rect 13804 45106 14084 45108
rect 13804 45054 14030 45106
rect 14082 45054 14084 45106
rect 13804 45052 14084 45054
rect 13580 44996 13636 45006
rect 13580 44902 13636 44940
rect 14028 44210 14084 45052
rect 14028 44158 14030 44210
rect 14082 44158 14084 44210
rect 13692 43764 13748 43774
rect 14028 43764 14084 44158
rect 13748 43708 14084 43764
rect 13692 43538 13748 43708
rect 13692 43486 13694 43538
rect 13746 43486 13748 43538
rect 13692 43474 13748 43486
rect 14140 43428 14196 46060
rect 14476 45780 14532 45790
rect 14476 45686 14532 45724
rect 14364 45108 14420 45118
rect 14364 43652 14420 45052
rect 14476 44996 14532 45006
rect 14700 44996 14756 45006
rect 14532 44994 14756 44996
rect 14532 44942 14702 44994
rect 14754 44942 14756 44994
rect 14532 44940 14756 44942
rect 14476 44930 14532 44940
rect 14700 44930 14756 44940
rect 14476 43652 14532 43662
rect 14364 43650 14532 43652
rect 14364 43598 14478 43650
rect 14530 43598 14532 43650
rect 14364 43596 14532 43598
rect 14476 43586 14532 43596
rect 14140 43372 14532 43428
rect 14028 43316 14084 43326
rect 13692 42756 13748 42766
rect 13468 42754 13748 42756
rect 13468 42702 13694 42754
rect 13746 42702 13748 42754
rect 13468 42700 13748 42702
rect 13692 42690 13748 42700
rect 14028 42754 14084 43260
rect 14028 42702 14030 42754
rect 14082 42702 14084 42754
rect 14028 42690 14084 42702
rect 13916 42644 13972 42654
rect 13916 42550 13972 42588
rect 13244 42082 13412 42084
rect 13244 42030 13246 42082
rect 13298 42030 13412 42082
rect 13244 42028 13412 42030
rect 13244 42018 13300 42028
rect 12572 41970 12852 41972
rect 12572 41918 12574 41970
rect 12626 41918 12852 41970
rect 12572 41916 12852 41918
rect 12572 41906 12628 41916
rect 11116 41804 11396 41860
rect 10892 41748 10948 41758
rect 10780 41412 10836 41422
rect 10892 41412 10948 41692
rect 11004 41412 11060 41422
rect 10892 41410 11060 41412
rect 10892 41358 11006 41410
rect 11058 41358 11060 41410
rect 10892 41356 11060 41358
rect 10780 41318 10836 41356
rect 11004 41346 11060 41356
rect 10668 40910 10670 40962
rect 10722 40910 10724 40962
rect 10668 40898 10724 40910
rect 11116 39730 11172 41804
rect 11676 41412 11732 41422
rect 11452 41410 11732 41412
rect 11452 41358 11678 41410
rect 11730 41358 11732 41410
rect 11452 41356 11732 41358
rect 11228 41188 11284 41198
rect 11452 41188 11508 41356
rect 11676 41346 11732 41356
rect 11228 41186 11508 41188
rect 11228 41134 11230 41186
rect 11282 41134 11508 41186
rect 11228 41132 11508 41134
rect 11228 41122 11284 41132
rect 11564 41076 11620 41086
rect 11564 40982 11620 41020
rect 12236 41076 12292 41086
rect 12236 40982 12292 41020
rect 12684 41076 12740 41086
rect 11788 40962 11844 40974
rect 11788 40910 11790 40962
rect 11842 40910 11844 40962
rect 11228 40404 11284 40414
rect 11788 40404 11844 40910
rect 11228 40402 11844 40404
rect 11228 40350 11230 40402
rect 11282 40350 11844 40402
rect 11228 40348 11844 40350
rect 12012 40962 12068 40974
rect 12012 40910 12014 40962
rect 12066 40910 12068 40962
rect 11228 39956 11284 40348
rect 11228 39890 11284 39900
rect 11116 39678 11118 39730
rect 11170 39678 11172 39730
rect 11116 39666 11172 39678
rect 11004 39620 11060 39630
rect 11004 39526 11060 39564
rect 11676 39618 11732 39630
rect 11676 39566 11678 39618
rect 11730 39566 11732 39618
rect 10556 39442 10612 39452
rect 11228 38834 11284 38846
rect 11228 38782 11230 38834
rect 11282 38782 11284 38834
rect 10668 38724 10724 38762
rect 10668 38658 10724 38668
rect 10780 38722 10836 38734
rect 10780 38670 10782 38722
rect 10834 38670 10836 38722
rect 10780 38276 10836 38670
rect 10780 38210 10836 38220
rect 11228 38052 11284 38782
rect 11228 37986 11284 37996
rect 11676 38164 11732 39566
rect 11900 39396 11956 39406
rect 11900 38946 11956 39340
rect 11900 38894 11902 38946
rect 11954 38894 11956 38946
rect 11900 38882 11956 38894
rect 10332 37154 10388 37166
rect 10332 37102 10334 37154
rect 10386 37102 10388 37154
rect 10220 37044 10276 37054
rect 10220 36950 10276 36988
rect 10220 35586 10276 35598
rect 10220 35534 10222 35586
rect 10274 35534 10276 35586
rect 10108 35476 10164 35486
rect 10108 35382 10164 35420
rect 10220 33908 10276 35534
rect 10332 35476 10388 37102
rect 11676 36932 11732 38108
rect 11900 38162 11956 38174
rect 11900 38110 11902 38162
rect 11954 38110 11956 38162
rect 11788 38052 11844 38062
rect 11788 37380 11844 37996
rect 11788 37286 11844 37324
rect 11900 37268 11956 38110
rect 11900 37202 11956 37212
rect 11676 36876 11844 36932
rect 11340 36594 11396 36606
rect 11340 36542 11342 36594
rect 11394 36542 11396 36594
rect 11004 35812 11060 35822
rect 10332 35410 10388 35420
rect 10556 35698 10612 35710
rect 10556 35646 10558 35698
rect 10610 35646 10612 35698
rect 10220 33842 10276 33852
rect 10556 34130 10612 35646
rect 10780 35700 10836 35710
rect 10780 35606 10836 35644
rect 10556 34078 10558 34130
rect 10610 34078 10612 34130
rect 9996 32620 10164 32676
rect 9996 32450 10052 32462
rect 9996 32398 9998 32450
rect 10050 32398 10052 32450
rect 9996 32340 10052 32398
rect 9996 32274 10052 32284
rect 10108 32116 10164 32620
rect 9548 31154 9604 31164
rect 9996 32060 10164 32116
rect 8988 30706 9044 30716
rect 9996 30660 10052 32060
rect 10108 31556 10164 31566
rect 10108 30994 10164 31500
rect 10108 30942 10110 30994
rect 10162 30942 10164 30994
rect 10108 30930 10164 30942
rect 10556 30996 10612 34078
rect 11004 34130 11060 35756
rect 11116 35476 11172 35486
rect 11116 35382 11172 35420
rect 11340 35476 11396 36542
rect 11340 35410 11396 35420
rect 11788 35698 11844 36876
rect 11788 35646 11790 35698
rect 11842 35646 11844 35698
rect 11228 35028 11284 35038
rect 11228 34934 11284 34972
rect 11004 34078 11006 34130
rect 11058 34078 11060 34130
rect 11004 34066 11060 34078
rect 11788 34132 11844 35646
rect 12012 34916 12068 40910
rect 12684 40962 12740 41020
rect 12684 40910 12686 40962
rect 12738 40910 12740 40962
rect 12684 40628 12740 40910
rect 12684 40562 12740 40572
rect 13916 40290 13972 40302
rect 13916 40238 13918 40290
rect 13970 40238 13972 40290
rect 12908 39842 12964 39854
rect 12908 39790 12910 39842
rect 12962 39790 12964 39842
rect 12908 39732 12964 39790
rect 13916 39844 13972 40238
rect 13916 39778 13972 39788
rect 12908 39666 12964 39676
rect 13580 39732 13636 39742
rect 13580 39638 13636 39676
rect 12684 39618 12740 39630
rect 12684 39566 12686 39618
rect 12738 39566 12740 39618
rect 12684 38724 12740 39566
rect 12684 38658 12740 38668
rect 12908 39506 12964 39518
rect 12908 39454 12910 39506
rect 12962 39454 12964 39506
rect 12908 37940 12964 39454
rect 13468 39396 13524 39406
rect 14028 39396 14084 39406
rect 13468 39302 13524 39340
rect 13580 39340 14028 39396
rect 13468 38276 13524 38286
rect 13468 38182 13524 38220
rect 13468 37940 13524 37950
rect 13580 37940 13636 39340
rect 14028 39302 14084 39340
rect 14028 38724 14084 38762
rect 14028 38658 14084 38668
rect 14364 38724 14420 38734
rect 14252 38612 14308 38622
rect 12908 37938 13636 37940
rect 12908 37886 13470 37938
rect 13522 37886 13636 37938
rect 12908 37884 13636 37886
rect 13692 38050 13748 38062
rect 13692 37998 13694 38050
rect 13746 37998 13748 38050
rect 12236 37268 12292 37278
rect 12236 35698 12292 37212
rect 12908 36258 12964 37884
rect 13468 37874 13524 37884
rect 12908 36206 12910 36258
rect 12962 36206 12964 36258
rect 12236 35646 12238 35698
rect 12290 35646 12292 35698
rect 12236 35634 12292 35646
rect 12684 35698 12740 35710
rect 12684 35646 12686 35698
rect 12738 35646 12740 35698
rect 12012 34850 12068 34860
rect 12348 35476 12404 35486
rect 12684 35476 12740 35646
rect 12908 35588 12964 36206
rect 13468 37380 13524 37390
rect 13468 36482 13524 37324
rect 13692 37268 13748 37998
rect 13692 37202 13748 37212
rect 14252 36594 14308 38556
rect 14364 38052 14420 38668
rect 14476 38388 14532 43372
rect 15036 39956 15092 48748
rect 15260 48242 15316 48972
rect 16492 49028 16548 49756
rect 16492 48962 16548 48972
rect 16716 49810 16772 49822
rect 16716 49758 16718 49810
rect 16770 49758 16772 49810
rect 16716 48466 16772 49758
rect 16828 49700 16884 49868
rect 16828 49644 17108 49700
rect 16716 48414 16718 48466
rect 16770 48414 16772 48466
rect 16716 48402 16772 48414
rect 16940 49476 16996 49486
rect 16828 48356 16884 48366
rect 16828 48262 16884 48300
rect 15260 48190 15262 48242
rect 15314 48190 15316 48242
rect 15260 48178 15316 48190
rect 16044 48242 16100 48254
rect 16044 48190 16046 48242
rect 16098 48190 16100 48242
rect 15708 48132 15764 48142
rect 15708 48038 15764 48076
rect 15820 48130 15876 48142
rect 15820 48078 15822 48130
rect 15874 48078 15876 48130
rect 15820 47684 15876 48078
rect 15820 47618 15876 47628
rect 16044 47348 16100 48190
rect 16044 47254 16100 47292
rect 16268 47572 16324 47582
rect 16268 47236 16324 47516
rect 16268 47170 16324 47180
rect 16940 46788 16996 49420
rect 17052 47068 17108 49644
rect 17388 49364 17444 49868
rect 18508 49810 18564 49822
rect 18508 49758 18510 49810
rect 18562 49758 18564 49810
rect 18060 49700 18116 49710
rect 18508 49700 18564 49758
rect 18060 49698 18564 49700
rect 18060 49646 18062 49698
rect 18114 49646 18564 49698
rect 18060 49644 18564 49646
rect 18060 49634 18116 49644
rect 17836 49588 17892 49598
rect 17836 49494 17892 49532
rect 17388 49308 17668 49364
rect 17500 49140 17556 49150
rect 17388 49138 17556 49140
rect 17388 49086 17502 49138
rect 17554 49086 17556 49138
rect 17388 49084 17556 49086
rect 17388 48356 17444 49084
rect 17500 49074 17556 49084
rect 17500 48468 17556 48478
rect 17612 48468 17668 49308
rect 18284 49028 18340 49038
rect 18284 48934 18340 48972
rect 17500 48466 17668 48468
rect 17500 48414 17502 48466
rect 17554 48414 17668 48466
rect 17500 48412 17668 48414
rect 17724 48916 17780 48926
rect 17724 48466 17780 48860
rect 17724 48414 17726 48466
rect 17778 48414 17780 48466
rect 17500 48402 17556 48412
rect 17724 48402 17780 48414
rect 17836 48914 17892 48926
rect 17836 48862 17838 48914
rect 17890 48862 17892 48914
rect 17388 48262 17444 48300
rect 17388 47236 17444 47246
rect 17276 47180 17388 47236
rect 17052 47012 17220 47068
rect 16940 46732 17108 46788
rect 16940 46562 16996 46574
rect 16940 46510 16942 46562
rect 16994 46510 16996 46562
rect 16604 46002 16660 46014
rect 16604 45950 16606 46002
rect 16658 45950 16660 46002
rect 16604 45332 16660 45950
rect 16604 45266 16660 45276
rect 16828 44994 16884 45006
rect 16828 44942 16830 44994
rect 16882 44942 16884 44994
rect 15932 43764 15988 43774
rect 15372 41858 15428 41870
rect 15372 41806 15374 41858
rect 15426 41806 15428 41858
rect 15372 41300 15428 41806
rect 15484 41300 15540 41310
rect 15372 41298 15540 41300
rect 15372 41246 15486 41298
rect 15538 41246 15540 41298
rect 15372 41244 15540 41246
rect 15484 41234 15540 41244
rect 15708 41186 15764 41198
rect 15708 41134 15710 41186
rect 15762 41134 15764 41186
rect 15708 41076 15764 41134
rect 15708 41010 15764 41020
rect 15036 39890 15092 39900
rect 15260 39620 15316 39630
rect 15932 39620 15988 43708
rect 16828 43540 16884 44942
rect 16940 43988 16996 46510
rect 16940 43922 16996 43932
rect 16828 43474 16884 43484
rect 16604 43426 16660 43438
rect 16604 43374 16606 43426
rect 16658 43374 16660 43426
rect 16604 43316 16660 43374
rect 16604 43250 16660 43260
rect 16044 41300 16100 41310
rect 16044 41298 16660 41300
rect 16044 41246 16046 41298
rect 16098 41246 16660 41298
rect 16044 41244 16660 41246
rect 16044 41234 16100 41244
rect 16604 41186 16660 41244
rect 16604 41134 16606 41186
rect 16658 41134 16660 41186
rect 16604 41122 16660 41134
rect 16380 40964 16436 40974
rect 16044 40962 16436 40964
rect 16044 40910 16382 40962
rect 16434 40910 16436 40962
rect 16044 40908 16436 40910
rect 16044 40514 16100 40908
rect 16380 40898 16436 40908
rect 16044 40462 16046 40514
rect 16098 40462 16100 40514
rect 16044 40450 16100 40462
rect 16828 40740 16884 40750
rect 16828 40402 16884 40684
rect 16828 40350 16830 40402
rect 16882 40350 16884 40402
rect 16828 40338 16884 40350
rect 17052 40292 17108 46732
rect 17164 46004 17220 47012
rect 17164 45910 17220 45948
rect 16268 40068 16324 40078
rect 16156 40012 16268 40068
rect 16044 39620 16100 39630
rect 15932 39618 16100 39620
rect 15932 39566 16046 39618
rect 16098 39566 16100 39618
rect 15932 39564 16100 39566
rect 15036 39172 15092 39182
rect 14588 39060 14644 39070
rect 14588 38966 14644 39004
rect 15036 38834 15092 39116
rect 15260 39060 15316 39564
rect 16044 39554 16100 39564
rect 15708 39508 15764 39518
rect 15708 39506 15876 39508
rect 15708 39454 15710 39506
rect 15762 39454 15876 39506
rect 15708 39452 15876 39454
rect 15708 39442 15764 39452
rect 15260 38966 15316 39004
rect 15372 39394 15428 39406
rect 15596 39396 15652 39406
rect 15372 39342 15374 39394
rect 15426 39342 15428 39394
rect 15036 38782 15038 38834
rect 15090 38782 15092 38834
rect 15036 38770 15092 38782
rect 14476 38322 14532 38332
rect 14588 38164 14644 38174
rect 14476 38052 14532 38062
rect 14364 38050 14532 38052
rect 14364 37998 14478 38050
rect 14530 37998 14532 38050
rect 14364 37996 14532 37998
rect 14476 37986 14532 37996
rect 14588 38050 14644 38108
rect 14588 37998 14590 38050
rect 14642 37998 14644 38050
rect 14588 37986 14644 37998
rect 14252 36542 14254 36594
rect 14306 36542 14308 36594
rect 14252 36530 14308 36542
rect 14364 37492 14420 37502
rect 13468 36430 13470 36482
rect 13522 36430 13524 36482
rect 13468 35700 13524 36430
rect 14364 35810 14420 37436
rect 15372 37492 15428 39342
rect 15484 39394 15652 39396
rect 15484 39342 15598 39394
rect 15650 39342 15652 39394
rect 15484 39340 15652 39342
rect 15484 37940 15540 39340
rect 15596 39330 15652 39340
rect 15708 38722 15764 38734
rect 15708 38670 15710 38722
rect 15762 38670 15764 38722
rect 15596 38612 15652 38622
rect 15596 38518 15652 38556
rect 15708 38276 15764 38670
rect 15708 38210 15764 38220
rect 15708 38052 15764 38062
rect 15708 37958 15764 37996
rect 15484 37874 15540 37884
rect 15372 37426 15428 37436
rect 15820 37492 15876 39452
rect 16156 39396 16212 40012
rect 16268 40002 16324 40012
rect 16828 39732 16884 39742
rect 16828 39638 16884 39676
rect 15820 37426 15876 37436
rect 15932 39340 16212 39396
rect 17052 39396 17108 40236
rect 15932 39172 15988 39340
rect 17052 39330 17108 39340
rect 14364 35758 14366 35810
rect 14418 35758 14420 35810
rect 14364 35746 14420 35758
rect 15372 36148 15428 36158
rect 13580 35700 13636 35710
rect 13468 35698 13636 35700
rect 13468 35646 13582 35698
rect 13634 35646 13636 35698
rect 13468 35644 13636 35646
rect 13132 35588 13188 35598
rect 12908 35586 13188 35588
rect 12908 35534 13134 35586
rect 13186 35534 13188 35586
rect 12908 35532 13188 35534
rect 13132 35522 13188 35532
rect 12404 35420 12740 35476
rect 12124 34692 12180 34702
rect 12124 34598 12180 34636
rect 11788 34038 11844 34076
rect 12236 34132 12292 34142
rect 12348 34132 12404 35420
rect 12236 34130 12404 34132
rect 12236 34078 12238 34130
rect 12290 34078 12404 34130
rect 12236 34076 12404 34078
rect 12460 35026 12516 35038
rect 12460 34974 12462 35026
rect 12514 34974 12516 35026
rect 12236 34066 12292 34076
rect 11116 33908 11172 33918
rect 11116 33814 11172 33852
rect 11116 33458 11172 33470
rect 11116 33406 11118 33458
rect 11170 33406 11172 33458
rect 11116 32564 11172 33406
rect 11116 32340 11172 32508
rect 11788 33124 11844 33134
rect 11788 32562 11844 33068
rect 11788 32510 11790 32562
rect 11842 32510 11844 32562
rect 11788 32498 11844 32510
rect 12124 32562 12180 32574
rect 12124 32510 12126 32562
rect 12178 32510 12180 32562
rect 10892 32284 11172 32340
rect 12012 32340 12068 32350
rect 10556 30902 10612 30940
rect 10780 31890 10836 31902
rect 10780 31838 10782 31890
rect 10834 31838 10836 31890
rect 10332 30772 10388 30782
rect 10332 30678 10388 30716
rect 10780 30772 10836 31838
rect 10892 30882 10948 32284
rect 12012 32246 12068 32284
rect 11340 32228 11396 32238
rect 11340 31780 11396 32172
rect 10892 30830 10894 30882
rect 10946 30830 10948 30882
rect 10892 30818 10948 30830
rect 11004 31778 11396 31780
rect 11004 31726 11342 31778
rect 11394 31726 11396 31778
rect 11004 31724 11396 31726
rect 10780 30706 10836 30716
rect 9996 30594 10052 30604
rect 10780 30322 10836 30334
rect 10780 30270 10782 30322
rect 10834 30270 10836 30322
rect 7980 30210 8484 30212
rect 7980 30158 7982 30210
rect 8034 30158 8484 30210
rect 7980 30156 8484 30158
rect 7980 30146 8036 30156
rect 2044 30046 2046 30098
rect 2098 30046 2100 30098
rect 2044 30034 2100 30046
rect 1708 29586 1764 29596
rect 2940 29986 2996 29998
rect 2940 29934 2942 29986
rect 2994 29934 2996 29986
rect 2940 29652 2996 29934
rect 2940 29586 2996 29596
rect 2044 29540 2100 29550
rect 2044 29446 2100 29484
rect 1708 29426 1764 29438
rect 1708 29374 1710 29426
rect 1762 29374 1764 29426
rect 1708 28980 1764 29374
rect 1708 28914 1764 28924
rect 2492 29314 2548 29326
rect 2492 29262 2494 29314
rect 2546 29262 2548 29314
rect 2492 28980 2548 29262
rect 4476 29036 4740 29046
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4476 28970 4740 28980
rect 2492 28914 2548 28924
rect 1708 28642 1764 28654
rect 1708 28590 1710 28642
rect 1762 28590 1764 28642
rect 1708 28308 1764 28590
rect 2044 28644 2100 28654
rect 2044 28418 2100 28588
rect 2044 28366 2046 28418
rect 2098 28366 2100 28418
rect 2044 28354 2100 28366
rect 2492 28642 2548 28654
rect 2492 28590 2494 28642
rect 2546 28590 2548 28642
rect 1708 28242 1764 28252
rect 2492 28308 2548 28590
rect 2492 28242 2548 28252
rect 8316 28644 8372 28654
rect 2044 27972 2100 27982
rect 2044 27878 2100 27916
rect 1708 27858 1764 27870
rect 1708 27806 1710 27858
rect 1762 27806 1764 27858
rect 1708 27636 1764 27806
rect 1708 27570 1764 27580
rect 2492 27746 2548 27758
rect 2492 27694 2494 27746
rect 2546 27694 2548 27746
rect 2492 27636 2548 27694
rect 2492 27570 2548 27580
rect 2716 27636 2772 27646
rect 1708 26964 1764 26974
rect 1708 26870 1764 26908
rect 2380 26962 2436 26974
rect 2380 26910 2382 26962
rect 2434 26910 2436 26962
rect 2044 26852 2100 26862
rect 2044 26758 2100 26796
rect 2380 26852 2436 26910
rect 2156 26740 2212 26750
rect 2044 26516 2100 26526
rect 2156 26516 2212 26684
rect 2044 26514 2212 26516
rect 2044 26462 2046 26514
rect 2098 26462 2212 26514
rect 2044 26460 2212 26462
rect 2044 26450 2100 26460
rect 1708 26290 1764 26302
rect 1708 26238 1710 26290
rect 1762 26238 1764 26290
rect 1708 26180 1764 26238
rect 2380 26292 2436 26796
rect 2492 26964 2548 26974
rect 2492 26514 2548 26908
rect 2716 26962 2772 27580
rect 4476 27468 4740 27478
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4476 27402 4740 27412
rect 8316 27412 8372 28588
rect 8316 27346 8372 27356
rect 8428 28530 8484 30156
rect 8652 30100 8708 30110
rect 10108 30100 10164 30110
rect 8652 30098 8932 30100
rect 8652 30046 8654 30098
rect 8706 30046 8932 30098
rect 8652 30044 8932 30046
rect 8652 30034 8708 30044
rect 8876 29650 8932 30044
rect 8876 29598 8878 29650
rect 8930 29598 8932 29650
rect 8876 29586 8932 29598
rect 10108 29426 10164 30044
rect 10108 29374 10110 29426
rect 10162 29374 10164 29426
rect 10108 29362 10164 29374
rect 10556 29428 10612 29438
rect 10556 29334 10612 29372
rect 8988 29314 9044 29326
rect 8988 29262 8990 29314
rect 9042 29262 9044 29314
rect 8988 29204 9044 29262
rect 10780 29316 10836 30270
rect 10780 29250 10836 29260
rect 8988 29138 9044 29148
rect 10332 29204 10388 29214
rect 10332 29110 10388 29148
rect 8428 28478 8430 28530
rect 8482 28478 8484 28530
rect 8428 27074 8484 28478
rect 9996 28868 10052 28878
rect 8428 27022 8430 27074
rect 8482 27022 8484 27074
rect 2716 26910 2718 26962
rect 2770 26910 2772 26962
rect 2716 26898 2772 26910
rect 3164 26962 3220 26974
rect 3164 26910 3166 26962
rect 3218 26910 3220 26962
rect 3164 26852 3220 26910
rect 3164 26786 3220 26796
rect 6524 26964 6580 26974
rect 2492 26462 2494 26514
rect 2546 26462 2548 26514
rect 2492 26450 2548 26462
rect 2380 26226 2436 26236
rect 1708 25620 1764 26124
rect 2940 26180 2996 26190
rect 2940 26086 2996 26124
rect 4476 25900 4740 25910
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4476 25834 4740 25844
rect 1708 25554 1764 25564
rect 2044 25508 2100 25518
rect 6524 25508 6580 26908
rect 8428 26964 8484 27022
rect 8428 26898 8484 26908
rect 8988 27972 9044 27982
rect 8316 26178 8372 26190
rect 8316 26126 8318 26178
rect 8370 26126 8372 26178
rect 8204 26068 8260 26078
rect 7196 26066 8260 26068
rect 7196 26014 8206 26066
rect 8258 26014 8260 26066
rect 7196 26012 8260 26014
rect 7196 25618 7252 26012
rect 8204 26002 8260 26012
rect 7196 25566 7198 25618
rect 7250 25566 7252 25618
rect 7196 25554 7252 25566
rect 1708 25394 1764 25406
rect 1708 25342 1710 25394
rect 1762 25342 1764 25394
rect 1708 24948 1764 25342
rect 2044 25394 2100 25452
rect 2044 25342 2046 25394
rect 2098 25342 2100 25394
rect 2044 25330 2100 25342
rect 5628 25506 6580 25508
rect 5628 25454 6526 25506
rect 6578 25454 6580 25506
rect 5628 25452 6580 25454
rect 1708 24882 1764 24892
rect 2492 25282 2548 25294
rect 2492 25230 2494 25282
rect 2546 25230 2548 25282
rect 2492 24948 2548 25230
rect 2492 24882 2548 24892
rect 2044 24836 2100 24846
rect 2044 24834 2212 24836
rect 2044 24782 2046 24834
rect 2098 24782 2212 24834
rect 2044 24780 2212 24782
rect 2044 24770 2100 24780
rect 1708 24722 1764 24734
rect 1708 24670 1710 24722
rect 1762 24670 1764 24722
rect 1708 24276 1764 24670
rect 1708 24210 1764 24220
rect 1708 23826 1764 23838
rect 1708 23774 1710 23826
rect 1762 23774 1764 23826
rect 1708 23604 1764 23774
rect 2044 23828 2100 23838
rect 2044 23734 2100 23772
rect 1708 23538 1764 23548
rect 2044 23266 2100 23278
rect 2044 23214 2046 23266
rect 2098 23214 2100 23266
rect 1708 23154 1764 23166
rect 1708 23102 1710 23154
rect 1762 23102 1764 23154
rect 1708 22932 1764 23102
rect 1708 22866 1764 22876
rect 2044 22372 2100 23214
rect 2156 23156 2212 24780
rect 5628 24722 5684 25452
rect 6524 25442 6580 25452
rect 8316 24836 8372 26126
rect 8316 24770 8372 24780
rect 5628 24670 5630 24722
rect 5682 24670 5684 24722
rect 5628 24658 5684 24670
rect 8988 24724 9044 27916
rect 9996 27970 10052 28812
rect 9996 27918 9998 27970
rect 10050 27918 10052 27970
rect 9996 27906 10052 27918
rect 9884 27636 9940 27646
rect 9100 27634 9940 27636
rect 9100 27582 9886 27634
rect 9938 27582 9940 27634
rect 9100 27580 9940 27582
rect 9100 27186 9156 27580
rect 9884 27570 9940 27580
rect 9100 27134 9102 27186
rect 9154 27134 9156 27186
rect 9100 27122 9156 27134
rect 11004 26292 11060 31724
rect 11340 31714 11396 31724
rect 11676 32004 11732 32014
rect 11676 31890 11732 31948
rect 11676 31838 11678 31890
rect 11730 31838 11732 31890
rect 11228 30996 11284 31006
rect 11676 30996 11732 31838
rect 12124 31778 12180 32510
rect 12124 31726 12126 31778
rect 12178 31726 12180 31778
rect 11228 30994 11732 30996
rect 11228 30942 11230 30994
rect 11282 30942 11732 30994
rect 11228 30940 11732 30942
rect 11900 30994 11956 31006
rect 11900 30942 11902 30994
rect 11954 30942 11956 30994
rect 11228 29652 11284 30940
rect 11676 30772 11732 30782
rect 11900 30772 11956 30942
rect 12124 30996 12180 31726
rect 12460 32452 12516 34974
rect 13020 35028 13076 35038
rect 12908 34692 12964 34702
rect 12908 34598 12964 34636
rect 13020 34130 13076 34972
rect 13468 34914 13524 35644
rect 13580 35634 13636 35644
rect 15260 35364 15316 35374
rect 13468 34862 13470 34914
rect 13522 34862 13524 34914
rect 13468 34850 13524 34862
rect 15148 35308 15260 35364
rect 14252 34804 14308 34814
rect 14252 34802 14644 34804
rect 14252 34750 14254 34802
rect 14306 34750 14644 34802
rect 14252 34748 14644 34750
rect 14252 34738 14308 34748
rect 13020 34078 13022 34130
rect 13074 34078 13076 34130
rect 12124 30930 12180 30940
rect 12348 31556 12404 31566
rect 11732 30716 11956 30772
rect 11228 29426 11284 29596
rect 11228 29374 11230 29426
rect 11282 29374 11284 29426
rect 11228 29362 11284 29374
rect 11340 30210 11396 30222
rect 11340 30158 11342 30210
rect 11394 30158 11396 30210
rect 11340 29428 11396 30158
rect 11340 29362 11396 29372
rect 11452 29428 11508 29438
rect 11676 29428 11732 30716
rect 11900 29988 11956 29998
rect 12348 29988 12404 31500
rect 11900 29986 12404 29988
rect 11900 29934 11902 29986
rect 11954 29934 12350 29986
rect 12402 29934 12404 29986
rect 11900 29932 12404 29934
rect 11900 29922 11956 29932
rect 11452 29426 11732 29428
rect 11452 29374 11454 29426
rect 11506 29374 11732 29426
rect 11452 29372 11732 29374
rect 12236 29426 12292 29438
rect 12236 29374 12238 29426
rect 12290 29374 12292 29426
rect 11452 29362 11508 29372
rect 12236 29316 12292 29374
rect 12236 29250 12292 29260
rect 11788 28644 11844 28654
rect 11788 27970 11844 28588
rect 11788 27918 11790 27970
rect 11842 27918 11844 27970
rect 11788 27906 11844 27918
rect 11116 27858 11172 27870
rect 11116 27806 11118 27858
rect 11170 27806 11172 27858
rect 11116 26516 11172 27806
rect 12348 27860 12404 29932
rect 12460 30882 12516 32396
rect 12684 32562 12740 32574
rect 12684 32510 12686 32562
rect 12738 32510 12740 32562
rect 12684 32004 12740 32510
rect 13020 32564 13076 34078
rect 13580 34132 13636 34142
rect 13580 34038 13636 34076
rect 14028 34130 14084 34142
rect 14028 34078 14030 34130
rect 14082 34078 14084 34130
rect 13244 34018 13300 34030
rect 13244 33966 13246 34018
rect 13298 33966 13300 34018
rect 13132 32564 13188 32574
rect 13020 32562 13188 32564
rect 13020 32510 13134 32562
rect 13186 32510 13188 32562
rect 13020 32508 13188 32510
rect 13244 32564 13300 33966
rect 13468 32564 13524 32574
rect 13244 32562 13524 32564
rect 13244 32510 13470 32562
rect 13522 32510 13524 32562
rect 13244 32508 13524 32510
rect 13132 32498 13188 32508
rect 13468 32452 13524 32508
rect 13580 32564 13636 32574
rect 13580 32470 13636 32508
rect 13468 32386 13524 32396
rect 14028 32228 14084 34078
rect 14588 33570 14644 34748
rect 15148 34354 15204 35308
rect 15260 35298 15316 35308
rect 15148 34302 15150 34354
rect 15202 34302 15204 34354
rect 14924 33908 14980 33918
rect 14588 33518 14590 33570
rect 14642 33518 14644 33570
rect 14588 33506 14644 33518
rect 14700 33572 14756 33582
rect 14700 33234 14756 33516
rect 14924 33346 14980 33852
rect 14924 33294 14926 33346
rect 14978 33294 14980 33346
rect 14924 33282 14980 33294
rect 15036 33460 15092 33470
rect 14700 33182 14702 33234
rect 14754 33182 14756 33234
rect 14700 33170 14756 33182
rect 14924 32788 14980 32798
rect 15036 32788 15092 33404
rect 15148 33346 15204 34302
rect 15260 33572 15316 33582
rect 15372 33572 15428 36092
rect 15932 35308 15988 39116
rect 17052 39172 17108 39182
rect 16044 39060 16100 39070
rect 16044 38052 16100 39004
rect 16604 38722 16660 38734
rect 16604 38670 16606 38722
rect 16658 38670 16660 38722
rect 16604 38668 16660 38670
rect 17052 38668 17108 39116
rect 17276 39060 17332 47180
rect 17388 47170 17444 47180
rect 17836 46898 17892 48862
rect 18060 48916 18116 48926
rect 18060 48822 18116 48860
rect 18172 48802 18228 48814
rect 18396 48804 18452 48814
rect 18172 48750 18174 48802
rect 18226 48750 18228 48802
rect 18172 48692 18228 48750
rect 18172 48626 18228 48636
rect 18284 48802 18452 48804
rect 18284 48750 18398 48802
rect 18450 48750 18452 48802
rect 18284 48748 18452 48750
rect 18060 48244 18116 48254
rect 18284 48244 18340 48748
rect 18396 48738 18452 48748
rect 18060 48242 18340 48244
rect 18060 48190 18062 48242
rect 18114 48190 18340 48242
rect 18060 48188 18340 48190
rect 18060 48178 18116 48188
rect 17948 48130 18004 48142
rect 17948 48078 17950 48130
rect 18002 48078 18004 48130
rect 17948 47572 18004 48078
rect 18508 48130 18564 49644
rect 18844 49698 18900 50372
rect 18844 49646 18846 49698
rect 18898 49646 18900 49698
rect 18844 48804 18900 49646
rect 18844 48738 18900 48748
rect 19068 48802 19124 48814
rect 19068 48750 19070 48802
rect 19122 48750 19124 48802
rect 18508 48078 18510 48130
rect 18562 48078 18564 48130
rect 18508 47908 18564 48078
rect 18508 47842 18564 47852
rect 18620 48692 18676 48702
rect 17948 47506 18004 47516
rect 18060 47796 18116 47806
rect 17836 46846 17838 46898
rect 17890 46846 17892 46898
rect 17836 46834 17892 46846
rect 17612 46674 17668 46686
rect 17612 46622 17614 46674
rect 17666 46622 17668 46674
rect 17612 45444 17668 46622
rect 17836 46674 17892 46686
rect 17836 46622 17838 46674
rect 17890 46622 17892 46674
rect 17724 45444 17780 45454
rect 17612 45388 17724 45444
rect 17724 45106 17780 45388
rect 17724 45054 17726 45106
rect 17778 45054 17780 45106
rect 17724 45042 17780 45054
rect 17612 44324 17668 44334
rect 17612 44230 17668 44268
rect 17836 44100 17892 46622
rect 18060 44996 18116 47740
rect 18620 47684 18676 48636
rect 19068 47908 19124 48750
rect 19068 47842 19124 47852
rect 19180 47684 19236 51436
rect 19404 51378 19460 51884
rect 19404 51326 19406 51378
rect 19458 51326 19460 51378
rect 19404 51314 19460 51326
rect 19292 51268 19348 51278
rect 19292 51174 19348 51212
rect 19516 50820 19572 54908
rect 19892 54852 19940 54908
rect 19996 54852 20044 54908
rect 19836 54842 20100 54852
rect 20188 54740 20244 55020
rect 20300 54982 20356 55020
rect 20076 54684 20244 54740
rect 20076 53508 20132 54684
rect 20412 53844 20468 55918
rect 20524 55412 20580 56924
rect 20524 55346 20580 55356
rect 20748 56084 20804 56094
rect 20636 55300 20692 55310
rect 20524 55188 20580 55198
rect 20524 55094 20580 55132
rect 20636 55186 20692 55244
rect 20636 55134 20638 55186
rect 20690 55134 20692 55186
rect 20076 53442 20132 53452
rect 20188 53788 20468 53844
rect 19836 53340 20100 53350
rect 19892 53284 19940 53340
rect 19996 53284 20044 53340
rect 19836 53274 20100 53284
rect 20188 53172 20244 53788
rect 20076 53116 20244 53172
rect 20076 52274 20132 53116
rect 20636 53060 20692 55134
rect 20748 53842 20804 56028
rect 20748 53790 20750 53842
rect 20802 53790 20804 53842
rect 20748 53778 20804 53790
rect 20076 52222 20078 52274
rect 20130 52222 20132 52274
rect 20076 52210 20132 52222
rect 20188 53004 20692 53060
rect 20748 53060 20804 53070
rect 19628 52162 19684 52174
rect 19628 52110 19630 52162
rect 19682 52110 19684 52162
rect 19628 51266 19684 52110
rect 19964 52164 20020 52174
rect 19964 52050 20020 52108
rect 20188 52162 20244 53004
rect 20748 52946 20804 53004
rect 20748 52894 20750 52946
rect 20802 52894 20804 52946
rect 20300 52836 20356 52846
rect 20524 52836 20580 52846
rect 20300 52834 20468 52836
rect 20300 52782 20302 52834
rect 20354 52782 20468 52834
rect 20300 52780 20468 52782
rect 20300 52770 20356 52780
rect 20188 52110 20190 52162
rect 20242 52110 20244 52162
rect 20188 52098 20244 52110
rect 20300 52388 20356 52398
rect 19964 51998 19966 52050
rect 20018 51998 20020 52050
rect 19964 51986 20020 51998
rect 19836 51772 20100 51782
rect 19892 51716 19940 51772
rect 19996 51716 20044 51772
rect 19836 51706 20100 51716
rect 19740 51604 19796 51614
rect 20300 51604 20356 52332
rect 19740 51510 19796 51548
rect 19964 51548 20356 51604
rect 19964 51492 20020 51548
rect 19964 51398 20020 51436
rect 19628 51214 19630 51266
rect 19682 51214 19684 51266
rect 19628 51202 19684 51214
rect 20300 51378 20356 51390
rect 20300 51326 20302 51378
rect 20354 51326 20356 51378
rect 20300 51268 20356 51326
rect 20412 51380 20468 52780
rect 20524 52386 20580 52780
rect 20748 52612 20804 52894
rect 20972 53060 21028 57484
rect 21420 57090 21476 57822
rect 21532 58324 21588 58334
rect 21532 57874 21588 58268
rect 21532 57822 21534 57874
rect 21586 57822 21588 57874
rect 21532 57810 21588 57822
rect 21420 57038 21422 57090
rect 21474 57038 21476 57090
rect 21420 57026 21476 57038
rect 21644 57650 21700 59164
rect 21644 57598 21646 57650
rect 21698 57598 21700 57650
rect 21644 57092 21700 57598
rect 21644 57026 21700 57036
rect 21308 56868 21364 56878
rect 21308 56774 21364 56812
rect 21644 56868 21700 56878
rect 21420 56756 21476 56766
rect 21420 56662 21476 56700
rect 21644 56306 21700 56812
rect 21756 56756 21812 59164
rect 21980 58548 22036 58558
rect 21868 58434 21924 58446
rect 21868 58382 21870 58434
rect 21922 58382 21924 58434
rect 21868 57204 21924 58382
rect 21980 57650 22036 58492
rect 21980 57598 21982 57650
rect 22034 57598 22036 57650
rect 21980 57586 22036 57598
rect 22092 57428 22148 59724
rect 22652 59686 22708 59724
rect 22428 59556 22484 59566
rect 21868 57138 21924 57148
rect 21980 57372 22148 57428
rect 22316 59500 22428 59556
rect 21756 56690 21812 56700
rect 21644 56254 21646 56306
rect 21698 56254 21700 56306
rect 21644 56242 21700 56254
rect 21980 55524 22036 57372
rect 22316 57316 22372 59500
rect 22428 59490 22484 59500
rect 22764 59220 22820 60732
rect 22988 61124 23044 61134
rect 22988 60786 23044 61068
rect 23100 61012 23156 61050
rect 23100 60946 23156 60956
rect 23212 60900 23268 60910
rect 23212 60806 23268 60844
rect 22988 60734 22990 60786
rect 23042 60734 23044 60786
rect 22988 60722 23044 60734
rect 23100 60788 23156 60798
rect 23100 60116 23156 60732
rect 22988 60114 23156 60116
rect 22988 60062 23102 60114
rect 23154 60062 23156 60114
rect 22988 60060 23156 60062
rect 22988 59556 23044 60060
rect 23100 60050 23156 60060
rect 23324 59892 23380 62132
rect 22988 59490 23044 59500
rect 23100 59836 23380 59892
rect 22764 59126 22820 59164
rect 22428 59106 22484 59118
rect 22428 59054 22430 59106
rect 22482 59054 22484 59106
rect 22428 57764 22484 59054
rect 22988 59108 23044 59118
rect 22876 58884 22932 58894
rect 22540 58324 22596 58334
rect 22540 58322 22820 58324
rect 22540 58270 22542 58322
rect 22594 58270 22820 58322
rect 22540 58268 22820 58270
rect 22540 58258 22596 58268
rect 22764 57874 22820 58268
rect 22764 57822 22766 57874
rect 22818 57822 22820 57874
rect 22764 57810 22820 57822
rect 22876 57874 22932 58828
rect 22876 57822 22878 57874
rect 22930 57822 22932 57874
rect 22876 57810 22932 57822
rect 22428 57698 22484 57708
rect 22652 57652 22708 57662
rect 22988 57652 23044 59052
rect 22652 57650 23044 57652
rect 22652 57598 22654 57650
rect 22706 57598 23044 57650
rect 22652 57596 23044 57598
rect 22652 57586 22708 57596
rect 22988 57428 23044 57438
rect 22316 57260 22596 57316
rect 22428 57092 22484 57102
rect 22092 56868 22148 56878
rect 22316 56868 22372 56878
rect 22092 56774 22148 56812
rect 22204 56866 22372 56868
rect 22204 56814 22318 56866
rect 22370 56814 22372 56866
rect 22204 56812 22372 56814
rect 22092 56308 22148 56318
rect 22204 56308 22260 56812
rect 22316 56802 22372 56812
rect 22092 56306 22260 56308
rect 22092 56254 22094 56306
rect 22146 56254 22260 56306
rect 22092 56252 22260 56254
rect 22092 56242 22148 56252
rect 21980 55458 22036 55468
rect 21308 55412 21364 55422
rect 21364 55356 21588 55412
rect 21308 55346 21364 55356
rect 21308 54402 21364 54414
rect 21308 54350 21310 54402
rect 21362 54350 21364 54402
rect 21308 53732 21364 54350
rect 21308 53638 21364 53676
rect 20972 52724 21028 53004
rect 21196 52948 21252 52958
rect 21196 52854 21252 52892
rect 20972 52658 21028 52668
rect 20748 52546 20804 52556
rect 21196 52388 21252 52398
rect 20524 52334 20526 52386
rect 20578 52334 20580 52386
rect 20524 52322 20580 52334
rect 20636 52386 21252 52388
rect 20636 52334 21198 52386
rect 21250 52334 21252 52386
rect 20636 52332 21252 52334
rect 20636 52274 20692 52332
rect 21196 52322 21252 52332
rect 20636 52222 20638 52274
rect 20690 52222 20692 52274
rect 20636 52210 20692 52222
rect 21420 52276 21476 52286
rect 21420 52182 21476 52220
rect 20524 51604 20580 51614
rect 20524 51510 20580 51548
rect 21196 51492 21252 51502
rect 21196 51398 21252 51436
rect 20636 51380 20692 51390
rect 20412 51378 20692 51380
rect 20412 51326 20638 51378
rect 20690 51326 20692 51378
rect 20412 51324 20692 51326
rect 20300 51202 20356 51212
rect 20636 51156 20692 51324
rect 20636 51090 20692 51100
rect 20748 51378 20804 51390
rect 20748 51326 20750 51378
rect 20802 51326 20804 51378
rect 18396 47628 18676 47684
rect 18732 47628 19236 47684
rect 19292 49810 19348 49822
rect 19292 49758 19294 49810
rect 19346 49758 19348 49810
rect 18396 47570 18452 47628
rect 18396 47518 18398 47570
rect 18450 47518 18452 47570
rect 18396 47506 18452 47518
rect 18508 47460 18564 47470
rect 18172 46674 18228 46686
rect 18172 46622 18174 46674
rect 18226 46622 18228 46674
rect 18172 45556 18228 46622
rect 18508 46562 18564 47404
rect 18508 46510 18510 46562
rect 18562 46510 18564 46562
rect 18508 46498 18564 46510
rect 18172 45500 18452 45556
rect 18284 45332 18340 45342
rect 18396 45332 18452 45500
rect 18396 45276 18676 45332
rect 18172 45220 18228 45230
rect 18284 45220 18340 45276
rect 18284 45164 18452 45220
rect 18172 45126 18228 45164
rect 18284 44996 18340 45006
rect 18060 44994 18340 44996
rect 18060 44942 18286 44994
rect 18338 44942 18340 44994
rect 18060 44940 18340 44942
rect 18284 44930 18340 44940
rect 17836 44034 17892 44044
rect 17500 43988 17556 43998
rect 17500 43426 17556 43932
rect 17500 43374 17502 43426
rect 17554 43374 17556 43426
rect 17500 42644 17556 43374
rect 17724 43652 17780 43662
rect 17724 42866 17780 43596
rect 18396 43652 18452 45164
rect 18172 43540 18228 43550
rect 18060 43484 18172 43540
rect 17948 42980 18004 42990
rect 18060 42980 18116 43484
rect 18172 43446 18228 43484
rect 18396 43538 18452 43596
rect 18396 43486 18398 43538
rect 18450 43486 18452 43538
rect 18396 43474 18452 43486
rect 18508 45106 18564 45118
rect 18508 45054 18510 45106
rect 18562 45054 18564 45106
rect 18508 43426 18564 45054
rect 18620 43988 18676 45276
rect 18732 45330 18788 47628
rect 19180 47460 19236 47470
rect 19292 47460 19348 49758
rect 19180 47458 19348 47460
rect 19180 47406 19182 47458
rect 19234 47406 19348 47458
rect 19180 47404 19348 47406
rect 19180 45668 19236 47404
rect 19180 45602 19236 45612
rect 19292 45778 19348 45790
rect 19292 45726 19294 45778
rect 19346 45726 19348 45778
rect 18732 45278 18734 45330
rect 18786 45278 18788 45330
rect 18732 45266 18788 45278
rect 18956 45332 19012 45342
rect 18956 45238 19012 45276
rect 19292 45332 19348 45726
rect 19516 45332 19572 50764
rect 20636 50932 20692 50942
rect 20188 50708 20244 50718
rect 20076 50594 20132 50606
rect 20076 50542 20078 50594
rect 20130 50542 20132 50594
rect 20076 50484 20132 50542
rect 20076 50418 20132 50428
rect 19836 50204 20100 50214
rect 19892 50148 19940 50204
rect 19996 50148 20044 50204
rect 19836 50138 20100 50148
rect 20076 49700 20132 49710
rect 20076 49606 20132 49644
rect 20188 48914 20244 50652
rect 20636 50482 20692 50876
rect 20748 50596 20804 51326
rect 21420 51378 21476 51390
rect 21420 51326 21422 51378
rect 21474 51326 21476 51378
rect 21308 51268 21364 51278
rect 20748 50502 20804 50540
rect 21196 51266 21364 51268
rect 21196 51214 21310 51266
rect 21362 51214 21364 51266
rect 21196 51212 21364 51214
rect 20636 50430 20638 50482
rect 20690 50430 20692 50482
rect 20636 50428 20692 50430
rect 20412 50372 20468 50382
rect 20636 50372 21028 50428
rect 20412 50370 20580 50372
rect 20412 50318 20414 50370
rect 20466 50318 20580 50370
rect 20412 50316 20580 50318
rect 20412 50306 20468 50316
rect 20412 49700 20468 49710
rect 20412 49026 20468 49644
rect 20412 48974 20414 49026
rect 20466 48974 20468 49026
rect 20412 48962 20468 48974
rect 20188 48862 20190 48914
rect 20242 48862 20244 48914
rect 20188 48850 20244 48862
rect 20524 48916 20580 50316
rect 20748 49364 20804 49374
rect 20748 49026 20804 49308
rect 20748 48974 20750 49026
rect 20802 48974 20804 49026
rect 20748 48962 20804 48974
rect 20636 48916 20692 48926
rect 20524 48914 20692 48916
rect 20524 48862 20638 48914
rect 20690 48862 20692 48914
rect 20524 48860 20692 48862
rect 20636 48850 20692 48860
rect 19628 48804 19684 48814
rect 19852 48804 19908 48814
rect 19628 48802 19908 48804
rect 19628 48750 19630 48802
rect 19682 48750 19854 48802
rect 19906 48750 19908 48802
rect 19628 48748 19908 48750
rect 19628 47236 19684 48748
rect 19852 48738 19908 48748
rect 19836 48636 20100 48646
rect 19892 48580 19940 48636
rect 19996 48580 20044 48636
rect 19836 48570 20100 48580
rect 20972 48468 21028 50372
rect 21196 49364 21252 51212
rect 21308 51202 21364 51212
rect 21420 51044 21476 51326
rect 21420 50978 21476 50988
rect 21420 50820 21476 50830
rect 21420 50484 21476 50764
rect 21308 50428 21476 50484
rect 21308 50370 21364 50428
rect 21308 50318 21310 50370
rect 21362 50318 21364 50370
rect 21308 50306 21364 50318
rect 21532 49364 21588 55356
rect 22092 53844 22148 53854
rect 22092 53750 22148 53788
rect 21868 53508 21924 53518
rect 21644 52946 21700 52958
rect 21644 52894 21646 52946
rect 21698 52894 21700 52946
rect 21644 52164 21700 52894
rect 21868 52948 21924 53452
rect 22204 52948 22260 56252
rect 22316 56194 22372 56206
rect 22316 56142 22318 56194
rect 22370 56142 22372 56194
rect 22316 55300 22372 56142
rect 22316 55234 22372 55244
rect 21868 52946 22036 52948
rect 21868 52894 21870 52946
rect 21922 52894 22036 52946
rect 21868 52892 22036 52894
rect 21868 52882 21924 52892
rect 21756 52834 21812 52846
rect 21756 52782 21758 52834
rect 21810 52782 21812 52834
rect 21756 52386 21812 52782
rect 21756 52334 21758 52386
rect 21810 52334 21812 52386
rect 21756 52322 21812 52334
rect 21868 52724 21924 52734
rect 21868 52164 21924 52668
rect 21644 52098 21700 52108
rect 21756 52108 21924 52164
rect 21756 50428 21812 52108
rect 21868 51380 21924 51390
rect 21868 51286 21924 51324
rect 21980 51156 22036 52892
rect 22204 52882 22260 52892
rect 22428 52274 22484 57036
rect 22540 56532 22596 57260
rect 22988 57090 23044 57372
rect 22988 57038 22990 57090
rect 23042 57038 23044 57090
rect 22988 57026 23044 57038
rect 22876 56868 22932 56878
rect 22652 56756 22708 56766
rect 22652 56662 22708 56700
rect 22876 56754 22932 56812
rect 22876 56702 22878 56754
rect 22930 56702 22932 56754
rect 22876 56690 22932 56702
rect 23100 56756 23156 59836
rect 23324 58996 23380 59006
rect 23212 57988 23268 57998
rect 23212 56866 23268 57932
rect 23324 57650 23380 58940
rect 23548 57762 23604 62132
rect 23772 61012 23828 63870
rect 23884 63922 24276 63924
rect 23884 63870 24222 63922
rect 24274 63870 24276 63922
rect 23884 63868 24276 63870
rect 23884 61124 23940 63868
rect 24220 63858 24276 63868
rect 24444 63924 24500 63934
rect 24444 63922 24612 63924
rect 24444 63870 24446 63922
rect 24498 63870 24612 63922
rect 24444 63868 24612 63870
rect 24444 63858 24500 63868
rect 24332 63812 24388 63822
rect 24332 63718 24388 63756
rect 24556 63476 24612 63868
rect 23884 61058 23940 61068
rect 23996 63420 24612 63476
rect 23772 60946 23828 60956
rect 23996 60900 24052 63420
rect 24556 63362 24612 63420
rect 24556 63310 24558 63362
rect 24610 63310 24612 63362
rect 24556 63298 24612 63310
rect 24220 63250 24276 63262
rect 24220 63198 24222 63250
rect 24274 63198 24276 63250
rect 24220 62916 24276 63198
rect 24220 62850 24276 62860
rect 24332 63140 24388 63150
rect 24220 62578 24276 62590
rect 24220 62526 24222 62578
rect 24274 62526 24276 62578
rect 24220 62354 24276 62526
rect 24220 62302 24222 62354
rect 24274 62302 24276 62354
rect 24220 62188 24276 62302
rect 23996 60834 24052 60844
rect 24108 62132 24276 62188
rect 23996 60674 24052 60686
rect 23996 60622 23998 60674
rect 24050 60622 24052 60674
rect 23660 60004 23716 60014
rect 23884 60004 23940 60014
rect 23660 60002 23884 60004
rect 23660 59950 23662 60002
rect 23714 59950 23884 60002
rect 23660 59948 23884 59950
rect 23660 59938 23716 59948
rect 23884 59910 23940 59948
rect 23996 59780 24052 60622
rect 23996 59714 24052 59724
rect 23996 59444 24052 59454
rect 23884 59388 23996 59444
rect 23660 59108 23716 59118
rect 23660 59106 23828 59108
rect 23660 59054 23662 59106
rect 23714 59054 23828 59106
rect 23660 59052 23828 59054
rect 23660 59042 23716 59052
rect 23772 58772 23828 59052
rect 23772 58706 23828 58716
rect 23548 57710 23550 57762
rect 23602 57710 23604 57762
rect 23548 57698 23604 57710
rect 23772 57876 23828 57886
rect 23324 57598 23326 57650
rect 23378 57598 23380 57650
rect 23324 57586 23380 57598
rect 23436 57652 23492 57662
rect 23212 56814 23214 56866
rect 23266 56814 23268 56866
rect 23212 56802 23268 56814
rect 23100 56690 23156 56700
rect 22540 56476 22708 56532
rect 22540 56084 22596 56094
rect 22540 55990 22596 56028
rect 22428 52222 22430 52274
rect 22482 52222 22484 52274
rect 22428 52210 22484 52222
rect 22204 52162 22260 52174
rect 22204 52110 22206 52162
rect 22258 52110 22260 52162
rect 22092 51604 22148 51614
rect 22092 51378 22148 51548
rect 22092 51326 22094 51378
rect 22146 51326 22148 51378
rect 22092 51314 22148 51326
rect 22204 51380 22260 52110
rect 22652 51604 22708 56476
rect 23100 55970 23156 55982
rect 23100 55918 23102 55970
rect 23154 55918 23156 55970
rect 22988 55300 23044 55310
rect 22988 53172 23044 55244
rect 23100 55188 23156 55918
rect 23436 55188 23492 57596
rect 23660 57428 23716 57438
rect 23548 57316 23604 57326
rect 23548 56866 23604 57260
rect 23660 56978 23716 57372
rect 23660 56926 23662 56978
rect 23714 56926 23716 56978
rect 23660 56914 23716 56926
rect 23548 56814 23550 56866
rect 23602 56814 23604 56866
rect 23548 56802 23604 56814
rect 23772 56866 23828 57820
rect 23884 57092 23940 59388
rect 23996 59378 24052 59388
rect 24108 59442 24164 62132
rect 24108 59390 24110 59442
rect 24162 59390 24164 59442
rect 23884 57026 23940 57036
rect 23996 57650 24052 57662
rect 23996 57598 23998 57650
rect 24050 57598 24052 57650
rect 23772 56814 23774 56866
rect 23826 56814 23828 56866
rect 23772 56802 23828 56814
rect 23996 56532 24052 57598
rect 24108 57652 24164 59390
rect 24220 61796 24276 61806
rect 24220 61682 24276 61740
rect 24220 61630 24222 61682
rect 24274 61630 24276 61682
rect 24220 59220 24276 61630
rect 24332 61572 24388 63084
rect 24556 62580 24612 62590
rect 24668 62580 24724 64988
rect 25004 63138 25060 65660
rect 25452 65660 25620 65716
rect 25788 65716 25844 65726
rect 25340 65604 25396 65614
rect 25228 65490 25284 65502
rect 25228 65438 25230 65490
rect 25282 65438 25284 65490
rect 25228 65380 25284 65438
rect 25228 65314 25284 65324
rect 25340 65156 25396 65548
rect 25228 65100 25396 65156
rect 25116 63700 25172 63710
rect 25116 63250 25172 63644
rect 25228 63588 25284 65100
rect 25452 63922 25508 65660
rect 25452 63870 25454 63922
rect 25506 63870 25508 63922
rect 25452 63858 25508 63870
rect 25564 65490 25620 65502
rect 25564 65438 25566 65490
rect 25618 65438 25620 65490
rect 25564 63812 25620 65438
rect 25228 63532 25508 63588
rect 25116 63198 25118 63250
rect 25170 63198 25172 63250
rect 25116 63186 25172 63198
rect 25228 63364 25284 63374
rect 25004 63086 25006 63138
rect 25058 63086 25060 63138
rect 25004 63074 25060 63086
rect 25228 63138 25284 63308
rect 25228 63086 25230 63138
rect 25282 63086 25284 63138
rect 24556 62578 24724 62580
rect 24556 62526 24558 62578
rect 24610 62526 24670 62578
rect 24722 62526 24724 62578
rect 24556 62524 24724 62526
rect 24556 62514 24612 62524
rect 24668 62514 24724 62524
rect 24780 62916 24836 62926
rect 24556 61572 24612 61582
rect 24332 61570 24612 61572
rect 24332 61518 24558 61570
rect 24610 61518 24612 61570
rect 24332 61516 24612 61518
rect 24556 61506 24612 61516
rect 24668 61012 24724 61022
rect 24780 61012 24836 62860
rect 25228 62188 25284 63086
rect 25116 62132 25284 62188
rect 25340 62242 25396 62254
rect 25340 62190 25342 62242
rect 25394 62190 25396 62242
rect 25116 61682 25172 62132
rect 25340 61796 25396 62190
rect 25340 61730 25396 61740
rect 25116 61630 25118 61682
rect 25170 61630 25172 61682
rect 25116 61618 25172 61630
rect 24668 61010 24836 61012
rect 24668 60958 24670 61010
rect 24722 60958 24836 61010
rect 24668 60956 24836 60958
rect 25340 61570 25396 61582
rect 25340 61518 25342 61570
rect 25394 61518 25396 61570
rect 24668 60946 24724 60956
rect 25340 60900 25396 61518
rect 25340 60834 25396 60844
rect 24332 60786 24388 60798
rect 24332 60734 24334 60786
rect 24386 60734 24388 60786
rect 24332 60114 24388 60734
rect 24332 60062 24334 60114
rect 24386 60062 24388 60114
rect 24332 59780 24388 60062
rect 25228 60674 25284 60686
rect 25228 60622 25230 60674
rect 25282 60622 25284 60674
rect 25228 60564 25284 60622
rect 24892 60004 24948 60014
rect 24332 59714 24388 59724
rect 24780 59948 24892 60004
rect 24556 59444 24612 59454
rect 24556 59350 24612 59388
rect 24444 59220 24500 59230
rect 24220 59164 24444 59220
rect 24108 57586 24164 57596
rect 24220 58772 24276 58782
rect 24220 56868 24276 58716
rect 24444 56980 24500 59164
rect 24668 59218 24724 59230
rect 24668 59166 24670 59218
rect 24722 59166 24724 59218
rect 24556 58996 24612 59006
rect 24556 58902 24612 58940
rect 24668 58772 24724 59166
rect 24668 58706 24724 58716
rect 24668 58546 24724 58558
rect 24668 58494 24670 58546
rect 24722 58494 24724 58546
rect 24668 58436 24724 58494
rect 24556 57876 24612 57886
rect 24556 57782 24612 57820
rect 24668 57650 24724 58380
rect 24668 57598 24670 57650
rect 24722 57598 24724 57650
rect 24668 57586 24724 57598
rect 24668 57092 24724 57102
rect 24444 56924 24612 56980
rect 23548 56194 23604 56206
rect 23548 56142 23550 56194
rect 23602 56142 23604 56194
rect 23548 56084 23604 56142
rect 23548 56018 23604 56028
rect 23996 56082 24052 56476
rect 23996 56030 23998 56082
rect 24050 56030 24052 56082
rect 23996 56018 24052 56030
rect 24108 56812 24220 56868
rect 23100 55186 23492 55188
rect 23100 55134 23438 55186
rect 23490 55134 23492 55186
rect 23100 55132 23492 55134
rect 23436 54514 23492 55132
rect 23436 54462 23438 54514
rect 23490 54462 23492 54514
rect 22988 53078 23044 53116
rect 23324 53732 23380 53742
rect 23324 53170 23380 53676
rect 23324 53118 23326 53170
rect 23378 53118 23380 53170
rect 23324 53106 23380 53118
rect 23212 53058 23268 53070
rect 23212 53006 23214 53058
rect 23266 53006 23268 53058
rect 22764 52948 22820 52958
rect 22764 52276 22820 52892
rect 22764 52210 22820 52220
rect 23212 52948 23268 53006
rect 22652 51538 22708 51548
rect 22876 52162 22932 52174
rect 22876 52110 22878 52162
rect 22930 52110 22932 52162
rect 22876 51492 22932 52110
rect 23100 52052 23156 52062
rect 23100 51958 23156 51996
rect 23212 51828 23268 52892
rect 23436 52500 23492 54462
rect 24108 53284 24164 56812
rect 24220 56774 24276 56812
rect 24332 56756 24388 56766
rect 24332 56662 24388 56700
rect 24444 56754 24500 56766
rect 24444 56702 24446 56754
rect 24498 56702 24500 56754
rect 24444 56644 24500 56702
rect 24444 56578 24500 56588
rect 24444 56308 24500 56318
rect 24444 56214 24500 56252
rect 24332 56084 24388 56094
rect 24556 56084 24612 56924
rect 24220 56082 24388 56084
rect 24220 56030 24334 56082
rect 24386 56030 24388 56082
rect 24220 56028 24388 56030
rect 24220 54740 24276 56028
rect 24332 56018 24388 56028
rect 24444 56028 24612 56084
rect 24444 54740 24500 56028
rect 24220 53842 24276 54684
rect 24220 53790 24222 53842
rect 24274 53790 24276 53842
rect 24220 53778 24276 53790
rect 24332 54684 24500 54740
rect 24556 54740 24612 54750
rect 24668 54740 24724 57036
rect 24556 54738 24724 54740
rect 24556 54686 24558 54738
rect 24610 54686 24724 54738
rect 24556 54684 24724 54686
rect 24780 54740 24836 59948
rect 24892 59938 24948 59948
rect 25228 59778 25284 60508
rect 25228 59726 25230 59778
rect 25282 59726 25284 59778
rect 25228 59220 25284 59726
rect 25452 59556 25508 63532
rect 25564 63364 25620 63756
rect 25564 63298 25620 63308
rect 25676 65378 25732 65390
rect 25676 65326 25678 65378
rect 25730 65326 25732 65378
rect 25564 63140 25620 63150
rect 25676 63140 25732 65326
rect 25788 64484 25844 65660
rect 25900 65604 25956 66220
rect 25900 65538 25956 65548
rect 26012 65380 26068 66892
rect 26124 66882 26180 66892
rect 26460 66946 26516 66958
rect 26460 66894 26462 66946
rect 26514 66894 26516 66946
rect 26460 66834 26516 66894
rect 26460 66782 26462 66834
rect 26514 66782 26516 66834
rect 26460 66770 26516 66782
rect 27020 66946 27076 66958
rect 27020 66894 27022 66946
rect 27074 66894 27076 66946
rect 26124 66500 26180 66510
rect 27020 66500 27076 66894
rect 26124 66498 26740 66500
rect 26124 66446 26126 66498
rect 26178 66446 26740 66498
rect 26124 66444 26740 66446
rect 26124 66434 26180 66444
rect 26236 66276 26292 66286
rect 26236 66182 26292 66220
rect 26124 66164 26180 66174
rect 26124 66070 26180 66108
rect 26012 65314 26068 65324
rect 26124 65716 26180 65726
rect 26124 65378 26180 65660
rect 26572 65492 26628 65502
rect 26572 65398 26628 65436
rect 26124 65326 26126 65378
rect 26178 65326 26180 65378
rect 26124 65156 26180 65326
rect 26236 65380 26292 65390
rect 26236 65378 26516 65380
rect 26236 65326 26238 65378
rect 26290 65326 26516 65378
rect 26236 65324 26516 65326
rect 26236 65314 26292 65324
rect 26124 65100 26292 65156
rect 25900 64818 25956 64830
rect 25900 64766 25902 64818
rect 25954 64766 25956 64818
rect 25900 64708 25956 64766
rect 26236 64708 26292 65100
rect 26460 64932 26516 65324
rect 26572 64932 26628 64942
rect 26460 64930 26628 64932
rect 26460 64878 26574 64930
rect 26626 64878 26628 64930
rect 26460 64876 26628 64878
rect 25900 64652 26292 64708
rect 25788 64428 26180 64484
rect 26124 64146 26180 64428
rect 26124 64094 26126 64146
rect 26178 64094 26180 64146
rect 26124 64082 26180 64094
rect 25900 63922 25956 63934
rect 25900 63870 25902 63922
rect 25954 63870 25956 63922
rect 25900 63812 25956 63870
rect 26012 63924 26068 63934
rect 26012 63830 26068 63868
rect 25900 63746 25956 63756
rect 26236 63588 26292 64652
rect 25564 63138 25732 63140
rect 25564 63086 25566 63138
rect 25618 63086 25732 63138
rect 25564 63084 25732 63086
rect 25900 63532 26292 63588
rect 26348 64482 26404 64494
rect 26348 64430 26350 64482
rect 26402 64430 26404 64482
rect 26348 64372 26404 64430
rect 26460 64484 26516 64494
rect 26460 64390 26516 64428
rect 25564 63074 25620 63084
rect 25676 61458 25732 61470
rect 25676 61406 25678 61458
rect 25730 61406 25732 61458
rect 25676 61124 25732 61406
rect 25676 61058 25732 61068
rect 25452 59490 25508 59500
rect 25788 59778 25844 59790
rect 25788 59726 25790 59778
rect 25842 59726 25844 59778
rect 25788 59332 25844 59726
rect 25788 59266 25844 59276
rect 25116 59164 25284 59220
rect 24892 58434 24948 58446
rect 24892 58382 24894 58434
rect 24946 58382 24948 58434
rect 24892 57540 24948 58382
rect 24892 57474 24948 57484
rect 24892 57316 24948 57326
rect 24892 57090 24948 57260
rect 24892 57038 24894 57090
rect 24946 57038 24948 57090
rect 24892 57026 24948 57038
rect 25116 55468 25172 59164
rect 25228 58994 25284 59006
rect 25228 58942 25230 58994
rect 25282 58942 25284 58994
rect 25228 58884 25284 58942
rect 25228 58818 25284 58828
rect 25340 58994 25396 59006
rect 25564 58996 25620 59006
rect 25340 58942 25342 58994
rect 25394 58942 25396 58994
rect 25340 57988 25396 58942
rect 25340 57922 25396 57932
rect 25452 58994 25620 58996
rect 25452 58942 25566 58994
rect 25618 58942 25620 58994
rect 25452 58940 25620 58942
rect 25228 57652 25284 57662
rect 25228 57558 25284 57596
rect 25452 57316 25508 58940
rect 25564 58930 25620 58940
rect 25676 58996 25732 59006
rect 25900 58996 25956 63532
rect 26012 62916 26068 62926
rect 26348 62916 26404 64316
rect 26460 64260 26516 64270
rect 26460 63924 26516 64204
rect 26572 64146 26628 64876
rect 26572 64094 26574 64146
rect 26626 64094 26628 64146
rect 26572 64082 26628 64094
rect 26684 64034 26740 66444
rect 27020 66434 27076 66444
rect 27804 66276 27860 66286
rect 28140 66276 28196 67116
rect 28364 67106 28420 67116
rect 28588 67618 28644 67630
rect 28588 67566 28590 67618
rect 28642 67566 28644 67618
rect 28588 67060 28644 67566
rect 29708 67508 29764 67518
rect 29260 67284 29316 67294
rect 29148 67172 29204 67182
rect 29148 67078 29204 67116
rect 28588 66994 28644 67004
rect 28700 66946 28756 66958
rect 28700 66894 28702 66946
rect 28754 66894 28756 66946
rect 27804 66182 27860 66220
rect 28028 66274 28196 66276
rect 28028 66222 28142 66274
rect 28194 66222 28196 66274
rect 28028 66220 28196 66222
rect 26908 66052 26964 66062
rect 26908 64930 26964 65996
rect 26908 64878 26910 64930
rect 26962 64878 26964 64930
rect 26908 64866 26964 64878
rect 27020 66050 27076 66062
rect 27020 65998 27022 66050
rect 27074 65998 27076 66050
rect 27020 64148 27076 65998
rect 27244 66052 27300 66062
rect 27244 65958 27300 65996
rect 27356 66050 27412 66062
rect 27356 65998 27358 66050
rect 27410 65998 27412 66050
rect 27356 65602 27412 65998
rect 27356 65550 27358 65602
rect 27410 65550 27412 65602
rect 27356 65538 27412 65550
rect 27468 66050 27524 66062
rect 27916 66052 27972 66062
rect 27468 65998 27470 66050
rect 27522 65998 27524 66050
rect 27468 65492 27524 65998
rect 27468 65426 27524 65436
rect 27580 66050 27972 66052
rect 27580 65998 27918 66050
rect 27970 65998 27972 66050
rect 27580 65996 27972 65998
rect 27244 64706 27300 64718
rect 27244 64654 27246 64706
rect 27298 64654 27300 64706
rect 27244 64372 27300 64654
rect 27468 64708 27524 64718
rect 27244 64306 27300 64316
rect 27356 64596 27412 64606
rect 27356 64260 27412 64540
rect 27356 64194 27412 64204
rect 27020 64082 27076 64092
rect 26684 63982 26686 64034
rect 26738 63982 26740 64034
rect 26684 63970 26740 63982
rect 27468 63924 27524 64652
rect 26460 63868 26628 63924
rect 26572 63698 26628 63868
rect 27468 63858 27524 63868
rect 27580 63810 27636 65996
rect 27916 65986 27972 65996
rect 27804 64706 27860 64718
rect 27804 64654 27806 64706
rect 27858 64654 27860 64706
rect 27804 64596 27860 64654
rect 28028 64706 28084 66220
rect 28140 66210 28196 66220
rect 28252 66276 28308 66286
rect 28028 64654 28030 64706
rect 28082 64654 28084 64706
rect 28028 64642 28084 64654
rect 27804 64530 27860 64540
rect 28140 64594 28196 64606
rect 28140 64542 28142 64594
rect 28194 64542 28196 64594
rect 28140 64148 28196 64542
rect 27580 63758 27582 63810
rect 27634 63758 27636 63810
rect 27580 63746 27636 63758
rect 27692 64092 28196 64148
rect 27692 63922 27748 64092
rect 27692 63870 27694 63922
rect 27746 63870 27748 63922
rect 26572 63646 26574 63698
rect 26626 63646 26628 63698
rect 26572 63634 26628 63646
rect 27692 63588 27748 63870
rect 28140 63812 28196 63822
rect 27804 63700 27860 63710
rect 28028 63700 28084 63710
rect 27804 63698 28084 63700
rect 27804 63646 27806 63698
rect 27858 63646 28030 63698
rect 28082 63646 28084 63698
rect 27804 63644 28084 63646
rect 27804 63634 27860 63644
rect 28028 63634 28084 63644
rect 27356 63532 27748 63588
rect 26068 62860 26404 62916
rect 27132 63028 27188 63038
rect 26012 62822 26068 62860
rect 26012 62242 26068 62254
rect 26012 62190 26014 62242
rect 26066 62190 26068 62242
rect 26012 62020 26068 62190
rect 26572 62132 26628 62142
rect 26012 61460 26068 61964
rect 26348 62076 26572 62132
rect 26236 61460 26292 61470
rect 26012 61458 26292 61460
rect 26012 61406 26238 61458
rect 26290 61406 26292 61458
rect 26012 61404 26292 61406
rect 26236 60564 26292 61404
rect 26348 61460 26404 62076
rect 26572 62066 26628 62076
rect 27132 62130 27188 62972
rect 27356 62188 27412 63532
rect 28140 62466 28196 63756
rect 28252 62916 28308 66220
rect 28700 66276 28756 66894
rect 28700 66210 28756 66220
rect 29260 66276 29316 67228
rect 29484 67284 29540 67294
rect 29484 67170 29540 67228
rect 29484 67118 29486 67170
rect 29538 67118 29540 67170
rect 29484 67106 29540 67118
rect 29708 67170 29764 67452
rect 29708 67118 29710 67170
rect 29762 67118 29764 67170
rect 29708 67106 29764 67118
rect 29260 66210 29316 66220
rect 28364 66162 28420 66174
rect 28364 66110 28366 66162
rect 28418 66110 28420 66162
rect 28364 65380 28420 66110
rect 28364 65314 28420 65324
rect 29260 66052 29316 66062
rect 28588 64596 28644 64606
rect 29148 64596 29204 64606
rect 28364 64594 29204 64596
rect 28364 64542 28590 64594
rect 28642 64542 29150 64594
rect 29202 64542 29204 64594
rect 28364 64540 29204 64542
rect 28364 63922 28420 64540
rect 28588 64530 28644 64540
rect 29148 64530 29204 64540
rect 28588 64372 28644 64382
rect 28364 63870 28366 63922
rect 28418 63870 28420 63922
rect 28364 63858 28420 63870
rect 28476 64316 28588 64372
rect 28364 63700 28420 63710
rect 28476 63700 28532 64316
rect 28588 64306 28644 64316
rect 28924 64260 28980 64270
rect 28588 64148 28644 64158
rect 28588 64054 28644 64092
rect 28812 64036 28868 64046
rect 28364 63698 28532 63700
rect 28364 63646 28366 63698
rect 28418 63646 28532 63698
rect 28364 63644 28532 63646
rect 28700 64034 28868 64036
rect 28700 63982 28814 64034
rect 28866 63982 28868 64034
rect 28700 63980 28868 63982
rect 28364 63634 28420 63644
rect 28476 62916 28532 62926
rect 28252 62914 28532 62916
rect 28252 62862 28478 62914
rect 28530 62862 28532 62914
rect 28252 62860 28532 62862
rect 28140 62414 28142 62466
rect 28194 62414 28196 62466
rect 28140 62402 28196 62414
rect 28252 62466 28308 62478
rect 28252 62414 28254 62466
rect 28306 62414 28308 62466
rect 27132 62078 27134 62130
rect 27186 62078 27188 62130
rect 26348 61458 26516 61460
rect 26348 61406 26350 61458
rect 26402 61406 26516 61458
rect 26348 61404 26516 61406
rect 26348 61394 26404 61404
rect 26236 60498 26292 60508
rect 26348 61124 26404 61134
rect 26012 60340 26068 60350
rect 26012 60002 26068 60284
rect 26236 60228 26292 60238
rect 26236 60134 26292 60172
rect 26012 59950 26014 60002
rect 26066 59950 26068 60002
rect 26012 59892 26068 59950
rect 26012 59220 26068 59836
rect 26236 59332 26292 59342
rect 26236 59238 26292 59276
rect 26012 59154 26068 59164
rect 26124 59218 26180 59230
rect 26124 59166 26126 59218
rect 26178 59166 26180 59218
rect 25676 58994 25844 58996
rect 25676 58942 25678 58994
rect 25730 58942 25844 58994
rect 25676 58940 25844 58942
rect 25900 58940 26068 58996
rect 25676 58930 25732 58940
rect 25788 58546 25844 58940
rect 25788 58494 25790 58546
rect 25842 58494 25844 58546
rect 25676 58434 25732 58446
rect 25676 58382 25678 58434
rect 25730 58382 25732 58434
rect 25676 57988 25732 58382
rect 25676 57922 25732 57932
rect 25788 57876 25844 58494
rect 25788 57810 25844 57820
rect 25452 57250 25508 57260
rect 25676 57204 25732 57214
rect 25676 56866 25732 57148
rect 25676 56814 25678 56866
rect 25730 56814 25732 56866
rect 25676 56802 25732 56814
rect 25340 56644 25396 56654
rect 25396 56588 25620 56644
rect 25340 56550 25396 56588
rect 25004 55412 25172 55468
rect 25228 56308 25284 56318
rect 24780 54684 24948 54740
rect 23884 53228 24164 53284
rect 23884 52724 23940 53228
rect 24220 53172 24276 53182
rect 24108 53116 24220 53172
rect 24108 53058 24164 53116
rect 24220 53106 24276 53116
rect 24108 53006 24110 53058
rect 24162 53006 24164 53058
rect 24108 52994 24164 53006
rect 23996 52948 24052 52958
rect 23996 52854 24052 52892
rect 24220 52946 24276 52958
rect 24220 52894 24222 52946
rect 24274 52894 24276 52946
rect 24220 52724 24276 52894
rect 23884 52668 24164 52724
rect 23996 52500 24052 52510
rect 23436 52444 23716 52500
rect 23548 52276 23604 52286
rect 23548 52182 23604 52220
rect 22876 51398 22932 51436
rect 23100 51772 23268 51828
rect 23436 52052 23492 52062
rect 22540 51380 22596 51390
rect 22204 51378 22596 51380
rect 22204 51326 22542 51378
rect 22594 51326 22596 51378
rect 22204 51324 22596 51326
rect 22204 51156 22260 51166
rect 21980 51100 22204 51156
rect 21196 49298 21252 49308
rect 21308 49308 21588 49364
rect 21644 50372 21812 50428
rect 22092 50596 22148 50606
rect 22092 50482 22148 50540
rect 22204 50594 22260 51100
rect 22204 50542 22206 50594
rect 22258 50542 22260 50594
rect 22204 50530 22260 50542
rect 22316 50820 22372 50830
rect 22540 50820 22596 51324
rect 22764 50820 22820 50830
rect 22540 50818 22820 50820
rect 22540 50766 22766 50818
rect 22818 50766 22820 50818
rect 22540 50764 22820 50766
rect 22316 50594 22372 50764
rect 22764 50754 22820 50764
rect 22316 50542 22318 50594
rect 22370 50542 22372 50594
rect 22316 50530 22372 50542
rect 22092 50430 22094 50482
rect 22146 50430 22148 50482
rect 22092 50428 22148 50430
rect 23100 50428 23156 51772
rect 23212 51492 23268 51502
rect 23212 51398 23268 51436
rect 23324 51380 23380 51390
rect 23324 51286 23380 51324
rect 23436 51378 23492 51996
rect 23436 51326 23438 51378
rect 23490 51326 23492 51378
rect 23436 51044 23492 51326
rect 23436 50978 23492 50988
rect 23324 50820 23380 50830
rect 23324 50706 23380 50764
rect 23324 50654 23326 50706
rect 23378 50654 23380 50706
rect 23324 50642 23380 50654
rect 23660 50484 23716 52444
rect 23996 52050 24052 52444
rect 23996 51998 23998 52050
rect 24050 51998 24052 52050
rect 23996 51986 24052 51998
rect 23772 51604 23828 51614
rect 23772 51380 23828 51548
rect 23772 51286 23828 51324
rect 23716 50428 23940 50484
rect 24108 50428 24164 52668
rect 24332 52724 24388 54684
rect 24556 54674 24612 54684
rect 24892 54628 24948 54684
rect 24444 54516 24500 54526
rect 24556 54516 24612 54526
rect 24444 54514 24556 54516
rect 24444 54462 24446 54514
rect 24498 54462 24556 54514
rect 24444 54460 24556 54462
rect 24444 54450 24500 54460
rect 24444 53732 24500 53742
rect 24444 53638 24500 53676
rect 24444 52948 24500 52958
rect 24556 52948 24612 54460
rect 24780 54514 24836 54526
rect 24780 54462 24782 54514
rect 24834 54462 24836 54514
rect 24668 54292 24724 54302
rect 24668 53170 24724 54236
rect 24780 53956 24836 54462
rect 24780 53890 24836 53900
rect 24668 53118 24670 53170
rect 24722 53118 24724 53170
rect 24668 53106 24724 53118
rect 24500 52892 24612 52948
rect 24444 52882 24500 52892
rect 24332 52668 24500 52724
rect 24220 52658 24276 52668
rect 24220 52164 24276 52174
rect 24220 52070 24276 52108
rect 24220 51380 24276 51390
rect 24220 51286 24276 51324
rect 22092 50372 22260 50428
rect 23100 50372 23380 50428
rect 23660 50390 23716 50428
rect 21644 50370 21700 50372
rect 21644 50318 21646 50370
rect 21698 50318 21700 50370
rect 21308 48916 21364 49308
rect 21420 49140 21476 49150
rect 21644 49140 21700 50318
rect 21420 49138 21700 49140
rect 21420 49086 21422 49138
rect 21474 49086 21700 49138
rect 21420 49084 21700 49086
rect 22204 49698 22260 50372
rect 22204 49646 22206 49698
rect 22258 49646 22260 49698
rect 21420 49074 21476 49084
rect 20860 48412 21028 48468
rect 21084 48860 21364 48916
rect 19628 47170 19684 47180
rect 20076 47348 20132 47358
rect 20076 47236 20132 47292
rect 20076 47234 20244 47236
rect 20076 47182 20078 47234
rect 20130 47182 20244 47234
rect 20076 47180 20244 47182
rect 20076 47170 20132 47180
rect 19836 47068 20100 47078
rect 19892 47012 19940 47068
rect 19996 47012 20044 47068
rect 19836 47002 20100 47012
rect 20076 45890 20132 45902
rect 20076 45838 20078 45890
rect 20130 45838 20132 45890
rect 20076 45668 20132 45838
rect 20188 45668 20244 47180
rect 20524 47234 20580 47246
rect 20524 47182 20526 47234
rect 20578 47182 20580 47234
rect 20524 47068 20580 47182
rect 20860 47068 20916 48412
rect 20972 48242 21028 48254
rect 20972 48190 20974 48242
rect 21026 48190 21028 48242
rect 20972 48132 21028 48190
rect 21084 48244 21140 48860
rect 21196 48468 21252 48478
rect 21196 48466 21700 48468
rect 21196 48414 21198 48466
rect 21250 48414 21700 48466
rect 21196 48412 21700 48414
rect 21196 48402 21252 48412
rect 21308 48244 21364 48254
rect 21084 48242 21364 48244
rect 21084 48190 21310 48242
rect 21362 48190 21364 48242
rect 21084 48188 21364 48190
rect 21308 48178 21364 48188
rect 21532 48244 21588 48254
rect 21532 48150 21588 48188
rect 20972 47348 21028 48076
rect 20972 47282 21028 47292
rect 21084 47684 21140 47694
rect 20524 47012 20804 47068
rect 20860 47012 21028 47068
rect 20636 46564 20692 46574
rect 20636 46470 20692 46508
rect 20748 46004 20804 47012
rect 20748 45780 20804 45948
rect 20748 45778 20916 45780
rect 20748 45726 20750 45778
rect 20802 45726 20916 45778
rect 20748 45724 20916 45726
rect 20748 45714 20804 45724
rect 20524 45668 20580 45678
rect 20188 45666 20580 45668
rect 20188 45614 20526 45666
rect 20578 45614 20580 45666
rect 20188 45612 20580 45614
rect 20076 45602 20132 45612
rect 19836 45500 20100 45510
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 19836 45434 20100 45444
rect 19516 45276 19908 45332
rect 19292 45266 19348 45276
rect 18844 45220 18900 45230
rect 18620 43922 18676 43932
rect 18732 44100 18788 44110
rect 18508 43374 18510 43426
rect 18562 43374 18564 43426
rect 17948 42978 18116 42980
rect 17948 42926 17950 42978
rect 18002 42926 18116 42978
rect 17948 42924 18116 42926
rect 18172 43316 18228 43326
rect 18508 43316 18564 43374
rect 18228 43260 18564 43316
rect 18172 42978 18228 43260
rect 18172 42926 18174 42978
rect 18226 42926 18228 42978
rect 17948 42914 18004 42924
rect 18172 42914 18228 42926
rect 17724 42814 17726 42866
rect 17778 42814 17780 42866
rect 17724 42802 17780 42814
rect 17500 42588 18228 42644
rect 17836 42084 17892 42094
rect 17836 40740 17892 42028
rect 17836 40402 17892 40684
rect 17836 40350 17838 40402
rect 17890 40350 17892 40402
rect 17836 40338 17892 40350
rect 17388 40290 17444 40302
rect 17388 40238 17390 40290
rect 17442 40238 17444 40290
rect 17388 39732 17444 40238
rect 17388 39666 17444 39676
rect 17500 40178 17556 40190
rect 17500 40126 17502 40178
rect 17554 40126 17556 40178
rect 17500 39620 17556 40126
rect 17500 39554 17556 39564
rect 17948 39956 18004 39966
rect 17500 39060 17556 39070
rect 17948 39060 18004 39900
rect 18060 39060 18116 39070
rect 17276 39058 17780 39060
rect 17276 39006 17502 39058
rect 17554 39006 17780 39058
rect 17276 39004 17780 39006
rect 17500 38994 17556 39004
rect 16604 38612 17108 38668
rect 16156 38052 16212 38062
rect 16716 38052 16772 38062
rect 16044 38050 16772 38052
rect 16044 37998 16158 38050
rect 16210 37998 16718 38050
rect 16770 37998 16772 38050
rect 16044 37996 16772 37998
rect 16156 37986 16212 37996
rect 16716 37986 16772 37996
rect 16492 37826 16548 37838
rect 16492 37774 16494 37826
rect 16546 37774 16548 37826
rect 16380 36708 16436 36718
rect 16380 36594 16436 36652
rect 16380 36542 16382 36594
rect 16434 36542 16436 36594
rect 16380 36530 16436 36542
rect 16492 36596 16548 37774
rect 16828 37492 16884 37502
rect 16492 36530 16548 36540
rect 16716 37266 16772 37278
rect 16716 37214 16718 37266
rect 16770 37214 16772 37266
rect 16716 36596 16772 37214
rect 16828 36706 16884 37436
rect 16828 36654 16830 36706
rect 16882 36654 16884 36706
rect 16828 36642 16884 36654
rect 16716 36530 16772 36540
rect 16716 36370 16772 36382
rect 16716 36318 16718 36370
rect 16770 36318 16772 36370
rect 16492 35700 16548 35710
rect 16492 35586 16548 35644
rect 16492 35534 16494 35586
rect 16546 35534 16548 35586
rect 16492 35522 16548 35534
rect 16716 35364 16772 36318
rect 16828 36258 16884 36270
rect 16828 36206 16830 36258
rect 16882 36206 16884 36258
rect 16828 35700 16884 36206
rect 16940 35700 16996 35710
rect 16828 35644 16940 35700
rect 15932 35252 16100 35308
rect 16716 35298 16772 35308
rect 15708 34356 15764 34366
rect 15708 34242 15764 34300
rect 15708 34190 15710 34242
rect 15762 34190 15764 34242
rect 15708 34178 15764 34190
rect 15316 33516 15428 33572
rect 15260 33506 15316 33516
rect 15148 33294 15150 33346
rect 15202 33294 15204 33346
rect 15148 33282 15204 33294
rect 14924 32786 15092 32788
rect 14924 32734 14926 32786
rect 14978 32734 15092 32786
rect 14924 32732 15092 32734
rect 14924 32722 14980 32732
rect 15148 32676 15204 32686
rect 15372 32676 15428 33516
rect 15484 33906 15540 33918
rect 15484 33854 15486 33906
rect 15538 33854 15540 33906
rect 15484 33572 15540 33854
rect 15484 33506 15540 33516
rect 15148 32674 15764 32676
rect 15148 32622 15150 32674
rect 15202 32622 15764 32674
rect 15148 32620 15764 32622
rect 15148 32610 15204 32620
rect 14588 32564 14644 32574
rect 14028 32162 14084 32172
rect 14140 32562 14644 32564
rect 14140 32510 14590 32562
rect 14642 32510 14644 32562
rect 14140 32508 14644 32510
rect 12684 31938 12740 31948
rect 14028 32004 14084 32014
rect 14140 32004 14196 32508
rect 14588 32498 14644 32508
rect 15596 32452 15652 32462
rect 15596 32358 15652 32396
rect 14028 32002 14196 32004
rect 14028 31950 14030 32002
rect 14082 31950 14196 32002
rect 14028 31948 14196 31950
rect 14700 32340 14756 32350
rect 14028 31938 14084 31948
rect 14700 31890 14756 32284
rect 14700 31838 14702 31890
rect 14754 31838 14756 31890
rect 14700 31826 14756 31838
rect 14812 32338 14868 32350
rect 14812 32286 14814 32338
rect 14866 32286 14868 32338
rect 14476 31780 14532 31790
rect 14476 31686 14532 31724
rect 14140 31668 14196 31678
rect 14140 31574 14196 31612
rect 12684 31556 12740 31566
rect 12684 31462 12740 31500
rect 13692 31556 13748 31566
rect 13692 31462 13748 31500
rect 14028 31554 14084 31566
rect 14028 31502 14030 31554
rect 14082 31502 14084 31554
rect 14028 31444 14084 31502
rect 12460 30830 12462 30882
rect 12514 30830 12516 30882
rect 12460 29538 12516 30830
rect 12796 30884 12852 30894
rect 12796 30790 12852 30828
rect 14028 30884 14084 31388
rect 14812 31108 14868 32286
rect 15372 31780 15428 31790
rect 15372 31686 15428 31724
rect 15596 31778 15652 31790
rect 15596 31726 15598 31778
rect 15650 31726 15652 31778
rect 15036 31556 15092 31566
rect 15036 31462 15092 31500
rect 15596 31444 15652 31726
rect 15708 31556 15764 32620
rect 16044 31892 16100 35252
rect 16828 35140 16884 35150
rect 16492 35084 16828 35140
rect 16380 35026 16436 35038
rect 16380 34974 16382 35026
rect 16434 34974 16436 35026
rect 16380 34916 16436 34974
rect 16156 34860 16380 34916
rect 16156 34356 16212 34860
rect 16380 34850 16436 34860
rect 16156 34262 16212 34300
rect 16268 34130 16324 34142
rect 16268 34078 16270 34130
rect 16322 34078 16324 34130
rect 16156 33908 16212 33918
rect 16156 33814 16212 33852
rect 16268 33572 16324 34078
rect 16156 32788 16212 32798
rect 16268 32788 16324 33516
rect 16156 32786 16324 32788
rect 16156 32734 16158 32786
rect 16210 32734 16324 32786
rect 16156 32732 16324 32734
rect 16156 32722 16212 32732
rect 16492 32564 16548 35084
rect 16828 35046 16884 35084
rect 16940 35138 16996 35644
rect 16940 35086 16942 35138
rect 16994 35086 16996 35138
rect 16940 35074 16996 35086
rect 16940 33236 16996 33246
rect 16716 33180 16940 33236
rect 16716 32674 16772 33180
rect 16940 33142 16996 33180
rect 17052 32788 17108 38612
rect 17500 38052 17556 38062
rect 17388 37940 17444 37978
rect 17500 37958 17556 37996
rect 17388 37874 17444 37884
rect 17276 37826 17332 37838
rect 17276 37774 17278 37826
rect 17330 37774 17332 37826
rect 17276 35138 17332 37774
rect 17612 37492 17668 37502
rect 17724 37492 17780 39004
rect 17948 39058 18116 39060
rect 17948 39006 18062 39058
rect 18114 39006 18116 39058
rect 17948 39004 18116 39006
rect 17612 37490 17780 37492
rect 17612 37438 17614 37490
rect 17666 37438 17780 37490
rect 17612 37436 17780 37438
rect 17836 38052 17892 38062
rect 17836 37490 17892 37996
rect 17948 38050 18004 39004
rect 18060 38994 18116 39004
rect 17948 37998 17950 38050
rect 18002 37998 18004 38050
rect 17948 37986 18004 37998
rect 18060 38050 18116 38062
rect 18060 37998 18062 38050
rect 18114 37998 18116 38050
rect 18060 37940 18116 37998
rect 18060 37874 18116 37884
rect 17836 37438 17838 37490
rect 17890 37438 17892 37490
rect 17500 36932 17556 36942
rect 17500 36594 17556 36876
rect 17500 36542 17502 36594
rect 17554 36542 17556 36594
rect 17500 36530 17556 36542
rect 17500 35810 17556 35822
rect 17500 35758 17502 35810
rect 17554 35758 17556 35810
rect 17388 35700 17444 35710
rect 17388 35606 17444 35644
rect 17500 35252 17556 35758
rect 17612 35476 17668 37436
rect 17612 35410 17668 35420
rect 17724 36596 17780 36606
rect 17276 35086 17278 35138
rect 17330 35086 17332 35138
rect 17276 35074 17332 35086
rect 17388 35196 17556 35252
rect 17164 34916 17220 34926
rect 17388 34916 17444 35196
rect 17724 35028 17780 36540
rect 17836 35308 17892 37438
rect 17948 37492 18004 37502
rect 17948 37154 18004 37436
rect 17948 37102 17950 37154
rect 18002 37102 18004 37154
rect 17948 35700 18004 37102
rect 18060 37266 18116 37278
rect 18060 37214 18062 37266
rect 18114 37214 18116 37266
rect 18060 37156 18116 37214
rect 18060 35922 18116 37100
rect 18060 35870 18062 35922
rect 18114 35870 18116 35922
rect 18060 35858 18116 35870
rect 17948 35644 18116 35700
rect 17836 35252 18004 35308
rect 17724 35026 17892 35028
rect 17724 34974 17726 35026
rect 17778 34974 17892 35026
rect 17724 34972 17892 34974
rect 17724 34962 17780 34972
rect 17220 34860 17444 34916
rect 17164 34822 17220 34860
rect 17612 33460 17668 33470
rect 17052 32732 17332 32788
rect 16716 32622 16718 32674
rect 16770 32622 16772 32674
rect 16716 32610 16772 32622
rect 16268 32562 16548 32564
rect 16268 32510 16494 32562
rect 16546 32510 16548 32562
rect 16268 32508 16548 32510
rect 16268 32002 16324 32508
rect 16492 32498 16548 32508
rect 16268 31950 16270 32002
rect 16322 31950 16324 32002
rect 16268 31938 16324 31950
rect 16716 31892 16772 31902
rect 16044 31836 16212 31892
rect 15820 31780 15876 31790
rect 15820 31686 15876 31724
rect 16044 31668 16100 31678
rect 15708 31500 15876 31556
rect 15596 31378 15652 31388
rect 14924 31108 14980 31118
rect 14812 31106 14980 31108
rect 14812 31054 14926 31106
rect 14978 31054 14980 31106
rect 14812 31052 14980 31054
rect 14924 31042 14980 31052
rect 15596 30996 15652 31006
rect 14028 30818 14084 30828
rect 15372 30994 15652 30996
rect 15372 30942 15598 30994
rect 15650 30942 15652 30994
rect 15372 30940 15652 30942
rect 12460 29486 12462 29538
rect 12514 29486 12516 29538
rect 12460 29474 12516 29486
rect 13020 30212 13076 30222
rect 12796 29428 12852 29438
rect 12852 29372 12964 29428
rect 12796 29334 12852 29372
rect 12796 28642 12852 28654
rect 12796 28590 12798 28642
rect 12850 28590 12852 28642
rect 12796 28084 12852 28590
rect 12796 28018 12852 28028
rect 12348 27794 12404 27804
rect 12572 27748 12628 27758
rect 12124 27300 12180 27310
rect 11228 27188 11284 27198
rect 11228 27094 11284 27132
rect 11116 26450 11172 26460
rect 12012 26516 12068 26526
rect 11676 26404 11732 26414
rect 11116 26292 11172 26302
rect 11004 26290 11172 26292
rect 11004 26238 11118 26290
rect 11170 26238 11172 26290
rect 11004 26236 11172 26238
rect 11116 25956 11172 26236
rect 11676 26290 11732 26348
rect 11676 26238 11678 26290
rect 11730 26238 11732 26290
rect 11340 26068 11396 26078
rect 11116 25900 11284 25956
rect 11116 25730 11172 25742
rect 11116 25678 11118 25730
rect 11170 25678 11172 25730
rect 8988 24658 9044 24668
rect 9324 25618 9380 25630
rect 9324 25566 9326 25618
rect 9378 25566 9380 25618
rect 2492 24610 2548 24622
rect 2492 24558 2494 24610
rect 2546 24558 2548 24610
rect 2492 24276 2548 24558
rect 6300 24612 6356 24622
rect 8428 24612 8484 24622
rect 6300 24518 6356 24556
rect 8204 24610 8484 24612
rect 8204 24558 8430 24610
rect 8482 24558 8484 24610
rect 8204 24556 8484 24558
rect 4476 24332 4740 24342
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4476 24266 4740 24276
rect 2492 24210 2548 24220
rect 7196 23938 7252 23950
rect 7196 23886 7198 23938
rect 7250 23886 7252 23938
rect 6972 23828 7028 23838
rect 6972 23734 7028 23772
rect 2492 23714 2548 23726
rect 2492 23662 2494 23714
rect 2546 23662 2548 23714
rect 2492 23604 2548 23662
rect 2492 23538 2548 23548
rect 7196 23492 7252 23886
rect 7644 23940 7700 23950
rect 7644 23846 7700 23884
rect 7756 23938 7812 23950
rect 7756 23886 7758 23938
rect 7810 23886 7812 23938
rect 7756 23604 7812 23886
rect 8092 23940 8148 23950
rect 8204 23940 8260 24556
rect 8428 24546 8484 24556
rect 8764 24612 8820 24622
rect 8764 24518 8820 24556
rect 8876 24610 8932 24622
rect 8876 24558 8878 24610
rect 8930 24558 8932 24610
rect 8316 24164 8372 24174
rect 8876 24164 8932 24558
rect 8316 24162 8932 24164
rect 8316 24110 8318 24162
rect 8370 24110 8932 24162
rect 8316 24108 8932 24110
rect 8316 24098 8372 24108
rect 8092 23938 8260 23940
rect 8092 23886 8094 23938
rect 8146 23886 8260 23938
rect 8092 23884 8260 23886
rect 9324 23940 9380 25566
rect 10444 25508 10500 25518
rect 10444 25414 10500 25452
rect 10220 25396 10276 25406
rect 10220 25394 10388 25396
rect 10220 25342 10222 25394
rect 10274 25342 10388 25394
rect 10220 25340 10388 25342
rect 10220 25330 10276 25340
rect 10220 24948 10276 24958
rect 10220 24854 10276 24892
rect 10108 24836 10164 24846
rect 8092 23828 8148 23884
rect 9324 23874 9380 23884
rect 9660 24610 9716 24622
rect 9660 24558 9662 24610
rect 9714 24558 9716 24610
rect 8092 23762 8148 23772
rect 8316 23826 8372 23838
rect 8316 23774 8318 23826
rect 8370 23774 8372 23826
rect 7756 23538 7812 23548
rect 7196 23426 7252 23436
rect 2156 23090 2212 23100
rect 5404 23156 5460 23166
rect 5404 23154 6020 23156
rect 5404 23102 5406 23154
rect 5458 23102 6020 23154
rect 5404 23100 6020 23102
rect 5404 23090 5460 23100
rect 2492 23042 2548 23054
rect 2492 22990 2494 23042
rect 2546 22990 2548 23042
rect 2492 22932 2548 22990
rect 2492 22866 2548 22876
rect 4476 22764 4740 22774
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4476 22698 4740 22708
rect 2044 22306 2100 22316
rect 1708 22260 1764 22270
rect 1708 22166 1764 22204
rect 2380 22258 2436 22270
rect 2380 22206 2382 22258
rect 2434 22206 2436 22258
rect 2044 22148 2100 22158
rect 2044 22146 2212 22148
rect 2044 22094 2046 22146
rect 2098 22094 2212 22146
rect 2044 22092 2212 22094
rect 2044 22082 2100 22092
rect 2044 21700 2100 21710
rect 2044 21606 2100 21644
rect 1708 21586 1764 21598
rect 1708 21534 1710 21586
rect 1762 21534 1764 21586
rect 1708 21476 1764 21534
rect 2156 21588 2212 22092
rect 2380 21812 2436 22206
rect 2380 21746 2436 21756
rect 2492 22260 2548 22270
rect 2492 21810 2548 22204
rect 2492 21758 2494 21810
rect 2546 21758 2548 21810
rect 2492 21746 2548 21758
rect 2716 22146 2772 22158
rect 2716 22094 2718 22146
rect 2770 22094 2772 22146
rect 2156 21522 2212 21532
rect 1708 20916 1764 21420
rect 1708 20850 1764 20860
rect 1708 20690 1764 20702
rect 1708 20638 1710 20690
rect 1762 20638 1764 20690
rect 1708 20244 1764 20638
rect 2044 20580 2100 20590
rect 2044 20578 2212 20580
rect 2044 20526 2046 20578
rect 2098 20526 2212 20578
rect 2044 20524 2212 20526
rect 2044 20514 2100 20524
rect 1708 20178 1764 20188
rect 2044 20132 2100 20142
rect 2044 20038 2100 20076
rect 1708 20018 1764 20030
rect 1708 19966 1710 20018
rect 1762 19966 1764 20018
rect 1708 19572 1764 19966
rect 1708 19506 1764 19516
rect 2044 18562 2100 18574
rect 2044 18510 2046 18562
rect 2098 18510 2100 18562
rect 1708 18450 1764 18462
rect 1708 18398 1710 18450
rect 1762 18398 1764 18450
rect 1708 18228 1764 18398
rect 2044 18340 2100 18510
rect 2044 18274 2100 18284
rect 1708 18162 1764 18172
rect 1708 17556 1764 17566
rect 1708 17462 1764 17500
rect 2044 17444 2100 17454
rect 2044 17350 2100 17388
rect 2156 17332 2212 20524
rect 2492 20578 2548 20590
rect 2492 20526 2494 20578
rect 2546 20526 2548 20578
rect 2492 20244 2548 20526
rect 2492 20178 2548 20188
rect 2492 19906 2548 19918
rect 2492 19854 2494 19906
rect 2546 19854 2548 19906
rect 2492 19572 2548 19854
rect 2716 19796 2772 22094
rect 3164 22146 3220 22158
rect 3164 22094 3166 22146
rect 3218 22094 3220 22146
rect 3164 21812 3220 22094
rect 3164 21746 3220 21756
rect 2940 21476 2996 21486
rect 2940 21382 2996 21420
rect 4476 21196 4740 21206
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4476 21130 4740 21140
rect 5964 20804 6020 23100
rect 6076 23044 6132 23054
rect 6076 22950 6132 22988
rect 6972 23044 7028 23054
rect 6972 22594 7028 22988
rect 8204 23042 8260 23054
rect 8204 22990 8206 23042
rect 8258 22990 8260 23042
rect 6972 22542 6974 22594
rect 7026 22542 7028 22594
rect 6972 22530 7028 22542
rect 7756 22594 7812 22606
rect 7756 22542 7758 22594
rect 7810 22542 7812 22594
rect 7084 22484 7140 22494
rect 7084 22390 7140 22428
rect 7756 22484 7812 22542
rect 7756 22418 7812 22428
rect 7980 22372 8036 22382
rect 8204 22372 8260 22990
rect 8316 22484 8372 23774
rect 8764 23828 8820 23838
rect 8428 22484 8484 22494
rect 8316 22428 8428 22484
rect 7980 22370 8260 22372
rect 7980 22318 7982 22370
rect 8034 22318 8260 22370
rect 7980 22316 8260 22318
rect 8428 22370 8484 22428
rect 8428 22318 8430 22370
rect 8482 22318 8484 22370
rect 6300 21586 6356 21598
rect 6300 21534 6302 21586
rect 6354 21534 6356 21586
rect 6076 20804 6132 20814
rect 5964 20802 6132 20804
rect 5964 20750 6078 20802
rect 6130 20750 6132 20802
rect 5964 20748 6132 20750
rect 2716 19730 2772 19740
rect 6076 20018 6132 20748
rect 6300 20692 6356 21534
rect 6524 21588 6580 21598
rect 6524 21494 6580 21532
rect 7868 21588 7924 21598
rect 7868 21494 7924 21532
rect 7980 21586 8036 22316
rect 8428 22306 8484 22318
rect 8764 22370 8820 23772
rect 9212 23604 9268 23614
rect 8764 22318 8766 22370
rect 8818 22318 8820 22370
rect 8764 22306 8820 22318
rect 8988 22484 9044 22494
rect 8988 21698 9044 22428
rect 8988 21646 8990 21698
rect 9042 21646 9044 21698
rect 8988 21634 9044 21646
rect 9212 22370 9268 23548
rect 9660 23604 9716 24558
rect 9996 24050 10052 24062
rect 9996 23998 9998 24050
rect 10050 23998 10052 24050
rect 9996 23716 10052 23998
rect 9996 23650 10052 23660
rect 9660 23538 9716 23548
rect 9772 23156 9828 23166
rect 9772 23062 9828 23100
rect 10108 22930 10164 24780
rect 10332 23492 10388 25340
rect 11116 24834 11172 25678
rect 11228 24948 11284 25900
rect 11340 25618 11396 26012
rect 11340 25566 11342 25618
rect 11394 25566 11396 25618
rect 11340 25554 11396 25566
rect 11228 24882 11284 24892
rect 11676 25506 11732 26238
rect 11676 25454 11678 25506
rect 11730 25454 11732 25506
rect 11116 24782 11118 24834
rect 11170 24782 11172 24834
rect 11116 24770 11172 24782
rect 10332 23156 10388 23436
rect 11116 24612 11172 24622
rect 10332 23154 10500 23156
rect 10332 23102 10334 23154
rect 10386 23102 10500 23154
rect 10332 23100 10500 23102
rect 10332 23090 10388 23100
rect 10108 22878 10110 22930
rect 10162 22878 10164 22930
rect 10108 22866 10164 22878
rect 10444 22484 10500 23100
rect 11116 23154 11172 24556
rect 11676 24612 11732 25454
rect 12012 26290 12068 26460
rect 12012 26238 12014 26290
rect 12066 26238 12068 26290
rect 11788 24724 11844 24734
rect 11788 24630 11844 24668
rect 11676 24546 11732 24556
rect 11228 24498 11284 24510
rect 11228 24446 11230 24498
rect 11282 24446 11284 24498
rect 11228 24052 11284 24446
rect 11228 23986 11284 23996
rect 11788 23940 11844 23950
rect 11116 23102 11118 23154
rect 11170 23102 11172 23154
rect 11116 23090 11172 23102
rect 11228 23716 11284 23726
rect 11228 23154 11284 23660
rect 11228 23102 11230 23154
rect 11282 23102 11284 23154
rect 11228 23090 11284 23102
rect 11788 23154 11844 23884
rect 12012 23828 12068 26238
rect 12124 24724 12180 27244
rect 12572 27188 12628 27692
rect 12796 27300 12852 27310
rect 12908 27300 12964 29372
rect 13020 29426 13076 30156
rect 13020 29374 13022 29426
rect 13074 29374 13076 29426
rect 13020 29362 13076 29374
rect 13580 30210 13636 30222
rect 13580 30158 13582 30210
rect 13634 30158 13636 30210
rect 13468 29202 13524 29214
rect 13468 29150 13470 29202
rect 13522 29150 13524 29202
rect 13468 28868 13524 29150
rect 13580 29204 13636 30158
rect 14252 30098 14308 30110
rect 14252 30046 14254 30098
rect 14306 30046 14308 30098
rect 14028 29652 14084 29662
rect 14028 29426 14084 29596
rect 14028 29374 14030 29426
rect 14082 29374 14084 29426
rect 14028 29362 14084 29374
rect 14252 29428 14308 30046
rect 14252 29362 14308 29372
rect 15148 29426 15204 29438
rect 15148 29374 15150 29426
rect 15202 29374 15204 29426
rect 13692 29316 13748 29326
rect 13692 29222 13748 29260
rect 13580 29138 13636 29148
rect 14252 29204 14308 29214
rect 13468 28802 13524 28812
rect 13468 28644 13524 28654
rect 13468 28550 13524 28588
rect 14252 28644 14308 29148
rect 14252 28550 14308 28588
rect 12852 27244 12964 27300
rect 13580 28530 13636 28542
rect 13580 28478 13582 28530
rect 13634 28478 13636 28530
rect 12796 27234 12852 27244
rect 13580 27188 13636 28478
rect 15036 28532 15092 28542
rect 15036 28438 15092 28476
rect 14364 28084 14420 28094
rect 14364 27990 14420 28028
rect 14924 28084 14980 28094
rect 13916 27746 13972 27758
rect 13916 27694 13918 27746
rect 13970 27694 13972 27746
rect 12348 25506 12404 25518
rect 12348 25454 12350 25506
rect 12402 25454 12404 25506
rect 12236 24724 12292 24734
rect 12124 24722 12292 24724
rect 12124 24670 12238 24722
rect 12290 24670 12292 24722
rect 12124 24668 12292 24670
rect 12236 24658 12292 24668
rect 12124 24052 12180 24062
rect 12124 23958 12180 23996
rect 12124 23828 12180 23838
rect 12012 23772 12124 23828
rect 12124 23762 12180 23772
rect 12348 23716 12404 25454
rect 12572 24610 12628 27132
rect 13468 27132 13636 27188
rect 13692 27636 13748 27646
rect 13468 27076 13524 27132
rect 13356 27020 13524 27076
rect 13692 27074 13748 27580
rect 13692 27022 13694 27074
rect 13746 27022 13748 27074
rect 13020 26404 13076 26414
rect 12796 26178 12852 26190
rect 12796 26126 12798 26178
rect 12850 26126 12852 26178
rect 12796 25732 12852 26126
rect 12796 25666 12852 25676
rect 12908 25394 12964 25406
rect 12908 25342 12910 25394
rect 12962 25342 12964 25394
rect 12908 25060 12964 25342
rect 12572 24558 12574 24610
rect 12626 24558 12628 24610
rect 12572 24546 12628 24558
rect 12684 25004 12908 25060
rect 12348 23650 12404 23660
rect 11788 23102 11790 23154
rect 11842 23102 11844 23154
rect 11788 23090 11844 23102
rect 12236 23156 12292 23166
rect 12124 23044 12180 23054
rect 11900 23042 12180 23044
rect 11900 22990 12126 23042
rect 12178 22990 12180 23042
rect 11900 22988 12180 22990
rect 10780 22484 10836 22494
rect 10444 22482 10836 22484
rect 10444 22430 10782 22482
rect 10834 22430 10836 22482
rect 10444 22428 10836 22430
rect 9212 22318 9214 22370
rect 9266 22318 9268 22370
rect 7980 21534 7982 21586
rect 8034 21534 8036 21586
rect 7980 21522 8036 21534
rect 8764 21586 8820 21598
rect 8764 21534 8766 21586
rect 8818 21534 8820 21586
rect 6860 21364 6916 21374
rect 6300 20626 6356 20636
rect 6748 21028 6804 21038
rect 6076 19966 6078 20018
rect 6130 19966 6132 20018
rect 4476 19628 4740 19638
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4476 19562 4740 19572
rect 2492 19506 2548 19516
rect 6076 18452 6132 19966
rect 6748 19346 6804 20972
rect 6860 20914 6916 21308
rect 6860 20862 6862 20914
rect 6914 20862 6916 20914
rect 6860 20850 6916 20862
rect 8764 20916 8820 21534
rect 9212 21588 9268 22318
rect 10108 22372 10164 22382
rect 10108 22278 10164 22316
rect 10444 22370 10500 22428
rect 10780 22418 10836 22428
rect 11788 22484 11844 22494
rect 11900 22484 11956 22988
rect 12124 22978 12180 22988
rect 11844 22428 11956 22484
rect 11788 22390 11844 22428
rect 10444 22318 10446 22370
rect 10498 22318 10500 22370
rect 10444 22306 10500 22318
rect 11228 22370 11284 22382
rect 11228 22318 11230 22370
rect 11282 22318 11284 22370
rect 11004 22148 11060 22158
rect 8988 21476 9044 21486
rect 8988 21362 9044 21420
rect 8988 21310 8990 21362
rect 9042 21310 9044 21362
rect 8988 21298 9044 21310
rect 8988 20916 9044 20926
rect 8764 20860 8988 20916
rect 8988 20822 9044 20860
rect 9212 20804 9268 21532
rect 9996 22036 10052 22046
rect 9660 21476 9716 21486
rect 9660 21382 9716 21420
rect 9548 21364 9604 21374
rect 9548 21270 9604 21308
rect 9212 20738 9268 20748
rect 9548 20802 9604 20814
rect 9548 20750 9550 20802
rect 9602 20750 9604 20802
rect 9324 20692 9380 20702
rect 6860 19906 6916 19918
rect 6860 19854 6862 19906
rect 6914 19854 6916 19906
rect 6860 19458 6916 19854
rect 7980 19908 8036 19918
rect 6860 19406 6862 19458
rect 6914 19406 6916 19458
rect 6860 19394 6916 19406
rect 7196 19684 7252 19694
rect 6748 19294 6750 19346
rect 6802 19294 6804 19346
rect 6748 19282 6804 19294
rect 7196 19234 7252 19628
rect 7196 19182 7198 19234
rect 7250 19182 7252 19234
rect 7196 19170 7252 19182
rect 7420 19234 7476 19246
rect 7420 19182 7422 19234
rect 7474 19182 7476 19234
rect 6076 18386 6132 18396
rect 6524 18450 6580 18462
rect 6524 18398 6526 18450
rect 6578 18398 6580 18450
rect 2492 18338 2548 18350
rect 2492 18286 2494 18338
rect 2546 18286 2548 18338
rect 2492 18228 2548 18286
rect 6524 18340 6580 18398
rect 6524 18274 6580 18284
rect 6972 18450 7028 18462
rect 6972 18398 6974 18450
rect 7026 18398 7028 18450
rect 2492 18162 2548 18172
rect 6972 18116 7028 18398
rect 4476 18060 4740 18070
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 6972 18050 7028 18060
rect 7084 18452 7140 18462
rect 4476 17994 4740 18004
rect 7084 17666 7140 18396
rect 7084 17614 7086 17666
rect 7138 17614 7140 17666
rect 7084 17602 7140 17614
rect 2156 17266 2212 17276
rect 2380 17554 2436 17566
rect 2380 17502 2382 17554
rect 2434 17502 2436 17554
rect 2044 16994 2100 17006
rect 2044 16942 2046 16994
rect 2098 16942 2100 16994
rect 1820 16882 1876 16894
rect 1820 16830 1822 16882
rect 1874 16830 1876 16882
rect 1820 16212 1876 16830
rect 2044 16772 2100 16942
rect 2380 16884 2436 17502
rect 2492 17556 2548 17566
rect 2492 17106 2548 17500
rect 2716 17556 2772 17566
rect 2716 17462 2772 17500
rect 7420 17556 7476 19182
rect 7868 19124 7924 19134
rect 7868 18450 7924 19068
rect 7868 18398 7870 18450
rect 7922 18398 7924 18450
rect 7868 18386 7924 18398
rect 7980 18450 8036 19852
rect 8988 19908 9044 19918
rect 8988 19814 9044 19852
rect 8764 19234 8820 19246
rect 8764 19182 8766 19234
rect 8818 19182 8820 19234
rect 8764 19124 8820 19182
rect 8876 19236 8932 19246
rect 8876 19234 9044 19236
rect 8876 19182 8878 19234
rect 8930 19182 9044 19234
rect 8876 19180 9044 19182
rect 8876 19170 8932 19180
rect 8764 19058 8820 19068
rect 8876 18676 8932 18686
rect 7980 18398 7982 18450
rect 8034 18398 8036 18450
rect 7980 18386 8036 18398
rect 8316 18452 8372 18462
rect 8372 18396 8484 18452
rect 8316 18386 8372 18396
rect 8204 18340 8260 18350
rect 7868 18228 7924 18238
rect 7868 17778 7924 18172
rect 8204 18226 8260 18284
rect 8204 18174 8206 18226
rect 8258 18174 8260 18226
rect 8204 18162 8260 18174
rect 7868 17726 7870 17778
rect 7922 17726 7924 17778
rect 7868 17714 7924 17726
rect 7420 17490 7476 17500
rect 2492 17054 2494 17106
rect 2546 17054 2548 17106
rect 2492 17042 2548 17054
rect 3164 17442 3220 17454
rect 3164 17390 3166 17442
rect 3218 17390 3220 17442
rect 2380 16818 2436 16828
rect 3164 16884 3220 17390
rect 3164 16818 3220 16828
rect 5180 17444 5236 17454
rect 2044 16706 2100 16716
rect 4476 16492 4740 16502
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4476 16426 4740 16436
rect 1820 16118 1876 16156
rect 4476 14924 4740 14934
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4476 14858 4740 14868
rect 5180 14532 5236 17388
rect 8428 16098 8484 18396
rect 8764 18450 8820 18462
rect 8764 18398 8766 18450
rect 8818 18398 8820 18450
rect 8764 16660 8820 18398
rect 8876 18338 8932 18620
rect 8876 18286 8878 18338
rect 8930 18286 8932 18338
rect 8876 18274 8932 18286
rect 8988 16884 9044 19180
rect 9324 18340 9380 20636
rect 9548 20132 9604 20750
rect 9548 20066 9604 20076
rect 9772 19458 9828 19470
rect 9772 19406 9774 19458
rect 9826 19406 9828 19458
rect 9660 19236 9716 19246
rect 9660 19142 9716 19180
rect 9548 18340 9604 18350
rect 9324 18338 9604 18340
rect 9324 18286 9550 18338
rect 9602 18286 9604 18338
rect 9324 18284 9604 18286
rect 8988 16818 9044 16828
rect 9548 18116 9604 18284
rect 8876 16772 8932 16782
rect 8876 16678 8932 16716
rect 8764 16594 8820 16604
rect 8988 16658 9044 16670
rect 8988 16606 8990 16658
rect 9042 16606 9044 16658
rect 8988 16212 9044 16606
rect 9100 16212 9156 16222
rect 8988 16210 9156 16212
rect 8988 16158 9102 16210
rect 9154 16158 9156 16210
rect 8988 16156 9156 16158
rect 9100 16146 9156 16156
rect 8428 16046 8430 16098
rect 8482 16046 8484 16098
rect 8428 16034 8484 16046
rect 5180 14466 5236 14476
rect 9548 14530 9604 18060
rect 9772 17780 9828 19406
rect 9884 19122 9940 19134
rect 9884 19070 9886 19122
rect 9938 19070 9940 19122
rect 9884 18676 9940 19070
rect 9884 18610 9940 18620
rect 9996 18564 10052 21980
rect 11004 21698 11060 22092
rect 11228 22036 11284 22318
rect 11228 21970 11284 21980
rect 12236 22146 12292 23100
rect 12684 23042 12740 25004
rect 12908 24994 12964 25004
rect 13020 24722 13076 26348
rect 13020 24670 13022 24722
rect 13074 24670 13076 24722
rect 13020 24658 13076 24670
rect 13356 24498 13412 27020
rect 13692 27010 13748 27022
rect 13580 26964 13636 26974
rect 13468 25732 13524 25742
rect 13468 25638 13524 25676
rect 13580 25618 13636 26908
rect 13916 26908 13972 27694
rect 14028 27298 14084 27310
rect 14028 27246 14030 27298
rect 14082 27246 14084 27298
rect 14028 27076 14084 27246
rect 14028 27010 14084 27020
rect 14140 27300 14196 27310
rect 14140 27074 14196 27244
rect 14140 27022 14142 27074
rect 14194 27022 14196 27074
rect 14140 27010 14196 27022
rect 14364 27186 14420 27198
rect 14364 27134 14366 27186
rect 14418 27134 14420 27186
rect 14364 26908 14420 27134
rect 13916 26852 14420 26908
rect 14476 27076 14532 27086
rect 13580 25566 13582 25618
rect 13634 25566 13636 25618
rect 13580 25554 13636 25566
rect 13356 24446 13358 24498
rect 13410 24446 13412 24498
rect 13356 24434 13412 24446
rect 13916 25282 13972 25294
rect 13916 25230 13918 25282
rect 13970 25230 13972 25282
rect 12908 23938 12964 23950
rect 12908 23886 12910 23938
rect 12962 23886 12964 23938
rect 12908 23828 12964 23886
rect 12908 23762 12964 23772
rect 13692 23828 13748 23838
rect 13468 23266 13524 23278
rect 13468 23214 13470 23266
rect 13522 23214 13524 23266
rect 13020 23156 13076 23166
rect 13020 23062 13076 23100
rect 13468 23156 13524 23214
rect 13468 23090 13524 23100
rect 12684 22990 12686 23042
rect 12738 22990 12740 23042
rect 12684 22978 12740 22990
rect 13692 22932 13748 23772
rect 13804 23380 13860 23390
rect 13804 23266 13860 23324
rect 13804 23214 13806 23266
rect 13858 23214 13860 23266
rect 13804 23202 13860 23214
rect 13468 22876 13748 22932
rect 13468 22372 13524 22876
rect 12236 22094 12238 22146
rect 12290 22094 12292 22146
rect 11004 21646 11006 21698
rect 11058 21646 11060 21698
rect 11004 21634 11060 21646
rect 10220 21586 10276 21598
rect 10220 21534 10222 21586
rect 10274 21534 10276 21586
rect 10108 21028 10164 21038
rect 10108 20934 10164 20972
rect 10220 19906 10276 21534
rect 10332 20916 10388 20926
rect 11900 20916 11956 20926
rect 10332 20822 10388 20860
rect 11788 20914 11956 20916
rect 11788 20862 11902 20914
rect 11954 20862 11956 20914
rect 11788 20860 11956 20862
rect 10556 20804 10612 20814
rect 10556 20710 10612 20748
rect 11452 20802 11508 20814
rect 11452 20750 11454 20802
rect 11506 20750 11508 20802
rect 10220 19854 10222 19906
rect 10274 19854 10276 19906
rect 9996 18508 10164 18564
rect 9772 17714 9828 17724
rect 9884 18452 9940 18462
rect 9884 18340 9940 18396
rect 10108 18450 10164 18508
rect 10108 18398 10110 18450
rect 10162 18398 10164 18450
rect 10108 18386 10164 18398
rect 9884 18284 10052 18340
rect 9884 16882 9940 18284
rect 9996 18228 10052 18284
rect 10220 18228 10276 19854
rect 11452 19908 11508 20750
rect 11452 19842 11508 19852
rect 11004 19684 11060 19694
rect 10444 19236 10500 19246
rect 9996 18172 10276 18228
rect 10332 19234 10500 19236
rect 10332 19182 10446 19234
rect 10498 19182 10500 19234
rect 10332 19180 10500 19182
rect 9996 17778 10052 17790
rect 9996 17726 9998 17778
rect 10050 17726 10052 17778
rect 9996 16996 10052 17726
rect 9996 16940 10276 16996
rect 9884 16830 9886 16882
rect 9938 16830 9940 16882
rect 9884 16818 9940 16830
rect 10108 16772 10164 16782
rect 10108 14754 10164 16716
rect 10108 14702 10110 14754
rect 10162 14702 10164 14754
rect 10108 14690 10164 14702
rect 10220 16660 10276 16940
rect 10220 14644 10276 16604
rect 10332 16548 10388 19180
rect 10444 19170 10500 19180
rect 11004 19234 11060 19628
rect 11004 19182 11006 19234
rect 11058 19182 11060 19234
rect 11004 19170 11060 19182
rect 11452 19234 11508 19246
rect 11452 19182 11454 19234
rect 11506 19182 11508 19234
rect 11452 19124 11508 19182
rect 11340 18452 11396 18462
rect 10556 18340 10612 18350
rect 10556 18246 10612 18284
rect 11340 18338 11396 18396
rect 11340 18286 11342 18338
rect 11394 18286 11396 18338
rect 10444 18228 10500 18238
rect 10444 18134 10500 18172
rect 11116 17780 11172 17790
rect 11116 17686 11172 17724
rect 11116 17556 11172 17566
rect 11004 17444 11060 17454
rect 10556 17442 11060 17444
rect 10556 17390 11006 17442
rect 11058 17390 11060 17442
rect 10556 17388 11060 17390
rect 10556 16994 10612 17388
rect 11004 17378 11060 17388
rect 10556 16942 10558 16994
rect 10610 16942 10612 16994
rect 10556 16930 10612 16942
rect 10332 16482 10388 16492
rect 10444 14644 10500 14654
rect 10220 14642 10500 14644
rect 10220 14590 10446 14642
rect 10498 14590 10500 14642
rect 10220 14588 10500 14590
rect 10444 14578 10500 14588
rect 9548 14478 9550 14530
rect 9602 14478 9604 14530
rect 9548 14466 9604 14478
rect 9772 14532 9828 14542
rect 9772 14438 9828 14476
rect 11116 14530 11172 17500
rect 11340 17220 11396 18286
rect 11452 17556 11508 19068
rect 11788 18900 11844 20860
rect 11900 20850 11956 20860
rect 12236 20468 12292 22094
rect 13356 22316 13524 22372
rect 13356 21924 13412 22316
rect 13580 22258 13636 22270
rect 13580 22206 13582 22258
rect 13634 22206 13636 22258
rect 13468 22148 13524 22158
rect 13468 22054 13524 22092
rect 13356 21868 13524 21924
rect 13468 21586 13524 21868
rect 13580 21812 13636 22206
rect 13916 22146 13972 25230
rect 14028 24722 14084 26852
rect 14252 25508 14308 25518
rect 14252 25414 14308 25452
rect 14252 25060 14308 25070
rect 14476 25060 14532 27020
rect 14700 27074 14756 27086
rect 14700 27022 14702 27074
rect 14754 27022 14756 27074
rect 14700 26404 14756 27022
rect 14924 26908 14980 28028
rect 15148 27748 15204 29374
rect 15148 27682 15204 27692
rect 15372 28644 15428 30940
rect 15596 30930 15652 30940
rect 15820 29540 15876 31500
rect 16044 31218 16100 31612
rect 16044 31166 16046 31218
rect 16098 31166 16100 31218
rect 16044 29650 16100 31166
rect 16044 29598 16046 29650
rect 16098 29598 16100 29650
rect 16044 29586 16100 29598
rect 15596 29538 15876 29540
rect 15596 29486 15822 29538
rect 15874 29486 15876 29538
rect 15596 29484 15876 29486
rect 15372 26908 15428 28588
rect 15484 29314 15540 29326
rect 15484 29262 15486 29314
rect 15538 29262 15540 29314
rect 15484 27076 15540 29262
rect 15596 28084 15652 29484
rect 15820 29474 15876 29484
rect 15932 29316 15988 29326
rect 15932 29222 15988 29260
rect 16044 29204 16100 29214
rect 16044 28644 16100 29148
rect 16156 28756 16212 31836
rect 16716 31798 16772 31836
rect 16604 31780 16660 31790
rect 16380 31556 16436 31566
rect 16380 30994 16436 31500
rect 16380 30942 16382 30994
rect 16434 30942 16436 30994
rect 16380 30930 16436 30942
rect 16604 31108 16660 31724
rect 16268 30772 16324 30782
rect 16268 29650 16324 30716
rect 16380 30324 16436 30334
rect 16604 30324 16660 31052
rect 16380 30322 16660 30324
rect 16380 30270 16382 30322
rect 16434 30270 16660 30322
rect 16380 30268 16660 30270
rect 16380 30258 16436 30268
rect 16268 29598 16270 29650
rect 16322 29598 16324 29650
rect 16268 29586 16324 29598
rect 16716 29540 16772 29550
rect 16716 29446 16772 29484
rect 16604 29204 16660 29214
rect 16604 29110 16660 29148
rect 16156 28690 16212 28700
rect 16604 28756 16660 28766
rect 17164 28756 17220 28766
rect 15932 28588 16100 28644
rect 15820 28532 15876 28542
rect 15708 28084 15764 28094
rect 15596 28082 15764 28084
rect 15596 28030 15710 28082
rect 15762 28030 15764 28082
rect 15596 28028 15764 28030
rect 15708 28018 15764 28028
rect 15820 28082 15876 28476
rect 15820 28030 15822 28082
rect 15874 28030 15876 28082
rect 15820 28018 15876 28030
rect 15932 28082 15988 28588
rect 15932 28030 15934 28082
rect 15986 28030 15988 28082
rect 15932 28018 15988 28030
rect 16492 27970 16548 27982
rect 16492 27918 16494 27970
rect 16546 27918 16548 27970
rect 15484 27010 15540 27020
rect 15596 27860 15652 27870
rect 14924 26852 15092 26908
rect 15372 26852 15540 26908
rect 14700 26338 14756 26348
rect 14924 26178 14980 26190
rect 14924 26126 14926 26178
rect 14978 26126 14980 26178
rect 14924 26068 14980 26126
rect 14924 26002 14980 26012
rect 14924 25732 14980 25742
rect 14700 25620 14756 25630
rect 14756 25564 14868 25620
rect 14700 25526 14756 25564
rect 14308 25004 14532 25060
rect 14252 24834 14308 25004
rect 14588 24948 14644 24958
rect 14588 24854 14644 24892
rect 14252 24782 14254 24834
rect 14306 24782 14308 24834
rect 14252 24770 14308 24782
rect 14028 24670 14030 24722
rect 14082 24670 14084 24722
rect 14028 24658 14084 24670
rect 14364 23380 14420 23390
rect 14364 23286 14420 23324
rect 14700 23042 14756 23054
rect 14700 22990 14702 23042
rect 14754 22990 14756 23042
rect 14588 22930 14644 22942
rect 14588 22878 14590 22930
rect 14642 22878 14644 22930
rect 14364 22482 14420 22494
rect 14364 22430 14366 22482
rect 14418 22430 14420 22482
rect 14364 22260 14420 22430
rect 13916 22094 13918 22146
rect 13970 22094 13972 22146
rect 13916 22036 13972 22094
rect 13916 21970 13972 21980
rect 14140 22204 14420 22260
rect 13580 21756 13972 21812
rect 13468 21534 13470 21586
rect 13522 21534 13524 21586
rect 13132 21474 13188 21486
rect 13132 21422 13134 21474
rect 13186 21422 13188 21474
rect 12908 20802 12964 20814
rect 12908 20750 12910 20802
rect 12962 20750 12964 20802
rect 12348 20578 12404 20590
rect 12348 20526 12350 20578
rect 12402 20526 12404 20578
rect 12348 20468 12404 20526
rect 12124 20412 12404 20468
rect 11900 19236 11956 19246
rect 11900 19142 11956 19180
rect 11676 18844 11844 18900
rect 11452 17490 11508 17500
rect 11564 18564 11620 18574
rect 11340 17154 11396 17164
rect 11116 14478 11118 14530
rect 11170 14478 11172 14530
rect 11116 14466 11172 14478
rect 11228 16884 11284 16894
rect 11228 16210 11284 16828
rect 11228 16158 11230 16210
rect 11282 16158 11284 16210
rect 11228 14532 11284 16158
rect 11564 15202 11620 18508
rect 11676 18452 11732 18844
rect 11788 18676 11844 18686
rect 12124 18676 12180 20412
rect 11788 18674 12180 18676
rect 11788 18622 11790 18674
rect 11842 18622 12180 18674
rect 11788 18620 12180 18622
rect 12236 20132 12292 20142
rect 11788 18610 11844 18620
rect 11676 18386 11732 18396
rect 12236 18450 12292 20076
rect 12348 19572 12404 19582
rect 12348 19234 12404 19516
rect 12796 19458 12852 19470
rect 12796 19406 12798 19458
rect 12850 19406 12852 19458
rect 12348 19182 12350 19234
rect 12402 19182 12404 19234
rect 12348 18564 12404 19182
rect 12348 18498 12404 18508
rect 12684 19236 12740 19246
rect 12236 18398 12238 18450
rect 12290 18398 12292 18450
rect 12236 18386 12292 18398
rect 12124 18116 12180 18126
rect 12124 17778 12180 18060
rect 12124 17726 12126 17778
rect 12178 17726 12180 17778
rect 12124 17714 12180 17726
rect 12348 17666 12404 17678
rect 12348 17614 12350 17666
rect 12402 17614 12404 17666
rect 12348 17556 12404 17614
rect 12348 17490 12404 17500
rect 11564 15150 11566 15202
rect 11618 15150 11620 15202
rect 11564 15138 11620 15150
rect 12124 17220 12180 17230
rect 12124 14642 12180 17164
rect 12684 16770 12740 19180
rect 12684 16718 12686 16770
rect 12738 16718 12740 16770
rect 12684 16706 12740 16718
rect 12684 16212 12740 16222
rect 12796 16212 12852 19406
rect 12908 19124 12964 20750
rect 13132 19348 13188 21422
rect 13468 20132 13524 21534
rect 13468 20066 13524 20076
rect 13692 20578 13748 20590
rect 13692 20526 13694 20578
rect 13746 20526 13748 20578
rect 13692 20132 13748 20526
rect 13132 19282 13188 19292
rect 13580 19460 13636 19470
rect 12908 19030 12964 19068
rect 12908 18340 12964 18350
rect 12908 18338 13412 18340
rect 12908 18286 12910 18338
rect 12962 18286 13412 18338
rect 12908 18284 13412 18286
rect 12908 18274 12964 18284
rect 12908 18116 12964 18126
rect 12908 17666 12964 18060
rect 12908 17614 12910 17666
rect 12962 17614 12964 17666
rect 12908 17602 12964 17614
rect 13356 17106 13412 18284
rect 13356 17054 13358 17106
rect 13410 17054 13412 17106
rect 13356 17042 13412 17054
rect 13468 16996 13524 17006
rect 13580 16996 13636 19404
rect 13692 18116 13748 20076
rect 13916 20020 13972 21756
rect 14028 20692 14084 20702
rect 14140 20692 14196 22204
rect 14588 22148 14644 22878
rect 14252 22092 14644 22148
rect 14252 21698 14308 22092
rect 14252 21646 14254 21698
rect 14306 21646 14308 21698
rect 14252 21634 14308 21646
rect 14252 21476 14308 21486
rect 14252 20802 14308 21420
rect 14252 20750 14254 20802
rect 14306 20750 14308 20802
rect 14252 20738 14308 20750
rect 14028 20690 14196 20692
rect 14028 20638 14030 20690
rect 14082 20638 14196 20690
rect 14028 20636 14196 20638
rect 14028 20626 14084 20636
rect 14140 20132 14196 20636
rect 14140 20076 14420 20132
rect 13916 19964 14084 20020
rect 13916 19796 13972 19806
rect 13916 19234 13972 19740
rect 13916 19182 13918 19234
rect 13970 19182 13972 19234
rect 13916 19170 13972 19182
rect 13692 18050 13748 18060
rect 14028 17890 14084 19964
rect 14028 17838 14030 17890
rect 14082 17838 14084 17890
rect 14028 17826 14084 17838
rect 14252 19684 14308 19694
rect 13692 17666 13748 17678
rect 13692 17614 13694 17666
rect 13746 17614 13748 17666
rect 13692 17332 13748 17614
rect 14252 17666 14308 19628
rect 14364 19234 14420 20076
rect 14588 19796 14644 19806
rect 14364 19182 14366 19234
rect 14418 19182 14420 19234
rect 14364 18228 14420 19182
rect 14476 19740 14588 19796
rect 14476 18228 14532 19740
rect 14588 19730 14644 19740
rect 14700 19458 14756 22990
rect 14812 22708 14868 25564
rect 14924 24946 14980 25676
rect 14924 24894 14926 24946
rect 14978 24894 14980 24946
rect 14924 24882 14980 24894
rect 15036 23940 15092 26852
rect 15372 26516 15428 26526
rect 15372 26290 15428 26460
rect 15372 26238 15374 26290
rect 15426 26238 15428 26290
rect 15148 25732 15204 25742
rect 15148 25506 15204 25676
rect 15148 25454 15150 25506
rect 15202 25454 15204 25506
rect 15148 25442 15204 25454
rect 15372 25508 15428 26238
rect 15372 24948 15428 25452
rect 15484 25506 15540 26852
rect 15484 25454 15486 25506
rect 15538 25454 15540 25506
rect 15484 25442 15540 25454
rect 15596 26402 15652 27804
rect 16380 27860 16436 27870
rect 16492 27860 16548 27918
rect 16380 27858 16548 27860
rect 16380 27806 16382 27858
rect 16434 27806 16548 27858
rect 16380 27804 16548 27806
rect 16380 27794 16436 27804
rect 16604 27186 16660 28700
rect 16828 28700 17164 28756
rect 16716 28084 16772 28094
rect 16716 27990 16772 28028
rect 16828 27970 16884 28700
rect 17164 28662 17220 28700
rect 16828 27918 16830 27970
rect 16882 27918 16884 27970
rect 16828 27906 16884 27918
rect 16604 27134 16606 27186
rect 16658 27134 16660 27186
rect 15596 26350 15598 26402
rect 15650 26350 15652 26402
rect 15484 24948 15540 24958
rect 15372 24946 15540 24948
rect 15372 24894 15486 24946
rect 15538 24894 15540 24946
rect 15372 24892 15540 24894
rect 15484 24882 15540 24892
rect 15036 23380 15092 23884
rect 15596 23716 15652 26350
rect 15820 27074 15876 27086
rect 15820 27022 15822 27074
rect 15874 27022 15876 27074
rect 15820 26068 15876 27022
rect 16268 26964 16324 26974
rect 15820 26002 15876 26012
rect 16156 26180 16212 26190
rect 15596 23650 15652 23660
rect 15148 23380 15204 23390
rect 14924 23378 15204 23380
rect 14924 23326 15150 23378
rect 15202 23326 15204 23378
rect 14924 23324 15204 23326
rect 14924 22932 14980 23324
rect 15148 23314 15204 23324
rect 16156 23380 16212 26124
rect 16268 25618 16324 26908
rect 16604 26516 16660 27134
rect 16940 26964 16996 27002
rect 16940 26898 16996 26908
rect 17052 26962 17108 26974
rect 17052 26910 17054 26962
rect 17106 26910 17108 26962
rect 16604 26450 16660 26460
rect 16828 26402 16884 26414
rect 16828 26350 16830 26402
rect 16882 26350 16884 26402
rect 16492 26290 16548 26302
rect 16492 26238 16494 26290
rect 16546 26238 16548 26290
rect 16492 26180 16548 26238
rect 16492 26114 16548 26124
rect 16268 25566 16270 25618
rect 16322 25566 16324 25618
rect 16268 25554 16324 25566
rect 16828 25508 16884 26350
rect 17052 26068 17108 26910
rect 17276 26964 17332 32732
rect 17612 32674 17668 33404
rect 17612 32622 17614 32674
rect 17666 32622 17668 32674
rect 17612 32610 17668 32622
rect 17724 32674 17780 32686
rect 17724 32622 17726 32674
rect 17778 32622 17780 32674
rect 17724 32564 17780 32622
rect 17500 31892 17556 31902
rect 17724 31892 17780 32508
rect 17556 31836 17780 31892
rect 17836 31892 17892 34972
rect 17948 34692 18004 35252
rect 18060 34914 18116 35644
rect 18172 35028 18228 42588
rect 18620 42532 18676 42542
rect 18620 42438 18676 42476
rect 18732 42084 18788 44044
rect 18844 42756 18900 45164
rect 19068 45108 19124 45118
rect 19068 45106 19684 45108
rect 19068 45054 19070 45106
rect 19122 45054 19684 45106
rect 19068 45052 19684 45054
rect 19068 45042 19124 45052
rect 19292 44548 19348 44558
rect 19628 44548 19684 45052
rect 19180 43540 19236 43550
rect 19180 43446 19236 43484
rect 19292 43428 19348 44492
rect 19516 44546 19684 44548
rect 19516 44494 19630 44546
rect 19682 44494 19684 44546
rect 19516 44492 19684 44494
rect 19404 44322 19460 44334
rect 19404 44270 19406 44322
rect 19458 44270 19460 44322
rect 19404 43988 19460 44270
rect 19404 43922 19460 43932
rect 19404 43428 19460 43438
rect 19292 43426 19460 43428
rect 19292 43374 19406 43426
rect 19458 43374 19460 43426
rect 19292 43372 19460 43374
rect 19404 43362 19460 43372
rect 19180 43204 19236 43214
rect 19180 42866 19236 43148
rect 19404 42980 19460 42990
rect 19516 42980 19572 44492
rect 19628 44482 19684 44492
rect 19852 44322 19908 45276
rect 19852 44270 19854 44322
rect 19906 44270 19908 44322
rect 19852 44258 19908 44270
rect 20188 44212 20244 44222
rect 20076 44100 20132 44138
rect 20076 44034 20132 44044
rect 19836 43932 20100 43942
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 19836 43866 20100 43876
rect 20188 43764 20244 44156
rect 20188 43698 20244 43708
rect 20524 43652 20580 45612
rect 20636 45666 20692 45678
rect 20636 45614 20638 45666
rect 20690 45614 20692 45666
rect 20636 45108 20692 45614
rect 20636 45042 20692 45052
rect 20748 44212 20804 44222
rect 20748 44118 20804 44156
rect 20524 43586 20580 43596
rect 20860 43316 20916 45724
rect 20972 45444 21028 47012
rect 20972 45378 21028 45388
rect 20636 43260 20916 43316
rect 19404 42978 19572 42980
rect 19404 42926 19406 42978
rect 19458 42926 19572 42978
rect 19404 42924 19572 42926
rect 19740 43204 19796 43214
rect 19740 42978 19796 43148
rect 19740 42926 19742 42978
rect 19794 42926 19796 42978
rect 19404 42914 19460 42924
rect 19740 42914 19796 42926
rect 20188 42980 20244 42990
rect 19180 42814 19182 42866
rect 19234 42814 19236 42866
rect 19180 42802 19236 42814
rect 18844 42308 18900 42700
rect 19964 42756 20020 42766
rect 19964 42662 20020 42700
rect 19836 42364 20100 42374
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 18844 42252 19124 42308
rect 19836 42298 20100 42308
rect 18844 42084 18900 42094
rect 18732 42082 18900 42084
rect 18732 42030 18846 42082
rect 18898 42030 18900 42082
rect 18732 42028 18900 42030
rect 18732 41074 18788 41086
rect 18732 41022 18734 41074
rect 18786 41022 18788 41074
rect 18620 40962 18676 40974
rect 18620 40910 18622 40962
rect 18674 40910 18676 40962
rect 18508 40628 18564 40638
rect 18284 40292 18340 40302
rect 18340 40236 18452 40292
rect 18284 40226 18340 40236
rect 18396 39060 18452 40236
rect 18508 39508 18564 40572
rect 18620 40514 18676 40910
rect 18620 40462 18622 40514
rect 18674 40462 18676 40514
rect 18620 40450 18676 40462
rect 18732 39732 18788 41022
rect 18732 39666 18788 39676
rect 18508 39452 18788 39508
rect 18508 39060 18564 39070
rect 18396 39058 18564 39060
rect 18396 39006 18510 39058
rect 18562 39006 18564 39058
rect 18396 39004 18564 39006
rect 18508 38994 18564 39004
rect 18284 38276 18340 38286
rect 18284 38162 18340 38220
rect 18284 38110 18286 38162
rect 18338 38110 18340 38162
rect 18284 38098 18340 38110
rect 18396 38050 18452 38062
rect 18396 37998 18398 38050
rect 18450 37998 18452 38050
rect 18396 37492 18452 37998
rect 18620 38050 18676 38062
rect 18620 37998 18622 38050
rect 18674 37998 18676 38050
rect 18620 37492 18676 37998
rect 18284 37436 18452 37492
rect 18508 37436 18676 37492
rect 18284 36708 18340 37436
rect 18396 37266 18452 37278
rect 18396 37214 18398 37266
rect 18450 37214 18452 37266
rect 18396 37156 18452 37214
rect 18396 37090 18452 37100
rect 18284 35700 18340 36652
rect 18396 35700 18452 35710
rect 18284 35698 18452 35700
rect 18284 35646 18398 35698
rect 18450 35646 18452 35698
rect 18284 35644 18452 35646
rect 18396 35634 18452 35644
rect 18172 34972 18452 35028
rect 18060 34862 18062 34914
rect 18114 34862 18116 34914
rect 18060 34850 18116 34862
rect 18284 34804 18340 34814
rect 18172 34802 18340 34804
rect 18172 34750 18286 34802
rect 18338 34750 18340 34802
rect 18172 34748 18340 34750
rect 18172 34692 18228 34748
rect 18284 34738 18340 34748
rect 17948 34636 18228 34692
rect 18396 33908 18452 34972
rect 18508 35026 18564 37436
rect 18620 37266 18676 37278
rect 18620 37214 18622 37266
rect 18674 37214 18676 37266
rect 18620 37156 18676 37214
rect 18620 37090 18676 37100
rect 18732 35812 18788 39452
rect 18844 38052 18900 42028
rect 19068 41970 19124 42252
rect 19068 41918 19070 41970
rect 19122 41918 19124 41970
rect 19068 41906 19124 41918
rect 20188 41858 20244 42924
rect 20188 41806 20190 41858
rect 20242 41806 20244 41858
rect 20188 41794 20244 41806
rect 19404 41188 19460 41198
rect 19964 41188 20020 41198
rect 19404 41186 19964 41188
rect 19404 41134 19406 41186
rect 19458 41134 19964 41186
rect 19404 41132 19964 41134
rect 19404 41122 19460 41132
rect 19964 41094 20020 41132
rect 19068 40962 19124 40974
rect 19068 40910 19070 40962
rect 19122 40910 19124 40962
rect 19068 40628 19124 40910
rect 19068 40562 19124 40572
rect 19628 40962 19684 40974
rect 19628 40910 19630 40962
rect 19682 40910 19684 40962
rect 19628 40068 19684 40910
rect 19852 40964 19908 41002
rect 19852 40898 19908 40908
rect 19836 40796 20100 40806
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 19836 40730 20100 40740
rect 19628 40002 19684 40012
rect 20412 40628 20468 40638
rect 20188 39844 20244 39854
rect 18956 39788 19684 39844
rect 18956 39730 19012 39788
rect 18956 39678 18958 39730
rect 19010 39678 19012 39730
rect 18956 39666 19012 39678
rect 19628 39732 19684 39788
rect 20076 39788 20188 39844
rect 19740 39732 19796 39742
rect 19628 39730 19796 39732
rect 19628 39678 19742 39730
rect 19794 39678 19796 39730
rect 19628 39676 19796 39678
rect 19740 39666 19796 39676
rect 19964 39732 20020 39742
rect 19964 39638 20020 39676
rect 19292 39618 19348 39630
rect 19292 39566 19294 39618
rect 19346 39566 19348 39618
rect 19292 39172 19348 39566
rect 19516 39620 19572 39630
rect 19516 39526 19572 39564
rect 19964 39508 20020 39518
rect 20076 39508 20132 39788
rect 20188 39778 20244 39788
rect 19964 39506 20132 39508
rect 19964 39454 19966 39506
rect 20018 39454 20132 39506
rect 19964 39452 20132 39454
rect 19964 39442 20020 39452
rect 20188 39394 20244 39406
rect 20188 39342 20190 39394
rect 20242 39342 20244 39394
rect 19836 39228 20100 39238
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 19836 39162 20100 39172
rect 19292 39106 19348 39116
rect 20188 39060 20244 39342
rect 20076 39004 20244 39060
rect 19852 38612 19908 38622
rect 18844 37986 18900 37996
rect 19516 38388 19572 38398
rect 19516 37940 19572 38332
rect 19852 38050 19908 38556
rect 19852 37998 19854 38050
rect 19906 37998 19908 38050
rect 19852 37986 19908 37998
rect 20076 38052 20132 39004
rect 20412 38834 20468 40572
rect 20412 38782 20414 38834
rect 20466 38782 20468 38834
rect 20412 38770 20468 38782
rect 20524 38500 20580 38510
rect 20188 38052 20244 38062
rect 20076 38050 20244 38052
rect 20076 37998 20190 38050
rect 20242 37998 20244 38050
rect 20076 37996 20244 37998
rect 19516 37938 19684 37940
rect 19516 37886 19518 37938
rect 19570 37886 19684 37938
rect 19516 37884 19684 37886
rect 19516 37874 19572 37884
rect 19292 37826 19348 37838
rect 19292 37774 19294 37826
rect 19346 37774 19348 37826
rect 19292 37716 19348 37774
rect 19292 37650 19348 37660
rect 18956 37492 19012 37502
rect 18956 37398 19012 37436
rect 18844 37266 18900 37278
rect 18844 37214 18846 37266
rect 18898 37214 18900 37266
rect 18844 36932 18900 37214
rect 18956 37156 19012 37166
rect 19404 37156 19460 37166
rect 18956 37154 19460 37156
rect 18956 37102 18958 37154
rect 19010 37102 19406 37154
rect 19458 37102 19460 37154
rect 18956 37100 19460 37102
rect 19628 37156 19684 37884
rect 19836 37660 20100 37670
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 19836 37594 20100 37604
rect 20076 37492 20132 37502
rect 20076 37268 20132 37436
rect 20076 37174 20132 37212
rect 19628 37100 19796 37156
rect 18956 37090 19012 37100
rect 19404 37090 19460 37100
rect 19516 37044 19572 37054
rect 19516 37042 19684 37044
rect 19516 36990 19518 37042
rect 19570 36990 19684 37042
rect 19516 36988 19684 36990
rect 19516 36978 19572 36988
rect 18844 36866 18900 36876
rect 19628 36594 19684 36988
rect 19628 36542 19630 36594
rect 19682 36542 19684 36594
rect 19628 36530 19684 36542
rect 19740 36260 19796 37100
rect 20188 37044 20244 37996
rect 20412 38052 20468 38062
rect 20412 37958 20468 37996
rect 20524 37828 20580 38444
rect 20188 36978 20244 36988
rect 20412 37772 20580 37828
rect 20412 36482 20468 37772
rect 20524 37492 20580 37502
rect 20524 37266 20580 37436
rect 20524 37214 20526 37266
rect 20578 37214 20580 37266
rect 20524 37202 20580 37214
rect 20412 36430 20414 36482
rect 20466 36430 20468 36482
rect 20412 36418 20468 36430
rect 20524 36932 20580 36942
rect 19628 36204 19796 36260
rect 18732 35756 18900 35812
rect 18508 34974 18510 35026
rect 18562 34974 18564 35026
rect 18508 34962 18564 34974
rect 18732 35588 18788 35598
rect 18732 34914 18788 35532
rect 18732 34862 18734 34914
rect 18786 34862 18788 34914
rect 18732 34850 18788 34862
rect 18060 33852 18452 33908
rect 18060 33460 18116 33852
rect 18060 33366 18116 33404
rect 18508 33572 18564 33582
rect 18844 33572 18900 35756
rect 18956 35810 19012 35822
rect 19404 35812 19460 35822
rect 18956 35758 18958 35810
rect 19010 35758 19012 35810
rect 18956 35140 19012 35758
rect 18956 35074 19012 35084
rect 19068 35756 19404 35812
rect 19068 35026 19124 35756
rect 19404 35718 19460 35756
rect 19068 34974 19070 35026
rect 19122 34974 19124 35026
rect 19068 34962 19124 34974
rect 19404 35476 19460 35486
rect 18844 33516 19012 33572
rect 18508 33460 18564 33516
rect 18508 33458 18788 33460
rect 18508 33406 18510 33458
rect 18562 33406 18788 33458
rect 18508 33404 18788 33406
rect 18508 33394 18564 33404
rect 18732 32786 18788 33404
rect 18732 32734 18734 32786
rect 18786 32734 18788 32786
rect 18732 32722 18788 32734
rect 18844 33348 18900 33358
rect 17948 32674 18004 32686
rect 17948 32622 17950 32674
rect 18002 32622 18004 32674
rect 17948 32564 18004 32622
rect 18060 32564 18116 32574
rect 17948 32562 18116 32564
rect 17948 32510 18062 32562
rect 18114 32510 18116 32562
rect 17948 32508 18116 32510
rect 18060 32498 18116 32508
rect 18508 32564 18564 32574
rect 18508 32470 18564 32508
rect 18620 32450 18676 32462
rect 18620 32398 18622 32450
rect 18674 32398 18676 32450
rect 18620 32004 18676 32398
rect 18844 32452 18900 33292
rect 18844 32386 18900 32396
rect 18620 31948 18900 32004
rect 17500 31826 17556 31836
rect 17836 31826 17892 31836
rect 18844 31890 18900 31948
rect 18844 31838 18846 31890
rect 18898 31838 18900 31890
rect 18844 31826 18900 31838
rect 18956 31668 19012 33516
rect 19292 33460 19348 33470
rect 19180 33124 19236 33134
rect 19292 33124 19348 33404
rect 19180 33122 19348 33124
rect 19180 33070 19182 33122
rect 19234 33070 19348 33122
rect 19180 33068 19348 33070
rect 19180 33058 19236 33068
rect 19180 32562 19236 32574
rect 19180 32510 19182 32562
rect 19234 32510 19236 32562
rect 19180 31780 19236 32510
rect 19180 31714 19236 31724
rect 18620 31612 19012 31668
rect 17612 31556 17668 31566
rect 17500 31108 17556 31118
rect 17500 31014 17556 31052
rect 17612 31106 17668 31500
rect 17612 31054 17614 31106
rect 17666 31054 17668 31106
rect 17612 31042 17668 31054
rect 17500 30772 17556 30782
rect 17500 30678 17556 30716
rect 18396 30098 18452 30110
rect 18396 30046 18398 30098
rect 18450 30046 18452 30098
rect 18284 29986 18340 29998
rect 18284 29934 18286 29986
rect 18338 29934 18340 29986
rect 17612 29314 17668 29326
rect 17612 29262 17614 29314
rect 17666 29262 17668 29314
rect 17500 28644 17556 28654
rect 17612 28644 17668 29262
rect 18284 28754 18340 29934
rect 18284 28702 18286 28754
rect 18338 28702 18340 28754
rect 18284 28690 18340 28702
rect 17556 28588 17668 28644
rect 17500 28550 17556 28588
rect 17500 28084 17556 28094
rect 17500 27990 17556 28028
rect 18284 27746 18340 27758
rect 18284 27694 18286 27746
rect 18338 27694 18340 27746
rect 17612 27412 17668 27422
rect 17612 27074 17668 27356
rect 17612 27022 17614 27074
rect 17666 27022 17668 27074
rect 17612 27010 17668 27022
rect 17388 26964 17444 26974
rect 17276 26962 17444 26964
rect 17276 26910 17390 26962
rect 17442 26910 17444 26962
rect 17276 26908 17444 26910
rect 17388 26292 17444 26908
rect 18284 26964 18340 27694
rect 18396 27298 18452 30046
rect 18396 27246 18398 27298
rect 18450 27246 18452 27298
rect 18396 27234 18452 27246
rect 18508 27634 18564 27646
rect 18508 27582 18510 27634
rect 18562 27582 18564 27634
rect 18284 26898 18340 26908
rect 18508 27186 18564 27582
rect 18508 27134 18510 27186
rect 18562 27134 18564 27186
rect 18508 26852 18564 27134
rect 18508 26786 18564 26796
rect 17388 26226 17444 26236
rect 17612 26628 17668 26638
rect 18620 26628 18676 31612
rect 19404 30324 19460 35420
rect 19628 33348 19684 36204
rect 19836 36092 20100 36102
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 19836 36026 20100 36036
rect 19740 35810 19796 35822
rect 20412 35812 20468 35822
rect 19740 35758 19742 35810
rect 19794 35758 19796 35810
rect 19740 35588 19796 35758
rect 19740 35522 19796 35532
rect 20300 35810 20468 35812
rect 20300 35758 20414 35810
rect 20466 35758 20468 35810
rect 20300 35756 20468 35758
rect 19836 34524 20100 34534
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 19836 34458 20100 34468
rect 19628 33254 19684 33292
rect 19852 33684 19908 33694
rect 19852 33124 19908 33628
rect 20300 33236 20356 35756
rect 20412 35746 20468 35756
rect 20412 34690 20468 34702
rect 20412 34638 20414 34690
rect 20466 34638 20468 34690
rect 20412 33684 20468 34638
rect 20412 33618 20468 33628
rect 20412 33236 20468 33246
rect 20300 33180 20412 33236
rect 20412 33170 20468 33180
rect 19628 33068 19908 33124
rect 19628 32788 19684 33068
rect 19836 32956 20100 32966
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20524 32900 20580 36876
rect 20636 36708 20692 43260
rect 20748 42980 20804 42990
rect 21084 42980 21140 47628
rect 21420 47572 21476 47582
rect 21644 47572 21700 48412
rect 22092 48466 22148 48478
rect 22092 48414 22094 48466
rect 22146 48414 22148 48466
rect 21756 48242 21812 48254
rect 21756 48190 21758 48242
rect 21810 48190 21812 48242
rect 21756 48132 21812 48190
rect 21756 48066 21812 48076
rect 21308 47516 21420 47572
rect 21308 47068 21364 47516
rect 21420 47506 21476 47516
rect 21532 47516 21700 47572
rect 21756 47684 21812 47694
rect 21532 47458 21588 47516
rect 21532 47406 21534 47458
rect 21586 47406 21588 47458
rect 21532 47394 21588 47406
rect 21756 47346 21812 47628
rect 21980 47572 22036 47582
rect 21980 47458 22036 47516
rect 21980 47406 21982 47458
rect 22034 47406 22036 47458
rect 21980 47394 22036 47406
rect 22092 47460 22148 48414
rect 22204 48354 22260 49646
rect 22204 48302 22206 48354
rect 22258 48302 22260 48354
rect 22204 48290 22260 48302
rect 22428 48244 22484 48254
rect 22428 47572 22484 48188
rect 22428 47506 22484 47516
rect 22876 48130 22932 48142
rect 22876 48078 22878 48130
rect 22930 48078 22932 48130
rect 22652 47460 22708 47470
rect 22876 47460 22932 48078
rect 22092 47404 22260 47460
rect 21756 47294 21758 47346
rect 21810 47294 21812 47346
rect 21756 47282 21812 47294
rect 21868 47236 21924 47246
rect 21868 47234 22036 47236
rect 21868 47182 21870 47234
rect 21922 47182 22036 47234
rect 21868 47180 22036 47182
rect 21868 47170 21924 47180
rect 21980 47068 22036 47180
rect 21308 47012 21588 47068
rect 21308 46674 21364 46686
rect 21308 46622 21310 46674
rect 21362 46622 21364 46674
rect 21308 45668 21364 46622
rect 21532 46114 21588 47012
rect 21756 47012 22036 47068
rect 22092 47234 22148 47246
rect 22092 47182 22094 47234
rect 22146 47182 22148 47234
rect 21756 46900 21812 47012
rect 21532 46062 21534 46114
rect 21586 46062 21588 46114
rect 21532 46050 21588 46062
rect 21644 46844 21812 46900
rect 22092 46900 22148 47182
rect 21420 45780 21476 45790
rect 21420 45778 21588 45780
rect 21420 45726 21422 45778
rect 21474 45726 21588 45778
rect 21420 45724 21588 45726
rect 21420 45714 21476 45724
rect 21308 45602 21364 45612
rect 21420 45332 21476 45342
rect 21308 45108 21364 45118
rect 21308 44546 21364 45052
rect 21308 44494 21310 44546
rect 21362 44494 21364 44546
rect 21308 44482 21364 44494
rect 21420 44434 21476 45276
rect 21532 44548 21588 45724
rect 21532 44482 21588 44492
rect 21420 44382 21422 44434
rect 21474 44382 21476 44434
rect 21420 44370 21476 44382
rect 21532 44100 21588 44110
rect 21532 44006 21588 44044
rect 21532 43652 21588 43662
rect 21644 43652 21700 46844
rect 22092 46834 22148 46844
rect 21756 46676 21812 46686
rect 21756 46562 21812 46620
rect 21756 46510 21758 46562
rect 21810 46510 21812 46562
rect 21756 46498 21812 46510
rect 21980 45892 22036 45902
rect 22204 45892 22260 47404
rect 22708 47404 22932 47460
rect 23324 47458 23380 50372
rect 23660 49026 23716 49038
rect 23660 48974 23662 49026
rect 23714 48974 23716 49026
rect 23660 48132 23716 48974
rect 23772 48468 23828 48478
rect 23772 48374 23828 48412
rect 23660 48066 23716 48076
rect 23324 47406 23326 47458
rect 23378 47406 23380 47458
rect 22652 47366 22708 47404
rect 23324 47394 23380 47406
rect 23100 47348 23156 47358
rect 22540 47236 22596 47246
rect 21980 45890 22260 45892
rect 21980 45838 21982 45890
rect 22034 45838 22260 45890
rect 21980 45836 22260 45838
rect 22316 47234 22596 47236
rect 22316 47182 22542 47234
rect 22594 47182 22596 47234
rect 22316 47180 22596 47182
rect 22316 45890 22372 47180
rect 22540 47170 22596 47180
rect 22428 46900 22484 46910
rect 22484 46844 22596 46900
rect 22428 46834 22484 46844
rect 22428 46564 22484 46574
rect 22428 46002 22484 46508
rect 22428 45950 22430 46002
rect 22482 45950 22484 46002
rect 22428 45938 22484 45950
rect 22316 45838 22318 45890
rect 22370 45838 22372 45890
rect 21980 45826 22036 45836
rect 22316 45826 22372 45838
rect 22540 45892 22596 46844
rect 21532 43650 21700 43652
rect 21532 43598 21534 43650
rect 21586 43598 21700 43650
rect 21532 43596 21700 43598
rect 21756 45668 21812 45678
rect 21756 44994 21812 45612
rect 22092 45668 22148 45678
rect 22092 45574 22148 45612
rect 21756 44942 21758 44994
rect 21810 44942 21812 44994
rect 21532 43586 21588 43596
rect 20748 42866 20804 42924
rect 20748 42814 20750 42866
rect 20802 42814 20804 42866
rect 20748 42802 20804 42814
rect 20972 42924 21140 42980
rect 21308 43316 21364 43326
rect 20748 40964 20804 40974
rect 20748 40290 20804 40908
rect 20748 40238 20750 40290
rect 20802 40238 20804 40290
rect 20748 40226 20804 40238
rect 20748 39844 20804 39854
rect 20748 39730 20804 39788
rect 20748 39678 20750 39730
rect 20802 39678 20804 39730
rect 20748 39666 20804 39678
rect 20748 39172 20804 39182
rect 20748 38274 20804 39116
rect 20860 38948 20916 38958
rect 20860 38834 20916 38892
rect 20860 38782 20862 38834
rect 20914 38782 20916 38834
rect 20860 38770 20916 38782
rect 20748 38222 20750 38274
rect 20802 38222 20804 38274
rect 20748 38210 20804 38222
rect 20860 38610 20916 38622
rect 20860 38558 20862 38610
rect 20914 38558 20916 38610
rect 20860 37828 20916 38558
rect 20972 38276 21028 42924
rect 21084 42756 21140 42766
rect 21084 40628 21140 42700
rect 21084 40534 21140 40572
rect 21308 42084 21364 43260
rect 21644 43316 21700 43326
rect 21756 43316 21812 44942
rect 21700 43260 21812 43316
rect 21868 45444 21924 45454
rect 21644 43250 21700 43260
rect 21868 43204 21924 45388
rect 22092 44548 22148 44558
rect 22092 44434 22148 44492
rect 22092 44382 22094 44434
rect 22146 44382 22148 44434
rect 22092 44370 22148 44382
rect 22204 43538 22260 43550
rect 22204 43486 22206 43538
rect 22258 43486 22260 43538
rect 22204 43316 22260 43486
rect 22540 43540 22596 45836
rect 22652 44324 22708 44334
rect 22652 44230 22708 44268
rect 23100 44100 23156 47292
rect 23660 47348 23716 47358
rect 23660 47254 23716 47292
rect 23212 47234 23268 47246
rect 23212 47182 23214 47234
rect 23266 47182 23268 47234
rect 23212 45890 23268 47182
rect 23884 47236 23940 50428
rect 23884 47170 23940 47180
rect 23996 50372 24164 50428
rect 23884 46564 23940 46574
rect 23660 46562 23940 46564
rect 23660 46510 23886 46562
rect 23938 46510 23940 46562
rect 23660 46508 23940 46510
rect 23212 45838 23214 45890
rect 23266 45838 23268 45890
rect 23212 45826 23268 45838
rect 23548 46452 23604 46462
rect 23548 45890 23604 46396
rect 23660 46002 23716 46508
rect 23884 46498 23940 46508
rect 23660 45950 23662 46002
rect 23714 45950 23716 46002
rect 23660 45938 23716 45950
rect 23548 45838 23550 45890
rect 23602 45838 23604 45890
rect 23548 45826 23604 45838
rect 23772 45892 23828 45902
rect 23772 45798 23828 45836
rect 23324 45668 23380 45678
rect 23324 45574 23380 45612
rect 23212 45108 23268 45118
rect 23212 44324 23268 45052
rect 23996 44324 24052 50372
rect 24332 49588 24388 49598
rect 24332 49138 24388 49532
rect 24332 49086 24334 49138
rect 24386 49086 24388 49138
rect 24332 49074 24388 49086
rect 24444 48580 24500 52668
rect 24892 52388 24948 54572
rect 24780 52332 24948 52388
rect 24444 48524 24612 48580
rect 24220 48468 24276 48478
rect 24220 48244 24276 48412
rect 24220 48242 24388 48244
rect 24220 48190 24222 48242
rect 24274 48190 24388 48242
rect 24220 48188 24388 48190
rect 24220 48178 24276 48188
rect 24220 47348 24276 47358
rect 23212 44258 23268 44268
rect 23884 44268 24052 44324
rect 24108 44436 24164 44446
rect 23100 44044 23268 44100
rect 22652 43540 22708 43550
rect 22876 43540 22932 43550
rect 22540 43538 22708 43540
rect 22540 43486 22654 43538
rect 22706 43486 22708 43538
rect 22540 43484 22708 43486
rect 22652 43474 22708 43484
rect 22764 43538 22932 43540
rect 22764 43486 22878 43538
rect 22930 43486 22932 43538
rect 22764 43484 22932 43486
rect 22204 43250 22260 43260
rect 21756 43148 21924 43204
rect 21644 42530 21700 42542
rect 21644 42478 21646 42530
rect 21698 42478 21700 42530
rect 21644 42420 21700 42478
rect 21756 42532 21812 43148
rect 22764 43092 22820 43484
rect 22876 43474 22932 43484
rect 23100 43538 23156 43550
rect 23100 43486 23102 43538
rect 23154 43486 23156 43538
rect 22092 43036 22820 43092
rect 22988 43426 23044 43438
rect 22988 43374 22990 43426
rect 23042 43374 23044 43426
rect 22092 42978 22148 43036
rect 22092 42926 22094 42978
rect 22146 42926 22148 42978
rect 22092 42914 22148 42926
rect 21980 42868 22036 42878
rect 22988 42868 23044 43374
rect 23100 42980 23156 43486
rect 23100 42914 23156 42924
rect 21980 42774 22036 42812
rect 22316 42812 23044 42868
rect 21756 42476 21924 42532
rect 21644 42354 21700 42364
rect 20972 38210 21028 38220
rect 21084 38948 21140 38958
rect 20860 37762 20916 37772
rect 20972 37378 21028 37390
rect 20972 37326 20974 37378
rect 21026 37326 21028 37378
rect 20860 37156 20916 37166
rect 20860 37062 20916 37100
rect 20972 37044 21028 37326
rect 20972 36978 21028 36988
rect 21084 36820 21140 38892
rect 21308 38834 21364 42028
rect 21868 41972 21924 42476
rect 22316 42082 22372 42812
rect 22428 42642 22484 42654
rect 22428 42590 22430 42642
rect 22482 42590 22484 42642
rect 22428 42420 22484 42590
rect 22764 42532 22820 42542
rect 23100 42532 23156 42542
rect 22764 42530 23156 42532
rect 22764 42478 22766 42530
rect 22818 42478 23102 42530
rect 23154 42478 23156 42530
rect 22764 42476 23156 42478
rect 22764 42466 22820 42476
rect 22540 42420 22596 42430
rect 22428 42364 22540 42420
rect 22540 42354 22596 42364
rect 22316 42030 22318 42082
rect 22370 42030 22372 42082
rect 22316 42018 22372 42030
rect 21980 41972 22036 41982
rect 21868 41916 21980 41972
rect 21980 41906 22036 41916
rect 22652 41860 22708 41870
rect 21532 41412 21588 41422
rect 21420 40964 21476 40974
rect 21420 40626 21476 40908
rect 21420 40574 21422 40626
rect 21474 40574 21476 40626
rect 21420 40562 21476 40574
rect 21532 40068 21588 41356
rect 21980 41300 22036 41310
rect 21980 41206 22036 41244
rect 21868 41074 21924 41086
rect 21868 41022 21870 41074
rect 21922 41022 21924 41074
rect 21868 40964 21924 41022
rect 22652 41076 22708 41804
rect 22876 41636 22932 42476
rect 23100 42466 23156 42476
rect 23212 42308 23268 44044
rect 23884 43876 23940 44268
rect 23996 44100 24052 44110
rect 24108 44100 24164 44380
rect 24220 44212 24276 47292
rect 24220 44146 24276 44156
rect 23996 44098 24164 44100
rect 23996 44046 23998 44098
rect 24050 44046 24164 44098
rect 23996 44044 24164 44046
rect 23996 44034 24052 44044
rect 23884 43820 24052 43876
rect 23324 43540 23380 43550
rect 23324 43446 23380 43484
rect 23772 43538 23828 43550
rect 23772 43486 23774 43538
rect 23826 43486 23828 43538
rect 22988 42252 23268 42308
rect 23324 42980 23380 42990
rect 22988 41860 23044 42252
rect 23100 41972 23156 41982
rect 23100 41970 23268 41972
rect 23100 41918 23102 41970
rect 23154 41918 23268 41970
rect 23100 41916 23268 41918
rect 23100 41906 23156 41916
rect 22988 41794 23044 41804
rect 22876 41580 23044 41636
rect 22652 40982 22708 41020
rect 22988 41076 23044 41580
rect 22988 40982 23044 41020
rect 23100 41188 23156 41198
rect 21868 40898 21924 40908
rect 23100 40628 23156 41132
rect 23100 40534 23156 40572
rect 22092 40514 22148 40526
rect 22092 40462 22094 40514
rect 22146 40462 22148 40514
rect 21308 38782 21310 38834
rect 21362 38782 21364 38834
rect 21308 38770 21364 38782
rect 21420 40012 21588 40068
rect 21868 40402 21924 40414
rect 21868 40350 21870 40402
rect 21922 40350 21924 40402
rect 21420 39730 21476 40012
rect 21420 39678 21422 39730
rect 21474 39678 21476 39730
rect 21420 38668 21476 39678
rect 21196 38612 21476 38668
rect 21532 39844 21588 39854
rect 21196 37378 21252 38612
rect 21196 37326 21198 37378
rect 21250 37326 21252 37378
rect 21196 37268 21252 37326
rect 21196 37202 21252 37212
rect 21308 37492 21364 37502
rect 20636 36642 20692 36652
rect 20748 36764 21140 36820
rect 20636 36260 20692 36270
rect 20636 34802 20692 36204
rect 20748 35922 20804 36764
rect 21308 36708 21364 37436
rect 20748 35870 20750 35922
rect 20802 35870 20804 35922
rect 20748 35858 20804 35870
rect 21196 36652 21364 36708
rect 20636 34750 20638 34802
rect 20690 34750 20692 34802
rect 20636 34738 20692 34750
rect 20748 34804 20804 34814
rect 20748 34710 20804 34748
rect 19836 32890 20100 32900
rect 20300 32844 20580 32900
rect 20636 33572 20692 33582
rect 19628 32732 19908 32788
rect 19852 32674 19908 32732
rect 19852 32622 19854 32674
rect 19906 32622 19908 32674
rect 19852 32610 19908 32622
rect 19628 31780 19684 31790
rect 19628 30996 19684 31724
rect 19836 31388 20100 31398
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 19836 31322 20100 31332
rect 20076 30996 20132 31006
rect 19628 30994 20132 30996
rect 19628 30942 20078 30994
rect 20130 30942 20132 30994
rect 19628 30940 20132 30942
rect 19460 30268 19796 30324
rect 19404 30230 19460 30268
rect 19740 30210 19796 30268
rect 19740 30158 19742 30210
rect 19794 30158 19796 30210
rect 19740 30146 19796 30158
rect 18956 30100 19012 30110
rect 18956 28756 19012 30044
rect 18844 27746 18900 27758
rect 18844 27694 18846 27746
rect 18898 27694 18900 27746
rect 18844 27634 18900 27694
rect 18844 27582 18846 27634
rect 18898 27582 18900 27634
rect 18844 27570 18900 27582
rect 18956 27412 19012 28700
rect 19068 29988 19124 29998
rect 19068 28644 19124 29932
rect 20076 29988 20132 30940
rect 20076 29922 20132 29932
rect 20300 30210 20356 32844
rect 20300 30158 20302 30210
rect 20354 30158 20356 30210
rect 19836 29820 20100 29830
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 19836 29754 20100 29764
rect 19068 27858 19124 28588
rect 19068 27806 19070 27858
rect 19122 27806 19124 27858
rect 19068 27794 19124 27806
rect 19628 28644 19684 28654
rect 18844 27356 19012 27412
rect 18844 27074 18900 27356
rect 18844 27022 18846 27074
rect 18898 27022 18900 27074
rect 18844 27010 18900 27022
rect 19628 27074 19684 28588
rect 19836 28252 20100 28262
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 19836 28186 20100 28196
rect 19852 27748 19908 27758
rect 19852 27654 19908 27692
rect 19628 27022 19630 27074
rect 19682 27022 19684 27074
rect 17612 26290 17668 26572
rect 18508 26572 18676 26628
rect 18732 26964 18788 26974
rect 17612 26238 17614 26290
rect 17666 26238 17668 26290
rect 17612 26226 17668 26238
rect 18060 26292 18116 26302
rect 18060 26198 18116 26236
rect 18508 26180 18564 26572
rect 17052 26002 17108 26012
rect 17948 26068 18004 26078
rect 18172 26068 18228 26078
rect 17948 25974 18004 26012
rect 18060 26012 18172 26068
rect 16828 25442 16884 25452
rect 18060 24834 18116 26012
rect 18172 26002 18228 26012
rect 18396 25620 18452 25630
rect 18396 25526 18452 25564
rect 18060 24782 18062 24834
rect 18114 24782 18116 24834
rect 18060 24770 18116 24782
rect 17724 24612 17780 24622
rect 17276 23940 17332 23950
rect 17276 23846 17332 23884
rect 17724 23940 17780 24556
rect 17724 23874 17780 23884
rect 18172 24498 18228 24510
rect 18172 24446 18174 24498
rect 18226 24446 18228 24498
rect 16156 23314 16212 23324
rect 18172 23266 18228 24446
rect 18508 24498 18564 26124
rect 18732 26068 18788 26908
rect 19068 26852 19124 26862
rect 18844 26628 18900 26638
rect 18844 26290 18900 26572
rect 18844 26238 18846 26290
rect 18898 26238 18900 26290
rect 18844 26226 18900 26238
rect 19068 26404 19124 26796
rect 19068 26290 19124 26348
rect 19068 26238 19070 26290
rect 19122 26238 19124 26290
rect 19068 26226 19124 26238
rect 19180 26740 19236 26750
rect 19180 26180 19236 26684
rect 19628 26628 19684 27022
rect 20076 26964 20132 27002
rect 20300 26908 20356 30158
rect 20524 32676 20580 32686
rect 20412 28756 20468 28766
rect 20412 28662 20468 28700
rect 20076 26852 20356 26908
rect 19836 26684 20100 26694
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 19836 26618 20100 26628
rect 19628 26562 19684 26572
rect 20188 26516 20244 26852
rect 20076 26460 20244 26516
rect 20076 26402 20132 26460
rect 20076 26350 20078 26402
rect 20130 26350 20132 26402
rect 20076 26338 20132 26350
rect 18732 26012 19124 26068
rect 19068 25618 19124 26012
rect 19068 25566 19070 25618
rect 19122 25566 19124 25618
rect 19068 25554 19124 25566
rect 18732 25508 18788 25518
rect 18732 24946 18788 25452
rect 18732 24894 18734 24946
rect 18786 24894 18788 24946
rect 18732 24882 18788 24894
rect 19180 24946 19236 26124
rect 19516 26290 19572 26302
rect 19516 26238 19518 26290
rect 19570 26238 19572 26290
rect 19516 25620 19572 26238
rect 20412 26292 20468 26302
rect 20412 26198 20468 26236
rect 19740 25844 19796 25854
rect 19740 25620 19796 25788
rect 19516 25554 19572 25564
rect 19628 25618 19796 25620
rect 19628 25566 19742 25618
rect 19794 25566 19796 25618
rect 19628 25564 19796 25566
rect 19404 25508 19460 25518
rect 19404 25414 19460 25452
rect 19180 24894 19182 24946
rect 19234 24894 19236 24946
rect 19180 24882 19236 24894
rect 19628 24610 19684 25564
rect 19740 25554 19796 25564
rect 20188 25284 20244 25294
rect 19836 25116 20100 25126
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 19836 25050 20100 25060
rect 19964 24948 20020 24958
rect 20188 24948 20244 25228
rect 19964 24946 20244 24948
rect 19964 24894 19966 24946
rect 20018 24894 20244 24946
rect 19964 24892 20244 24894
rect 19964 24882 20020 24892
rect 19628 24558 19630 24610
rect 19682 24558 19684 24610
rect 18508 24446 18510 24498
rect 18562 24446 18564 24498
rect 18508 24434 18564 24446
rect 19292 24498 19348 24510
rect 19292 24446 19294 24498
rect 19346 24446 19348 24498
rect 19068 23940 19124 23950
rect 19068 23826 19124 23884
rect 19292 23938 19348 24446
rect 19292 23886 19294 23938
rect 19346 23886 19348 23938
rect 19292 23874 19348 23886
rect 19068 23774 19070 23826
rect 19122 23774 19124 23826
rect 18172 23214 18174 23266
rect 18226 23214 18228 23266
rect 18172 23202 18228 23214
rect 18508 23268 18564 23278
rect 17500 23154 17556 23166
rect 17500 23102 17502 23154
rect 17554 23102 17556 23154
rect 16716 23044 16772 23054
rect 14924 22866 14980 22876
rect 16604 23042 16772 23044
rect 16604 22990 16718 23042
rect 16770 22990 16772 23042
rect 16604 22988 16772 22990
rect 14812 22652 15092 22708
rect 14812 22482 14868 22494
rect 14812 22430 14814 22482
rect 14866 22430 14868 22482
rect 14812 20804 14868 22430
rect 14812 20738 14868 20748
rect 14924 22484 14980 22494
rect 14812 20020 14868 20030
rect 14924 20020 14980 22428
rect 15036 20132 15092 22652
rect 15148 22036 15204 22046
rect 15148 20242 15204 21980
rect 16380 21474 16436 21486
rect 16380 21422 16382 21474
rect 16434 21422 16436 21474
rect 16380 21028 16436 21422
rect 15932 20972 16436 21028
rect 16604 21026 16660 22988
rect 16716 22978 16772 22988
rect 16828 22932 16884 22942
rect 16828 22930 16996 22932
rect 16828 22878 16830 22930
rect 16882 22878 16996 22930
rect 16828 22876 16996 22878
rect 16828 22866 16884 22876
rect 16940 22482 16996 22876
rect 16940 22430 16942 22482
rect 16994 22430 16996 22482
rect 16940 22418 16996 22430
rect 17500 22372 17556 23102
rect 17724 22372 17780 22382
rect 17500 22370 17780 22372
rect 17500 22318 17726 22370
rect 17778 22318 17780 22370
rect 17500 22316 17780 22318
rect 17724 21700 17780 22316
rect 18396 22372 18452 22382
rect 18396 22278 18452 22316
rect 18172 21812 18228 21822
rect 17724 21634 17780 21644
rect 17948 21756 18172 21812
rect 16604 20974 16606 21026
rect 16658 20974 16660 21026
rect 15148 20190 15150 20242
rect 15202 20190 15204 20242
rect 15148 20178 15204 20190
rect 15372 20802 15428 20814
rect 15372 20750 15374 20802
rect 15426 20750 15428 20802
rect 15036 20066 15092 20076
rect 15372 20020 15428 20750
rect 15708 20804 15764 20814
rect 15932 20804 15988 20972
rect 16604 20962 16660 20974
rect 16716 21474 16772 21486
rect 16716 21422 16718 21474
rect 16770 21422 16772 21474
rect 15708 20802 15988 20804
rect 15708 20750 15710 20802
rect 15762 20750 15988 20802
rect 15708 20748 15988 20750
rect 16044 20802 16100 20814
rect 16044 20750 16046 20802
rect 16098 20750 16100 20802
rect 15708 20738 15764 20748
rect 14812 20018 14980 20020
rect 14812 19966 14814 20018
rect 14866 19966 14980 20018
rect 14812 19964 14980 19966
rect 15260 19964 15372 20020
rect 14812 19954 14868 19964
rect 15260 19460 15316 19964
rect 15372 19954 15428 19964
rect 15708 19908 15764 19918
rect 15708 19684 15764 19852
rect 15708 19618 15764 19628
rect 14700 19406 14702 19458
rect 14754 19406 14756 19458
rect 14700 19394 14756 19406
rect 14924 19404 15316 19460
rect 14588 19348 14644 19358
rect 14588 19254 14644 19292
rect 14924 19236 14980 19404
rect 15484 19348 15540 19358
rect 14812 19234 14980 19236
rect 14812 19182 14926 19234
rect 14978 19182 14980 19234
rect 14812 19180 14980 19182
rect 14476 18172 14756 18228
rect 14364 18162 14420 18172
rect 14252 17614 14254 17666
rect 14306 17614 14308 17666
rect 14252 17602 14308 17614
rect 13692 17266 13748 17276
rect 13468 16994 13636 16996
rect 13468 16942 13470 16994
rect 13522 16942 13636 16994
rect 13468 16940 13636 16942
rect 14700 16994 14756 18172
rect 14812 17666 14868 19180
rect 14924 19170 14980 19180
rect 15036 19236 15092 19246
rect 15036 18340 15092 19180
rect 14812 17614 14814 17666
rect 14866 17614 14868 17666
rect 14812 17602 14868 17614
rect 14924 18338 15092 18340
rect 14924 18286 15038 18338
rect 15090 18286 15092 18338
rect 14924 18284 15092 18286
rect 14924 17668 14980 18284
rect 15036 18274 15092 18284
rect 15372 18338 15428 18350
rect 15372 18286 15374 18338
rect 15426 18286 15428 18338
rect 15148 17668 15204 17678
rect 14924 17666 15204 17668
rect 14924 17614 15150 17666
rect 15202 17614 15204 17666
rect 14924 17612 15204 17614
rect 15148 17602 15204 17612
rect 14700 16942 14702 16994
rect 14754 16942 14756 16994
rect 13468 16930 13524 16940
rect 14700 16930 14756 16942
rect 12684 16210 12852 16212
rect 12684 16158 12686 16210
rect 12738 16158 12852 16210
rect 12684 16156 12852 16158
rect 14028 16882 14084 16894
rect 14028 16830 14030 16882
rect 14082 16830 14084 16882
rect 12684 16146 12740 16156
rect 14028 16100 14084 16830
rect 14476 16100 14532 16110
rect 14028 16098 14532 16100
rect 14028 16046 14478 16098
rect 14530 16046 14532 16098
rect 14028 16044 14532 16046
rect 12796 15876 12852 15886
rect 12796 15782 12852 15820
rect 13692 15876 13748 15886
rect 13692 15426 13748 15820
rect 13692 15374 13694 15426
rect 13746 15374 13748 15426
rect 13692 15362 13748 15374
rect 14476 15316 14532 16044
rect 15148 15988 15204 15998
rect 15148 15894 15204 15932
rect 14476 15222 14532 15260
rect 12124 14590 12126 14642
rect 12178 14590 12180 14642
rect 12124 14578 12180 14590
rect 11228 14466 11284 14476
rect 11900 14532 11956 14542
rect 11900 14438 11956 14476
rect 4476 13356 4740 13366
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4476 13290 4740 13300
rect 4476 11788 4740 11798
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4476 11722 4740 11732
rect 4476 10220 4740 10230
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4476 10154 4740 10164
rect 4476 8652 4740 8662
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4476 8586 4740 8596
rect 15372 8428 15428 18286
rect 15484 18004 15540 19292
rect 15820 19234 15876 20748
rect 16044 20692 16100 20750
rect 15820 19182 15822 19234
rect 15874 19182 15876 19234
rect 15820 19170 15876 19182
rect 15932 20636 16044 20692
rect 15596 18228 15652 18238
rect 15596 18134 15652 18172
rect 15932 18116 15988 20636
rect 16044 20598 16100 20636
rect 16156 20804 16212 20814
rect 16044 20132 16100 20142
rect 16044 20038 16100 20076
rect 16156 19796 16212 20748
rect 16716 20244 16772 21422
rect 17612 21474 17668 21486
rect 17612 21422 17614 21474
rect 17666 21422 17668 21474
rect 16828 21362 16884 21374
rect 16828 21310 16830 21362
rect 16882 21310 16884 21362
rect 16828 20916 16884 21310
rect 16828 20850 16884 20860
rect 17164 20804 17220 20814
rect 17164 20802 17332 20804
rect 17164 20750 17166 20802
rect 17218 20750 17332 20802
rect 17164 20748 17332 20750
rect 17164 20738 17220 20748
rect 16716 20178 16772 20188
rect 16044 19740 16212 19796
rect 16604 20020 16660 20030
rect 16604 19906 16660 19964
rect 16604 19854 16606 19906
rect 16658 19854 16660 19906
rect 16044 18450 16100 19740
rect 16604 19684 16660 19854
rect 16604 19618 16660 19628
rect 16828 19460 16884 19470
rect 16828 19366 16884 19404
rect 16940 19236 16996 19246
rect 16940 19142 16996 19180
rect 16044 18398 16046 18450
rect 16098 18398 16100 18450
rect 16044 18386 16100 18398
rect 16156 19124 16212 19134
rect 16380 19124 16436 19134
rect 16716 19124 16772 19134
rect 16212 19122 16772 19124
rect 16212 19070 16382 19122
rect 16434 19070 16718 19122
rect 16770 19070 16772 19122
rect 16212 19068 16772 19070
rect 15932 18050 15988 18060
rect 15484 17948 15652 18004
rect 15596 17666 15652 17948
rect 16156 17778 16212 19068
rect 16380 19058 16436 19068
rect 16716 19058 16772 19068
rect 16828 19012 16884 19022
rect 16380 18620 16772 18676
rect 16268 18450 16324 18462
rect 16268 18398 16270 18450
rect 16322 18398 16324 18450
rect 16268 18340 16324 18398
rect 16268 18274 16324 18284
rect 16156 17726 16158 17778
rect 16210 17726 16212 17778
rect 16156 17714 16212 17726
rect 16380 18116 16436 18620
rect 16492 18452 16548 18490
rect 16548 18396 16660 18452
rect 16492 18386 16548 18396
rect 15596 17614 15598 17666
rect 15650 17614 15652 17666
rect 15596 17602 15652 17614
rect 16380 17444 16436 18060
rect 16492 18228 16548 18238
rect 16492 17666 16548 18172
rect 16492 17614 16494 17666
rect 16546 17614 16548 17666
rect 16492 17602 16548 17614
rect 16492 17444 16548 17454
rect 16380 17388 16492 17444
rect 16492 17378 16548 17388
rect 16604 16884 16660 18396
rect 16716 18450 16772 18620
rect 16716 18398 16718 18450
rect 16770 18398 16772 18450
rect 16716 18386 16772 18398
rect 16716 18228 16772 18238
rect 16828 18228 16884 18956
rect 16716 18226 16884 18228
rect 16716 18174 16718 18226
rect 16770 18174 16884 18226
rect 16716 18172 16884 18174
rect 16716 18162 16772 18172
rect 17052 17892 17108 17902
rect 16828 17890 17108 17892
rect 16828 17838 17054 17890
rect 17106 17838 17108 17890
rect 16828 17836 17108 17838
rect 16828 16996 16884 17836
rect 17052 17826 17108 17836
rect 16940 17668 16996 17678
rect 16940 17666 17108 17668
rect 16940 17614 16942 17666
rect 16994 17614 17108 17666
rect 16940 17612 17108 17614
rect 16940 17602 16996 17612
rect 16828 16940 16996 16996
rect 16604 16828 16884 16884
rect 16828 16770 16884 16828
rect 16828 16718 16830 16770
rect 16882 16718 16884 16770
rect 16828 16706 16884 16718
rect 16604 15988 16660 15998
rect 16660 15932 16772 15988
rect 16604 15922 16660 15932
rect 16380 15540 16436 15550
rect 15372 8372 16100 8428
rect 4476 7084 4740 7094
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4476 7018 4740 7028
rect 4476 5516 4740 5526
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4476 5450 4740 5460
rect 4476 3948 4740 3958
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4476 3882 4740 3892
rect 12684 3444 12740 3454
rect 13132 3444 13188 3454
rect 12684 3442 13188 3444
rect 12684 3390 12686 3442
rect 12738 3390 13134 3442
rect 13186 3390 13188 3442
rect 12684 3388 13188 3390
rect 12684 3378 12740 3388
rect 12796 800 12852 3388
rect 13132 3378 13188 3388
rect 13468 3444 13524 3454
rect 13468 3350 13524 3388
rect 15820 3442 15876 3454
rect 15820 3390 15822 3442
rect 15874 3390 15876 3442
rect 15820 3220 15876 3390
rect 16044 3442 16100 8372
rect 16268 3556 16324 3566
rect 16044 3390 16046 3442
rect 16098 3390 16100 3442
rect 16044 3378 16100 3390
rect 16156 3554 16324 3556
rect 16156 3502 16270 3554
rect 16322 3502 16324 3554
rect 16156 3500 16324 3502
rect 16156 3220 16212 3500
rect 16268 3490 16324 3500
rect 16380 3444 16436 15484
rect 16716 15538 16772 15932
rect 16716 15486 16718 15538
rect 16770 15486 16772 15538
rect 16716 15474 16772 15486
rect 16828 15428 16884 15438
rect 16940 15428 16996 16940
rect 16828 15426 16996 15428
rect 16828 15374 16830 15426
rect 16882 15374 16996 15426
rect 16828 15372 16996 15374
rect 16828 15362 16884 15372
rect 17052 8428 17108 17612
rect 17276 17108 17332 20748
rect 17612 20692 17668 21422
rect 17724 20916 17780 20926
rect 17780 20860 17892 20916
rect 17724 20850 17780 20860
rect 17836 20802 17892 20860
rect 17836 20750 17838 20802
rect 17890 20750 17892 20802
rect 17836 20738 17892 20750
rect 17612 20626 17668 20636
rect 17948 20242 18004 21756
rect 18172 21718 18228 21756
rect 17948 20190 17950 20242
rect 18002 20190 18004 20242
rect 17612 20132 17668 20142
rect 17500 19906 17556 19918
rect 17500 19854 17502 19906
rect 17554 19854 17556 19906
rect 17388 19796 17444 19806
rect 17388 19702 17444 19740
rect 17500 19012 17556 19854
rect 17500 18946 17556 18956
rect 17388 18452 17444 18462
rect 17612 18452 17668 20076
rect 17836 19684 17892 19694
rect 17724 19572 17780 19582
rect 17724 19234 17780 19516
rect 17724 19182 17726 19234
rect 17778 19182 17780 19234
rect 17724 19170 17780 19182
rect 17836 19234 17892 19628
rect 17948 19348 18004 20190
rect 18508 21586 18564 23212
rect 18508 21534 18510 21586
rect 18562 21534 18564 21586
rect 18508 20242 18564 21534
rect 18844 22370 18900 22382
rect 18844 22318 18846 22370
rect 18898 22318 18900 22370
rect 18844 21476 18900 22318
rect 19068 21812 19124 23774
rect 19628 23044 19684 24558
rect 20300 24610 20356 24622
rect 20300 24558 20302 24610
rect 20354 24558 20356 24610
rect 19852 24498 19908 24510
rect 19852 24446 19854 24498
rect 19906 24446 19908 24498
rect 19852 24050 19908 24446
rect 20300 24500 20356 24558
rect 20300 24434 20356 24444
rect 19852 23998 19854 24050
rect 19906 23998 19908 24050
rect 19852 23986 19908 23998
rect 20524 23828 20580 32620
rect 20636 28420 20692 33516
rect 21196 33572 21252 36652
rect 21308 36484 21364 36494
rect 21308 36390 21364 36428
rect 21420 36260 21476 36270
rect 21196 33506 21252 33516
rect 21308 36258 21476 36260
rect 21308 36206 21422 36258
rect 21474 36206 21476 36258
rect 21308 36204 21476 36206
rect 21308 32228 21364 36204
rect 21420 36194 21476 36204
rect 21420 35700 21476 35710
rect 21420 35606 21476 35644
rect 21532 32676 21588 39788
rect 21868 39172 21924 40350
rect 21868 39106 21924 39116
rect 22092 38946 22148 40462
rect 22764 40516 22820 40526
rect 22764 40422 22820 40460
rect 23212 39732 23268 41916
rect 23212 39638 23268 39676
rect 22092 38894 22094 38946
rect 22146 38894 22148 38946
rect 22092 38882 22148 38894
rect 21756 38388 21812 38398
rect 21756 38162 21812 38332
rect 22988 38388 23044 38398
rect 22092 38276 22148 38286
rect 22092 38182 22148 38220
rect 21756 38110 21758 38162
rect 21810 38110 21812 38162
rect 21756 38098 21812 38110
rect 21868 38164 21924 38174
rect 21644 38052 21700 38062
rect 21644 37156 21700 37996
rect 21868 37490 21924 38108
rect 22988 38050 23044 38332
rect 22988 37998 22990 38050
rect 23042 37998 23044 38050
rect 22988 37986 23044 37998
rect 23100 38052 23156 38062
rect 22204 37938 22260 37950
rect 22204 37886 22206 37938
rect 22258 37886 22260 37938
rect 22092 37826 22148 37838
rect 22092 37774 22094 37826
rect 22146 37774 22148 37826
rect 22092 37604 22148 37774
rect 22092 37538 22148 37548
rect 21868 37438 21870 37490
rect 21922 37438 21924 37490
rect 21868 37426 21924 37438
rect 22092 37380 22148 37390
rect 21644 37062 21700 37100
rect 21980 37378 22148 37380
rect 21980 37326 22094 37378
rect 22146 37326 22148 37378
rect 21980 37324 22148 37326
rect 21868 36370 21924 36382
rect 21868 36318 21870 36370
rect 21922 36318 21924 36370
rect 21644 36258 21700 36270
rect 21644 36206 21646 36258
rect 21698 36206 21700 36258
rect 21644 35586 21700 36206
rect 21644 35534 21646 35586
rect 21698 35534 21700 35586
rect 21644 35522 21700 35534
rect 21868 35588 21924 36318
rect 21980 35700 22036 37324
rect 22092 37314 22148 37324
rect 22204 37268 22260 37886
rect 22652 37828 22708 37838
rect 22204 36370 22260 37212
rect 22540 37826 22708 37828
rect 22540 37774 22654 37826
rect 22706 37774 22708 37826
rect 22540 37772 22708 37774
rect 22540 37156 22596 37772
rect 22652 37762 22708 37772
rect 22988 37492 23044 37502
rect 23100 37492 23156 37996
rect 23324 38052 23380 42924
rect 23772 42754 23828 43486
rect 23884 43540 23940 43550
rect 23884 43446 23940 43484
rect 23772 42702 23774 42754
rect 23826 42702 23828 42754
rect 23772 42644 23828 42702
rect 23436 42532 23492 42542
rect 23772 42532 23828 42588
rect 23996 42754 24052 43820
rect 24108 43650 24164 44044
rect 24332 43988 24388 48188
rect 24444 47236 24500 47246
rect 24444 45108 24500 47180
rect 24444 45042 24500 45052
rect 24556 44436 24612 48524
rect 24780 48468 24836 52332
rect 24780 48402 24836 48412
rect 24892 52164 24948 52174
rect 24668 48130 24724 48142
rect 24668 48078 24670 48130
rect 24722 48078 24724 48130
rect 24668 47908 24724 48078
rect 24668 47842 24724 47852
rect 24780 48132 24836 48142
rect 24780 47458 24836 48076
rect 24780 47406 24782 47458
rect 24834 47406 24836 47458
rect 24668 46676 24724 46686
rect 24780 46676 24836 47406
rect 24668 46674 24836 46676
rect 24668 46622 24670 46674
rect 24722 46622 24836 46674
rect 24668 46620 24836 46622
rect 24668 45332 24724 46620
rect 24892 46116 24948 52108
rect 25004 46228 25060 55412
rect 25228 54292 25284 56252
rect 25452 56082 25508 56094
rect 25452 56030 25454 56082
rect 25506 56030 25508 56082
rect 25340 55970 25396 55982
rect 25340 55918 25342 55970
rect 25394 55918 25396 55970
rect 25340 54964 25396 55918
rect 25340 54898 25396 54908
rect 25340 54292 25396 54302
rect 25228 54290 25396 54292
rect 25228 54238 25342 54290
rect 25394 54238 25396 54290
rect 25228 54236 25396 54238
rect 25340 53842 25396 54236
rect 25452 54292 25508 56030
rect 25564 55412 25620 56588
rect 25564 55346 25620 55356
rect 25900 56082 25956 56094
rect 25900 56030 25902 56082
rect 25954 56030 25956 56082
rect 25900 55188 25956 56030
rect 25676 54516 25732 54526
rect 25900 54516 25956 55132
rect 25452 54198 25508 54236
rect 25564 54514 25956 54516
rect 25564 54462 25678 54514
rect 25730 54462 25956 54514
rect 25564 54460 25956 54462
rect 25340 53790 25342 53842
rect 25394 53790 25396 53842
rect 25340 53778 25396 53790
rect 25564 53730 25620 54460
rect 25676 54450 25732 54460
rect 25564 53678 25566 53730
rect 25618 53678 25620 53730
rect 25564 53666 25620 53678
rect 25788 54290 25844 54302
rect 25788 54238 25790 54290
rect 25842 54238 25844 54290
rect 25228 53618 25284 53630
rect 25228 53566 25230 53618
rect 25282 53566 25284 53618
rect 25228 53060 25284 53566
rect 25788 53508 25844 54238
rect 25788 53442 25844 53452
rect 26012 53284 26068 58940
rect 26124 57428 26180 59166
rect 26236 59108 26292 59118
rect 26236 58994 26292 59052
rect 26236 58942 26238 58994
rect 26290 58942 26292 58994
rect 26236 58930 26292 58942
rect 26348 58322 26404 61068
rect 26460 59444 26516 61404
rect 26572 61346 26628 61358
rect 26572 61294 26574 61346
rect 26626 61294 26628 61346
rect 26572 61012 26628 61294
rect 26572 60946 26628 60956
rect 26796 61346 26852 61358
rect 26796 61294 26798 61346
rect 26850 61294 26852 61346
rect 26572 60788 26628 60798
rect 26572 60226 26628 60732
rect 26572 60174 26574 60226
rect 26626 60174 26628 60226
rect 26572 60162 26628 60174
rect 26796 60228 26852 61294
rect 26908 61348 26964 61358
rect 26908 61254 26964 61292
rect 27020 61346 27076 61358
rect 27020 61294 27022 61346
rect 27074 61294 27076 61346
rect 26460 59378 26516 59388
rect 26796 59218 26852 60172
rect 26908 60564 26964 60574
rect 26908 60002 26964 60508
rect 27020 60340 27076 61294
rect 27020 60274 27076 60284
rect 26908 59950 26910 60002
rect 26962 59950 26964 60002
rect 26908 59938 26964 59950
rect 27132 60002 27188 62078
rect 27132 59950 27134 60002
rect 27186 59950 27188 60002
rect 27132 59938 27188 59950
rect 27244 62132 27412 62188
rect 27468 62242 27524 62254
rect 27468 62190 27470 62242
rect 27522 62190 27524 62242
rect 27468 62188 27524 62190
rect 27916 62242 27972 62254
rect 27916 62190 27918 62242
rect 27970 62190 27972 62242
rect 27468 62132 27748 62188
rect 27244 59890 27300 62132
rect 27468 62020 27524 62132
rect 27468 61954 27524 61964
rect 27580 61908 27636 61918
rect 27468 61572 27524 61582
rect 27580 61572 27636 61852
rect 27468 61570 27636 61572
rect 27468 61518 27470 61570
rect 27522 61518 27636 61570
rect 27468 61516 27636 61518
rect 27692 61570 27748 62132
rect 27692 61518 27694 61570
rect 27746 61518 27748 61570
rect 27468 61506 27524 61516
rect 27692 61506 27748 61518
rect 27804 62130 27860 62142
rect 27804 62078 27806 62130
rect 27858 62078 27860 62130
rect 27804 61572 27860 62078
rect 27916 62020 27972 62190
rect 27916 61954 27972 61964
rect 28252 61796 28308 62414
rect 28252 61730 28308 61740
rect 27916 61572 27972 61582
rect 27804 61570 27972 61572
rect 27804 61518 27918 61570
rect 27970 61518 27972 61570
rect 27804 61516 27972 61518
rect 27916 61506 27972 61516
rect 28364 61570 28420 62860
rect 28476 62850 28532 62860
rect 28476 62356 28532 62366
rect 28476 62262 28532 62300
rect 28700 62132 28756 63980
rect 28812 63970 28868 63980
rect 28924 64034 28980 64204
rect 28924 63982 28926 64034
rect 28978 63982 28980 64034
rect 28924 63970 28980 63982
rect 28700 62066 28756 62076
rect 28812 63252 28868 63262
rect 28812 62354 28868 63196
rect 28812 62302 28814 62354
rect 28866 62302 28868 62354
rect 28364 61518 28366 61570
rect 28418 61518 28420 61570
rect 28140 61346 28196 61358
rect 28140 61294 28142 61346
rect 28194 61294 28196 61346
rect 28140 61012 28196 61294
rect 28252 61348 28308 61358
rect 28364 61348 28420 61518
rect 28476 61348 28532 61358
rect 28364 61292 28476 61348
rect 28252 61124 28308 61292
rect 28476 61282 28532 61292
rect 28252 61068 28532 61124
rect 28140 60956 28420 61012
rect 28140 60786 28196 60798
rect 28140 60734 28142 60786
rect 28194 60734 28196 60786
rect 27356 60676 27412 60686
rect 27356 60582 27412 60620
rect 28140 60564 28196 60734
rect 28252 60564 28308 60574
rect 28140 60508 28252 60564
rect 28252 60498 28308 60508
rect 28028 60228 28084 60238
rect 28028 60134 28084 60172
rect 28364 60226 28420 60956
rect 28476 60898 28532 61068
rect 28476 60846 28478 60898
rect 28530 60846 28532 60898
rect 28476 60834 28532 60846
rect 28700 60788 28756 60798
rect 28700 60694 28756 60732
rect 28588 60676 28644 60686
rect 28588 60582 28644 60620
rect 28812 60564 28868 62302
rect 29260 62188 29316 65996
rect 29372 66050 29428 66062
rect 29372 65998 29374 66050
rect 29426 65998 29428 66050
rect 29372 65380 29428 65998
rect 29484 65380 29540 65390
rect 29428 65378 29540 65380
rect 29428 65326 29486 65378
rect 29538 65326 29540 65378
rect 29428 65324 29540 65326
rect 29372 65286 29428 65324
rect 29372 64708 29428 64718
rect 29372 64614 29428 64652
rect 29484 64260 29540 65324
rect 29932 64930 29988 67788
rect 30044 67396 30100 68796
rect 30044 67330 30100 67340
rect 30044 67058 30100 67070
rect 30044 67006 30046 67058
rect 30098 67006 30100 67058
rect 30044 66948 30100 67006
rect 30156 67060 30212 69020
rect 30268 67956 30324 70364
rect 31052 70354 31108 70364
rect 32396 70354 32452 70364
rect 31164 70196 31220 70206
rect 30828 70194 31220 70196
rect 30828 70142 31166 70194
rect 31218 70142 31220 70194
rect 30828 70140 31220 70142
rect 30716 70084 30772 70094
rect 30716 69990 30772 70028
rect 30380 69636 30436 69646
rect 30380 69410 30436 69580
rect 30828 69524 30884 70140
rect 31164 70130 31220 70140
rect 33180 70194 33236 70476
rect 33964 70306 34020 70700
rect 34748 70690 34804 70700
rect 33964 70254 33966 70306
rect 34018 70254 34020 70306
rect 33964 70242 34020 70254
rect 33180 70142 33182 70194
rect 33234 70142 33236 70194
rect 33180 70130 33236 70142
rect 32508 70084 32564 70094
rect 32508 70082 33012 70084
rect 32508 70030 32510 70082
rect 32562 70030 33012 70082
rect 32508 70028 33012 70030
rect 32508 70018 32564 70028
rect 31276 69636 31332 69646
rect 31276 69542 31332 69580
rect 30380 69358 30382 69410
rect 30434 69358 30436 69410
rect 30380 69346 30436 69358
rect 30492 69468 30884 69524
rect 30940 69522 30996 69534
rect 30940 69470 30942 69522
rect 30994 69470 30996 69522
rect 30380 67956 30436 67966
rect 30268 67954 30436 67956
rect 30268 67902 30382 67954
rect 30434 67902 30436 67954
rect 30268 67900 30436 67902
rect 30380 67890 30436 67900
rect 30380 67396 30436 67406
rect 30380 67170 30436 67340
rect 30380 67118 30382 67170
rect 30434 67118 30436 67170
rect 30380 67106 30436 67118
rect 30492 67170 30548 69468
rect 30604 69298 30660 69310
rect 30604 69246 30606 69298
rect 30658 69246 30660 69298
rect 30604 67284 30660 69246
rect 30828 69188 30884 69198
rect 30828 69094 30884 69132
rect 30604 67218 30660 67228
rect 30828 68964 30884 68974
rect 30492 67118 30494 67170
rect 30546 67118 30548 67170
rect 30492 67106 30548 67118
rect 30156 66994 30212 67004
rect 30604 67060 30660 67070
rect 30604 66966 30660 67004
rect 30044 66882 30100 66892
rect 30716 66948 30772 66958
rect 30268 66162 30324 66174
rect 30268 66110 30270 66162
rect 30322 66110 30324 66162
rect 30044 66052 30100 66062
rect 30268 66052 30324 66110
rect 30604 66164 30660 66174
rect 30716 66164 30772 66892
rect 30604 66162 30772 66164
rect 30604 66110 30606 66162
rect 30658 66110 30772 66162
rect 30604 66108 30772 66110
rect 30828 66164 30884 68908
rect 30940 67058 30996 69470
rect 32956 69522 33012 70028
rect 34860 69972 34916 70814
rect 32956 69470 32958 69522
rect 33010 69470 33012 69522
rect 32956 69458 33012 69470
rect 34300 69916 34916 69972
rect 34972 69972 35028 71036
rect 36428 70532 36484 70542
rect 36428 70194 36484 70476
rect 36428 70142 36430 70194
rect 36482 70142 36484 70194
rect 36428 70130 36484 70142
rect 36092 70082 36148 70094
rect 36092 70030 36094 70082
rect 36146 70030 36148 70082
rect 34972 69916 35140 69972
rect 34300 69522 34356 69916
rect 34300 69470 34302 69522
rect 34354 69470 34356 69522
rect 34300 69458 34356 69470
rect 31164 69356 31444 69412
rect 31052 69188 31108 69198
rect 31164 69188 31220 69356
rect 31388 69298 31444 69356
rect 33404 69410 33460 69422
rect 33404 69358 33406 69410
rect 33458 69358 33460 69410
rect 31388 69246 31390 69298
rect 31442 69246 31444 69298
rect 31388 69234 31444 69246
rect 31836 69300 31892 69310
rect 31836 69206 31892 69244
rect 33292 69300 33348 69310
rect 31052 69186 31220 69188
rect 31052 69134 31054 69186
rect 31106 69134 31220 69186
rect 31052 69132 31220 69134
rect 31052 69122 31108 69132
rect 30940 67006 30942 67058
rect 30994 67006 30996 67058
rect 30940 66994 30996 67006
rect 31052 68628 31108 68638
rect 31052 66498 31108 68572
rect 31164 67508 31220 69132
rect 31164 67442 31220 67452
rect 31276 69188 31332 69198
rect 31276 67170 31332 69132
rect 31612 69188 31668 69198
rect 31612 69094 31668 69132
rect 32844 69186 32900 69198
rect 32844 69134 32846 69186
rect 32898 69134 32900 69186
rect 32844 68964 32900 69134
rect 33068 69186 33124 69198
rect 33068 69134 33070 69186
rect 33122 69134 33124 69186
rect 33068 69076 33124 69134
rect 33068 69010 33124 69020
rect 32844 68898 32900 68908
rect 33292 68850 33348 69244
rect 33292 68798 33294 68850
rect 33346 68798 33348 68850
rect 33292 68786 33348 68798
rect 32956 68628 33012 68638
rect 32956 68534 33012 68572
rect 33404 68514 33460 69358
rect 34412 69412 34468 69422
rect 34412 69318 34468 69356
rect 34972 69300 35028 69310
rect 33964 69188 34020 69226
rect 34972 69206 35028 69244
rect 33964 69122 34020 69132
rect 34188 69186 34244 69198
rect 34188 69134 34190 69186
rect 34242 69134 34244 69186
rect 34188 69076 34244 69134
rect 34636 69188 34692 69198
rect 34636 69094 34692 69132
rect 34748 69186 34804 69198
rect 34748 69134 34750 69186
rect 34802 69134 34804 69186
rect 34748 69076 34804 69134
rect 34748 69020 35028 69076
rect 34188 69010 34244 69020
rect 33516 68852 33572 68862
rect 33516 68758 33572 68796
rect 34972 68852 35028 69020
rect 34972 68786 35028 68796
rect 35084 68964 35140 69916
rect 35196 69804 35460 69814
rect 35252 69748 35300 69804
rect 35356 69748 35404 69804
rect 35196 69738 35460 69748
rect 35644 69636 35700 69646
rect 35308 69634 35700 69636
rect 35308 69582 35646 69634
rect 35698 69582 35700 69634
rect 35308 69580 35700 69582
rect 35308 69410 35364 69580
rect 35644 69570 35700 69580
rect 35308 69358 35310 69410
rect 35362 69358 35364 69410
rect 35308 69346 35364 69358
rect 36092 69412 36148 70030
rect 36428 69636 36484 69646
rect 36428 69542 36484 69580
rect 34412 68740 34468 68750
rect 34412 68646 34468 68684
rect 33404 68462 33406 68514
rect 33458 68462 33460 68514
rect 33404 68450 33460 68462
rect 34748 68626 34804 68638
rect 34748 68574 34750 68626
rect 34802 68574 34804 68626
rect 31276 67118 31278 67170
rect 31330 67118 31332 67170
rect 31276 67106 31332 67118
rect 31500 68180 31556 68190
rect 31500 67172 31556 68124
rect 32508 67954 32564 67966
rect 32508 67902 32510 67954
rect 32562 67902 32564 67954
rect 32060 67172 32116 67182
rect 31500 67170 32116 67172
rect 31500 67118 32062 67170
rect 32114 67118 32116 67170
rect 31500 67116 32116 67118
rect 31500 67058 31556 67116
rect 31500 67006 31502 67058
rect 31554 67006 31556 67058
rect 31500 66994 31556 67006
rect 32060 67060 32116 67116
rect 32508 67172 32564 67902
rect 32508 67106 32564 67116
rect 33068 67618 33124 67630
rect 33068 67566 33070 67618
rect 33122 67566 33124 67618
rect 33068 67396 33124 67566
rect 32060 66994 32116 67004
rect 31052 66446 31054 66498
rect 31106 66446 31108 66498
rect 31052 66434 31108 66446
rect 31052 66276 31108 66286
rect 30940 66164 30996 66174
rect 30828 66162 30996 66164
rect 30828 66110 30942 66162
rect 30994 66110 30996 66162
rect 30828 66108 30996 66110
rect 30604 66098 30660 66108
rect 30100 65996 30324 66052
rect 30044 65958 30100 65996
rect 30268 65602 30324 65614
rect 30268 65550 30270 65602
rect 30322 65550 30324 65602
rect 29932 64878 29934 64930
rect 29986 64878 29988 64930
rect 29932 64866 29988 64878
rect 30044 65490 30100 65502
rect 30044 65438 30046 65490
rect 30098 65438 30100 65490
rect 29820 64708 29876 64718
rect 30044 64708 30100 65438
rect 30156 65492 30212 65502
rect 30156 65398 30212 65436
rect 29820 64706 30100 64708
rect 29820 64654 29822 64706
rect 29874 64654 30100 64706
rect 29820 64652 30100 64654
rect 30268 64708 30324 65550
rect 29484 64194 29540 64204
rect 29596 64482 29652 64494
rect 29596 64430 29598 64482
rect 29650 64430 29652 64482
rect 29596 64148 29652 64430
rect 29820 64372 29876 64652
rect 30268 64642 30324 64652
rect 30716 65490 30772 65502
rect 30716 65438 30718 65490
rect 30770 65438 30772 65490
rect 29820 64306 29876 64316
rect 30156 64484 30212 64494
rect 30604 64484 30660 64494
rect 30156 64482 30660 64484
rect 30156 64430 30158 64482
rect 30210 64430 30606 64482
rect 30658 64430 30660 64482
rect 30156 64428 30660 64430
rect 30156 64260 30212 64428
rect 30604 64418 30660 64428
rect 30156 64194 30212 64204
rect 30716 64372 30772 65438
rect 29596 64092 29764 64148
rect 29372 64036 29428 64046
rect 29372 63942 29428 63980
rect 29596 63922 29652 63934
rect 29596 63870 29598 63922
rect 29650 63870 29652 63922
rect 29484 63812 29540 63822
rect 29484 63718 29540 63756
rect 29484 62356 29540 62366
rect 29484 62262 29540 62300
rect 29148 62132 29316 62188
rect 29036 61796 29092 61806
rect 29036 61570 29092 61740
rect 29036 61518 29038 61570
rect 29090 61518 29092 61570
rect 29036 61506 29092 61518
rect 28924 61012 28980 61022
rect 28924 60918 28980 60956
rect 29036 60564 29092 60574
rect 28812 60508 29036 60564
rect 28364 60174 28366 60226
rect 28418 60174 28420 60226
rect 28364 60162 28420 60174
rect 27244 59838 27246 59890
rect 27298 59838 27300 59890
rect 27132 59444 27188 59482
rect 27132 59378 27188 59388
rect 26908 59332 26964 59342
rect 26964 59276 27076 59332
rect 26908 59266 26964 59276
rect 26796 59166 26798 59218
rect 26850 59166 26852 59218
rect 26796 59154 26852 59166
rect 26348 58270 26350 58322
rect 26402 58270 26404 58322
rect 26348 58258 26404 58270
rect 26684 58772 26740 58782
rect 26684 58322 26740 58716
rect 26908 58436 26964 58446
rect 26908 58342 26964 58380
rect 26684 58270 26686 58322
rect 26738 58270 26740 58322
rect 26684 58258 26740 58270
rect 26124 57362 26180 57372
rect 26460 58212 26516 58222
rect 26460 56978 26516 58156
rect 26460 56926 26462 56978
rect 26514 56926 26516 56978
rect 26460 56914 26516 56926
rect 26572 57204 26628 57214
rect 26572 56082 26628 57148
rect 26572 56030 26574 56082
rect 26626 56030 26628 56082
rect 26572 56018 26628 56030
rect 26348 55970 26404 55982
rect 26348 55918 26350 55970
rect 26402 55918 26404 55970
rect 26236 55412 26292 55422
rect 26124 54626 26180 54638
rect 26124 54574 26126 54626
rect 26178 54574 26180 54626
rect 26124 54516 26180 54574
rect 26124 54450 26180 54460
rect 26124 53956 26180 53966
rect 26124 53730 26180 53900
rect 26124 53678 26126 53730
rect 26178 53678 26180 53730
rect 26124 53666 26180 53678
rect 26012 53228 26180 53284
rect 25116 53004 25284 53060
rect 26012 53060 26068 53070
rect 25116 52052 25172 53004
rect 26012 52966 26068 53004
rect 25676 52946 25732 52958
rect 25676 52894 25678 52946
rect 25730 52894 25732 52946
rect 25228 52836 25284 52846
rect 25228 52274 25284 52780
rect 25340 52834 25396 52846
rect 25340 52782 25342 52834
rect 25394 52782 25396 52834
rect 25340 52724 25396 52782
rect 25340 52658 25396 52668
rect 25676 52612 25732 52894
rect 25676 52546 25732 52556
rect 25340 52388 25396 52398
rect 25340 52386 26068 52388
rect 25340 52334 25342 52386
rect 25394 52334 26068 52386
rect 25340 52332 26068 52334
rect 25340 52322 25396 52332
rect 25228 52222 25230 52274
rect 25282 52222 25284 52274
rect 25228 52210 25284 52222
rect 25116 51986 25172 51996
rect 25676 52162 25732 52174
rect 25676 52110 25678 52162
rect 25730 52110 25732 52162
rect 25228 51380 25284 51390
rect 25676 51380 25732 52110
rect 26012 51490 26068 52332
rect 26012 51438 26014 51490
rect 26066 51438 26068 51490
rect 26012 51426 26068 51438
rect 25116 51378 25732 51380
rect 25116 51326 25230 51378
rect 25282 51326 25732 51378
rect 25116 51324 25732 51326
rect 25116 48132 25172 51324
rect 25228 51314 25284 51324
rect 25340 50372 25396 50382
rect 25340 49922 25396 50316
rect 25340 49870 25342 49922
rect 25394 49870 25396 49922
rect 25340 49858 25396 49870
rect 25228 49588 25284 49598
rect 25228 49494 25284 49532
rect 26124 49476 26180 53228
rect 26236 52724 26292 55356
rect 26348 55300 26404 55918
rect 27020 55468 27076 59276
rect 27132 59220 27188 59230
rect 27132 59126 27188 59164
rect 27244 58772 27300 59838
rect 28028 60002 28084 60014
rect 28028 59950 28030 60002
rect 28082 59950 28084 60002
rect 27692 59780 27748 59790
rect 28028 59780 28084 59950
rect 27580 59778 28084 59780
rect 27580 59726 27694 59778
rect 27746 59726 28084 59778
rect 27580 59724 28084 59726
rect 27468 59332 27524 59342
rect 27580 59332 27636 59724
rect 27692 59714 27748 59724
rect 27468 59330 27636 59332
rect 27468 59278 27470 59330
rect 27522 59278 27636 59330
rect 27468 59276 27636 59278
rect 27692 59444 27748 59454
rect 27468 59266 27524 59276
rect 27244 58706 27300 58716
rect 27692 58658 27748 59388
rect 27692 58606 27694 58658
rect 27746 58606 27748 58658
rect 27692 58594 27748 58606
rect 27804 59332 27860 59342
rect 27244 57540 27300 57550
rect 27244 57446 27300 57484
rect 27356 55972 27412 55982
rect 27356 55878 27412 55916
rect 26348 55206 26404 55244
rect 26908 55412 27076 55468
rect 27804 55524 27860 59276
rect 29036 59218 29092 60508
rect 29148 60004 29204 62132
rect 29260 62020 29316 62030
rect 29260 61460 29316 61964
rect 29260 61366 29316 61404
rect 29372 61458 29428 61470
rect 29372 61406 29374 61458
rect 29426 61406 29428 61458
rect 29372 60788 29428 61406
rect 29596 61460 29652 63870
rect 29596 61394 29652 61404
rect 29708 60900 29764 64092
rect 30380 64146 30436 64158
rect 30380 64094 30382 64146
rect 30434 64094 30436 64146
rect 30380 64036 30436 64094
rect 30380 63970 30436 63980
rect 30044 63922 30100 63934
rect 30044 63870 30046 63922
rect 30098 63870 30100 63922
rect 30044 63028 30100 63870
rect 30492 63922 30548 63934
rect 30492 63870 30494 63922
rect 30546 63870 30548 63922
rect 30044 62962 30100 62972
rect 30380 63810 30436 63822
rect 30380 63758 30382 63810
rect 30434 63758 30436 63810
rect 30044 62244 30100 62254
rect 29932 62020 29988 62030
rect 29932 61570 29988 61964
rect 29932 61518 29934 61570
rect 29986 61518 29988 61570
rect 29932 61506 29988 61518
rect 29372 60722 29428 60732
rect 29484 60844 29764 60900
rect 29820 61458 29876 61470
rect 29820 61406 29822 61458
rect 29874 61406 29876 61458
rect 29148 59938 29204 59948
rect 29036 59166 29038 59218
rect 29090 59166 29092 59218
rect 29036 59154 29092 59166
rect 27916 59106 27972 59118
rect 27916 59054 27918 59106
rect 27970 59054 27972 59106
rect 27916 58772 27972 59054
rect 27916 57988 27972 58716
rect 28812 59106 28868 59118
rect 28812 59054 28814 59106
rect 28866 59054 28868 59106
rect 28028 58436 28084 58446
rect 28028 58342 28084 58380
rect 28812 58436 28868 59054
rect 29484 58658 29540 60844
rect 29820 60788 29876 61406
rect 29820 60722 29876 60732
rect 30044 61458 30100 62188
rect 30044 61406 30046 61458
rect 30098 61406 30100 61458
rect 29596 60676 29652 60686
rect 29596 60114 29652 60620
rect 29596 60062 29598 60114
rect 29650 60062 29652 60114
rect 29596 60050 29652 60062
rect 29708 60674 29764 60686
rect 29708 60622 29710 60674
rect 29762 60622 29764 60674
rect 29708 60564 29764 60622
rect 30044 60564 30100 61406
rect 30268 62020 30324 62030
rect 30268 60898 30324 61964
rect 30380 61010 30436 63758
rect 30492 61796 30548 63870
rect 30716 62132 30772 64316
rect 30716 62066 30772 62076
rect 30828 62020 30884 66108
rect 30940 66098 30996 66108
rect 31052 66162 31108 66220
rect 31052 66110 31054 66162
rect 31106 66110 31108 66162
rect 31052 66098 31108 66110
rect 31612 66052 31668 66062
rect 30940 64932 30996 64942
rect 30940 64930 31220 64932
rect 30940 64878 30942 64930
rect 30994 64878 31220 64930
rect 30940 64876 31220 64878
rect 30940 64866 30996 64876
rect 31164 64706 31220 64876
rect 31164 64654 31166 64706
rect 31218 64654 31220 64706
rect 31164 63252 31220 64654
rect 31164 63158 31220 63196
rect 31388 64036 31444 64046
rect 31164 62356 31220 62366
rect 31052 62244 31108 62254
rect 30828 61954 30884 61964
rect 30940 62132 30996 62142
rect 30492 61794 30884 61796
rect 30492 61742 30494 61794
rect 30546 61742 30884 61794
rect 30492 61740 30884 61742
rect 30492 61730 30548 61740
rect 30380 60958 30382 61010
rect 30434 60958 30436 61010
rect 30380 60946 30436 60958
rect 30604 61572 30660 61582
rect 30604 61012 30660 61516
rect 30828 61570 30884 61740
rect 30828 61518 30830 61570
rect 30882 61518 30884 61570
rect 30828 61506 30884 61518
rect 30268 60846 30270 60898
rect 30322 60846 30324 60898
rect 30268 60834 30324 60846
rect 30604 60898 30660 60956
rect 30604 60846 30606 60898
rect 30658 60846 30660 60898
rect 30604 60834 30660 60846
rect 30156 60788 30212 60798
rect 30156 60694 30212 60732
rect 29708 60508 30100 60564
rect 29484 58606 29486 58658
rect 29538 58606 29540 58658
rect 29484 58594 29540 58606
rect 28812 58370 28868 58380
rect 27916 57922 27972 57932
rect 28140 58324 28196 58334
rect 27804 55458 27860 55468
rect 28028 55972 28084 55982
rect 27244 55412 27300 55422
rect 26460 54964 26516 54974
rect 26516 54908 26852 54964
rect 26460 54898 26516 54908
rect 26460 54740 26516 54750
rect 26460 54646 26516 54684
rect 26796 54626 26852 54908
rect 26796 54574 26798 54626
rect 26850 54574 26852 54626
rect 26796 54562 26852 54574
rect 26908 54626 26964 55412
rect 26908 54574 26910 54626
rect 26962 54574 26964 54626
rect 26908 54516 26964 54574
rect 26908 54450 26964 54460
rect 27020 55298 27076 55310
rect 27020 55246 27022 55298
rect 27074 55246 27076 55298
rect 27020 54852 27076 55246
rect 27244 55186 27300 55356
rect 28028 55410 28084 55916
rect 28028 55358 28030 55410
rect 28082 55358 28084 55410
rect 28028 55346 28084 55358
rect 28140 55298 28196 58268
rect 28252 58212 28308 58222
rect 28252 58118 28308 58156
rect 28364 58210 28420 58222
rect 28364 58158 28366 58210
rect 28418 58158 28420 58210
rect 28364 57876 28420 58158
rect 28364 57810 28420 57820
rect 28588 57652 28644 57662
rect 28588 56978 28644 57596
rect 29708 57204 29764 60508
rect 30940 59890 30996 62076
rect 31052 60788 31108 62188
rect 31052 60674 31108 60732
rect 31052 60622 31054 60674
rect 31106 60622 31108 60674
rect 31052 60116 31108 60622
rect 31052 60050 31108 60060
rect 30940 59838 30942 59890
rect 30994 59838 30996 59890
rect 30940 59826 30996 59838
rect 29820 59108 29876 59118
rect 30268 59108 30324 59118
rect 29820 59106 30100 59108
rect 29820 59054 29822 59106
rect 29874 59054 30100 59106
rect 29820 59052 30100 59054
rect 29820 59042 29876 59052
rect 30044 58546 30100 59052
rect 30044 58494 30046 58546
rect 30098 58494 30100 58546
rect 30044 58482 30100 58494
rect 29820 58436 29876 58446
rect 29820 57540 29876 58380
rect 30156 58436 30212 58446
rect 30156 58342 30212 58380
rect 29932 58324 29988 58334
rect 29932 58212 29988 58268
rect 30268 58212 30324 59052
rect 30940 58548 30996 58558
rect 31164 58548 31220 62300
rect 31388 61572 31444 63980
rect 31612 64034 31668 65996
rect 32732 66052 32788 66062
rect 32732 66050 32900 66052
rect 32732 65998 32734 66050
rect 32786 65998 32900 66050
rect 32732 65996 32900 65998
rect 32732 65986 32788 65996
rect 32172 65602 32228 65614
rect 32172 65550 32174 65602
rect 32226 65550 32228 65602
rect 31948 65492 32004 65502
rect 31948 65398 32004 65436
rect 31948 64820 32004 64830
rect 32172 64820 32228 65550
rect 32620 65604 32676 65614
rect 31948 64818 32228 64820
rect 31948 64766 31950 64818
rect 32002 64766 32228 64818
rect 31948 64764 32228 64766
rect 32284 65492 32340 65502
rect 31948 64754 32004 64764
rect 32172 64484 32228 64494
rect 32284 64484 32340 65436
rect 32508 65492 32564 65502
rect 32508 65398 32564 65436
rect 32228 64428 32340 64484
rect 32396 64484 32452 64494
rect 31724 64260 31780 64270
rect 31724 64146 31780 64204
rect 31724 64094 31726 64146
rect 31778 64094 31780 64146
rect 31724 64082 31780 64094
rect 31612 63982 31614 64034
rect 31666 63982 31668 64034
rect 31612 63970 31668 63982
rect 31948 64036 32004 64046
rect 31948 63942 32004 63980
rect 31836 63924 31892 63934
rect 31612 62244 31668 62282
rect 31612 62178 31668 62188
rect 31836 61682 31892 63868
rect 32172 63924 32228 64428
rect 32172 63922 32340 63924
rect 32172 63870 32174 63922
rect 32226 63870 32340 63922
rect 32172 63868 32340 63870
rect 32172 63858 32228 63868
rect 32284 63588 32340 63868
rect 32396 63810 32452 64428
rect 32508 64036 32564 64046
rect 32620 64036 32676 65548
rect 32508 64034 32676 64036
rect 32508 63982 32510 64034
rect 32562 63982 32676 64034
rect 32508 63980 32676 63982
rect 32844 65492 32900 65996
rect 32956 65492 33012 65502
rect 32844 65490 33012 65492
rect 32844 65438 32958 65490
rect 33010 65438 33012 65490
rect 32844 65436 33012 65438
rect 32844 65380 32900 65436
rect 32956 65426 33012 65436
rect 32508 63970 32564 63980
rect 32396 63758 32398 63810
rect 32450 63758 32452 63810
rect 32396 63746 32452 63758
rect 32284 63532 32564 63588
rect 32396 63028 32452 63038
rect 32284 62244 32340 62282
rect 32284 62178 32340 62188
rect 31836 61630 31838 61682
rect 31890 61630 31892 61682
rect 31836 61618 31892 61630
rect 32396 61682 32452 62972
rect 32508 62132 32564 63532
rect 32844 62244 32900 65324
rect 33068 64820 33124 67340
rect 33404 67618 33460 67630
rect 33404 67566 33406 67618
rect 33458 67566 33460 67618
rect 33404 67172 33460 67566
rect 33292 66052 33348 66062
rect 33292 65958 33348 65996
rect 33404 65940 33460 67116
rect 34412 66948 34468 66958
rect 34300 66946 34468 66948
rect 34300 66894 34414 66946
rect 34466 66894 34468 66946
rect 34300 66892 34468 66894
rect 33628 66164 33684 66174
rect 34076 66164 34132 66174
rect 34300 66164 34356 66892
rect 34412 66882 34468 66892
rect 34748 66948 34804 68574
rect 34748 66882 34804 66892
rect 34524 66500 34580 66510
rect 34524 66386 34580 66444
rect 34524 66334 34526 66386
rect 34578 66334 34580 66386
rect 34524 66322 34580 66334
rect 33628 66162 33908 66164
rect 33628 66110 33630 66162
rect 33682 66110 33908 66162
rect 33628 66108 33908 66110
rect 33628 66098 33684 66108
rect 33404 65874 33460 65884
rect 33516 66052 33572 66062
rect 32956 64764 33124 64820
rect 33404 65716 33460 65726
rect 33404 65490 33460 65660
rect 33516 65604 33572 65996
rect 33516 65538 33572 65548
rect 33740 65940 33796 65950
rect 33404 65438 33406 65490
rect 33458 65438 33460 65490
rect 32956 63700 33012 64764
rect 33404 64708 33460 65438
rect 33628 65490 33684 65502
rect 33628 65438 33630 65490
rect 33682 65438 33684 65490
rect 33068 64652 33460 64708
rect 33516 65378 33572 65390
rect 33516 65326 33518 65378
rect 33570 65326 33572 65378
rect 33068 63924 33124 64652
rect 33516 64596 33572 65326
rect 33068 63858 33124 63868
rect 33180 64540 33572 64596
rect 33628 65380 33684 65438
rect 33180 63922 33236 64540
rect 33516 64148 33572 64158
rect 33516 64054 33572 64092
rect 33628 64036 33684 65324
rect 33628 63942 33684 63980
rect 33180 63870 33182 63922
rect 33234 63870 33236 63922
rect 33180 63858 33236 63870
rect 33292 63924 33348 63934
rect 33292 63830 33348 63868
rect 32956 63644 33348 63700
rect 33068 62692 33124 62702
rect 33068 62578 33124 62636
rect 33068 62526 33070 62578
rect 33122 62526 33124 62578
rect 33068 62514 33124 62526
rect 33292 62580 33348 63644
rect 33292 62578 33460 62580
rect 33292 62526 33294 62578
rect 33346 62526 33460 62578
rect 33292 62524 33460 62526
rect 33292 62514 33348 62524
rect 32844 62178 32900 62188
rect 33180 62356 33236 62366
rect 33180 62188 33236 62300
rect 32508 62066 32564 62076
rect 32956 62130 33012 62142
rect 33180 62132 33348 62188
rect 32956 62078 32958 62130
rect 33010 62078 33012 62130
rect 32396 61630 32398 61682
rect 32450 61630 32452 61682
rect 32396 61618 32452 61630
rect 32732 61796 32788 61806
rect 31388 61478 31444 61516
rect 32172 61572 32228 61582
rect 32172 61478 32228 61516
rect 32508 61570 32564 61582
rect 32508 61518 32510 61570
rect 32562 61518 32564 61570
rect 31500 61460 31556 61470
rect 31500 61366 31556 61404
rect 32508 61460 32564 61518
rect 32508 61394 32564 61404
rect 32732 61570 32788 61740
rect 32732 61518 32734 61570
rect 32786 61518 32788 61570
rect 31724 61236 31780 61246
rect 31500 61012 31556 61022
rect 31500 60918 31556 60956
rect 30996 58492 31220 58548
rect 31276 59778 31332 59790
rect 31276 59726 31278 59778
rect 31330 59726 31332 59778
rect 30940 58454 30996 58492
rect 29932 58210 30324 58212
rect 29932 58158 29934 58210
rect 29986 58158 30324 58210
rect 29932 58156 30324 58158
rect 31276 58212 31332 59726
rect 31500 58212 31556 58222
rect 31276 58156 31500 58212
rect 29932 58146 29988 58156
rect 29820 57474 29876 57484
rect 28588 56926 28590 56978
rect 28642 56926 28644 56978
rect 28588 56914 28644 56926
rect 29036 57148 29764 57204
rect 28588 55412 28644 55422
rect 28140 55246 28142 55298
rect 28194 55246 28196 55298
rect 28140 55234 28196 55246
rect 28364 55298 28420 55310
rect 28364 55246 28366 55298
rect 28418 55246 28420 55298
rect 27244 55134 27246 55186
rect 27298 55134 27300 55186
rect 27244 55122 27300 55134
rect 28364 55188 28420 55246
rect 28364 55122 28420 55132
rect 28588 55298 28644 55356
rect 28588 55246 28590 55298
rect 28642 55246 28644 55298
rect 27916 55076 27972 55086
rect 27916 54982 27972 55020
rect 27020 54404 27076 54796
rect 27916 54516 27972 54526
rect 27468 54404 27524 54414
rect 27020 54338 27076 54348
rect 27244 54402 27524 54404
rect 27244 54350 27470 54402
rect 27522 54350 27524 54402
rect 27244 54348 27524 54350
rect 26908 54292 26964 54302
rect 26796 54290 26964 54292
rect 26796 54238 26910 54290
rect 26962 54238 26964 54290
rect 26796 54236 26964 54238
rect 26684 53844 26740 53854
rect 26684 53750 26740 53788
rect 26796 53730 26852 54236
rect 26908 54226 26964 54236
rect 27244 54180 27300 54348
rect 27468 54338 27524 54348
rect 27916 54402 27972 54460
rect 27916 54350 27918 54402
rect 27970 54350 27972 54402
rect 27132 53844 27188 53854
rect 26796 53678 26798 53730
rect 26850 53678 26852 53730
rect 26796 53666 26852 53678
rect 27020 53788 27132 53844
rect 26572 53508 26628 53518
rect 26572 53414 26628 53452
rect 26684 53284 26740 53294
rect 26684 53170 26740 53228
rect 26684 53118 26686 53170
rect 26738 53118 26740 53170
rect 26684 53106 26740 53118
rect 26236 52658 26292 52668
rect 26348 52946 26404 52958
rect 26348 52894 26350 52946
rect 26402 52894 26404 52946
rect 26348 52164 26404 52894
rect 26348 52098 26404 52108
rect 26908 52948 26964 52958
rect 26460 52052 26516 52062
rect 26460 51958 26516 51996
rect 26908 50708 26964 52892
rect 26908 50642 26964 50652
rect 26348 50596 26404 50606
rect 26348 50594 26740 50596
rect 26348 50542 26350 50594
rect 26402 50542 26740 50594
rect 26348 50540 26740 50542
rect 26348 50530 26404 50540
rect 26236 50372 26292 50382
rect 26460 50372 26516 50382
rect 26292 50370 26516 50372
rect 26292 50318 26462 50370
rect 26514 50318 26516 50370
rect 26292 50316 26516 50318
rect 26236 50306 26292 50316
rect 26460 50306 26516 50316
rect 26572 50372 26628 50382
rect 26572 50278 26628 50316
rect 26348 49812 26404 49822
rect 26348 49718 26404 49756
rect 26572 49810 26628 49822
rect 26572 49758 26574 49810
rect 26626 49758 26628 49810
rect 26012 49420 26180 49476
rect 26460 49698 26516 49710
rect 26460 49646 26462 49698
rect 26514 49646 26516 49698
rect 25116 48066 25172 48076
rect 25228 48242 25284 48254
rect 25228 48190 25230 48242
rect 25282 48190 25284 48242
rect 25228 47236 25284 48190
rect 25228 47170 25284 47180
rect 25564 47346 25620 47358
rect 25564 47294 25566 47346
rect 25618 47294 25620 47346
rect 25340 46676 25396 46686
rect 25340 46582 25396 46620
rect 25564 46564 25620 47294
rect 25788 46676 25844 46686
rect 25788 46582 25844 46620
rect 25564 46498 25620 46508
rect 25228 46452 25284 46462
rect 25228 46358 25284 46396
rect 25788 46228 25844 46238
rect 25004 46172 25172 46228
rect 24892 46060 25060 46116
rect 24668 45266 24724 45276
rect 24892 45892 24948 45902
rect 24108 43598 24110 43650
rect 24162 43598 24164 43650
rect 24108 43586 24164 43598
rect 24220 43932 24388 43988
rect 24444 44380 24612 44436
rect 24220 43428 24276 43932
rect 24332 43764 24388 43774
rect 24332 43650 24388 43708
rect 24332 43598 24334 43650
rect 24386 43598 24388 43650
rect 24332 43586 24388 43598
rect 23996 42702 23998 42754
rect 24050 42702 24052 42754
rect 23436 42530 23828 42532
rect 23436 42478 23438 42530
rect 23490 42478 23828 42530
rect 23436 42476 23828 42478
rect 23436 42466 23492 42476
rect 23772 42308 23828 42476
rect 23884 42532 23940 42542
rect 23884 42438 23940 42476
rect 23772 42252 23940 42308
rect 23660 41972 23716 41982
rect 23548 40964 23604 40974
rect 23436 40962 23604 40964
rect 23436 40910 23550 40962
rect 23602 40910 23604 40962
rect 23436 40908 23604 40910
rect 23436 40516 23492 40908
rect 23548 40898 23604 40908
rect 23660 40964 23716 41916
rect 23884 41970 23940 42252
rect 23884 41918 23886 41970
rect 23938 41918 23940 41970
rect 23884 41906 23940 41918
rect 23772 41858 23828 41870
rect 23772 41806 23774 41858
rect 23826 41806 23828 41858
rect 23772 41748 23828 41806
rect 23996 41748 24052 42702
rect 24108 43372 24276 43428
rect 24108 42084 24164 43372
rect 24332 42756 24388 42766
rect 24332 42662 24388 42700
rect 24108 42028 24276 42084
rect 23772 41692 24052 41748
rect 24108 41858 24164 41870
rect 24108 41806 24110 41858
rect 24162 41806 24164 41858
rect 24108 41412 24164 41806
rect 23660 40740 23716 40908
rect 23436 40422 23492 40460
rect 23548 40684 23716 40740
rect 23772 41356 24164 41412
rect 23324 37986 23380 37996
rect 22988 37490 23156 37492
rect 22988 37438 22990 37490
rect 23042 37438 23156 37490
rect 22988 37436 23156 37438
rect 23324 37828 23380 37838
rect 22988 37426 23044 37436
rect 22764 37380 22820 37390
rect 22764 37378 22932 37380
rect 22764 37326 22766 37378
rect 22818 37326 22932 37378
rect 22764 37324 22932 37326
rect 22764 37314 22820 37324
rect 22652 37268 22708 37278
rect 22652 37174 22708 37212
rect 22540 37090 22596 37100
rect 22204 36318 22206 36370
rect 22258 36318 22260 36370
rect 22204 36306 22260 36318
rect 22652 36596 22708 36606
rect 22652 36370 22708 36540
rect 22652 36318 22654 36370
rect 22706 36318 22708 36370
rect 22652 36306 22708 36318
rect 22764 36370 22820 36382
rect 22764 36318 22766 36370
rect 22818 36318 22820 36370
rect 22428 36260 22484 36270
rect 22428 36166 22484 36204
rect 22428 35756 22708 35812
rect 21980 35634 22036 35644
rect 22316 35698 22372 35710
rect 22316 35646 22318 35698
rect 22370 35646 22372 35698
rect 21868 35522 21924 35532
rect 22092 35588 22148 35598
rect 22316 35588 22372 35646
rect 22092 35586 22372 35588
rect 22092 35534 22094 35586
rect 22146 35534 22372 35586
rect 22092 35532 22372 35534
rect 22092 35364 22148 35532
rect 22428 35476 22484 35756
rect 22652 35698 22708 35756
rect 22652 35646 22654 35698
rect 22706 35646 22708 35698
rect 22652 35634 22708 35646
rect 22764 35700 22820 36318
rect 21644 35308 22148 35364
rect 22204 35420 22484 35476
rect 22540 35586 22596 35598
rect 22540 35534 22542 35586
rect 22594 35534 22596 35586
rect 21644 34914 21700 35308
rect 21644 34862 21646 34914
rect 21698 34862 21700 34914
rect 21644 34850 21700 34862
rect 21756 34804 21812 34814
rect 21756 34710 21812 34748
rect 21532 32610 21588 32620
rect 21868 34692 21924 34702
rect 22204 34692 22260 35420
rect 22540 35140 22596 35534
rect 22316 35084 22596 35140
rect 22316 34914 22372 35084
rect 22316 34862 22318 34914
rect 22370 34862 22372 34914
rect 22316 34850 22372 34862
rect 22652 35026 22708 35038
rect 22652 34974 22654 35026
rect 22706 34974 22708 35026
rect 21868 34690 22260 34692
rect 21868 34638 21870 34690
rect 21922 34638 22260 34690
rect 21868 34636 22260 34638
rect 21868 32564 21924 34636
rect 22652 34020 22708 34974
rect 22652 33954 22708 33964
rect 21980 33460 22036 33470
rect 21980 32676 22036 33404
rect 22428 33348 22484 33358
rect 22316 33292 22428 33348
rect 22316 32788 22372 33292
rect 22428 33282 22484 33292
rect 22764 33124 22820 35644
rect 22876 33348 22932 37324
rect 23100 37156 23156 37166
rect 22988 35924 23044 35934
rect 22988 35810 23044 35868
rect 22988 35758 22990 35810
rect 23042 35758 23044 35810
rect 22988 35746 23044 35758
rect 23100 33796 23156 37100
rect 23212 36260 23268 36270
rect 23324 36260 23380 37772
rect 23548 36596 23604 40684
rect 23660 38948 23716 38958
rect 23660 38724 23716 38892
rect 23660 37266 23716 38668
rect 23660 37214 23662 37266
rect 23714 37214 23716 37266
rect 23660 37202 23716 37214
rect 23660 36596 23716 36606
rect 23604 36594 23716 36596
rect 23604 36542 23662 36594
rect 23714 36542 23716 36594
rect 23604 36540 23716 36542
rect 23548 36502 23604 36540
rect 23660 36530 23716 36540
rect 23212 36258 23380 36260
rect 23212 36206 23214 36258
rect 23266 36206 23380 36258
rect 23212 36204 23380 36206
rect 23212 35028 23268 36204
rect 23548 35924 23604 35934
rect 23548 35830 23604 35868
rect 23212 34962 23268 34972
rect 23772 34244 23828 41356
rect 24108 41188 24164 41198
rect 24220 41188 24276 42028
rect 24332 41972 24388 41982
rect 24444 41972 24500 44380
rect 24556 44212 24612 44222
rect 24556 44210 24836 44212
rect 24556 44158 24558 44210
rect 24610 44158 24836 44210
rect 24556 44156 24836 44158
rect 24556 44146 24612 44156
rect 24556 42754 24612 42766
rect 24556 42702 24558 42754
rect 24610 42702 24612 42754
rect 24556 42644 24612 42702
rect 24780 42756 24836 44156
rect 24892 44210 24948 45836
rect 24892 44158 24894 44210
rect 24946 44158 24948 44210
rect 24892 44146 24948 44158
rect 25004 43428 25060 46060
rect 25116 44548 25172 46172
rect 25564 45332 25620 45342
rect 25340 45108 25396 45118
rect 25340 45014 25396 45052
rect 25116 44482 25172 44492
rect 25116 44322 25172 44334
rect 25116 44270 25118 44322
rect 25170 44270 25172 44322
rect 25116 43652 25172 44270
rect 25116 43586 25172 43596
rect 25564 43538 25620 45276
rect 25564 43486 25566 43538
rect 25618 43486 25620 43538
rect 25564 43474 25620 43486
rect 25004 43372 25172 43428
rect 25004 43204 25060 43214
rect 24780 42700 24948 42756
rect 24556 42578 24612 42588
rect 24668 42532 24724 42542
rect 24556 42084 24612 42094
rect 24556 41990 24612 42028
rect 24332 41970 24500 41972
rect 24332 41918 24334 41970
rect 24386 41918 24500 41970
rect 24332 41916 24500 41918
rect 24332 41906 24388 41916
rect 24444 41860 24500 41916
rect 24444 41794 24500 41804
rect 24668 41748 24724 42476
rect 24780 42530 24836 42542
rect 24780 42478 24782 42530
rect 24834 42478 24836 42530
rect 24780 42196 24836 42478
rect 24780 42130 24836 42140
rect 24892 41860 24948 42700
rect 25004 42754 25060 43148
rect 25004 42702 25006 42754
rect 25058 42702 25060 42754
rect 25004 42690 25060 42702
rect 24892 41804 25060 41860
rect 25004 41748 25060 41804
rect 24668 41692 24948 41748
rect 24780 41524 24836 41534
rect 24108 41186 24276 41188
rect 24108 41134 24110 41186
rect 24162 41134 24276 41186
rect 24108 41132 24276 41134
rect 24444 41300 24500 41310
rect 24108 41122 24164 41132
rect 23884 40628 23940 40638
rect 23884 40534 23940 40572
rect 24332 40628 24388 40638
rect 24332 40514 24388 40572
rect 24444 40626 24500 41244
rect 24444 40574 24446 40626
rect 24498 40574 24500 40626
rect 24444 40562 24500 40574
rect 24668 41076 24724 41086
rect 24668 40626 24724 41020
rect 24780 41074 24836 41468
rect 24780 41022 24782 41074
rect 24834 41022 24836 41074
rect 24780 41010 24836 41022
rect 24668 40574 24670 40626
rect 24722 40574 24724 40626
rect 24668 40562 24724 40574
rect 24332 40462 24334 40514
rect 24386 40462 24388 40514
rect 24332 40450 24388 40462
rect 23996 40404 24052 40414
rect 23996 40402 24276 40404
rect 23996 40350 23998 40402
rect 24050 40350 24276 40402
rect 23996 40348 24276 40350
rect 23996 40338 24052 40348
rect 23884 40292 23940 40302
rect 23884 40178 23940 40236
rect 23884 40126 23886 40178
rect 23938 40126 23940 40178
rect 23884 40114 23940 40126
rect 24220 38722 24276 40348
rect 24220 38670 24222 38722
rect 24274 38670 24276 38722
rect 24220 38658 24276 38670
rect 24332 39732 24388 39742
rect 24332 38836 24388 39676
rect 24668 39060 24724 39070
rect 24668 38946 24724 39004
rect 24668 38894 24670 38946
rect 24722 38894 24724 38946
rect 24668 38882 24724 38894
rect 23884 38388 23940 38398
rect 23884 38162 23940 38332
rect 23884 38110 23886 38162
rect 23938 38110 23940 38162
rect 23884 38098 23940 38110
rect 24220 38052 24276 38062
rect 24108 37604 24164 37614
rect 24108 37266 24164 37548
rect 24220 37492 24276 37996
rect 24332 38050 24388 38780
rect 24556 38724 24612 38762
rect 24556 38658 24612 38668
rect 24892 38668 24948 41692
rect 25004 41682 25060 41692
rect 25116 41300 25172 43372
rect 25788 42980 25844 46172
rect 26012 43204 26068 49420
rect 26460 49364 26516 49646
rect 26348 49308 26516 49364
rect 26348 43764 26404 49308
rect 26460 49140 26516 49150
rect 26460 49046 26516 49084
rect 26572 47012 26628 49758
rect 26684 49140 26740 50540
rect 27020 50594 27076 53788
rect 27132 53778 27188 53788
rect 27132 53618 27188 53630
rect 27132 53566 27134 53618
rect 27186 53566 27188 53618
rect 27132 53172 27188 53566
rect 27244 53618 27300 54124
rect 27916 54068 27972 54350
rect 28364 54404 28420 54414
rect 28364 54310 28420 54348
rect 27916 54012 28196 54068
rect 27916 53844 27972 53854
rect 27916 53750 27972 53788
rect 27468 53732 27524 53742
rect 27692 53732 27748 53742
rect 27468 53730 27748 53732
rect 27468 53678 27470 53730
rect 27522 53678 27694 53730
rect 27746 53678 27748 53730
rect 27468 53676 27748 53678
rect 27468 53666 27524 53676
rect 27692 53666 27748 53676
rect 28028 53732 28084 53742
rect 28028 53638 28084 53676
rect 27244 53566 27246 53618
rect 27298 53566 27300 53618
rect 27244 53554 27300 53566
rect 27244 53172 27300 53182
rect 27132 53170 27300 53172
rect 27132 53118 27246 53170
rect 27298 53118 27300 53170
rect 27132 53116 27300 53118
rect 27244 52500 27300 53116
rect 27468 52948 27524 52958
rect 27468 52854 27524 52892
rect 27916 52948 27972 52958
rect 27916 52854 27972 52892
rect 27356 52836 27412 52846
rect 27356 52742 27412 52780
rect 27244 52434 27300 52444
rect 27916 52500 27972 52510
rect 27972 52444 28084 52500
rect 27916 52434 27972 52444
rect 27020 50542 27022 50594
rect 27074 50542 27076 50594
rect 27020 50530 27076 50542
rect 27244 52276 27300 52286
rect 26908 49812 26964 49822
rect 26908 49252 26964 49756
rect 27020 49810 27076 49822
rect 27020 49758 27022 49810
rect 27074 49758 27076 49810
rect 27020 49588 27076 49758
rect 27244 49812 27300 52220
rect 28028 51268 28084 52444
rect 28140 52388 28196 54012
rect 28588 53956 28644 55246
rect 29036 54404 29092 57148
rect 30156 57092 30212 57102
rect 29148 56980 29204 56990
rect 29148 56866 29204 56924
rect 29148 56814 29150 56866
rect 29202 56814 29204 56866
rect 29148 56802 29204 56814
rect 30156 56754 30212 57036
rect 30156 56702 30158 56754
rect 30210 56702 30212 56754
rect 30156 56690 30212 56702
rect 29484 56644 29540 56654
rect 29484 56642 29652 56644
rect 29484 56590 29486 56642
rect 29538 56590 29652 56642
rect 29484 56588 29652 56590
rect 29484 56578 29540 56588
rect 29484 55972 29540 55982
rect 29260 55970 29540 55972
rect 29260 55918 29486 55970
rect 29538 55918 29540 55970
rect 29260 55916 29540 55918
rect 29260 55298 29316 55916
rect 29484 55906 29540 55916
rect 29260 55246 29262 55298
rect 29314 55246 29316 55298
rect 29260 55234 29316 55246
rect 29148 55076 29204 55086
rect 29148 54982 29204 55020
rect 29596 54964 29652 56588
rect 29932 55970 29988 55982
rect 29932 55918 29934 55970
rect 29986 55918 29988 55970
rect 29932 55412 29988 55918
rect 29932 55346 29988 55356
rect 30044 55524 30100 55534
rect 29932 55074 29988 55086
rect 29932 55022 29934 55074
rect 29986 55022 29988 55074
rect 29820 54964 29876 54974
rect 29596 54908 29820 54964
rect 29148 54628 29204 54638
rect 29148 54534 29204 54572
rect 29484 54626 29540 54638
rect 29484 54574 29486 54626
rect 29538 54574 29540 54626
rect 29036 54348 29204 54404
rect 28588 53890 28644 53900
rect 28252 53508 28308 53518
rect 28252 52612 28308 53452
rect 28364 53172 28420 53182
rect 28364 53078 28420 53116
rect 29036 53060 29092 53070
rect 29036 52966 29092 53004
rect 28476 52946 28532 52958
rect 28476 52894 28478 52946
rect 28530 52894 28532 52946
rect 28364 52724 28420 52734
rect 28364 52630 28420 52668
rect 28252 52546 28308 52556
rect 28140 52332 28308 52388
rect 28252 51380 28308 52332
rect 28476 52276 28532 52894
rect 28812 52946 28868 52958
rect 28812 52894 28814 52946
rect 28866 52894 28868 52946
rect 28588 52276 28644 52286
rect 28476 52220 28588 52276
rect 28588 52182 28644 52220
rect 28812 52276 28868 52894
rect 28812 52210 28868 52220
rect 28924 52834 28980 52846
rect 28924 52782 28926 52834
rect 28978 52782 28980 52834
rect 28476 52052 28532 52062
rect 28924 52052 28980 52782
rect 29036 52724 29092 52734
rect 29036 52162 29092 52668
rect 29148 52500 29204 54348
rect 29484 53732 29540 54574
rect 29820 54626 29876 54908
rect 29820 54574 29822 54626
rect 29874 54574 29876 54626
rect 29820 54562 29876 54574
rect 29932 54852 29988 55022
rect 29372 53676 29484 53732
rect 29148 52434 29204 52444
rect 29260 52948 29316 52958
rect 29260 52386 29316 52892
rect 29260 52334 29262 52386
rect 29314 52334 29316 52386
rect 29260 52322 29316 52334
rect 29036 52110 29038 52162
rect 29090 52110 29092 52162
rect 29036 52098 29092 52110
rect 29148 52276 29204 52286
rect 28476 51602 28532 51996
rect 28476 51550 28478 51602
rect 28530 51550 28532 51602
rect 28476 51538 28532 51550
rect 28588 51996 28980 52052
rect 28588 51490 28644 51996
rect 28588 51438 28590 51490
rect 28642 51438 28644 51490
rect 28588 51426 28644 51438
rect 28252 51324 28532 51380
rect 28140 51268 28196 51278
rect 28028 51266 28196 51268
rect 28028 51214 28142 51266
rect 28194 51214 28196 51266
rect 28028 51212 28196 51214
rect 27468 50036 27524 50046
rect 27468 49942 27524 49980
rect 28140 50036 28196 51212
rect 28476 51156 28532 51324
rect 29036 51378 29092 51390
rect 29036 51326 29038 51378
rect 29090 51326 29092 51378
rect 28476 51100 28868 51156
rect 28140 49942 28196 49980
rect 28252 50596 28308 50606
rect 27244 49718 27300 49756
rect 27692 49922 27748 49934
rect 27692 49870 27694 49922
rect 27746 49870 27748 49922
rect 27356 49588 27412 49598
rect 27020 49586 27412 49588
rect 27020 49534 27358 49586
rect 27410 49534 27412 49586
rect 27020 49532 27412 49534
rect 27356 49522 27412 49532
rect 26684 49074 26740 49084
rect 26796 49196 26964 49252
rect 26572 46674 26628 46956
rect 26572 46622 26574 46674
rect 26626 46622 26628 46674
rect 26572 46610 26628 46622
rect 26796 47460 26852 49196
rect 26908 49140 26964 49196
rect 27244 49140 27300 49150
rect 26908 49138 27300 49140
rect 26908 49086 27246 49138
rect 27298 49086 27300 49138
rect 26908 49084 27300 49086
rect 27244 49074 27300 49084
rect 27692 49026 27748 49870
rect 28252 49922 28308 50540
rect 28252 49870 28254 49922
rect 28306 49870 28308 49922
rect 28252 49858 28308 49870
rect 28700 49812 28756 49822
rect 28700 49698 28756 49756
rect 28700 49646 28702 49698
rect 28754 49646 28756 49698
rect 28140 49586 28196 49598
rect 28140 49534 28142 49586
rect 28194 49534 28196 49586
rect 28140 49138 28196 49534
rect 28140 49086 28142 49138
rect 28194 49086 28196 49138
rect 28140 49074 28196 49086
rect 27692 48974 27694 49026
rect 27746 48974 27748 49026
rect 26796 46674 26852 47404
rect 26796 46622 26798 46674
rect 26850 46622 26852 46674
rect 26796 46610 26852 46622
rect 26908 48804 26964 48814
rect 26684 44210 26740 44222
rect 26684 44158 26686 44210
rect 26738 44158 26740 44210
rect 26460 44100 26516 44110
rect 26684 44100 26740 44158
rect 26516 44044 26740 44100
rect 26460 44006 26516 44044
rect 26348 43708 26628 43764
rect 26348 43428 26404 43466
rect 26348 43362 26404 43372
rect 26012 43138 26068 43148
rect 26348 43204 26404 43214
rect 26404 43148 26516 43204
rect 26348 43138 26404 43148
rect 25788 42924 26292 42980
rect 25788 42866 25844 42924
rect 25788 42814 25790 42866
rect 25842 42814 25844 42866
rect 25788 42802 25844 42814
rect 26236 42754 26292 42924
rect 26236 42702 26238 42754
rect 26290 42702 26292 42754
rect 26236 42690 26292 42702
rect 25228 42644 25284 42654
rect 25228 42194 25284 42588
rect 26012 42644 26068 42654
rect 26012 42550 26068 42588
rect 26348 42532 26404 42542
rect 26348 42438 26404 42476
rect 25228 42142 25230 42194
rect 25282 42142 25284 42194
rect 25228 42084 25284 42142
rect 25228 42018 25284 42028
rect 25788 42308 25844 42318
rect 26460 42308 26516 43148
rect 25452 41970 25508 41982
rect 25452 41918 25454 41970
rect 25506 41918 25508 41970
rect 25116 41234 25172 41244
rect 25340 41860 25396 41870
rect 25116 40962 25172 40974
rect 25116 40910 25118 40962
rect 25170 40910 25172 40962
rect 25116 40740 25172 40910
rect 25116 40292 25172 40684
rect 25340 40626 25396 41804
rect 25452 41748 25508 41918
rect 25452 41682 25508 41692
rect 25452 41300 25508 41310
rect 25452 40964 25508 41244
rect 25564 41186 25620 41198
rect 25564 41134 25566 41186
rect 25618 41134 25620 41186
rect 25564 41076 25620 41134
rect 25564 41010 25620 41020
rect 25788 41074 25844 42252
rect 26124 42252 26516 42308
rect 26124 41970 26180 42252
rect 26572 42196 26628 43708
rect 26796 43428 26852 43438
rect 26124 41918 26126 41970
rect 26178 41918 26180 41970
rect 26124 41906 26180 41918
rect 26236 42140 26628 42196
rect 26684 42754 26740 42766
rect 26684 42702 26686 42754
rect 26738 42702 26740 42754
rect 26684 42644 26740 42702
rect 26796 42754 26852 43372
rect 26796 42702 26798 42754
rect 26850 42702 26852 42754
rect 26796 42690 26852 42702
rect 26684 42194 26740 42588
rect 26908 42532 26964 48748
rect 27244 48132 27300 48142
rect 27244 48038 27300 48076
rect 27244 47796 27300 47806
rect 27132 46900 27188 46910
rect 27132 46806 27188 46844
rect 27020 45780 27076 45790
rect 27020 44322 27076 45724
rect 27132 45218 27188 45230
rect 27132 45166 27134 45218
rect 27186 45166 27188 45218
rect 27132 44434 27188 45166
rect 27132 44382 27134 44434
rect 27186 44382 27188 44434
rect 27132 44370 27188 44382
rect 27020 44270 27022 44322
rect 27074 44270 27076 44322
rect 27020 44258 27076 44270
rect 27132 44212 27188 44222
rect 27132 42754 27188 44156
rect 27244 44100 27300 47740
rect 27692 47570 27748 48974
rect 28700 48804 28756 49646
rect 27692 47518 27694 47570
rect 27746 47518 27748 47570
rect 27580 47348 27636 47358
rect 27468 46900 27524 46910
rect 27580 46900 27636 47292
rect 27692 47068 27748 47518
rect 28364 48748 28756 48804
rect 28028 47460 28084 47470
rect 28028 47366 28084 47404
rect 28140 47348 28196 47358
rect 28140 47234 28196 47292
rect 28140 47182 28142 47234
rect 28194 47182 28196 47234
rect 28140 47170 28196 47182
rect 28252 47236 28308 47246
rect 28252 47142 28308 47180
rect 27692 47012 27860 47068
rect 28364 47012 28420 48748
rect 28700 47458 28756 47470
rect 28700 47406 28702 47458
rect 28754 47406 28756 47458
rect 27468 46898 27636 46900
rect 27468 46846 27470 46898
rect 27522 46846 27636 46898
rect 27468 46844 27636 46846
rect 27692 46900 27748 46910
rect 27468 46834 27524 46844
rect 27692 46806 27748 46844
rect 27580 46564 27636 46574
rect 27580 46470 27636 46508
rect 27804 46340 27860 47012
rect 28028 46956 28420 47012
rect 28476 47012 28532 47022
rect 28028 46452 28084 46956
rect 28140 46676 28196 46686
rect 28364 46676 28420 46686
rect 28140 46674 28420 46676
rect 28140 46622 28142 46674
rect 28194 46622 28366 46674
rect 28418 46622 28420 46674
rect 28140 46620 28420 46622
rect 28140 46610 28196 46620
rect 28364 46610 28420 46620
rect 28028 46396 28196 46452
rect 27916 46340 27972 46350
rect 27804 46284 27916 46340
rect 27916 46274 27972 46284
rect 27580 46060 28084 46116
rect 27356 45780 27412 45790
rect 27356 45330 27412 45724
rect 27356 45278 27358 45330
rect 27410 45278 27412 45330
rect 27356 45266 27412 45278
rect 27580 45330 27636 46060
rect 27692 45892 27748 45902
rect 27692 45890 27972 45892
rect 27692 45838 27694 45890
rect 27746 45838 27972 45890
rect 27692 45836 27972 45838
rect 27692 45826 27748 45836
rect 27580 45278 27582 45330
rect 27634 45278 27636 45330
rect 27468 44994 27524 45006
rect 27468 44942 27470 44994
rect 27522 44942 27524 44994
rect 27468 44548 27524 44942
rect 27468 44482 27524 44492
rect 27580 44434 27636 45278
rect 27580 44382 27582 44434
rect 27634 44382 27636 44434
rect 27356 44324 27412 44334
rect 27580 44324 27636 44382
rect 27356 44322 27636 44324
rect 27356 44270 27358 44322
rect 27410 44270 27636 44322
rect 27356 44268 27636 44270
rect 27916 45332 27972 45836
rect 28028 45890 28084 46060
rect 28028 45838 28030 45890
rect 28082 45838 28084 45890
rect 28028 45826 28084 45838
rect 28028 45332 28084 45342
rect 27916 45330 28084 45332
rect 27916 45278 28030 45330
rect 28082 45278 28084 45330
rect 27916 45276 28084 45278
rect 27916 44322 27972 45276
rect 28028 45266 28084 45276
rect 27916 44270 27918 44322
rect 27970 44270 27972 44322
rect 27356 44258 27412 44268
rect 27916 44258 27972 44270
rect 28140 44100 28196 46396
rect 28476 46002 28532 46956
rect 28700 46900 28756 47406
rect 28700 46834 28756 46844
rect 28588 46786 28644 46798
rect 28588 46734 28590 46786
rect 28642 46734 28644 46786
rect 28588 46116 28644 46734
rect 28700 46674 28756 46686
rect 28700 46622 28702 46674
rect 28754 46622 28756 46674
rect 28700 46340 28756 46622
rect 28700 46274 28756 46284
rect 28588 46060 28756 46116
rect 28476 45950 28478 46002
rect 28530 45950 28532 46002
rect 28476 45938 28532 45950
rect 28476 45780 28532 45790
rect 28476 45686 28532 45724
rect 28700 45332 28756 46060
rect 28700 45266 28756 45276
rect 28588 45220 28644 45230
rect 28588 45126 28644 45164
rect 28476 45106 28532 45118
rect 28476 45054 28478 45106
rect 28530 45054 28532 45106
rect 28364 44996 28420 45006
rect 28364 44322 28420 44940
rect 28364 44270 28366 44322
rect 28418 44270 28420 44322
rect 28364 44258 28420 44270
rect 28476 44100 28532 45054
rect 27244 44044 27412 44100
rect 28140 44044 28420 44100
rect 27132 42702 27134 42754
rect 27186 42702 27188 42754
rect 27132 42690 27188 42702
rect 26908 42466 26964 42476
rect 27020 42530 27076 42542
rect 27020 42478 27022 42530
rect 27074 42478 27076 42530
rect 26684 42142 26686 42194
rect 26738 42142 26740 42194
rect 26236 41748 26292 42140
rect 26684 42130 26740 42142
rect 26908 42196 26964 42206
rect 27020 42196 27076 42478
rect 26908 42194 27076 42196
rect 26908 42142 26910 42194
rect 26962 42142 27076 42194
rect 26908 42140 27076 42142
rect 26908 42130 26964 42140
rect 27132 42082 27188 42094
rect 27132 42030 27134 42082
rect 27186 42030 27188 42082
rect 25788 41022 25790 41074
rect 25842 41022 25844 41074
rect 25788 41010 25844 41022
rect 25900 41692 26292 41748
rect 26460 41970 26516 41982
rect 26460 41918 26462 41970
rect 26514 41918 26516 41970
rect 25452 40898 25508 40908
rect 25340 40574 25342 40626
rect 25394 40574 25396 40626
rect 25340 40562 25396 40574
rect 25116 40226 25172 40236
rect 25452 40516 25508 40526
rect 25452 39060 25508 40460
rect 25788 40516 25844 40526
rect 25788 40422 25844 40460
rect 25452 38966 25508 39004
rect 25564 39396 25620 39406
rect 24892 38612 25172 38668
rect 24332 37998 24334 38050
rect 24386 37998 24388 38050
rect 24332 37986 24388 37998
rect 25004 37940 25060 37950
rect 25004 37846 25060 37884
rect 24332 37492 24388 37502
rect 24220 37490 24388 37492
rect 24220 37438 24334 37490
rect 24386 37438 24388 37490
rect 24220 37436 24388 37438
rect 24332 37426 24388 37436
rect 24444 37492 24500 37502
rect 24108 37214 24110 37266
rect 24162 37214 24164 37266
rect 24108 37202 24164 37214
rect 24444 36594 24500 37436
rect 24444 36542 24446 36594
rect 24498 36542 24500 36594
rect 24444 36530 24500 36542
rect 24556 37378 24612 37390
rect 24556 37326 24558 37378
rect 24610 37326 24612 37378
rect 23996 35924 24052 35934
rect 23996 35830 24052 35868
rect 24556 35140 24612 37326
rect 24668 37268 24724 37278
rect 24668 37174 24724 37212
rect 24892 36260 24948 36270
rect 24892 35364 24948 36204
rect 24892 35298 24948 35308
rect 24556 35074 24612 35084
rect 24780 34804 24836 34814
rect 24332 34802 24836 34804
rect 24332 34750 24782 34802
rect 24834 34750 24836 34802
rect 24332 34748 24836 34750
rect 24332 34354 24388 34748
rect 24780 34738 24836 34748
rect 24332 34302 24334 34354
rect 24386 34302 24388 34354
rect 24332 34290 24388 34302
rect 23996 34244 24052 34254
rect 23772 34242 24052 34244
rect 23772 34190 23998 34242
rect 24050 34190 24052 34242
rect 23772 34188 24052 34190
rect 25116 34244 25172 38612
rect 25340 37380 25396 37390
rect 25228 37378 25396 37380
rect 25228 37326 25342 37378
rect 25394 37326 25396 37378
rect 25228 37324 25396 37326
rect 25228 36260 25284 37324
rect 25340 37314 25396 37324
rect 25452 37268 25508 37278
rect 25452 37174 25508 37212
rect 25340 37156 25396 37166
rect 25340 37042 25396 37100
rect 25340 36990 25342 37042
rect 25394 36990 25396 37042
rect 25340 36978 25396 36990
rect 25564 36932 25620 39340
rect 25676 37266 25732 37278
rect 25676 37214 25678 37266
rect 25730 37214 25732 37266
rect 25676 37156 25732 37214
rect 25676 37090 25732 37100
rect 25788 37268 25844 37278
rect 25452 36876 25620 36932
rect 25452 36820 25508 36876
rect 25228 36194 25284 36204
rect 25340 36764 25508 36820
rect 25340 35308 25396 36764
rect 25676 36372 25732 36382
rect 25788 36372 25844 37212
rect 25900 36482 25956 41692
rect 26460 41188 26516 41918
rect 27132 41972 27188 42030
rect 27244 42084 27300 42094
rect 27244 41990 27300 42028
rect 26460 41122 26516 41132
rect 26572 41300 26628 41310
rect 27132 41300 27188 41916
rect 26572 41298 27188 41300
rect 26572 41246 26574 41298
rect 26626 41246 27188 41298
rect 26572 41244 27188 41246
rect 26124 40964 26180 40974
rect 26124 40870 26180 40908
rect 25900 36430 25902 36482
rect 25954 36430 25956 36482
rect 25900 36418 25956 36430
rect 26012 40740 26068 40750
rect 25676 36370 25844 36372
rect 25676 36318 25678 36370
rect 25730 36318 25844 36370
rect 25676 36316 25844 36318
rect 25676 36306 25732 36316
rect 26012 36260 26068 40684
rect 26460 40404 26516 40414
rect 26460 40310 26516 40348
rect 26236 37940 26292 37950
rect 26124 37492 26180 37502
rect 26124 37398 26180 37436
rect 26236 37490 26292 37884
rect 26236 37438 26238 37490
rect 26290 37438 26292 37490
rect 26236 37426 26292 37438
rect 26348 37266 26404 37278
rect 26348 37214 26350 37266
rect 26402 37214 26404 37266
rect 26348 36596 26404 37214
rect 26348 36530 26404 36540
rect 26460 36708 26516 36718
rect 25788 36204 26068 36260
rect 25788 35698 25844 36204
rect 26460 36036 26516 36652
rect 26012 35924 26068 35934
rect 26068 35868 26292 35924
rect 26012 35830 26068 35868
rect 25788 35646 25790 35698
rect 25842 35646 25844 35698
rect 25788 35634 25844 35646
rect 25228 35252 25396 35308
rect 25228 34468 25284 35252
rect 25564 34916 25620 34926
rect 25564 34914 26180 34916
rect 25564 34862 25566 34914
rect 25618 34862 26180 34914
rect 25564 34860 26180 34862
rect 25564 34850 25620 34860
rect 25228 34402 25284 34412
rect 25900 34690 25956 34702
rect 25900 34638 25902 34690
rect 25954 34638 25956 34690
rect 25228 34244 25284 34254
rect 25116 34242 25284 34244
rect 25116 34190 25230 34242
rect 25282 34190 25284 34242
rect 25116 34188 25284 34190
rect 23996 34178 24052 34188
rect 25228 34178 25284 34188
rect 23660 34132 23716 34142
rect 23660 34038 23716 34076
rect 24220 34130 24276 34142
rect 24220 34078 24222 34130
rect 24274 34078 24276 34130
rect 23212 34020 23268 34030
rect 23548 34020 23604 34030
rect 23268 34018 23604 34020
rect 23268 33966 23550 34018
rect 23602 33966 23604 34018
rect 23268 33964 23604 33966
rect 23212 33926 23268 33964
rect 23548 33954 23604 33964
rect 23100 33740 23380 33796
rect 23100 33458 23156 33470
rect 23100 33406 23102 33458
rect 23154 33406 23156 33458
rect 22932 33292 23044 33348
rect 22876 33282 22932 33292
rect 22540 33068 22820 33124
rect 22540 32900 22596 33068
rect 22540 32844 22708 32900
rect 22428 32788 22484 32798
rect 22316 32786 22484 32788
rect 22316 32734 22430 32786
rect 22482 32734 22484 32786
rect 22316 32732 22484 32734
rect 22428 32722 22484 32732
rect 21980 32610 22036 32620
rect 22540 32676 22596 32686
rect 22540 32582 22596 32620
rect 21308 32162 21364 32172
rect 21756 32508 21924 32564
rect 21644 32004 21700 32014
rect 20860 32002 21700 32004
rect 20860 31950 21646 32002
rect 21698 31950 21700 32002
rect 20860 31948 21700 31950
rect 20860 31106 20916 31948
rect 21644 31938 21700 31948
rect 21756 31780 21812 32508
rect 21980 32452 22036 32462
rect 22428 32452 22484 32462
rect 20860 31054 20862 31106
rect 20914 31054 20916 31106
rect 20860 31042 20916 31054
rect 21644 31724 21812 31780
rect 21868 32450 22036 32452
rect 21868 32398 21982 32450
rect 22034 32398 22036 32450
rect 21868 32396 22036 32398
rect 21532 30884 21588 30894
rect 21644 30884 21700 31724
rect 21588 30828 21700 30884
rect 21756 31554 21812 31566
rect 21756 31502 21758 31554
rect 21810 31502 21812 31554
rect 21532 30210 21588 30828
rect 21532 30158 21534 30210
rect 21586 30158 21588 30210
rect 21532 30146 21588 30158
rect 21756 30212 21812 31502
rect 21868 30884 21924 32396
rect 21980 32386 22036 32396
rect 22092 32450 22484 32452
rect 22092 32398 22430 32450
rect 22482 32398 22484 32450
rect 22092 32396 22484 32398
rect 21980 32004 22036 32014
rect 22092 32004 22148 32396
rect 22428 32386 22484 32396
rect 21980 32002 22148 32004
rect 21980 31950 21982 32002
rect 22034 31950 22148 32002
rect 21980 31948 22148 31950
rect 21980 31938 22036 31948
rect 22652 31666 22708 32844
rect 22988 32788 23044 33292
rect 23100 33124 23156 33406
rect 23100 33058 23156 33068
rect 22876 32732 23044 32788
rect 22764 32562 22820 32574
rect 22764 32510 22766 32562
rect 22818 32510 22820 32562
rect 22764 32228 22820 32510
rect 22764 32162 22820 32172
rect 22652 31614 22654 31666
rect 22706 31614 22708 31666
rect 22316 31554 22372 31566
rect 22540 31556 22596 31566
rect 22316 31502 22318 31554
rect 22370 31502 22372 31554
rect 22316 30884 22372 31502
rect 21868 30828 22372 30884
rect 22428 31500 22540 31556
rect 21756 30146 21812 30156
rect 21868 30210 21924 30222
rect 21868 30158 21870 30210
rect 21922 30158 21924 30210
rect 20860 29988 20916 29998
rect 20860 29986 21252 29988
rect 20860 29934 20862 29986
rect 20914 29934 21252 29986
rect 20860 29932 21252 29934
rect 20860 29922 20916 29932
rect 21196 28644 21252 29932
rect 21308 29986 21364 29998
rect 21308 29934 21310 29986
rect 21362 29934 21364 29986
rect 21308 29204 21364 29934
rect 21420 29986 21476 29998
rect 21420 29934 21422 29986
rect 21474 29934 21476 29986
rect 21420 29428 21476 29934
rect 21868 29876 21924 30158
rect 21868 29810 21924 29820
rect 21756 29652 21812 29662
rect 21812 29596 21924 29652
rect 21756 29586 21812 29596
rect 21420 29372 21812 29428
rect 21308 29148 21700 29204
rect 21644 28754 21700 29148
rect 21644 28702 21646 28754
rect 21698 28702 21700 28754
rect 21644 28690 21700 28702
rect 21420 28644 21476 28654
rect 21196 28642 21476 28644
rect 21196 28590 21422 28642
rect 21474 28590 21476 28642
rect 21196 28588 21476 28590
rect 20636 28364 21252 28420
rect 21084 28196 21140 28206
rect 20748 27412 20804 27422
rect 20636 26290 20692 26302
rect 20636 26238 20638 26290
rect 20690 26238 20692 26290
rect 20636 26180 20692 26238
rect 20636 26114 20692 26124
rect 20636 25732 20692 25742
rect 20748 25732 20804 27356
rect 20860 27188 20916 27198
rect 20860 27094 20916 27132
rect 20972 26068 21028 26078
rect 20972 25974 21028 26012
rect 20636 25730 20804 25732
rect 20636 25678 20638 25730
rect 20690 25678 20804 25730
rect 20636 25676 20804 25678
rect 20636 25666 20692 25676
rect 20748 25394 20804 25406
rect 20748 25342 20750 25394
rect 20802 25342 20804 25394
rect 20636 25282 20692 25294
rect 20636 25230 20638 25282
rect 20690 25230 20692 25282
rect 20636 24052 20692 25230
rect 20748 24500 20804 25342
rect 20748 24434 20804 24444
rect 21084 24052 21140 28140
rect 21196 24276 21252 28364
rect 21308 26964 21364 27002
rect 21308 26898 21364 26908
rect 21420 24724 21476 28588
rect 21756 28308 21812 29372
rect 21868 28644 21924 29596
rect 21868 28550 21924 28588
rect 21980 28642 22036 30828
rect 22316 30212 22372 30222
rect 22316 30118 22372 30156
rect 22204 30098 22260 30110
rect 22204 30046 22206 30098
rect 22258 30046 22260 30098
rect 22204 29988 22260 30046
rect 21980 28590 21982 28642
rect 22034 28590 22036 28642
rect 21980 28578 22036 28590
rect 22092 29092 22148 29102
rect 21532 28252 21812 28308
rect 21980 28420 22036 28430
rect 21532 27972 21588 28252
rect 21532 26962 21588 27916
rect 21980 27746 22036 28364
rect 21980 27694 21982 27746
rect 22034 27694 22036 27746
rect 21644 27636 21700 27646
rect 21644 27074 21700 27580
rect 21980 27524 22036 27694
rect 21980 27458 22036 27468
rect 21644 27022 21646 27074
rect 21698 27022 21700 27074
rect 21644 27010 21700 27022
rect 21532 26910 21534 26962
rect 21586 26910 21588 26962
rect 21532 26898 21588 26910
rect 21532 26404 21588 26414
rect 21532 26178 21588 26348
rect 21532 26126 21534 26178
rect 21586 26126 21588 26178
rect 21532 25284 21588 26126
rect 21644 26292 21700 26302
rect 21644 25620 21700 26236
rect 21644 25554 21700 25564
rect 21868 25394 21924 25406
rect 21868 25342 21870 25394
rect 21922 25342 21924 25394
rect 21588 25228 21812 25284
rect 21532 25190 21588 25228
rect 21420 24658 21476 24668
rect 21196 24220 21700 24276
rect 21532 24052 21588 24062
rect 20636 24050 21588 24052
rect 20636 23998 21534 24050
rect 21586 23998 21588 24050
rect 20636 23996 21588 23998
rect 21532 23986 21588 23996
rect 20748 23828 20804 23838
rect 20524 23826 20804 23828
rect 20524 23774 20750 23826
rect 20802 23774 20804 23826
rect 20524 23772 20804 23774
rect 20300 23714 20356 23726
rect 20300 23662 20302 23714
rect 20354 23662 20356 23714
rect 20300 23604 20356 23662
rect 19836 23548 20100 23558
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20300 23538 20356 23548
rect 19836 23482 20100 23492
rect 19068 21746 19124 21756
rect 19292 22988 19684 23044
rect 20300 23156 20356 23166
rect 20300 23042 20356 23100
rect 20300 22990 20302 23042
rect 20354 22990 20356 23042
rect 18956 21476 19012 21486
rect 18844 21474 19012 21476
rect 18844 21422 18958 21474
rect 19010 21422 19012 21474
rect 18844 21420 19012 21422
rect 18956 21028 19012 21420
rect 18508 20190 18510 20242
rect 18562 20190 18564 20242
rect 18508 20178 18564 20190
rect 18732 20972 19012 21028
rect 19292 21028 19348 22988
rect 19628 22820 19684 22830
rect 19516 22764 19628 22820
rect 19516 22372 19572 22764
rect 19628 22754 19684 22764
rect 19740 22372 19796 22382
rect 19404 22370 19572 22372
rect 19404 22318 19518 22370
rect 19570 22318 19572 22370
rect 19404 22316 19572 22318
rect 19404 21140 19460 22316
rect 19516 22306 19572 22316
rect 19628 22370 19796 22372
rect 19628 22318 19742 22370
rect 19794 22318 19796 22370
rect 19628 22316 19796 22318
rect 19516 21700 19572 21710
rect 19516 21586 19572 21644
rect 19516 21534 19518 21586
rect 19570 21534 19572 21586
rect 19516 21522 19572 21534
rect 19628 21140 19684 22316
rect 19740 22306 19796 22316
rect 19836 21980 20100 21990
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 19836 21914 20100 21924
rect 20300 21700 20356 22990
rect 20524 22820 20580 23772
rect 20748 23762 20804 23772
rect 20524 22754 20580 22764
rect 20636 23604 20692 23614
rect 20636 23154 20692 23548
rect 21644 23492 21700 24220
rect 21644 23426 21700 23436
rect 20972 23268 21028 23278
rect 20972 23174 21028 23212
rect 20636 23102 20638 23154
rect 20690 23102 20692 23154
rect 20524 22594 20580 22606
rect 20524 22542 20526 22594
rect 20578 22542 20580 22594
rect 20076 21644 20356 21700
rect 20412 22370 20468 22382
rect 20412 22318 20414 22370
rect 20466 22318 20468 22370
rect 19404 21084 19572 21140
rect 19292 20972 19460 21028
rect 18732 20018 18788 20972
rect 19292 20244 19348 20254
rect 18732 19966 18734 20018
rect 18786 19966 18788 20018
rect 17948 19282 18004 19292
rect 18620 19908 18676 19918
rect 17836 19182 17838 19234
rect 17890 19182 17892 19234
rect 17836 19170 17892 19182
rect 18620 19234 18676 19852
rect 18620 19182 18622 19234
rect 18674 19182 18676 19234
rect 18620 19170 18676 19182
rect 17724 18452 17780 18462
rect 17612 18450 17780 18452
rect 17612 18398 17726 18450
rect 17778 18398 17780 18450
rect 17612 18396 17780 18398
rect 18732 18452 18788 19966
rect 19180 20018 19236 20030
rect 19180 19966 19182 20018
rect 19234 19966 19236 20018
rect 19068 19234 19124 19246
rect 19068 19182 19070 19234
rect 19122 19182 19124 19234
rect 18956 18452 19012 18462
rect 18732 18450 19012 18452
rect 18732 18398 18958 18450
rect 19010 18398 19012 18450
rect 18732 18396 19012 18398
rect 17388 17778 17444 18396
rect 17388 17726 17390 17778
rect 17442 17726 17444 17778
rect 17388 17714 17444 17726
rect 17724 17780 17780 18396
rect 18060 18340 18116 18350
rect 17724 17714 17780 17724
rect 17948 17892 18004 17902
rect 17276 17052 17668 17108
rect 17500 16884 17556 16894
rect 17276 16324 17332 16334
rect 17276 16210 17332 16268
rect 17276 16158 17278 16210
rect 17330 16158 17332 16210
rect 17276 16146 17332 16158
rect 16940 8372 17108 8428
rect 17500 8428 17556 16828
rect 17612 16772 17668 17052
rect 17612 16770 17892 16772
rect 17612 16718 17614 16770
rect 17666 16718 17892 16770
rect 17612 16716 17892 16718
rect 17612 16706 17668 16716
rect 17836 16098 17892 16716
rect 17836 16046 17838 16098
rect 17890 16046 17892 16098
rect 17724 15316 17780 15326
rect 17836 15316 17892 16046
rect 17724 15314 17836 15316
rect 17724 15262 17726 15314
rect 17778 15262 17836 15314
rect 17724 15260 17836 15262
rect 17724 15250 17780 15260
rect 17836 15222 17892 15260
rect 17948 14530 18004 17836
rect 18060 17668 18116 18284
rect 18060 17574 18116 17612
rect 18284 18340 18340 18350
rect 18284 16884 18340 18284
rect 18620 18340 18676 18350
rect 18620 18338 18788 18340
rect 18620 18286 18622 18338
rect 18674 18286 18788 18338
rect 18620 18284 18788 18286
rect 18620 18274 18676 18284
rect 18508 18228 18564 18238
rect 18284 16818 18340 16828
rect 18396 18226 18564 18228
rect 18396 18174 18510 18226
rect 18562 18174 18564 18226
rect 18396 18172 18564 18174
rect 18396 15202 18452 18172
rect 18508 18162 18564 18172
rect 18508 17666 18564 17678
rect 18508 17614 18510 17666
rect 18562 17614 18564 17666
rect 18508 17444 18564 17614
rect 18620 17444 18676 17454
rect 18508 17388 18620 17444
rect 18620 17378 18676 17388
rect 18620 16212 18676 16222
rect 18620 16118 18676 16156
rect 18396 15150 18398 15202
rect 18450 15150 18452 15202
rect 18396 15138 18452 15150
rect 18508 15316 18564 15326
rect 17948 14478 17950 14530
rect 18002 14478 18004 14530
rect 17948 14466 18004 14478
rect 18172 14530 18228 14542
rect 18172 14478 18174 14530
rect 18226 14478 18228 14530
rect 17500 8372 17780 8428
rect 16380 3378 16436 3388
rect 16828 4226 16884 4238
rect 16828 4174 16830 4226
rect 16882 4174 16884 4226
rect 15820 3164 16212 3220
rect 16156 800 16212 3164
rect 16828 2548 16884 4174
rect 16940 3444 16996 8372
rect 17276 3554 17332 3566
rect 17276 3502 17278 3554
rect 17330 3502 17332 3554
rect 17052 3444 17108 3454
rect 16940 3442 17108 3444
rect 16940 3390 17054 3442
rect 17106 3390 17108 3442
rect 16940 3388 17108 3390
rect 17052 3378 17108 3388
rect 17276 2548 17332 3502
rect 17724 3444 17780 8372
rect 17724 3378 17780 3388
rect 17948 3554 18004 3566
rect 17948 3502 17950 3554
rect 18002 3502 18004 3554
rect 16828 2492 17332 2548
rect 17948 2548 18004 3502
rect 18172 3442 18228 14478
rect 18508 13746 18564 15260
rect 18732 14754 18788 18284
rect 18956 17892 19012 18396
rect 18956 17826 19012 17836
rect 18956 17666 19012 17678
rect 18956 17614 18958 17666
rect 19010 17614 19012 17666
rect 18956 16324 19012 17614
rect 18956 15652 19012 16268
rect 18956 15586 19012 15596
rect 19068 15540 19124 19182
rect 19180 18676 19236 19966
rect 19292 19794 19348 20188
rect 19292 19742 19294 19794
rect 19346 19742 19348 19794
rect 19292 19730 19348 19742
rect 19180 18620 19348 18676
rect 19068 15474 19124 15484
rect 19180 18450 19236 18462
rect 19180 18398 19182 18450
rect 19234 18398 19236 18450
rect 19180 14756 19236 18398
rect 19292 18340 19348 18620
rect 19292 18274 19348 18284
rect 18732 14702 18734 14754
rect 18786 14702 18788 14754
rect 18732 14690 18788 14702
rect 18844 14700 19236 14756
rect 19292 17668 19348 17678
rect 18508 13694 18510 13746
rect 18562 13694 18564 13746
rect 18508 13682 18564 13694
rect 18396 11508 18452 11518
rect 18396 11394 18452 11452
rect 18396 11342 18398 11394
rect 18450 11342 18452 11394
rect 18396 11330 18452 11342
rect 18732 11396 18788 11406
rect 18732 11302 18788 11340
rect 18172 3390 18174 3442
rect 18226 3390 18228 3442
rect 18172 3378 18228 3390
rect 18396 4226 18452 4238
rect 18396 4174 18398 4226
rect 18450 4174 18452 4226
rect 18396 2548 18452 4174
rect 17948 2492 18452 2548
rect 18620 3554 18676 3566
rect 18620 3502 18622 3554
rect 18674 3502 18676 3554
rect 18620 2548 18676 3502
rect 18844 3442 18900 14700
rect 19292 14530 19348 17612
rect 19292 14478 19294 14530
rect 19346 14478 19348 14530
rect 19292 14466 19348 14478
rect 19292 14308 19348 14318
rect 19292 13858 19348 14252
rect 19292 13806 19294 13858
rect 19346 13806 19348 13858
rect 19292 13794 19348 13806
rect 19404 12180 19460 20972
rect 19516 20020 19572 21084
rect 19628 21084 20020 21140
rect 19628 20132 19684 21084
rect 19964 20914 20020 21084
rect 19964 20862 19966 20914
rect 20018 20862 20020 20914
rect 19964 20850 20020 20862
rect 20076 20916 20132 21644
rect 20188 21474 20244 21486
rect 20188 21422 20190 21474
rect 20242 21422 20244 21474
rect 20188 21028 20244 21422
rect 20412 21476 20468 22318
rect 20412 21410 20468 21420
rect 20300 21028 20356 21038
rect 20188 21026 20356 21028
rect 20188 20974 20302 21026
rect 20354 20974 20356 21026
rect 20188 20972 20356 20974
rect 20300 20962 20356 20972
rect 20412 20916 20468 20926
rect 20524 20916 20580 22542
rect 20076 20860 20244 20916
rect 20188 20804 20244 20860
rect 20412 20914 20580 20916
rect 20412 20862 20414 20914
rect 20466 20862 20580 20914
rect 20412 20860 20580 20862
rect 20412 20850 20468 20860
rect 20188 20748 20356 20804
rect 19836 20412 20100 20422
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 19836 20346 20100 20356
rect 19628 20066 19684 20076
rect 19516 19954 19572 19964
rect 19964 20020 20020 20030
rect 19964 19926 20020 19964
rect 19628 19906 19684 19918
rect 19628 19854 19630 19906
rect 19682 19854 19684 19906
rect 19628 18676 19684 19854
rect 19852 19348 19908 19358
rect 19852 19254 19908 19292
rect 19836 18844 20100 18854
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 19836 18778 20100 18788
rect 19628 18620 19796 18676
rect 19740 18452 19796 18620
rect 19740 18386 19796 18396
rect 20188 18450 20244 18462
rect 20188 18398 20190 18450
rect 20242 18398 20244 18450
rect 19628 18226 19684 18238
rect 19628 18174 19630 18226
rect 19682 18174 19684 18226
rect 19628 17778 19684 18174
rect 19628 17726 19630 17778
rect 19682 17726 19684 17778
rect 19628 17714 19684 17726
rect 20076 17780 20132 17790
rect 20076 17686 20132 17724
rect 20188 17668 20244 18398
rect 20188 17602 20244 17612
rect 19516 17554 19572 17566
rect 19516 17502 19518 17554
rect 19570 17502 19572 17554
rect 19516 16212 19572 17502
rect 20188 17444 20244 17454
rect 19836 17276 20100 17286
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 19836 17210 20100 17220
rect 19516 16146 19572 16156
rect 19836 15708 20100 15718
rect 19628 15652 19684 15662
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 19836 15642 20100 15652
rect 19628 14530 19684 15596
rect 19628 14478 19630 14530
rect 19682 14478 19684 14530
rect 19628 14466 19684 14478
rect 19964 14532 20020 14542
rect 20188 14532 20244 17388
rect 19964 14530 20244 14532
rect 19964 14478 19966 14530
rect 20018 14478 20244 14530
rect 19964 14476 20244 14478
rect 19964 14466 20020 14476
rect 20300 14308 20356 20748
rect 20412 20020 20468 20030
rect 20412 19346 20468 19964
rect 20636 19796 20692 23102
rect 21420 23042 21476 23054
rect 21420 22990 21422 23042
rect 21474 22990 21476 23042
rect 21420 22372 21476 22990
rect 21756 23044 21812 25228
rect 21868 25172 21924 25342
rect 21868 24612 21924 25116
rect 21868 24546 21924 24556
rect 22092 24948 22148 29036
rect 22204 28420 22260 29932
rect 22428 28868 22484 31500
rect 22540 31490 22596 31500
rect 22540 30212 22596 30222
rect 22540 30118 22596 30156
rect 22652 29988 22708 31614
rect 22876 31332 22932 32732
rect 22876 30884 22932 31276
rect 22988 32562 23044 32574
rect 22988 32510 22990 32562
rect 23042 32510 23044 32562
rect 22988 31108 23044 32510
rect 23324 32004 23380 33740
rect 24220 32788 24276 34078
rect 24444 34132 24500 34142
rect 24444 34038 24500 34076
rect 24668 34130 24724 34142
rect 24668 34078 24670 34130
rect 24722 34078 24724 34130
rect 24668 34020 24724 34078
rect 24668 33954 24724 33964
rect 24780 34132 24836 34142
rect 24220 32722 24276 32732
rect 24780 32786 24836 34076
rect 25452 34132 25508 34142
rect 25452 34038 25508 34076
rect 25676 34132 25732 34142
rect 25676 34038 25732 34076
rect 25788 34132 25844 34142
rect 25900 34132 25956 34638
rect 25788 34130 25956 34132
rect 25788 34078 25790 34130
rect 25842 34078 25956 34130
rect 25788 34076 25956 34078
rect 25564 34018 25620 34030
rect 25564 33966 25566 34018
rect 25618 33966 25620 34018
rect 25228 33796 25284 33806
rect 25228 33684 25284 33740
rect 25004 33628 25284 33684
rect 24780 32734 24782 32786
rect 24834 32734 24836 32786
rect 24780 32722 24836 32734
rect 24892 33236 24948 33246
rect 24556 32676 24612 32686
rect 24892 32676 24948 33180
rect 24556 32674 24724 32676
rect 24556 32622 24558 32674
rect 24610 32622 24724 32674
rect 24556 32620 24724 32622
rect 24556 32610 24612 32620
rect 24444 32564 24500 32574
rect 23436 32450 23492 32462
rect 23436 32398 23438 32450
rect 23490 32398 23492 32450
rect 23436 32228 23492 32398
rect 23436 32162 23492 32172
rect 24220 32450 24276 32462
rect 24220 32398 24222 32450
rect 24274 32398 24276 32450
rect 24220 32004 24276 32398
rect 23324 31948 23492 32004
rect 22988 31042 23044 31052
rect 23100 31892 23156 31902
rect 22988 30884 23044 30894
rect 22764 30882 23044 30884
rect 22764 30830 22990 30882
rect 23042 30830 23044 30882
rect 22764 30828 23044 30830
rect 22764 30210 22820 30828
rect 22988 30818 23044 30828
rect 22764 30158 22766 30210
rect 22818 30158 22820 30210
rect 22764 30146 22820 30158
rect 22652 29932 23044 29988
rect 22540 29876 22596 29886
rect 22596 29820 22932 29876
rect 22540 29810 22596 29820
rect 22652 29650 22708 29662
rect 22652 29598 22654 29650
rect 22706 29598 22708 29650
rect 22652 29428 22708 29598
rect 22652 29426 22820 29428
rect 22652 29374 22654 29426
rect 22706 29374 22820 29426
rect 22652 29372 22820 29374
rect 22652 29362 22708 29372
rect 22652 29204 22708 29214
rect 22540 28868 22596 28878
rect 22428 28866 22596 28868
rect 22428 28814 22542 28866
rect 22594 28814 22596 28866
rect 22428 28812 22596 28814
rect 22540 28802 22596 28812
rect 22652 28642 22708 29148
rect 22652 28590 22654 28642
rect 22706 28590 22708 28642
rect 22652 28578 22708 28590
rect 22540 28420 22596 28430
rect 22204 28354 22260 28364
rect 22428 28418 22596 28420
rect 22428 28366 22542 28418
rect 22594 28366 22596 28418
rect 22428 28364 22596 28366
rect 22428 28084 22484 28364
rect 22540 28354 22596 28364
rect 21868 23714 21924 23726
rect 21868 23662 21870 23714
rect 21922 23662 21924 23714
rect 21868 23548 21924 23662
rect 22092 23548 22148 24892
rect 22204 28028 22484 28084
rect 22540 28084 22596 28094
rect 22204 27188 22260 28028
rect 22540 27990 22596 28028
rect 22204 23604 22260 27132
rect 22316 27858 22372 27870
rect 22316 27806 22318 27858
rect 22370 27806 22372 27858
rect 22316 26292 22372 27806
rect 22428 27748 22484 27758
rect 22428 27654 22484 27692
rect 22540 27636 22596 27646
rect 22428 27524 22484 27534
rect 22428 27074 22484 27468
rect 22540 27298 22596 27580
rect 22540 27246 22542 27298
rect 22594 27246 22596 27298
rect 22540 27234 22596 27246
rect 22652 27188 22708 27198
rect 22652 27094 22708 27132
rect 22428 27022 22430 27074
rect 22482 27022 22484 27074
rect 22428 27010 22484 27022
rect 22316 26226 22372 26236
rect 22428 26852 22484 26862
rect 22428 24834 22484 26796
rect 22428 24782 22430 24834
rect 22482 24782 22484 24834
rect 22428 24770 22484 24782
rect 22540 26290 22596 26302
rect 22540 26238 22542 26290
rect 22594 26238 22596 26290
rect 22204 23548 22484 23604
rect 21868 23492 22148 23548
rect 21868 23380 21924 23492
rect 21868 23314 21924 23324
rect 22204 23380 22260 23390
rect 22204 23286 22260 23324
rect 21756 22988 22036 23044
rect 21420 22306 21476 22316
rect 21980 22932 22036 22988
rect 22092 22932 22148 22942
rect 21980 22930 22148 22932
rect 21980 22878 22094 22930
rect 22146 22878 22148 22930
rect 21980 22876 22148 22878
rect 20748 22260 20804 22270
rect 20748 22258 21364 22260
rect 20748 22206 20750 22258
rect 20802 22206 21364 22258
rect 20748 22204 21364 22206
rect 20748 22194 20804 22204
rect 21308 20914 21364 22204
rect 21308 20862 21310 20914
rect 21362 20862 21364 20914
rect 20860 20132 20916 20142
rect 20860 20018 20916 20076
rect 20860 19966 20862 20018
rect 20914 19966 20916 20018
rect 20860 19954 20916 19966
rect 21308 19906 21364 20862
rect 21868 21700 21924 21710
rect 21532 20802 21588 20814
rect 21532 20750 21534 20802
rect 21586 20750 21588 20802
rect 21308 19854 21310 19906
rect 21362 19854 21364 19906
rect 20636 19740 20916 19796
rect 20412 19294 20414 19346
rect 20466 19294 20468 19346
rect 20412 19282 20468 19294
rect 20748 19124 20804 19134
rect 20748 19030 20804 19068
rect 20636 18452 20692 18462
rect 20524 18450 20692 18452
rect 20524 18398 20638 18450
rect 20690 18398 20692 18450
rect 20524 18396 20692 18398
rect 20524 15202 20580 18396
rect 20636 18386 20692 18396
rect 20748 18452 20804 18462
rect 20748 16210 20804 18396
rect 20748 16158 20750 16210
rect 20802 16158 20804 16210
rect 20748 16146 20804 16158
rect 20524 15150 20526 15202
rect 20578 15150 20580 15202
rect 20412 14532 20468 14542
rect 20524 14532 20580 15150
rect 20412 14530 20580 14532
rect 20412 14478 20414 14530
rect 20466 14478 20580 14530
rect 20412 14476 20580 14478
rect 20412 14466 20468 14476
rect 20300 14252 20804 14308
rect 19836 14140 20100 14150
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 19836 14074 20100 14084
rect 20748 13076 20804 14252
rect 20748 12982 20804 13020
rect 19836 12572 20100 12582
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 19836 12506 20100 12516
rect 19964 12404 20020 12414
rect 19964 12310 20020 12348
rect 20860 12404 20916 19740
rect 21308 19348 21364 19854
rect 20972 19346 21364 19348
rect 20972 19294 21310 19346
rect 21362 19294 21364 19346
rect 20972 19292 21364 19294
rect 20972 18450 21028 19292
rect 21308 19282 21364 19292
rect 21420 20020 21476 20030
rect 20972 18398 20974 18450
rect 21026 18398 21028 18450
rect 20972 18386 21028 18398
rect 21084 18452 21140 18462
rect 21084 18358 21140 18396
rect 21420 17666 21476 19964
rect 21532 18116 21588 20750
rect 21868 20020 21924 21644
rect 21868 19926 21924 19964
rect 21756 19348 21812 19358
rect 21756 19234 21812 19292
rect 21756 19182 21758 19234
rect 21810 19182 21812 19234
rect 21756 19170 21812 19182
rect 21868 19236 21924 19246
rect 21532 18050 21588 18060
rect 21420 17614 21422 17666
rect 21474 17614 21476 17666
rect 21420 17602 21476 17614
rect 21868 16882 21924 19180
rect 21868 16830 21870 16882
rect 21922 16830 21924 16882
rect 21868 16212 21924 16830
rect 21868 16146 21924 16156
rect 21868 15314 21924 15326
rect 21868 15262 21870 15314
rect 21922 15262 21924 15314
rect 21868 15090 21924 15262
rect 21868 15038 21870 15090
rect 21922 15038 21924 15090
rect 21868 15026 21924 15038
rect 21868 14644 21924 14654
rect 21980 14644 22036 22876
rect 22092 22866 22148 22876
rect 22428 21588 22484 23548
rect 22540 23156 22596 26238
rect 22764 25172 22820 29372
rect 22876 28866 22932 29820
rect 22876 28814 22878 28866
rect 22930 28814 22932 28866
rect 22876 28802 22932 28814
rect 22988 28530 23044 29932
rect 23100 29650 23156 31836
rect 23212 30884 23268 30894
rect 23212 30790 23268 30828
rect 23324 30098 23380 30110
rect 23324 30046 23326 30098
rect 23378 30046 23380 30098
rect 23212 29988 23268 29998
rect 23324 29988 23380 30046
rect 23268 29932 23380 29988
rect 23212 29922 23268 29932
rect 23100 29598 23102 29650
rect 23154 29598 23156 29650
rect 23100 29586 23156 29598
rect 23324 29314 23380 29326
rect 23324 29262 23326 29314
rect 23378 29262 23380 29314
rect 23324 28980 23380 29262
rect 23436 29092 23492 31948
rect 24220 31938 24276 31948
rect 24444 32002 24500 32508
rect 24444 31950 24446 32002
rect 24498 31950 24500 32002
rect 24444 31938 24500 31950
rect 23996 31892 24052 31902
rect 23548 31556 23604 31566
rect 23548 31554 23716 31556
rect 23548 31502 23550 31554
rect 23602 31502 23716 31554
rect 23548 31500 23716 31502
rect 23548 31490 23604 31500
rect 23548 31332 23604 31342
rect 23548 31106 23604 31276
rect 23548 31054 23550 31106
rect 23602 31054 23604 31106
rect 23548 31042 23604 31054
rect 23660 30996 23716 31500
rect 23996 31554 24052 31836
rect 23996 31502 23998 31554
rect 24050 31502 24052 31554
rect 23996 31332 24052 31502
rect 23996 31266 24052 31276
rect 24556 31554 24612 31566
rect 24556 31502 24558 31554
rect 24610 31502 24612 31554
rect 24556 31444 24612 31502
rect 24108 31106 24164 31118
rect 24108 31054 24110 31106
rect 24162 31054 24164 31106
rect 23772 30996 23828 31006
rect 23660 30940 23772 30996
rect 23772 30930 23828 30940
rect 23772 30322 23828 30334
rect 23772 30270 23774 30322
rect 23826 30270 23828 30322
rect 23772 29988 23828 30270
rect 24108 30212 24164 31054
rect 24444 30996 24500 31006
rect 24444 30902 24500 30940
rect 24108 30146 24164 30156
rect 23772 29922 23828 29932
rect 24556 29988 24612 31388
rect 24668 30548 24724 32620
rect 24668 30482 24724 30492
rect 24780 32002 24836 32014
rect 24780 31950 24782 32002
rect 24834 31950 24836 32002
rect 24556 29922 24612 29932
rect 24780 29764 24836 31950
rect 24892 31890 24948 32620
rect 24892 31838 24894 31890
rect 24946 31838 24948 31890
rect 24892 31826 24948 31838
rect 25004 30884 25060 33628
rect 25228 33460 25284 33470
rect 25564 33460 25620 33966
rect 25228 33458 25620 33460
rect 25228 33406 25230 33458
rect 25282 33406 25620 33458
rect 25228 33404 25620 33406
rect 25788 34020 25844 34076
rect 25228 33394 25284 33404
rect 25116 32788 25172 32798
rect 25116 32694 25172 32732
rect 25788 32788 25844 33964
rect 25788 32722 25844 32732
rect 25900 33346 25956 33358
rect 25900 33294 25902 33346
rect 25954 33294 25956 33346
rect 25340 32674 25396 32686
rect 25340 32622 25342 32674
rect 25394 32622 25396 32674
rect 25340 32004 25396 32622
rect 25452 32564 25508 32574
rect 25452 32470 25508 32508
rect 25900 32004 25956 33294
rect 26012 32452 26068 32462
rect 26012 32358 26068 32396
rect 26012 32004 26068 32014
rect 25900 31948 26012 32004
rect 25340 31938 25396 31948
rect 26012 31938 26068 31948
rect 25676 31890 25732 31902
rect 25676 31838 25678 31890
rect 25730 31838 25732 31890
rect 25676 31780 25732 31838
rect 25676 31714 25732 31724
rect 25900 31780 25956 31790
rect 25228 31668 25284 31678
rect 25228 31666 25396 31668
rect 25228 31614 25230 31666
rect 25282 31614 25396 31666
rect 25228 31612 25396 31614
rect 25228 31602 25284 31612
rect 25228 31332 25284 31342
rect 25228 30994 25284 31276
rect 25228 30942 25230 30994
rect 25282 30942 25284 30994
rect 25228 30930 25284 30942
rect 25004 30828 25172 30884
rect 25116 30772 25172 30828
rect 25116 30716 25284 30772
rect 24444 29708 24836 29764
rect 23436 29026 23492 29036
rect 23548 29426 23604 29438
rect 23548 29374 23550 29426
rect 23602 29374 23604 29426
rect 22988 28478 22990 28530
rect 23042 28478 23044 28530
rect 22988 28466 23044 28478
rect 23100 28924 23380 28980
rect 23100 28532 23156 28924
rect 23100 28466 23156 28476
rect 23212 28756 23268 28766
rect 23548 28756 23604 29374
rect 24444 29426 24500 29708
rect 24444 29374 24446 29426
rect 24498 29374 24500 29426
rect 23268 28700 23604 28756
rect 24108 29314 24164 29326
rect 24108 29262 24110 29314
rect 24162 29262 24164 29314
rect 24108 28756 24164 29262
rect 24444 29204 24500 29374
rect 24444 29138 24500 29148
rect 24556 29538 24612 29550
rect 24556 29486 24558 29538
rect 24610 29486 24612 29538
rect 23212 28530 23268 28700
rect 24108 28690 24164 28700
rect 23996 28644 24052 28654
rect 23996 28550 24052 28588
rect 23212 28478 23214 28530
rect 23266 28478 23268 28530
rect 23212 28466 23268 28478
rect 23436 28532 23492 28542
rect 23436 28438 23492 28476
rect 24556 28308 24612 29486
rect 24780 29428 24836 29438
rect 24780 29334 24836 29372
rect 24668 29316 24724 29326
rect 24668 28754 24724 29260
rect 24668 28702 24670 28754
rect 24722 28702 24724 28754
rect 24668 28690 24724 28702
rect 24556 28252 25060 28308
rect 23324 28084 23380 28094
rect 23324 27990 23380 28028
rect 24668 28084 24724 28094
rect 24668 27990 24724 28028
rect 23548 27972 23604 27982
rect 24108 27972 24164 27982
rect 22988 27860 23044 27870
rect 22988 27766 23044 27804
rect 23548 27858 23604 27916
rect 23548 27806 23550 27858
rect 23602 27806 23604 27858
rect 23548 27794 23604 27806
rect 23660 27970 24164 27972
rect 23660 27918 24110 27970
rect 24162 27918 24164 27970
rect 23660 27916 24164 27918
rect 23212 27636 23268 27646
rect 23212 27542 23268 27580
rect 23324 27412 23380 27422
rect 23324 27074 23380 27356
rect 23436 27300 23492 27310
rect 23436 27188 23492 27244
rect 23436 27132 23548 27188
rect 23324 27022 23326 27074
rect 23378 27022 23380 27074
rect 23324 27010 23380 27022
rect 23492 27086 23548 27132
rect 23492 27076 23604 27086
rect 23492 27020 23548 27076
rect 23548 27010 23604 27020
rect 23660 26908 23716 27916
rect 24108 27906 24164 27916
rect 24220 27858 24276 27870
rect 24220 27806 24222 27858
rect 24274 27806 24276 27858
rect 24108 27634 24164 27646
rect 24108 27582 24110 27634
rect 24162 27582 24164 27634
rect 23996 27300 24052 27310
rect 23996 27074 24052 27244
rect 24108 27188 24164 27582
rect 24220 27300 24276 27806
rect 24220 27234 24276 27244
rect 24108 27122 24164 27132
rect 24668 27186 24724 27198
rect 24668 27134 24670 27186
rect 24722 27134 24724 27186
rect 23996 27022 23998 27074
rect 24050 27022 24052 27074
rect 23996 27010 24052 27022
rect 24220 27076 24276 27086
rect 24220 26982 24276 27020
rect 23324 26852 23716 26908
rect 24108 26964 24164 26974
rect 23324 26404 23380 26852
rect 23492 26796 23604 26852
rect 23772 26850 23828 26862
rect 23772 26798 23774 26850
rect 23826 26798 23828 26850
rect 23324 26338 23380 26348
rect 23436 26516 23492 26526
rect 23436 26290 23492 26460
rect 23660 26516 23716 26526
rect 23660 26402 23716 26460
rect 23660 26350 23662 26402
rect 23714 26350 23716 26402
rect 23660 26338 23716 26350
rect 23436 26238 23438 26290
rect 23490 26238 23492 26290
rect 23100 26178 23156 26190
rect 23100 26126 23102 26178
rect 23154 26126 23156 26178
rect 23100 25844 23156 26126
rect 23100 25778 23156 25788
rect 23436 25620 23492 26238
rect 23772 26180 23828 26798
rect 23884 26852 23940 26862
rect 23884 26758 23940 26796
rect 24108 26628 24164 26908
rect 23996 26572 24164 26628
rect 24556 26964 24612 26974
rect 23996 26402 24052 26572
rect 23996 26350 23998 26402
rect 24050 26350 24052 26402
rect 23996 26338 24052 26350
rect 24444 26402 24500 26414
rect 24444 26350 24446 26402
rect 24498 26350 24500 26402
rect 24220 26292 24276 26302
rect 24220 26198 24276 26236
rect 23884 26180 23940 26190
rect 23772 26178 24052 26180
rect 23772 26126 23886 26178
rect 23938 26126 24052 26178
rect 23772 26124 24052 26126
rect 23884 26114 23940 26124
rect 22652 24500 22708 24510
rect 22652 23938 22708 24444
rect 22652 23886 22654 23938
rect 22706 23886 22708 23938
rect 22652 23874 22708 23886
rect 22652 23268 22708 23278
rect 22652 23174 22708 23212
rect 22540 23090 22596 23100
rect 22764 22372 22820 25116
rect 23100 25564 23492 25620
rect 22988 24052 23044 24062
rect 23100 24052 23156 25564
rect 23772 24946 23828 24958
rect 23772 24894 23774 24946
rect 23826 24894 23828 24946
rect 23212 24724 23268 24734
rect 23212 24722 23380 24724
rect 23212 24670 23214 24722
rect 23266 24670 23380 24722
rect 23212 24668 23380 24670
rect 23212 24658 23268 24668
rect 23212 24052 23268 24062
rect 23100 24050 23268 24052
rect 23100 23998 23214 24050
rect 23266 23998 23268 24050
rect 23100 23996 23268 23998
rect 22988 23938 23044 23996
rect 23212 23986 23268 23996
rect 22988 23886 22990 23938
rect 23042 23886 23044 23938
rect 22988 23874 23044 23886
rect 22988 23380 23044 23390
rect 22764 22306 22820 22316
rect 22876 23044 22932 23054
rect 22876 21810 22932 22988
rect 22876 21758 22878 21810
rect 22930 21758 22932 21810
rect 22876 21746 22932 21758
rect 22988 21812 23044 23324
rect 23100 23042 23156 23054
rect 23100 22990 23102 23042
rect 23154 22990 23156 23042
rect 23100 22930 23156 22990
rect 23100 22878 23102 22930
rect 23154 22878 23156 22930
rect 23100 22866 23156 22878
rect 23212 22708 23268 22718
rect 23100 21812 23156 21822
rect 22988 21756 23100 21812
rect 23100 21718 23156 21756
rect 22428 21532 22596 21588
rect 22316 21476 22372 21486
rect 22372 21420 22484 21476
rect 22316 21382 22372 21420
rect 22428 20802 22484 21420
rect 22540 20916 22596 21532
rect 22540 20850 22596 20860
rect 22988 21474 23044 21486
rect 22988 21422 22990 21474
rect 23042 21422 23044 21474
rect 22428 20750 22430 20802
rect 22482 20750 22484 20802
rect 22428 20738 22484 20750
rect 22988 20692 23044 21422
rect 23100 20916 23156 20926
rect 23212 20916 23268 22652
rect 23324 22482 23380 24668
rect 23548 24722 23604 24734
rect 23548 24670 23550 24722
rect 23602 24670 23604 24722
rect 23548 24162 23604 24670
rect 23548 24110 23550 24162
rect 23602 24110 23604 24162
rect 23548 24098 23604 24110
rect 23660 24052 23716 24062
rect 23660 23958 23716 23996
rect 23548 23156 23604 23166
rect 23548 23062 23604 23100
rect 23772 23044 23828 24894
rect 23884 24836 23940 24846
rect 23884 24500 23940 24780
rect 23996 24722 24052 26124
rect 24444 25844 24500 26350
rect 24556 26402 24612 26908
rect 24556 26350 24558 26402
rect 24610 26350 24612 26402
rect 24556 26338 24612 26350
rect 24332 25620 24388 25630
rect 24332 24946 24388 25564
rect 24332 24894 24334 24946
rect 24386 24894 24388 24946
rect 24332 24882 24388 24894
rect 24444 24948 24500 25788
rect 24556 24948 24612 24958
rect 24444 24892 24556 24948
rect 24556 24854 24612 24892
rect 24668 24834 24724 27134
rect 24780 26850 24836 26862
rect 24780 26798 24782 26850
rect 24834 26798 24836 26850
rect 24780 26516 24836 26798
rect 24780 26450 24836 26460
rect 24668 24782 24670 24834
rect 24722 24782 24724 24834
rect 24668 24770 24724 24782
rect 23996 24670 23998 24722
rect 24050 24670 24052 24722
rect 23996 24658 24052 24670
rect 23884 24434 23940 24444
rect 24892 23938 24948 23950
rect 24892 23886 24894 23938
rect 24946 23886 24948 23938
rect 24332 23826 24388 23838
rect 24332 23774 24334 23826
rect 24386 23774 24388 23826
rect 24108 23044 24164 23054
rect 23772 22978 23828 22988
rect 23996 23042 24164 23044
rect 23996 22990 24110 23042
rect 24162 22990 24164 23042
rect 23996 22988 24164 22990
rect 23324 22430 23326 22482
rect 23378 22430 23380 22482
rect 23324 21700 23380 22430
rect 23324 21634 23380 21644
rect 23436 22484 23492 22494
rect 23436 21026 23492 22428
rect 23772 21700 23828 21710
rect 23660 21698 23828 21700
rect 23660 21646 23774 21698
rect 23826 21646 23828 21698
rect 23660 21644 23828 21646
rect 23548 21588 23604 21598
rect 23548 21494 23604 21532
rect 23436 20974 23438 21026
rect 23490 20974 23492 21026
rect 23436 20962 23492 20974
rect 23100 20914 23268 20916
rect 23100 20862 23102 20914
rect 23154 20862 23268 20914
rect 23100 20860 23268 20862
rect 23324 20916 23380 20926
rect 23100 20850 23156 20860
rect 22540 20636 23044 20692
rect 22540 20130 22596 20636
rect 22540 20078 22542 20130
rect 22594 20078 22596 20130
rect 22540 20066 22596 20078
rect 22316 19516 22820 19572
rect 22316 19458 22372 19516
rect 22316 19406 22318 19458
rect 22370 19406 22372 19458
rect 22316 19394 22372 19406
rect 22764 19234 22820 19516
rect 23324 19460 23380 20860
rect 22764 19182 22766 19234
rect 22818 19182 22820 19234
rect 22764 19170 22820 19182
rect 23212 19404 23380 19460
rect 22204 19124 22260 19134
rect 22428 19124 22484 19134
rect 22260 19068 22372 19124
rect 22204 19058 22260 19068
rect 22092 19012 22148 19022
rect 22092 17778 22148 18956
rect 22316 19010 22372 19068
rect 22428 19030 22484 19068
rect 22316 18958 22318 19010
rect 22370 18958 22372 19010
rect 22316 18946 22372 18958
rect 22876 19012 22932 19022
rect 22876 18918 22932 18956
rect 22988 19010 23044 19022
rect 22988 18958 22990 19010
rect 23042 18958 23044 19010
rect 22988 18788 23044 18958
rect 22428 18732 23044 18788
rect 22428 18674 22484 18732
rect 22428 18622 22430 18674
rect 22482 18622 22484 18674
rect 22428 18610 22484 18622
rect 22540 18564 22596 18574
rect 22204 18450 22260 18462
rect 22204 18398 22206 18450
rect 22258 18398 22260 18450
rect 22204 18116 22260 18398
rect 22540 18450 22596 18508
rect 23100 18564 23156 18574
rect 22540 18398 22542 18450
rect 22594 18398 22596 18450
rect 22540 18386 22596 18398
rect 22764 18450 22820 18462
rect 22764 18398 22766 18450
rect 22818 18398 22820 18450
rect 22764 18340 22820 18398
rect 22764 18274 22820 18284
rect 22204 18050 22260 18060
rect 22092 17726 22094 17778
rect 22146 17726 22148 17778
rect 22092 17714 22148 17726
rect 22204 16772 22260 16782
rect 22204 15092 22260 16716
rect 22652 16212 22708 16222
rect 22876 16212 22932 16222
rect 22708 16210 22932 16212
rect 22708 16158 22878 16210
rect 22930 16158 22932 16210
rect 22708 16156 22932 16158
rect 22652 16146 22708 16156
rect 22652 15652 22708 15662
rect 22316 15428 22372 15438
rect 22652 15428 22708 15596
rect 22316 15426 22708 15428
rect 22316 15374 22318 15426
rect 22370 15374 22654 15426
rect 22706 15374 22708 15426
rect 22316 15372 22708 15374
rect 22316 15362 22372 15372
rect 22652 15362 22708 15372
rect 22764 15426 22820 15438
rect 22764 15374 22766 15426
rect 22818 15374 22820 15426
rect 22316 15092 22372 15102
rect 22204 15090 22372 15092
rect 22204 15038 22318 15090
rect 22370 15038 22372 15090
rect 22204 15036 22372 15038
rect 21868 14642 22260 14644
rect 21868 14590 21870 14642
rect 21922 14590 22260 14642
rect 21868 14588 22260 14590
rect 21868 14578 21924 14588
rect 21420 14420 21476 14430
rect 21420 14418 21588 14420
rect 21420 14366 21422 14418
rect 21474 14366 21588 14418
rect 21420 14364 21588 14366
rect 21420 14354 21476 14364
rect 21308 14308 21364 14318
rect 21308 14214 21364 14252
rect 21420 13636 21476 13646
rect 21420 13542 21476 13580
rect 21532 13188 21588 14364
rect 21532 13122 21588 13132
rect 21868 13746 21924 13758
rect 21868 13694 21870 13746
rect 21922 13694 21924 13746
rect 21756 12964 21812 12974
rect 19404 12114 19460 12124
rect 19516 12292 19572 12302
rect 19516 11394 19572 12236
rect 20300 12180 20356 12190
rect 19740 11620 19796 11630
rect 19516 11342 19518 11394
rect 19570 11342 19572 11394
rect 19516 11330 19572 11342
rect 19628 11618 19796 11620
rect 19628 11566 19742 11618
rect 19794 11566 19796 11618
rect 19628 11564 19796 11566
rect 19628 9156 19684 11564
rect 19740 11554 19796 11564
rect 19852 11506 19908 11518
rect 19852 11454 19854 11506
rect 19906 11454 19908 11506
rect 19852 11172 19908 11454
rect 20300 11396 20356 12124
rect 20748 12180 20804 12190
rect 20860 12180 20916 12348
rect 21644 12908 21756 12964
rect 20972 12292 21028 12302
rect 20972 12290 21140 12292
rect 20972 12238 20974 12290
rect 21026 12238 21140 12290
rect 20972 12236 21140 12238
rect 20972 12226 21028 12236
rect 20748 12178 20916 12180
rect 20748 12126 20750 12178
rect 20802 12126 20916 12178
rect 20748 12124 20916 12126
rect 20748 12114 20804 12124
rect 20972 11844 21028 11854
rect 20300 11330 20356 11340
rect 20524 11394 20580 11406
rect 20524 11342 20526 11394
rect 20578 11342 20580 11394
rect 19852 11106 19908 11116
rect 19836 11004 20100 11014
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 19836 10938 20100 10948
rect 19836 9436 20100 9446
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 19836 9370 20100 9380
rect 19628 9090 19684 9100
rect 20524 8932 20580 11342
rect 20748 11284 20804 11294
rect 20972 11284 21028 11788
rect 21084 11620 21140 12236
rect 21532 12180 21588 12190
rect 21308 12178 21588 12180
rect 21308 12126 21534 12178
rect 21586 12126 21588 12178
rect 21308 12124 21588 12126
rect 21196 11620 21252 11630
rect 21084 11618 21252 11620
rect 21084 11566 21198 11618
rect 21250 11566 21252 11618
rect 21084 11564 21252 11566
rect 21196 11554 21252 11564
rect 20748 11282 21028 11284
rect 20748 11230 20750 11282
rect 20802 11230 21028 11282
rect 20748 11228 21028 11230
rect 20748 11218 20804 11228
rect 20972 10498 21028 11228
rect 20972 10446 20974 10498
rect 21026 10446 21028 10498
rect 20972 10434 21028 10446
rect 20524 8866 20580 8876
rect 19836 7868 20100 7878
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 19836 7802 20100 7812
rect 19836 6300 20100 6310
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 19836 6234 20100 6244
rect 19836 4732 20100 4742
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 19836 4666 20100 4676
rect 18844 3390 18846 3442
rect 18898 3390 18900 3442
rect 18844 3378 18900 3390
rect 19068 4226 19124 4238
rect 19068 4174 19070 4226
rect 19122 4174 19124 4226
rect 19068 2548 19124 4174
rect 19740 4226 19796 4238
rect 19740 4174 19742 4226
rect 19794 4174 19796 4226
rect 19180 3444 19236 3454
rect 19180 3350 19236 3388
rect 19516 3444 19572 3454
rect 19740 3444 19796 4174
rect 20860 4226 20916 4238
rect 20860 4174 20862 4226
rect 20914 4174 20916 4226
rect 19516 3442 19796 3444
rect 19516 3390 19518 3442
rect 19570 3390 19796 3442
rect 19516 3388 19796 3390
rect 19852 3444 19908 3454
rect 18620 2492 19124 2548
rect 16828 800 16884 2492
rect 18172 800 18228 2492
rect 18844 800 18900 2492
rect 19516 800 19572 3388
rect 19852 3350 19908 3388
rect 20188 3444 20244 3454
rect 19836 3164 20100 3174
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 19836 3098 20100 3108
rect 20188 800 20244 3388
rect 20860 3444 20916 4174
rect 21084 3444 21140 3454
rect 20860 3442 21140 3444
rect 20860 3390 21086 3442
rect 21138 3390 21140 3442
rect 20860 3388 21140 3390
rect 21308 3444 21364 12124
rect 21532 12114 21588 12124
rect 21644 12180 21700 12908
rect 21756 12898 21812 12908
rect 21868 12180 21924 13694
rect 22092 13188 22148 13198
rect 21420 11618 21476 11630
rect 21420 11566 21422 11618
rect 21474 11566 21476 11618
rect 21420 10610 21476 11566
rect 21532 11508 21588 11518
rect 21644 11508 21700 12124
rect 21756 12124 21924 12180
rect 21980 12178 22036 12190
rect 21980 12126 21982 12178
rect 22034 12126 22036 12178
rect 21756 11788 21812 12124
rect 21980 11844 22036 12126
rect 22092 11954 22148 13132
rect 22204 12068 22260 14588
rect 22316 14306 22372 15036
rect 22316 14254 22318 14306
rect 22370 14254 22372 14306
rect 22316 12852 22372 14254
rect 22540 14308 22596 14318
rect 22540 13858 22596 14252
rect 22540 13806 22542 13858
rect 22594 13806 22596 13858
rect 22540 13794 22596 13806
rect 22652 14308 22708 14318
rect 22764 14308 22820 15374
rect 22652 14306 22820 14308
rect 22652 14254 22654 14306
rect 22706 14254 22820 14306
rect 22652 14252 22820 14254
rect 22652 13636 22708 14252
rect 22652 13570 22708 13580
rect 22316 12786 22372 12796
rect 22540 13076 22596 13086
rect 22540 12178 22596 13020
rect 22540 12126 22542 12178
rect 22594 12126 22596 12178
rect 22540 12114 22596 12126
rect 22204 12066 22484 12068
rect 22204 12014 22206 12066
rect 22258 12014 22484 12066
rect 22204 12012 22484 12014
rect 22204 12002 22260 12012
rect 22092 11902 22094 11954
rect 22146 11902 22148 11954
rect 22092 11890 22148 11902
rect 21756 11732 21924 11788
rect 21980 11778 22036 11788
rect 21532 11506 21700 11508
rect 21532 11454 21534 11506
rect 21586 11454 21700 11506
rect 21532 11452 21700 11454
rect 21532 11442 21588 11452
rect 21420 10558 21422 10610
rect 21474 10558 21476 10610
rect 21420 9604 21476 10558
rect 21868 11284 21924 11732
rect 22428 11284 22484 12012
rect 22652 11508 22708 11518
rect 22876 11508 22932 16156
rect 22988 15540 23044 15550
rect 22988 15446 23044 15484
rect 23100 14642 23156 18508
rect 23212 18228 23268 19404
rect 23660 19348 23716 21644
rect 23772 21634 23828 21644
rect 23996 21252 24052 22988
rect 24108 22978 24164 22988
rect 24332 22484 24388 23774
rect 24444 23828 24500 23838
rect 24444 23734 24500 23772
rect 24556 23268 24612 23278
rect 24556 23154 24612 23212
rect 24556 23102 24558 23154
rect 24610 23102 24612 23154
rect 24556 22596 24612 23102
rect 24556 22530 24612 22540
rect 24332 22418 24388 22428
rect 24892 21924 24948 23886
rect 24892 21858 24948 21868
rect 25004 22932 25060 28252
rect 25228 28084 25284 30716
rect 25340 30660 25396 31612
rect 25452 31556 25508 31566
rect 25452 31462 25508 31500
rect 25676 31556 25732 31566
rect 25676 31462 25732 31500
rect 25788 31554 25844 31566
rect 25788 31502 25790 31554
rect 25842 31502 25844 31554
rect 25788 31332 25844 31502
rect 25340 30594 25396 30604
rect 25452 31276 25788 31332
rect 25452 29650 25508 31276
rect 25788 31238 25844 31276
rect 25788 30436 25844 30446
rect 25452 29598 25454 29650
rect 25506 29598 25508 29650
rect 25452 29586 25508 29598
rect 25564 30380 25788 30436
rect 25564 29650 25620 30380
rect 25788 30370 25844 30380
rect 25900 30322 25956 31724
rect 26124 30884 26180 34860
rect 26236 34914 26292 35868
rect 26460 35922 26516 35980
rect 26460 35870 26462 35922
rect 26514 35870 26516 35922
rect 26460 35858 26516 35870
rect 26572 35476 26628 41244
rect 27020 41076 27076 41086
rect 26908 41020 27020 41076
rect 26908 40626 26964 41020
rect 27020 40982 27076 41020
rect 26908 40574 26910 40626
rect 26962 40574 26964 40626
rect 26908 40404 26964 40574
rect 26236 34862 26238 34914
rect 26290 34862 26292 34914
rect 26236 34850 26292 34862
rect 26460 35420 26628 35476
rect 26684 40348 26964 40404
rect 27244 40404 27300 40414
rect 26236 34244 26292 34254
rect 26236 34242 26404 34244
rect 26236 34190 26238 34242
rect 26290 34190 26404 34242
rect 26236 34188 26404 34190
rect 26236 34178 26292 34188
rect 26236 32676 26292 32686
rect 26236 32582 26292 32620
rect 26348 32564 26404 34188
rect 26460 33796 26516 35420
rect 26572 35252 26628 35262
rect 26572 34354 26628 35196
rect 26572 34302 26574 34354
rect 26626 34302 26628 34354
rect 26572 34290 26628 34302
rect 26460 33730 26516 33740
rect 26684 33348 26740 40348
rect 27244 40310 27300 40348
rect 26796 39620 26852 39630
rect 26796 39526 26852 39564
rect 27244 38722 27300 38734
rect 27244 38670 27246 38722
rect 27298 38670 27300 38722
rect 27132 38162 27188 38174
rect 27132 38110 27134 38162
rect 27186 38110 27188 38162
rect 26908 37828 26964 37838
rect 26908 35924 26964 37772
rect 27132 37492 27188 38110
rect 27132 37426 27188 37436
rect 27244 37716 27300 38670
rect 27020 37380 27076 37390
rect 27020 37154 27076 37324
rect 27020 37102 27022 37154
rect 27074 37102 27076 37154
rect 27020 37090 27076 37102
rect 27244 36708 27300 37660
rect 27132 36652 27300 36708
rect 26908 35830 26964 35868
rect 27020 36036 27076 36046
rect 26908 34916 26964 34926
rect 26908 34822 26964 34860
rect 27020 34914 27076 35980
rect 27020 34862 27022 34914
rect 27074 34862 27076 34914
rect 27020 34850 27076 34862
rect 27132 34468 27188 36652
rect 27244 36484 27300 36494
rect 27244 36370 27300 36428
rect 27244 36318 27246 36370
rect 27298 36318 27300 36370
rect 27244 36306 27300 36318
rect 27356 36260 27412 44044
rect 27580 43540 27636 43550
rect 27580 42754 27636 43484
rect 27916 42868 27972 42878
rect 27916 42774 27972 42812
rect 27580 42702 27582 42754
rect 27634 42702 27636 42754
rect 27580 42308 27636 42702
rect 27580 42242 27636 42252
rect 28252 42532 28308 42542
rect 27692 41972 27748 41982
rect 27692 41878 27748 41916
rect 27468 41300 27524 41310
rect 27468 41206 27524 41244
rect 28028 41300 28084 41310
rect 28028 41206 28084 41244
rect 27580 41188 27636 41198
rect 27468 39396 27524 39406
rect 27468 39302 27524 39340
rect 27468 38724 27524 38762
rect 27468 38658 27524 38668
rect 27580 38274 27636 41132
rect 27580 38222 27582 38274
rect 27634 38222 27636 38274
rect 27580 38210 27636 38222
rect 27916 38164 27972 38174
rect 27916 38070 27972 38108
rect 28252 38052 28308 42476
rect 28364 38668 28420 44044
rect 28476 44034 28532 44044
rect 28700 45108 28756 45118
rect 28476 43428 28532 43438
rect 28700 43428 28756 45052
rect 28476 43426 28756 43428
rect 28476 43374 28478 43426
rect 28530 43374 28756 43426
rect 28476 43372 28756 43374
rect 28476 42084 28532 43372
rect 28476 42018 28532 42028
rect 28700 41412 28756 41422
rect 28700 41298 28756 41356
rect 28700 41246 28702 41298
rect 28754 41246 28756 41298
rect 28700 38724 28756 41246
rect 28364 38612 28532 38668
rect 28700 38658 28756 38668
rect 28476 38276 28532 38612
rect 28476 38220 28644 38276
rect 28476 38052 28532 38062
rect 28252 38050 28532 38052
rect 28252 37998 28478 38050
rect 28530 37998 28532 38050
rect 28252 37996 28532 37998
rect 28476 37986 28532 37996
rect 27804 37828 27860 37838
rect 27692 37826 27860 37828
rect 27692 37774 27806 37826
rect 27858 37774 27860 37826
rect 27692 37772 27860 37774
rect 27468 37492 27524 37502
rect 27468 37044 27524 37436
rect 27468 36978 27524 36988
rect 27468 36596 27524 36606
rect 27468 36502 27524 36540
rect 27356 36204 27524 36260
rect 27356 36036 27412 36046
rect 27356 35922 27412 35980
rect 27356 35870 27358 35922
rect 27410 35870 27412 35922
rect 27356 35858 27412 35870
rect 27356 35140 27412 35150
rect 27244 34692 27300 34702
rect 27244 34598 27300 34636
rect 27132 34412 27300 34468
rect 26908 34132 26964 34142
rect 26908 34038 26964 34076
rect 27020 34018 27076 34030
rect 27020 33966 27022 34018
rect 27074 33966 27076 34018
rect 27020 33348 27076 33966
rect 26348 32498 26404 32508
rect 26460 33292 26740 33348
rect 26796 33292 27076 33348
rect 26460 32676 26516 33292
rect 26572 33124 26628 33134
rect 26796 33124 26852 33292
rect 27132 33236 27188 33246
rect 27132 33142 27188 33180
rect 26628 33068 26852 33124
rect 26908 33124 26964 33134
rect 26572 33030 26628 33068
rect 26572 32676 26628 32686
rect 26460 32674 26628 32676
rect 26460 32622 26574 32674
rect 26626 32622 26628 32674
rect 26460 32620 26628 32622
rect 26348 31666 26404 31678
rect 26348 31614 26350 31666
rect 26402 31614 26404 31666
rect 26236 31556 26292 31566
rect 26236 31462 26292 31500
rect 26348 31444 26404 31614
rect 26348 31378 26404 31388
rect 26348 30884 26404 30894
rect 26124 30828 26348 30884
rect 26348 30818 26404 30828
rect 26460 30660 26516 32620
rect 26572 32610 26628 32620
rect 26908 32450 26964 33068
rect 26908 32398 26910 32450
rect 26962 32398 26964 32450
rect 26908 32386 26964 32398
rect 27020 32452 27076 32462
rect 27244 32452 27300 34412
rect 27076 32396 27300 32452
rect 26684 32004 26740 32014
rect 25900 30270 25902 30322
rect 25954 30270 25956 30322
rect 25900 30258 25956 30270
rect 26124 30604 26516 30660
rect 26572 30884 26628 30894
rect 25564 29598 25566 29650
rect 25618 29598 25620 29650
rect 25564 29586 25620 29598
rect 25900 29540 25956 29550
rect 25788 29428 25844 29438
rect 25788 29334 25844 29372
rect 25900 29426 25956 29484
rect 25900 29374 25902 29426
rect 25954 29374 25956 29426
rect 25900 29362 25956 29374
rect 25676 29316 25732 29326
rect 25676 29222 25732 29260
rect 25452 28532 25508 28542
rect 25340 28084 25396 28094
rect 25284 28082 25396 28084
rect 25284 28030 25342 28082
rect 25394 28030 25396 28082
rect 25284 28028 25396 28030
rect 25228 27990 25284 28028
rect 25340 28018 25396 28028
rect 25228 27858 25284 27870
rect 25228 27806 25230 27858
rect 25282 27806 25284 27858
rect 25228 27524 25284 27806
rect 25116 27300 25172 27310
rect 25116 27074 25172 27244
rect 25116 27022 25118 27074
rect 25170 27022 25172 27074
rect 25116 27010 25172 27022
rect 25116 26516 25172 26526
rect 25116 26422 25172 26460
rect 25228 26514 25284 27468
rect 25452 27188 25508 28476
rect 25900 28084 25956 28094
rect 25564 27860 25620 27870
rect 25564 27766 25620 27804
rect 25900 27858 25956 28028
rect 25900 27806 25902 27858
rect 25954 27806 25956 27858
rect 25900 27794 25956 27806
rect 25452 26962 25508 27132
rect 25900 27300 25956 27310
rect 25900 27186 25956 27244
rect 25900 27134 25902 27186
rect 25954 27134 25956 27186
rect 25900 27122 25956 27134
rect 25452 26910 25454 26962
rect 25506 26910 25508 26962
rect 25452 26898 25508 26910
rect 25228 26462 25230 26514
rect 25282 26462 25284 26514
rect 25228 26450 25284 26462
rect 26012 26516 26068 26526
rect 26012 26422 26068 26460
rect 25452 26404 25508 26414
rect 25452 26310 25508 26348
rect 25788 26404 25844 26414
rect 25788 26290 25844 26348
rect 25788 26238 25790 26290
rect 25842 26238 25844 26290
rect 25788 26226 25844 26238
rect 25452 25060 25508 25070
rect 25340 24834 25396 24846
rect 25340 24782 25342 24834
rect 25394 24782 25396 24834
rect 25116 24722 25172 24734
rect 25116 24670 25118 24722
rect 25170 24670 25172 24722
rect 25116 24052 25172 24670
rect 25116 23986 25172 23996
rect 25340 23156 25396 24782
rect 25452 24834 25508 25004
rect 25452 24782 25454 24834
rect 25506 24782 25508 24834
rect 25452 24770 25508 24782
rect 25788 24834 25844 24846
rect 25788 24782 25790 24834
rect 25842 24782 25844 24834
rect 25564 23828 25620 23838
rect 25564 23734 25620 23772
rect 25340 23062 25396 23100
rect 25676 23154 25732 23166
rect 25676 23102 25678 23154
rect 25730 23102 25732 23154
rect 25676 22932 25732 23102
rect 25004 22876 25732 22932
rect 24444 21700 24500 21710
rect 24108 21586 24164 21598
rect 24108 21534 24110 21586
rect 24162 21534 24164 21586
rect 24108 21476 24164 21534
rect 24332 21588 24388 21598
rect 24332 21494 24388 21532
rect 24108 21410 24164 21420
rect 23436 19292 23716 19348
rect 23772 20802 23828 20814
rect 23772 20750 23774 20802
rect 23826 20750 23828 20802
rect 23772 19348 23828 20750
rect 23996 20802 24052 21196
rect 24332 20916 24388 20926
rect 24444 20916 24500 21644
rect 24332 20914 24500 20916
rect 24332 20862 24334 20914
rect 24386 20862 24500 20914
rect 24332 20860 24500 20862
rect 24556 21698 24612 21710
rect 24556 21646 24558 21698
rect 24610 21646 24612 21698
rect 24332 20850 24388 20860
rect 23996 20750 23998 20802
rect 24050 20750 24052 20802
rect 23996 20738 24052 20750
rect 24556 20244 24612 21646
rect 25004 21700 25060 22876
rect 25788 22596 25844 24782
rect 26124 24722 26180 30604
rect 26572 30210 26628 30828
rect 26572 30158 26574 30210
rect 26626 30158 26628 30210
rect 26572 28644 26628 30158
rect 26684 29426 26740 31948
rect 27020 31780 27076 32396
rect 27132 31780 27188 31790
rect 27020 31778 27188 31780
rect 27020 31726 27134 31778
rect 27186 31726 27188 31778
rect 27020 31724 27188 31726
rect 26908 31668 26964 31678
rect 26796 31554 26852 31566
rect 26796 31502 26798 31554
rect 26850 31502 26852 31554
rect 26796 30436 26852 31502
rect 26796 30370 26852 30380
rect 26684 29374 26686 29426
rect 26738 29374 26740 29426
rect 26684 29362 26740 29374
rect 26572 28578 26628 28588
rect 26684 29204 26740 29214
rect 26124 24670 26126 24722
rect 26178 24670 26180 24722
rect 26124 24052 26180 24670
rect 26124 23986 26180 23996
rect 26236 28420 26292 28430
rect 26236 27746 26292 28364
rect 26236 27694 26238 27746
rect 26290 27694 26292 27746
rect 26236 23380 26292 27694
rect 26348 27300 26404 27310
rect 26348 27186 26404 27244
rect 26348 27134 26350 27186
rect 26402 27134 26404 27186
rect 26348 26964 26404 27134
rect 26348 26898 26404 26908
rect 26348 26402 26404 26414
rect 26348 26350 26350 26402
rect 26402 26350 26404 26402
rect 26348 25956 26404 26350
rect 26572 26068 26628 26078
rect 26404 25900 26516 25956
rect 26348 25890 26404 25900
rect 26460 23492 26516 25900
rect 26572 25506 26628 26012
rect 26572 25454 26574 25506
rect 26626 25454 26628 25506
rect 26572 25442 26628 25454
rect 26572 25060 26628 25070
rect 26572 24722 26628 25004
rect 26572 24670 26574 24722
rect 26626 24670 26628 24722
rect 26572 24658 26628 24670
rect 25564 22540 25844 22596
rect 25900 23324 26292 23380
rect 26348 23380 26404 23390
rect 25228 22372 25284 22382
rect 25228 22278 25284 22316
rect 25564 21924 25620 22540
rect 25340 21868 25620 21924
rect 25676 22372 25732 22382
rect 25340 21812 25396 21868
rect 25004 21634 25060 21644
rect 25228 21810 25396 21812
rect 25228 21758 25342 21810
rect 25394 21758 25396 21810
rect 25228 21756 25396 21758
rect 24556 20178 24612 20188
rect 24668 21586 24724 21598
rect 24668 21534 24670 21586
rect 24722 21534 24724 21586
rect 24668 19908 24724 21534
rect 25116 21586 25172 21598
rect 25116 21534 25118 21586
rect 25170 21534 25172 21586
rect 24444 19906 24724 19908
rect 24444 19854 24670 19906
rect 24722 19854 24724 19906
rect 24444 19852 24724 19854
rect 23772 19292 24276 19348
rect 23324 19234 23380 19246
rect 23324 19182 23326 19234
rect 23378 19182 23380 19234
rect 23324 18452 23380 19182
rect 23436 18900 23492 19292
rect 23548 19124 23604 19134
rect 23548 19030 23604 19068
rect 24108 19122 24164 19134
rect 24108 19070 24110 19122
rect 24162 19070 24164 19122
rect 23660 19012 23716 19022
rect 23660 19010 23828 19012
rect 23660 18958 23662 19010
rect 23714 18958 23828 19010
rect 23660 18956 23828 18958
rect 23660 18946 23716 18956
rect 23436 18844 23604 18900
rect 23324 18386 23380 18396
rect 23212 18172 23380 18228
rect 23212 18004 23268 18014
rect 23212 17106 23268 17948
rect 23212 17054 23214 17106
rect 23266 17054 23268 17106
rect 23212 17042 23268 17054
rect 23324 15316 23380 18172
rect 23548 17444 23604 18844
rect 23660 18788 23716 18798
rect 23660 18450 23716 18732
rect 23772 18564 23828 18956
rect 23772 18498 23828 18508
rect 23884 19010 23940 19022
rect 23884 18958 23886 19010
rect 23938 18958 23940 19010
rect 23660 18398 23662 18450
rect 23714 18398 23716 18450
rect 23660 18386 23716 18398
rect 23884 17780 23940 18958
rect 23996 18450 24052 18462
rect 23996 18398 23998 18450
rect 24050 18398 24052 18450
rect 23996 18004 24052 18398
rect 24108 18340 24164 19070
rect 24108 18246 24164 18284
rect 24220 18228 24276 19292
rect 24332 18452 24388 18462
rect 24332 18358 24388 18396
rect 24220 18162 24276 18172
rect 24444 18004 24500 19852
rect 24668 19842 24724 19852
rect 24780 20020 24836 20030
rect 24780 19346 24836 19964
rect 24780 19294 24782 19346
rect 24834 19294 24836 19346
rect 24780 19236 24836 19294
rect 24780 19170 24836 19180
rect 25116 19234 25172 21534
rect 25116 19182 25118 19234
rect 25170 19182 25172 19234
rect 25116 19170 25172 19182
rect 24668 18788 24724 18798
rect 24556 18676 24612 18686
rect 24556 18582 24612 18620
rect 24668 18564 24724 18732
rect 25228 18676 25284 21756
rect 25340 21746 25396 21756
rect 25452 21700 25508 21710
rect 25452 21606 25508 21644
rect 25564 21476 25620 21486
rect 25452 21420 25564 21476
rect 25340 20244 25396 20254
rect 25340 20130 25396 20188
rect 25340 20078 25342 20130
rect 25394 20078 25396 20130
rect 25340 20066 25396 20078
rect 25452 19348 25508 21420
rect 25564 21410 25620 21420
rect 25676 20020 25732 22316
rect 25676 19926 25732 19964
rect 25900 19908 25956 23324
rect 26012 23154 26068 23166
rect 26012 23102 26014 23154
rect 26066 23102 26068 23154
rect 26012 22708 26068 23102
rect 26348 23154 26404 23324
rect 26348 23102 26350 23154
rect 26402 23102 26404 23154
rect 26348 23090 26404 23102
rect 26124 23044 26180 23054
rect 26124 22950 26180 22988
rect 26012 22652 26292 22708
rect 26012 21700 26068 21710
rect 26012 21586 26068 21644
rect 26012 21534 26014 21586
rect 26066 21534 26068 21586
rect 26012 21522 26068 21534
rect 26236 21586 26292 22652
rect 26348 22484 26404 22494
rect 26348 21698 26404 22428
rect 26348 21646 26350 21698
rect 26402 21646 26404 21698
rect 26348 21634 26404 21646
rect 26236 21534 26238 21586
rect 26290 21534 26292 21586
rect 26236 21252 26292 21534
rect 26460 21588 26516 23436
rect 26572 23042 26628 23054
rect 26572 22990 26574 23042
rect 26626 22990 26628 23042
rect 26572 22708 26628 22990
rect 26572 22642 26628 22652
rect 26460 21522 26516 21532
rect 26684 21476 26740 29148
rect 26796 28756 26852 28766
rect 26908 28756 26964 31612
rect 26796 28754 26964 28756
rect 26796 28702 26798 28754
rect 26850 28702 26964 28754
rect 26796 28700 26964 28702
rect 26796 28690 26852 28700
rect 26796 28084 26852 28094
rect 26796 27990 26852 28028
rect 26796 26516 26852 26526
rect 26796 26178 26852 26460
rect 26796 26126 26798 26178
rect 26850 26126 26852 26178
rect 26796 24834 26852 26126
rect 26796 24782 26798 24834
rect 26850 24782 26852 24834
rect 26796 22484 26852 24782
rect 26908 23548 26964 28700
rect 27020 26908 27076 31724
rect 27132 31714 27188 31724
rect 27356 31668 27412 35084
rect 27468 34914 27524 36204
rect 27468 34862 27470 34914
rect 27522 34862 27524 34914
rect 27468 34356 27524 34862
rect 27468 34290 27524 34300
rect 27580 34916 27636 34926
rect 27692 34916 27748 37772
rect 27804 37762 27860 37772
rect 28140 37826 28196 37838
rect 28140 37774 28142 37826
rect 28194 37774 28196 37826
rect 28140 36484 28196 37774
rect 28364 37826 28420 37838
rect 28588 37828 28644 38220
rect 28364 37774 28366 37826
rect 28418 37774 28420 37826
rect 28252 37716 28308 37726
rect 28364 37716 28420 37774
rect 28308 37660 28420 37716
rect 28476 37772 28644 37828
rect 28252 37650 28308 37660
rect 28140 36418 28196 36428
rect 27636 34914 27748 34916
rect 27636 34862 27694 34914
rect 27746 34862 27748 34914
rect 27636 34860 27748 34862
rect 27468 33572 27524 33582
rect 27468 33478 27524 33516
rect 27580 33348 27636 34860
rect 27692 34850 27748 34860
rect 27916 36036 27972 36046
rect 27916 34914 27972 35980
rect 27916 34862 27918 34914
rect 27970 34862 27972 34914
rect 27916 34850 27972 34862
rect 28140 35700 28196 35710
rect 28028 34804 28084 34814
rect 28028 34710 28084 34748
rect 27692 34356 27748 34366
rect 27692 34262 27748 34300
rect 28028 34242 28084 34254
rect 28028 34190 28030 34242
rect 28082 34190 28084 34242
rect 28028 33572 28084 34190
rect 27580 33282 27636 33292
rect 27692 33516 28084 33572
rect 27692 33346 27748 33516
rect 27692 33294 27694 33346
rect 27746 33294 27748 33346
rect 27692 31892 27748 33294
rect 27916 33346 27972 33358
rect 27916 33294 27918 33346
rect 27970 33294 27972 33346
rect 27916 32900 27972 33294
rect 27916 32834 27972 32844
rect 27692 31826 27748 31836
rect 28140 31780 28196 35644
rect 28476 35140 28532 37772
rect 28588 36258 28644 36270
rect 28588 36206 28590 36258
rect 28642 36206 28644 36258
rect 28588 36148 28644 36206
rect 28588 36082 28644 36092
rect 28476 35074 28532 35084
rect 28476 34690 28532 34702
rect 28476 34638 28478 34690
rect 28530 34638 28532 34690
rect 28476 34356 28532 34638
rect 28476 34290 28532 34300
rect 28364 34244 28420 34254
rect 28364 34132 28420 34188
rect 28364 34130 28532 34132
rect 28364 34078 28366 34130
rect 28418 34078 28532 34130
rect 28364 34076 28532 34078
rect 28364 34066 28420 34076
rect 28476 33572 28532 34076
rect 28588 34020 28644 34030
rect 28588 33926 28644 33964
rect 28476 33348 28532 33516
rect 28588 33348 28644 33358
rect 28476 33346 28644 33348
rect 28476 33294 28590 33346
rect 28642 33294 28644 33346
rect 28476 33292 28644 33294
rect 28588 33282 28644 33292
rect 28364 33122 28420 33134
rect 28364 33070 28366 33122
rect 28418 33070 28420 33122
rect 28364 31892 28420 33070
rect 28476 33124 28532 33134
rect 28476 33030 28532 33068
rect 28364 31826 28420 31836
rect 28140 31714 28196 31724
rect 27244 31612 27412 31668
rect 28588 31668 28644 31678
rect 27244 31556 27300 31612
rect 28588 31574 28644 31612
rect 27468 31556 27524 31566
rect 27132 31500 27300 31556
rect 27356 31554 27524 31556
rect 27356 31502 27470 31554
rect 27522 31502 27524 31554
rect 27356 31500 27524 31502
rect 27132 30996 27188 31500
rect 27132 28754 27188 30940
rect 27356 31444 27412 31500
rect 27468 31490 27524 31500
rect 27692 31554 27748 31566
rect 27692 31502 27694 31554
rect 27746 31502 27748 31554
rect 27244 30884 27300 30894
rect 27244 30790 27300 30828
rect 27244 30100 27300 30110
rect 27244 30006 27300 30044
rect 27356 29764 27412 31388
rect 27692 31332 27748 31502
rect 27804 31556 27860 31566
rect 27804 31462 27860 31500
rect 28140 31554 28196 31566
rect 28140 31502 28142 31554
rect 28194 31502 28196 31554
rect 28140 31444 28196 31502
rect 28140 31378 28196 31388
rect 27692 31266 27748 31276
rect 28700 30996 28756 31006
rect 27468 30212 27524 30222
rect 27468 30118 27524 30156
rect 27580 30212 27636 30222
rect 28028 30212 28084 30222
rect 27580 30210 28084 30212
rect 27580 30158 27582 30210
rect 27634 30158 28030 30210
rect 28082 30158 28084 30210
rect 27580 30156 28084 30158
rect 27580 30146 27636 30156
rect 28028 30146 28084 30156
rect 28588 30212 28644 30222
rect 27692 29988 27748 29998
rect 28140 29988 28196 29998
rect 27692 29894 27748 29932
rect 28028 29986 28196 29988
rect 28028 29934 28142 29986
rect 28194 29934 28196 29986
rect 28028 29932 28196 29934
rect 27132 28702 27134 28754
rect 27186 28702 27188 28754
rect 27132 28690 27188 28702
rect 27244 29708 27412 29764
rect 27132 28084 27188 28094
rect 27132 27188 27188 28028
rect 27244 27748 27300 29708
rect 27356 29316 27412 29326
rect 28028 29316 28084 29932
rect 28140 29922 28196 29932
rect 28252 29986 28308 29998
rect 28252 29934 28254 29986
rect 28306 29934 28308 29986
rect 27356 29314 28084 29316
rect 27356 29262 27358 29314
rect 27410 29262 28084 29314
rect 27356 29260 28084 29262
rect 27356 29250 27412 29260
rect 28028 28868 28084 28878
rect 28252 28868 28308 29934
rect 28028 28866 28308 28868
rect 28028 28814 28030 28866
rect 28082 28814 28308 28866
rect 28028 28812 28308 28814
rect 28364 29988 28420 29998
rect 28364 28866 28420 29932
rect 28364 28814 28366 28866
rect 28418 28814 28420 28866
rect 28028 28802 28084 28812
rect 28364 28802 28420 28814
rect 28588 28754 28644 30156
rect 28700 30210 28756 30940
rect 28812 30772 28868 51100
rect 29036 49028 29092 51326
rect 29036 48962 29092 48972
rect 29036 48802 29092 48814
rect 29036 48750 29038 48802
rect 29090 48750 29092 48802
rect 28924 47572 28980 47582
rect 28924 47012 28980 47516
rect 29036 47236 29092 48750
rect 29036 47170 29092 47180
rect 28924 46956 29092 47012
rect 28924 43652 28980 43662
rect 28924 43558 28980 43596
rect 29036 38668 29092 46956
rect 29148 46452 29204 52220
rect 29372 52050 29428 53676
rect 29484 53666 29540 53676
rect 29708 53620 29764 53630
rect 29708 53506 29764 53564
rect 29708 53454 29710 53506
rect 29762 53454 29764 53506
rect 29484 52946 29540 52958
rect 29484 52894 29486 52946
rect 29538 52894 29540 52946
rect 29484 52834 29540 52894
rect 29484 52782 29486 52834
rect 29538 52782 29540 52834
rect 29484 52770 29540 52782
rect 29596 52612 29652 52622
rect 29372 51998 29374 52050
rect 29426 51998 29428 52050
rect 29372 51986 29428 51998
rect 29484 52500 29540 52510
rect 29484 50820 29540 52444
rect 29596 52050 29652 52556
rect 29596 51998 29598 52050
rect 29650 51998 29652 52050
rect 29596 51986 29652 51998
rect 29708 51828 29764 53454
rect 29932 53508 29988 54796
rect 30044 53620 30100 55468
rect 30268 55186 30324 58156
rect 31500 58118 31556 58156
rect 30828 57876 30884 57886
rect 30828 57782 30884 57820
rect 30940 57652 30996 57662
rect 30940 57558 30996 57596
rect 31276 57540 31332 57550
rect 31388 57540 31444 57550
rect 31332 57538 31444 57540
rect 31332 57486 31390 57538
rect 31442 57486 31444 57538
rect 31332 57484 31444 57486
rect 30380 56980 30436 56990
rect 30380 56306 30436 56924
rect 31052 56868 31108 56878
rect 30492 56644 30548 56654
rect 30940 56644 30996 56654
rect 31052 56644 31108 56812
rect 30492 56642 31108 56644
rect 30492 56590 30494 56642
rect 30546 56590 30942 56642
rect 30994 56590 31108 56642
rect 30492 56588 31108 56590
rect 30492 56578 30548 56588
rect 30940 56578 30996 56588
rect 30380 56254 30382 56306
rect 30434 56254 30436 56306
rect 30380 56242 30436 56254
rect 30268 55134 30270 55186
rect 30322 55134 30324 55186
rect 30268 55122 30324 55134
rect 30380 55412 30436 55422
rect 30156 54628 30212 54638
rect 30156 54534 30212 54572
rect 30044 53526 30100 53564
rect 30268 53732 30324 53742
rect 29932 53442 29988 53452
rect 30044 53172 30100 53182
rect 30044 53078 30100 53116
rect 30268 53170 30324 53676
rect 30380 53618 30436 55356
rect 30492 55300 30548 55310
rect 30548 55244 30660 55300
rect 30492 55234 30548 55244
rect 30492 54626 30548 54638
rect 30492 54574 30494 54626
rect 30546 54574 30548 54626
rect 30492 54516 30548 54574
rect 30492 54450 30548 54460
rect 30380 53566 30382 53618
rect 30434 53566 30436 53618
rect 30380 53554 30436 53566
rect 30604 53284 30660 55244
rect 30716 55076 30772 55086
rect 30716 54982 30772 55020
rect 30268 53118 30270 53170
rect 30322 53118 30324 53170
rect 30268 53106 30324 53118
rect 30492 53228 30660 53284
rect 30828 54740 30884 54750
rect 30156 53060 30212 53070
rect 29820 52834 29876 52846
rect 29820 52782 29822 52834
rect 29874 52782 29876 52834
rect 29820 52724 29876 52782
rect 29932 52724 29988 52734
rect 29820 52722 29988 52724
rect 29820 52670 29934 52722
rect 29986 52670 29988 52722
rect 29820 52668 29988 52670
rect 29932 52658 29988 52668
rect 30156 52162 30212 53004
rect 30156 52110 30158 52162
rect 30210 52110 30212 52162
rect 30156 52098 30212 52110
rect 30380 52724 30436 52734
rect 30380 52050 30436 52668
rect 30380 51998 30382 52050
rect 30434 51998 30436 52050
rect 30380 51986 30436 51998
rect 29932 51940 29988 51950
rect 29932 51846 29988 51884
rect 30044 51938 30100 51950
rect 30044 51886 30046 51938
rect 30098 51886 30100 51938
rect 29484 50754 29540 50764
rect 29596 51772 29764 51828
rect 29596 50596 29652 51772
rect 29708 51268 29764 51278
rect 29708 51266 29988 51268
rect 29708 51214 29710 51266
rect 29762 51214 29988 51266
rect 29708 51212 29988 51214
rect 29708 51202 29764 51212
rect 29932 50818 29988 51212
rect 29932 50766 29934 50818
rect 29986 50766 29988 50818
rect 29932 50754 29988 50766
rect 30044 50706 30100 51886
rect 30044 50654 30046 50706
rect 30098 50654 30100 50706
rect 30044 50642 30100 50654
rect 29484 50540 29652 50596
rect 29372 49588 29428 49598
rect 29260 49586 29428 49588
rect 29260 49534 29374 49586
rect 29426 49534 29428 49586
rect 29260 49532 29428 49534
rect 29260 48804 29316 49532
rect 29372 49522 29428 49532
rect 29260 48710 29316 48748
rect 29372 48914 29428 48926
rect 29372 48862 29374 48914
rect 29426 48862 29428 48914
rect 29260 47234 29316 47246
rect 29260 47182 29262 47234
rect 29314 47182 29316 47234
rect 29260 46900 29316 47182
rect 29372 47124 29428 48862
rect 29372 47058 29428 47068
rect 29260 46834 29316 46844
rect 29260 46676 29316 46686
rect 29484 46676 29540 50540
rect 30380 49924 30436 49934
rect 30380 49830 30436 49868
rect 30156 49812 30212 49822
rect 30156 49718 30212 49756
rect 29596 49698 29652 49710
rect 29596 49646 29598 49698
rect 29650 49646 29652 49698
rect 29596 49586 29652 49646
rect 29596 49534 29598 49586
rect 29650 49534 29652 49586
rect 29596 49522 29652 49534
rect 30268 49588 30324 49598
rect 30268 49586 30436 49588
rect 30268 49534 30270 49586
rect 30322 49534 30436 49586
rect 30268 49532 30436 49534
rect 30268 49522 30324 49532
rect 29820 49028 29876 49038
rect 29820 48804 29876 48972
rect 29820 48748 30324 48804
rect 29932 48244 29988 48254
rect 29820 47460 29876 47470
rect 29820 47366 29876 47404
rect 29596 47348 29652 47358
rect 29596 47254 29652 47292
rect 29708 47234 29764 47246
rect 29708 47182 29710 47234
rect 29762 47182 29764 47234
rect 29708 47124 29764 47182
rect 29708 47058 29764 47068
rect 29932 46786 29988 48188
rect 30156 47458 30212 47470
rect 30156 47406 30158 47458
rect 30210 47406 30212 47458
rect 30156 47124 30212 47406
rect 30156 47058 30212 47068
rect 29932 46734 29934 46786
rect 29986 46734 29988 46786
rect 29708 46676 29764 46686
rect 29260 46674 29764 46676
rect 29260 46622 29262 46674
rect 29314 46622 29710 46674
rect 29762 46622 29764 46674
rect 29260 46620 29764 46622
rect 29260 46610 29316 46620
rect 29148 46396 29428 46452
rect 29260 46228 29316 46238
rect 29148 45108 29204 45118
rect 29148 45014 29204 45052
rect 29260 44884 29316 46172
rect 29372 45220 29428 46396
rect 29372 45126 29428 45164
rect 29596 44996 29652 45006
rect 29596 44902 29652 44940
rect 29148 44828 29316 44884
rect 29708 44884 29764 46620
rect 29820 45108 29876 45118
rect 29932 45108 29988 46734
rect 29820 45106 29988 45108
rect 29820 45054 29822 45106
rect 29874 45054 29988 45106
rect 29820 45052 29988 45054
rect 30268 45778 30324 48748
rect 30380 46674 30436 49532
rect 30492 49140 30548 53228
rect 30828 53172 30884 54684
rect 30940 54516 30996 54526
rect 31052 54516 31108 56588
rect 31164 55074 31220 55086
rect 31164 55022 31166 55074
rect 31218 55022 31220 55074
rect 31164 54852 31220 55022
rect 31276 55076 31332 57484
rect 31388 57474 31444 57484
rect 31612 56644 31668 56654
rect 31276 55010 31332 55020
rect 31500 56196 31556 56206
rect 31164 54738 31220 54796
rect 31164 54686 31166 54738
rect 31218 54686 31220 54738
rect 31164 54674 31220 54686
rect 31052 54460 31220 54516
rect 30940 54422 30996 54460
rect 31052 53732 31108 53742
rect 30828 53078 30884 53116
rect 30940 53284 30996 53294
rect 30604 52946 30660 52958
rect 30604 52894 30606 52946
rect 30658 52894 30660 52946
rect 30604 52164 30660 52894
rect 30716 52724 30772 52734
rect 30716 52630 30772 52668
rect 30716 52164 30772 52174
rect 30604 52162 30772 52164
rect 30604 52110 30718 52162
rect 30770 52110 30772 52162
rect 30604 52108 30772 52110
rect 30716 52098 30772 52108
rect 30940 52052 30996 53228
rect 31052 53170 31108 53676
rect 31052 53118 31054 53170
rect 31106 53118 31108 53170
rect 31052 53106 31108 53118
rect 30940 51958 30996 51996
rect 31052 52050 31108 52062
rect 31052 51998 31054 52050
rect 31106 51998 31108 52050
rect 31052 51940 31108 51998
rect 30940 50370 30996 50382
rect 30940 50318 30942 50370
rect 30994 50318 30996 50370
rect 30940 50148 30996 50318
rect 31052 50148 31108 51884
rect 31164 50372 31220 54460
rect 31388 52948 31444 52958
rect 31388 52854 31444 52892
rect 31388 52724 31444 52734
rect 31388 51492 31444 52668
rect 31500 51828 31556 56140
rect 31612 54404 31668 56588
rect 31612 54338 31668 54348
rect 31724 55410 31780 61180
rect 32732 61012 32788 61518
rect 32732 60946 32788 60956
rect 32060 60900 32116 60910
rect 31836 59778 31892 59790
rect 31836 59726 31838 59778
rect 31890 59726 31892 59778
rect 31836 58212 31892 59726
rect 32060 59444 32116 60844
rect 32284 60786 32340 60798
rect 32284 60734 32286 60786
rect 32338 60734 32340 60786
rect 32172 60002 32228 60014
rect 32172 59950 32174 60002
rect 32226 59950 32228 60002
rect 32172 59668 32228 59950
rect 32284 60004 32340 60734
rect 32508 60788 32564 60798
rect 32284 59938 32340 59948
rect 32396 60674 32452 60686
rect 32396 60622 32398 60674
rect 32450 60622 32452 60674
rect 32396 59892 32452 60622
rect 32396 59826 32452 59836
rect 32172 59602 32228 59612
rect 32508 59556 32564 60732
rect 32956 60786 33012 62078
rect 32956 60734 32958 60786
rect 33010 60734 33012 60786
rect 32956 60722 33012 60734
rect 33180 61460 33236 61470
rect 32844 60676 32900 60686
rect 32844 60114 32900 60620
rect 33180 60674 33236 61404
rect 33180 60622 33182 60674
rect 33234 60622 33236 60674
rect 33180 60610 33236 60622
rect 32844 60062 32846 60114
rect 32898 60062 32900 60114
rect 32844 60050 32900 60062
rect 33068 60004 33124 60014
rect 33124 59948 33236 60004
rect 33068 59938 33124 59948
rect 32508 59500 33012 59556
rect 32060 59388 32452 59444
rect 32284 59220 32340 59230
rect 31948 59218 32340 59220
rect 31948 59166 32286 59218
rect 32338 59166 32340 59218
rect 31948 59164 32340 59166
rect 31948 59106 32004 59164
rect 32284 59154 32340 59164
rect 31948 59054 31950 59106
rect 32002 59054 32004 59106
rect 31948 59042 32004 59054
rect 32396 58994 32452 59388
rect 32396 58942 32398 58994
rect 32450 58942 32452 58994
rect 32396 58436 32452 58942
rect 32396 58370 32452 58380
rect 32620 59332 32676 59342
rect 31948 58212 32004 58222
rect 31836 58156 31948 58212
rect 31836 57652 31892 57662
rect 31836 56866 31892 57596
rect 31948 57316 32004 58156
rect 32620 57874 32676 59276
rect 32844 58884 32900 58894
rect 32732 58660 32788 58670
rect 32732 58546 32788 58604
rect 32732 58494 32734 58546
rect 32786 58494 32788 58546
rect 32732 58482 32788 58494
rect 32620 57822 32622 57874
rect 32674 57822 32676 57874
rect 32620 57810 32676 57822
rect 31948 57260 32228 57316
rect 31836 56814 31838 56866
rect 31890 56814 31892 56866
rect 31836 56196 31892 56814
rect 31836 56130 31892 56140
rect 31836 55970 31892 55982
rect 31836 55918 31838 55970
rect 31890 55918 31892 55970
rect 31836 55524 31892 55918
rect 32060 55524 32116 55534
rect 31836 55468 32060 55524
rect 31724 55358 31726 55410
rect 31778 55358 31780 55410
rect 31612 53842 31668 53854
rect 31612 53790 31614 53842
rect 31666 53790 31668 53842
rect 31612 53508 31668 53790
rect 31612 53442 31668 53452
rect 31724 52724 31780 55358
rect 32060 55298 32116 55468
rect 32060 55246 32062 55298
rect 32114 55246 32116 55298
rect 32060 55234 32116 55246
rect 32172 55076 32228 57260
rect 32844 56866 32900 58828
rect 32956 58434 33012 59500
rect 33068 59444 33124 59454
rect 33180 59444 33236 59948
rect 33068 59442 33236 59444
rect 33068 59390 33070 59442
rect 33122 59390 33236 59442
rect 33068 59388 33236 59390
rect 33292 59556 33348 62132
rect 33404 60340 33460 62524
rect 33516 62468 33572 62478
rect 33516 62374 33572 62412
rect 33628 61682 33684 61694
rect 33628 61630 33630 61682
rect 33682 61630 33684 61682
rect 33628 60788 33684 61630
rect 33740 61458 33796 65884
rect 33852 64146 33908 66108
rect 34076 66162 34356 66164
rect 34076 66110 34078 66162
rect 34130 66110 34356 66162
rect 34076 66108 34356 66110
rect 34076 66098 34132 66108
rect 33964 66052 34020 66062
rect 33964 65958 34020 65996
rect 34188 65604 34244 65614
rect 34188 65510 34244 65548
rect 33964 65490 34020 65502
rect 33964 65438 33966 65490
rect 34018 65438 34020 65490
rect 33964 65380 34020 65438
rect 33964 65314 34020 65324
rect 34076 65378 34132 65390
rect 34076 65326 34078 65378
rect 34130 65326 34132 65378
rect 34076 65268 34132 65326
rect 34076 65202 34132 65212
rect 34076 64820 34132 64830
rect 34300 64820 34356 66108
rect 34076 64818 34356 64820
rect 34076 64766 34078 64818
rect 34130 64766 34356 64818
rect 34076 64764 34356 64766
rect 34076 64754 34132 64764
rect 34076 64596 34132 64606
rect 33852 64094 33854 64146
rect 33906 64094 33908 64146
rect 33852 64082 33908 64094
rect 33964 64260 34020 64270
rect 33852 62356 33908 62366
rect 33852 62262 33908 62300
rect 33964 62130 34020 64204
rect 34076 64034 34132 64540
rect 34076 63982 34078 64034
rect 34130 63982 34132 64034
rect 34076 62578 34132 63982
rect 34188 64036 34244 64046
rect 34188 63942 34244 63980
rect 34076 62526 34078 62578
rect 34130 62526 34132 62578
rect 34076 62514 34132 62526
rect 34300 62916 34356 64764
rect 34524 65490 34580 65502
rect 34524 65438 34526 65490
rect 34578 65438 34580 65490
rect 34412 64594 34468 64606
rect 34412 64542 34414 64594
rect 34466 64542 34468 64594
rect 34412 64484 34468 64542
rect 34412 64418 34468 64428
rect 34524 64260 34580 65438
rect 34972 65492 35028 65502
rect 34972 64930 35028 65436
rect 34972 64878 34974 64930
rect 35026 64878 35028 64930
rect 34972 64866 35028 64878
rect 34524 64194 34580 64204
rect 34636 64706 34692 64718
rect 34636 64654 34638 64706
rect 34690 64654 34692 64706
rect 34636 64148 34692 64654
rect 34972 64596 35028 64606
rect 35084 64596 35140 68908
rect 35532 69298 35588 69310
rect 35532 69246 35534 69298
rect 35586 69246 35588 69298
rect 35532 68964 35588 69246
rect 35644 69188 35700 69198
rect 35644 69186 35812 69188
rect 35644 69134 35646 69186
rect 35698 69134 35812 69186
rect 35644 69132 35812 69134
rect 35644 69122 35700 69132
rect 35532 68898 35588 68908
rect 35644 68626 35700 68638
rect 35644 68574 35646 68626
rect 35698 68574 35700 68626
rect 35308 68516 35364 68526
rect 35644 68516 35700 68574
rect 35756 68628 35812 69132
rect 35756 68562 35812 68572
rect 35980 68738 36036 68750
rect 35980 68686 35982 68738
rect 36034 68686 36036 68738
rect 35308 68514 35700 68516
rect 35308 68462 35310 68514
rect 35362 68462 35700 68514
rect 35308 68460 35700 68462
rect 35980 68516 36036 68686
rect 35308 68450 35364 68460
rect 35196 68236 35460 68246
rect 35252 68180 35300 68236
rect 35356 68180 35404 68236
rect 35196 68170 35460 68180
rect 35532 67060 35588 68460
rect 35980 68450 36036 68460
rect 36092 68516 36148 69356
rect 36988 69412 37044 71598
rect 37212 70866 37268 70878
rect 37212 70814 37214 70866
rect 37266 70814 37268 70866
rect 37212 70532 37268 70814
rect 37212 70466 37268 70476
rect 38444 70644 38500 70654
rect 37212 70082 37268 70094
rect 37212 70030 37214 70082
rect 37266 70030 37268 70082
rect 37212 69636 37268 70030
rect 37212 69570 37268 69580
rect 38444 69522 38500 70588
rect 39564 70532 39620 70542
rect 39340 70084 39396 70094
rect 39340 70082 39508 70084
rect 39340 70030 39342 70082
rect 39394 70030 39508 70082
rect 39340 70028 39508 70030
rect 39340 70018 39396 70028
rect 38444 69470 38446 69522
rect 38498 69470 38500 69522
rect 38444 69458 38500 69470
rect 36988 69346 37044 69356
rect 38556 69412 38612 69422
rect 36316 69300 36372 69310
rect 36316 69206 36372 69244
rect 37548 69300 37604 69310
rect 37548 69206 37604 69244
rect 37212 69186 37268 69198
rect 37212 69134 37214 69186
rect 37266 69134 37268 69186
rect 36428 68738 36484 68750
rect 36428 68686 36430 68738
rect 36482 68686 36484 68738
rect 36316 68626 36372 68638
rect 36316 68574 36318 68626
rect 36370 68574 36372 68626
rect 36316 68516 36372 68574
rect 36092 68460 36372 68516
rect 36428 68628 36484 68686
rect 36652 68740 36708 68750
rect 36652 68738 36820 68740
rect 36652 68686 36654 68738
rect 36706 68686 36820 68738
rect 36652 68684 36820 68686
rect 36652 68674 36708 68684
rect 35644 67620 35700 67630
rect 35868 67620 35924 67630
rect 35644 67618 35868 67620
rect 35644 67566 35646 67618
rect 35698 67566 35868 67618
rect 35644 67564 35868 67566
rect 35644 67554 35700 67564
rect 35868 67526 35924 67564
rect 36092 67396 36148 68460
rect 36428 68404 36484 68572
rect 36764 68626 36820 68684
rect 36764 68574 36766 68626
rect 36818 68574 36820 68626
rect 36764 68562 36820 68574
rect 37100 68626 37156 68638
rect 37100 68574 37102 68626
rect 37154 68574 37156 68626
rect 37100 68516 37156 68574
rect 37100 68450 37156 68460
rect 37212 68514 37268 69134
rect 37436 69188 37492 69198
rect 37436 69094 37492 69132
rect 37660 69186 37716 69198
rect 37660 69134 37662 69186
rect 37714 69134 37716 69186
rect 37324 68852 37380 68890
rect 37324 68786 37380 68796
rect 37212 68462 37214 68514
rect 37266 68462 37268 68514
rect 37212 68450 37268 68462
rect 37324 68628 37380 68638
rect 37548 68628 37604 68638
rect 36204 68348 36484 68404
rect 36204 67730 36260 68348
rect 36204 67678 36206 67730
rect 36258 67678 36260 67730
rect 36204 67666 36260 67678
rect 37324 67732 37380 68572
rect 37436 68626 37604 68628
rect 37436 68574 37550 68626
rect 37602 68574 37604 68626
rect 37436 68572 37604 68574
rect 37436 68066 37492 68572
rect 37548 68562 37604 68572
rect 37436 68014 37438 68066
rect 37490 68014 37492 68066
rect 37436 68002 37492 68014
rect 37548 67844 37604 67854
rect 37660 67844 37716 69134
rect 38108 69188 38164 69198
rect 38332 69188 38388 69198
rect 38108 69186 38276 69188
rect 38108 69134 38110 69186
rect 38162 69134 38276 69186
rect 38108 69132 38276 69134
rect 38108 69122 38164 69132
rect 38108 68852 38164 68862
rect 38108 68758 38164 68796
rect 38220 68850 38276 69132
rect 38220 68798 38222 68850
rect 38274 68798 38276 68850
rect 38220 68786 38276 68798
rect 37884 68626 37940 68638
rect 37884 68574 37886 68626
rect 37938 68574 37940 68626
rect 37884 68516 37940 68574
rect 37884 68450 37940 68460
rect 37548 67842 37660 67844
rect 37548 67790 37550 67842
rect 37602 67790 37660 67842
rect 37548 67788 37660 67790
rect 37548 67778 37604 67788
rect 37660 67750 37716 67788
rect 37436 67732 37492 67742
rect 37324 67730 37492 67732
rect 37324 67678 37438 67730
rect 37490 67678 37492 67730
rect 37324 67676 37492 67678
rect 38332 67732 38388 69132
rect 38556 69186 38612 69356
rect 39228 69300 39284 69310
rect 38556 69134 38558 69186
rect 38610 69134 38612 69186
rect 38444 68964 38500 68974
rect 38556 68964 38612 69134
rect 39116 69298 39284 69300
rect 39116 69246 39230 69298
rect 39282 69246 39284 69298
rect 39116 69244 39284 69246
rect 38556 68908 38948 68964
rect 38444 68628 38500 68908
rect 38780 68738 38836 68750
rect 38780 68686 38782 68738
rect 38834 68686 38836 68738
rect 38556 68628 38612 68638
rect 38444 68626 38612 68628
rect 38444 68574 38558 68626
rect 38610 68574 38612 68626
rect 38444 68572 38612 68574
rect 38444 67732 38500 67742
rect 38332 67730 38500 67732
rect 38332 67678 38446 67730
rect 38498 67678 38500 67730
rect 38332 67676 38500 67678
rect 37436 67666 37492 67676
rect 38444 67666 38500 67676
rect 38108 67618 38164 67630
rect 38108 67566 38110 67618
rect 38162 67566 38164 67618
rect 38108 67508 38164 67566
rect 38108 67442 38164 67452
rect 35532 66994 35588 67004
rect 35644 67340 36148 67396
rect 35196 66668 35460 66678
rect 35252 66612 35300 66668
rect 35356 66612 35404 66668
rect 35196 66602 35460 66612
rect 35196 66274 35252 66286
rect 35196 66222 35198 66274
rect 35250 66222 35252 66274
rect 35196 65492 35252 66222
rect 35420 66274 35476 66286
rect 35420 66222 35422 66274
rect 35474 66222 35476 66274
rect 35420 66052 35476 66222
rect 35420 65986 35476 65996
rect 35196 65426 35252 65436
rect 35196 65100 35460 65110
rect 35252 65044 35300 65100
rect 35356 65044 35404 65100
rect 35196 65034 35460 65044
rect 35028 64540 35140 64596
rect 34972 64530 35028 64540
rect 35644 64372 35700 67340
rect 36764 66948 36820 66958
rect 36652 66946 36820 66948
rect 36652 66894 36766 66946
rect 36818 66894 36820 66946
rect 36652 66892 36820 66894
rect 36204 66164 36260 66174
rect 35756 66052 35812 66062
rect 35756 66050 36148 66052
rect 35756 65998 35758 66050
rect 35810 65998 36148 66050
rect 35756 65996 36148 65998
rect 35756 65986 35812 65996
rect 35756 64708 35812 64746
rect 35756 64642 35812 64652
rect 35868 64706 35924 64718
rect 35868 64654 35870 64706
rect 35922 64654 35924 64706
rect 35868 64372 35924 64654
rect 35644 64316 35924 64372
rect 35980 64594 36036 64606
rect 35980 64542 35982 64594
rect 36034 64542 36036 64594
rect 35980 64372 36036 64542
rect 34636 64082 34692 64092
rect 34524 63812 34580 63822
rect 34524 63718 34580 63756
rect 35196 63532 35460 63542
rect 35252 63476 35300 63532
rect 35356 63476 35404 63532
rect 35196 63466 35460 63476
rect 35756 63252 35812 64316
rect 35980 64306 36036 64316
rect 36092 64148 36148 65996
rect 36204 64932 36260 66108
rect 36428 66162 36484 66174
rect 36428 66110 36430 66162
rect 36482 66110 36484 66162
rect 36316 66052 36372 66062
rect 36316 65958 36372 65996
rect 36428 65268 36484 66110
rect 36428 65202 36484 65212
rect 36428 64932 36484 64942
rect 36204 64930 36484 64932
rect 36204 64878 36430 64930
rect 36482 64878 36484 64930
rect 36204 64876 36484 64878
rect 36428 64866 36484 64876
rect 36652 64372 36708 66892
rect 36764 66882 36820 66892
rect 38556 66612 38612 68572
rect 38780 67844 38836 68686
rect 38892 68628 38948 68908
rect 39116 68852 39172 69244
rect 39228 69234 39284 69244
rect 39340 69300 39396 69310
rect 39340 69206 39396 69244
rect 39340 68964 39396 68974
rect 39452 68964 39508 70028
rect 39564 69412 39620 70476
rect 39900 70308 39956 71710
rect 40236 71652 40292 71662
rect 40236 70418 40292 71596
rect 40348 71650 40404 71662
rect 40348 71598 40350 71650
rect 40402 71598 40404 71650
rect 40348 70644 40404 71598
rect 40908 71652 40964 71662
rect 40908 71558 40964 71596
rect 41020 71540 41076 71550
rect 41020 71538 41748 71540
rect 41020 71486 41022 71538
rect 41074 71486 41748 71538
rect 41020 71484 41748 71486
rect 41020 71474 41076 71484
rect 40348 70578 40404 70588
rect 40236 70366 40238 70418
rect 40290 70366 40292 70418
rect 40236 70354 40292 70366
rect 39900 70242 39956 70252
rect 40908 70308 40964 70318
rect 39788 70194 39844 70206
rect 39788 70142 39790 70194
rect 39842 70142 39844 70194
rect 39676 69412 39732 69422
rect 39564 69410 39732 69412
rect 39564 69358 39678 69410
rect 39730 69358 39732 69410
rect 39564 69356 39732 69358
rect 39676 69346 39732 69356
rect 39788 69300 39844 70142
rect 40124 70194 40180 70206
rect 40124 70142 40126 70194
rect 40178 70142 40180 70194
rect 39788 69244 39956 69300
rect 39396 68908 39508 68964
rect 39340 68898 39396 68908
rect 39116 68786 39172 68796
rect 39228 68740 39284 68750
rect 39228 68646 39284 68684
rect 39116 68628 39172 68638
rect 38892 68626 39172 68628
rect 38892 68574 39118 68626
rect 39170 68574 39172 68626
rect 38892 68572 39172 68574
rect 39004 67844 39060 67854
rect 38780 67788 39004 67844
rect 38780 67618 38836 67630
rect 38780 67566 38782 67618
rect 38834 67566 38836 67618
rect 38780 67508 38836 67566
rect 38780 67442 38836 67452
rect 38108 66556 38612 66612
rect 37324 66276 37380 66286
rect 37324 66274 37492 66276
rect 37324 66222 37326 66274
rect 37378 66222 37492 66274
rect 37324 66220 37492 66222
rect 37324 66210 37380 66220
rect 36988 66164 37044 66174
rect 36988 66070 37044 66108
rect 37324 66050 37380 66062
rect 37324 65998 37326 66050
rect 37378 65998 37380 66050
rect 37324 65716 37380 65998
rect 36652 64306 36708 64316
rect 36764 65660 37380 65716
rect 35756 63186 35812 63196
rect 35868 64092 36148 64148
rect 34300 62466 34356 62860
rect 34748 63138 34804 63150
rect 34748 63086 34750 63138
rect 34802 63086 34804 63138
rect 34748 62580 34804 63086
rect 35868 63138 35924 64092
rect 36652 63812 36708 63822
rect 35980 63810 36708 63812
rect 35980 63758 36654 63810
rect 36706 63758 36708 63810
rect 35980 63756 36708 63758
rect 35980 63250 36036 63756
rect 36652 63746 36708 63756
rect 35980 63198 35982 63250
rect 36034 63198 36036 63250
rect 35980 63186 36036 63198
rect 36092 63364 36148 63374
rect 35868 63086 35870 63138
rect 35922 63086 35924 63138
rect 35868 63074 35924 63086
rect 36092 63138 36148 63308
rect 36092 63086 36094 63138
rect 36146 63086 36148 63138
rect 36092 63074 36148 63086
rect 35196 62916 35252 62926
rect 35196 62822 35252 62860
rect 35644 62916 35700 62926
rect 35644 62822 35700 62860
rect 34748 62514 34804 62524
rect 35644 62692 35700 62702
rect 34300 62414 34302 62466
rect 34354 62414 34356 62466
rect 34300 62356 34356 62414
rect 33964 62078 33966 62130
rect 34018 62078 34020 62130
rect 33964 62066 34020 62078
rect 34076 62300 34356 62356
rect 35196 62356 35252 62366
rect 34076 61908 34132 62300
rect 35196 62262 35252 62300
rect 34748 62242 34804 62254
rect 34748 62190 34750 62242
rect 34802 62190 34804 62242
rect 33740 61406 33742 61458
rect 33794 61406 33796 61458
rect 33740 61394 33796 61406
rect 33852 61852 34132 61908
rect 34188 62020 34244 62030
rect 33628 60674 33684 60732
rect 33740 60900 33796 60910
rect 33740 60786 33796 60844
rect 33740 60734 33742 60786
rect 33794 60734 33796 60786
rect 33740 60722 33796 60734
rect 33628 60622 33630 60674
rect 33682 60622 33684 60674
rect 33628 60610 33684 60622
rect 33404 60284 33684 60340
rect 33068 58660 33124 59388
rect 33180 58884 33236 58894
rect 33292 58884 33348 59500
rect 33516 59332 33572 59342
rect 33236 58828 33348 58884
rect 33404 59276 33516 59332
rect 33180 58818 33236 58828
rect 33404 58772 33460 59276
rect 33516 59238 33572 59276
rect 33628 59330 33684 60284
rect 33628 59278 33630 59330
rect 33682 59278 33684 59330
rect 33628 59266 33684 59278
rect 33740 59218 33796 59230
rect 33740 59166 33742 59218
rect 33794 59166 33796 59218
rect 33292 58716 33460 58772
rect 33516 58884 33572 58894
rect 33180 58660 33236 58670
rect 33068 58658 33236 58660
rect 33068 58606 33182 58658
rect 33234 58606 33236 58658
rect 33068 58604 33236 58606
rect 33180 58594 33236 58604
rect 32956 58382 32958 58434
rect 33010 58382 33012 58434
rect 32956 58370 33012 58382
rect 33180 58436 33236 58446
rect 32844 56814 32846 56866
rect 32898 56814 32900 56866
rect 32284 56642 32340 56654
rect 32284 56590 32286 56642
rect 32338 56590 32340 56642
rect 32284 56532 32340 56590
rect 32284 56466 32340 56476
rect 32508 56644 32564 56654
rect 32508 56306 32564 56588
rect 32508 56254 32510 56306
rect 32562 56254 32564 56306
rect 32508 56242 32564 56254
rect 32396 56084 32452 56094
rect 32396 55186 32452 56028
rect 32396 55134 32398 55186
rect 32450 55134 32452 55186
rect 32396 55122 32452 55134
rect 31948 55020 32228 55076
rect 31836 54740 31892 54750
rect 31836 54646 31892 54684
rect 31724 52658 31780 52668
rect 31836 52834 31892 52846
rect 31836 52782 31838 52834
rect 31890 52782 31892 52834
rect 31836 52164 31892 52782
rect 31836 52098 31892 52108
rect 31500 51772 31892 51828
rect 31836 51492 31892 51772
rect 31388 51436 31556 51492
rect 31388 51268 31444 51278
rect 31164 50306 31220 50316
rect 31276 51212 31388 51268
rect 31276 50594 31332 51212
rect 31388 51202 31444 51212
rect 31276 50542 31278 50594
rect 31330 50542 31332 50594
rect 30940 50092 31220 50148
rect 30604 49922 30660 49934
rect 30604 49870 30606 49922
rect 30658 49870 30660 49922
rect 30604 49364 30660 49870
rect 31164 49924 31220 50092
rect 30604 49298 30660 49308
rect 30716 49812 30772 49822
rect 30492 49084 30660 49140
rect 30492 48916 30548 48926
rect 30492 48822 30548 48860
rect 30492 47460 30548 47470
rect 30492 47366 30548 47404
rect 30380 46622 30382 46674
rect 30434 46622 30436 46674
rect 30380 46610 30436 46622
rect 30268 45726 30270 45778
rect 30322 45726 30324 45778
rect 29820 45042 29876 45052
rect 29708 44828 29876 44884
rect 29148 43650 29204 44828
rect 29260 44100 29316 44110
rect 29260 44006 29316 44044
rect 29148 43598 29150 43650
rect 29202 43598 29204 43650
rect 29148 43586 29204 43598
rect 29596 43652 29652 43662
rect 29484 43538 29540 43550
rect 29484 43486 29486 43538
rect 29538 43486 29540 43538
rect 29372 43428 29428 43438
rect 29260 43426 29428 43428
rect 29260 43374 29374 43426
rect 29426 43374 29428 43426
rect 29260 43372 29428 43374
rect 29260 42644 29316 43372
rect 29372 43362 29428 43372
rect 29148 42588 29316 42644
rect 29148 41970 29204 42588
rect 29484 42532 29540 43486
rect 29596 42756 29652 43596
rect 29596 42662 29652 42700
rect 29708 42642 29764 42654
rect 29708 42590 29710 42642
rect 29762 42590 29764 42642
rect 29596 42532 29652 42542
rect 29484 42476 29596 42532
rect 29596 42466 29652 42476
rect 29708 42084 29764 42590
rect 29708 42018 29764 42028
rect 29148 41918 29150 41970
rect 29202 41918 29204 41970
rect 29148 41906 29204 41918
rect 29260 41970 29316 41982
rect 29260 41918 29262 41970
rect 29314 41918 29316 41970
rect 29148 41412 29204 41422
rect 29260 41412 29316 41918
rect 29484 41970 29540 41982
rect 29484 41918 29486 41970
rect 29538 41918 29540 41970
rect 29372 41860 29428 41870
rect 29372 41766 29428 41804
rect 29484 41636 29540 41918
rect 29484 41570 29540 41580
rect 29596 41970 29652 41982
rect 29596 41918 29598 41970
rect 29650 41918 29652 41970
rect 29260 41356 29428 41412
rect 29148 41298 29204 41356
rect 29148 41246 29150 41298
rect 29202 41246 29204 41298
rect 29148 41234 29204 41246
rect 29260 41188 29316 41198
rect 29260 41094 29316 41132
rect 29372 39396 29428 41356
rect 29596 39620 29652 41918
rect 29596 39554 29652 39564
rect 29708 41186 29764 41198
rect 29708 41134 29710 41186
rect 29762 41134 29764 41186
rect 29372 39330 29428 39340
rect 29596 38948 29652 38958
rect 29596 38854 29652 38892
rect 28924 38612 29092 38668
rect 29708 38612 29764 41134
rect 29820 40628 29876 44828
rect 30268 44324 30324 45726
rect 30380 46450 30436 46462
rect 30380 46398 30382 46450
rect 30434 46398 30436 46450
rect 30380 45780 30436 46398
rect 30380 45714 30436 45724
rect 30492 44324 30548 44334
rect 30268 44322 30548 44324
rect 30268 44270 30494 44322
rect 30546 44270 30548 44322
rect 30268 44268 30548 44270
rect 29932 43540 29988 43550
rect 29932 43446 29988 43484
rect 30156 42754 30212 42766
rect 30156 42702 30158 42754
rect 30210 42702 30212 42754
rect 29932 42530 29988 42542
rect 29932 42478 29934 42530
rect 29986 42478 29988 42530
rect 29932 40852 29988 42478
rect 30156 42532 30212 42702
rect 30156 42466 30212 42476
rect 29932 40786 29988 40796
rect 29820 40572 29988 40628
rect 29820 39508 29876 39518
rect 29820 39414 29876 39452
rect 28924 36932 28980 38612
rect 29484 38556 29708 38612
rect 29372 38164 29428 38174
rect 29372 38050 29428 38108
rect 29372 37998 29374 38050
rect 29426 37998 29428 38050
rect 29372 37986 29428 37998
rect 29148 37828 29204 37838
rect 29036 37826 29204 37828
rect 29036 37774 29150 37826
rect 29202 37774 29204 37826
rect 29036 37772 29204 37774
rect 29036 37044 29092 37772
rect 29148 37762 29204 37772
rect 29260 37826 29316 37838
rect 29260 37774 29262 37826
rect 29314 37774 29316 37826
rect 29148 37380 29204 37390
rect 29260 37380 29316 37774
rect 29148 37378 29316 37380
rect 29148 37326 29150 37378
rect 29202 37326 29316 37378
rect 29148 37324 29316 37326
rect 29372 37492 29428 37502
rect 29148 37314 29204 37324
rect 29036 36988 29316 37044
rect 28924 36876 29092 36932
rect 28924 34356 28980 34366
rect 28924 34130 28980 34300
rect 28924 34078 28926 34130
rect 28978 34078 28980 34130
rect 28924 34066 28980 34078
rect 29036 32900 29092 36876
rect 29260 36594 29316 36988
rect 29260 36542 29262 36594
rect 29314 36542 29316 36594
rect 29260 36530 29316 36542
rect 29372 36482 29428 37436
rect 29484 37268 29540 38556
rect 29708 38546 29764 38556
rect 29932 38052 29988 40572
rect 30044 39508 30100 39518
rect 30044 38668 30100 39452
rect 30156 39394 30212 39406
rect 30156 39342 30158 39394
rect 30210 39342 30212 39394
rect 30156 39284 30212 39342
rect 30156 39218 30212 39228
rect 30268 38834 30324 44268
rect 30492 44258 30548 44268
rect 30380 43428 30436 43438
rect 30380 41748 30436 43372
rect 30492 41972 30548 41982
rect 30492 41878 30548 41916
rect 30380 41692 30548 41748
rect 30380 41076 30436 41086
rect 30380 40982 30436 41020
rect 30380 40852 30436 40862
rect 30380 39956 30436 40796
rect 30492 40180 30548 41692
rect 30604 40516 30660 49084
rect 30716 48244 30772 49756
rect 30940 48244 30996 48254
rect 30772 48242 30996 48244
rect 30772 48190 30942 48242
rect 30994 48190 30996 48242
rect 30772 48188 30996 48190
rect 30716 48178 30772 48188
rect 30940 48178 30996 48188
rect 31164 47908 31220 49868
rect 31276 48354 31332 50542
rect 31388 49812 31444 49822
rect 31388 49718 31444 49756
rect 31276 48302 31278 48354
rect 31330 48302 31332 48354
rect 31276 48290 31332 48302
rect 31388 49364 31444 49374
rect 31388 48356 31444 49308
rect 31052 47852 31220 47908
rect 30716 47572 30772 47582
rect 30772 47516 30884 47572
rect 30716 47506 30772 47516
rect 30828 47348 30884 47516
rect 31052 47458 31108 47852
rect 31276 47460 31332 47470
rect 31388 47460 31444 48300
rect 31052 47406 31054 47458
rect 31106 47406 31108 47458
rect 31052 47394 31108 47406
rect 31164 47458 31444 47460
rect 31164 47406 31278 47458
rect 31330 47406 31444 47458
rect 31164 47404 31444 47406
rect 30940 47348 30996 47358
rect 30828 47346 30996 47348
rect 30828 47294 30942 47346
rect 30994 47294 30996 47346
rect 30828 47292 30996 47294
rect 30940 47282 30996 47292
rect 31052 45108 31108 45118
rect 31164 45108 31220 47404
rect 31276 47394 31332 47404
rect 31276 47124 31332 47134
rect 31276 46674 31332 47068
rect 31500 46900 31556 51436
rect 31724 51436 31892 51492
rect 31724 49924 31780 51436
rect 31836 51268 31892 51278
rect 31836 51174 31892 51212
rect 31612 49922 31780 49924
rect 31612 49870 31726 49922
rect 31778 49870 31780 49922
rect 31612 49868 31780 49870
rect 31612 49028 31668 49868
rect 31724 49858 31780 49868
rect 31836 50260 31892 50270
rect 31836 49252 31892 50204
rect 31612 48962 31668 48972
rect 31724 49196 31892 49252
rect 31276 46622 31278 46674
rect 31330 46622 31332 46674
rect 31276 45220 31332 46622
rect 31388 46844 31556 46900
rect 31612 48130 31668 48142
rect 31612 48078 31614 48130
rect 31666 48078 31668 48130
rect 31612 47458 31668 48078
rect 31612 47406 31614 47458
rect 31666 47406 31668 47458
rect 31612 47348 31668 47406
rect 31388 45332 31444 46844
rect 31500 46676 31556 46686
rect 31612 46676 31668 47292
rect 31724 46900 31780 49196
rect 31836 47460 31892 47470
rect 31836 47366 31892 47404
rect 31724 46844 31892 46900
rect 31500 46674 31668 46676
rect 31500 46622 31502 46674
rect 31554 46622 31668 46674
rect 31500 46620 31668 46622
rect 31500 46610 31556 46620
rect 31500 45332 31556 45342
rect 31388 45330 31556 45332
rect 31388 45278 31502 45330
rect 31554 45278 31556 45330
rect 31388 45276 31556 45278
rect 31276 45126 31332 45164
rect 31108 45052 31220 45108
rect 30940 44996 30996 45006
rect 30940 43428 30996 44940
rect 30940 43362 30996 43372
rect 30716 42756 30772 42766
rect 30716 42662 30772 42700
rect 31052 42754 31108 45052
rect 31388 44994 31444 45006
rect 31388 44942 31390 44994
rect 31442 44942 31444 44994
rect 31276 44436 31332 44446
rect 31388 44436 31444 44942
rect 31276 44434 31444 44436
rect 31276 44382 31278 44434
rect 31330 44382 31444 44434
rect 31276 44380 31444 44382
rect 31500 44884 31556 45276
rect 31612 45106 31668 45118
rect 31612 45054 31614 45106
rect 31666 45054 31668 45106
rect 31612 44996 31668 45054
rect 31612 44930 31668 44940
rect 31276 44370 31332 44380
rect 31500 43764 31556 44828
rect 31500 43698 31556 43708
rect 31052 42702 31054 42754
rect 31106 42702 31108 42754
rect 31052 42690 31108 42702
rect 31388 42754 31444 42766
rect 31388 42702 31390 42754
rect 31442 42702 31444 42754
rect 31164 42530 31220 42542
rect 31164 42478 31166 42530
rect 31218 42478 31220 42530
rect 30828 42082 30884 42094
rect 30828 42030 30830 42082
rect 30882 42030 30884 42082
rect 30828 41860 30884 42030
rect 30828 41794 30884 41804
rect 30604 40422 30660 40460
rect 30492 40114 30548 40124
rect 30380 39900 30772 39956
rect 30716 39618 30772 39900
rect 31164 39620 31220 42478
rect 31388 42532 31444 42702
rect 31612 42756 31668 42766
rect 31612 42642 31668 42700
rect 31612 42590 31614 42642
rect 31666 42590 31668 42642
rect 31612 42578 31668 42590
rect 31388 42466 31444 42476
rect 31276 41076 31332 41086
rect 31276 39730 31332 41020
rect 31276 39678 31278 39730
rect 31330 39678 31332 39730
rect 31276 39666 31332 39678
rect 31836 39732 31892 46844
rect 31948 46676 32004 55020
rect 32172 54516 32228 54526
rect 32172 53172 32228 54460
rect 32284 53172 32340 53182
rect 32172 53116 32284 53172
rect 32284 53078 32340 53116
rect 32396 52948 32452 52958
rect 32396 52162 32452 52892
rect 32396 52110 32398 52162
rect 32450 52110 32452 52162
rect 32396 52098 32452 52110
rect 32732 52050 32788 52062
rect 32732 51998 32734 52050
rect 32786 51998 32788 52050
rect 32620 51940 32676 51950
rect 32620 51846 32676 51884
rect 32732 51716 32788 51998
rect 32732 51650 32788 51660
rect 32620 49140 32676 49150
rect 32620 49138 32788 49140
rect 32620 49086 32622 49138
rect 32674 49086 32788 49138
rect 32620 49084 32788 49086
rect 32620 49074 32676 49084
rect 32620 48916 32676 48926
rect 32060 48244 32116 48254
rect 32060 48150 32116 48188
rect 32508 48130 32564 48142
rect 32508 48078 32510 48130
rect 32562 48078 32564 48130
rect 32508 47684 32564 48078
rect 32508 47618 32564 47628
rect 32620 47570 32676 48860
rect 32732 48244 32788 49084
rect 32732 48178 32788 48188
rect 32620 47518 32622 47570
rect 32674 47518 32676 47570
rect 32620 47506 32676 47518
rect 32844 47572 32900 56814
rect 32956 57988 33012 57998
rect 32956 50428 33012 57932
rect 33180 57538 33236 58380
rect 33180 57486 33182 57538
rect 33234 57486 33236 57538
rect 33180 57474 33236 57486
rect 33292 57428 33348 58716
rect 33516 58658 33572 58828
rect 33516 58606 33518 58658
rect 33570 58606 33572 58658
rect 33516 58594 33572 58606
rect 33404 58548 33460 58558
rect 33404 58454 33460 58492
rect 33740 58548 33796 59166
rect 33740 58482 33796 58492
rect 33516 57652 33572 57662
rect 33516 57558 33572 57596
rect 33292 57372 33572 57428
rect 33516 56754 33572 57372
rect 33516 56702 33518 56754
rect 33570 56702 33572 56754
rect 33516 56690 33572 56702
rect 33180 56644 33236 56654
rect 33180 56550 33236 56588
rect 33068 56532 33124 56542
rect 33068 56082 33124 56476
rect 33068 56030 33070 56082
rect 33122 56030 33124 56082
rect 33068 56018 33124 56030
rect 33516 56084 33572 56094
rect 33516 55990 33572 56028
rect 33292 55412 33348 55422
rect 33180 55356 33292 55412
rect 33180 53844 33236 55356
rect 33292 55346 33348 55356
rect 33292 54404 33348 54414
rect 33292 54310 33348 54348
rect 33404 54292 33460 54302
rect 33404 54290 33572 54292
rect 33404 54238 33406 54290
rect 33458 54238 33572 54290
rect 33404 54236 33572 54238
rect 33404 54226 33460 54236
rect 33180 53788 33348 53844
rect 33180 53620 33236 53630
rect 33068 53172 33124 53182
rect 33068 53078 33124 53116
rect 33180 51378 33236 53564
rect 33292 52836 33348 53788
rect 33516 53732 33572 54236
rect 33740 53732 33796 53742
rect 33516 53730 33796 53732
rect 33516 53678 33742 53730
rect 33794 53678 33796 53730
rect 33516 53676 33796 53678
rect 33740 53666 33796 53676
rect 33852 53508 33908 61852
rect 34188 61796 34244 61964
rect 34076 61740 34244 61796
rect 34748 61796 34804 62190
rect 35644 62242 35700 62636
rect 36540 62580 36596 62590
rect 36540 62486 36596 62524
rect 35644 62190 35646 62242
rect 35698 62190 35700 62242
rect 35196 61964 35460 61974
rect 35252 61908 35300 61964
rect 35356 61908 35404 61964
rect 35196 61898 35460 61908
rect 33964 61570 34020 61582
rect 33964 61518 33966 61570
rect 34018 61518 34020 61570
rect 33964 61348 34020 61518
rect 33964 58212 34020 61292
rect 34076 58436 34132 61740
rect 34748 61730 34804 61740
rect 34636 61572 34692 61582
rect 35084 61572 35140 61582
rect 34636 61570 35140 61572
rect 34636 61518 34638 61570
rect 34690 61518 35086 61570
rect 35138 61518 35140 61570
rect 34636 61516 35140 61518
rect 34636 61506 34692 61516
rect 34748 60788 34804 60798
rect 34524 60786 34804 60788
rect 34524 60734 34750 60786
rect 34802 60734 34804 60786
rect 34524 60732 34804 60734
rect 34188 59780 34244 59790
rect 34188 59386 34244 59724
rect 34188 59334 34190 59386
rect 34242 59334 34244 59386
rect 34524 59442 34580 60732
rect 34748 60722 34804 60732
rect 34972 60786 35028 60798
rect 34972 60734 34974 60786
rect 35026 60734 35028 60786
rect 34860 60676 34916 60686
rect 34860 60582 34916 60620
rect 34972 60340 35028 60734
rect 34748 60284 35028 60340
rect 34524 59390 34526 59442
rect 34578 59390 34580 59442
rect 34524 59378 34580 59390
rect 34636 60004 34692 60014
rect 34188 59322 34244 59334
rect 34300 59330 34356 59342
rect 34300 59278 34302 59330
rect 34354 59278 34356 59330
rect 34300 59220 34356 59278
rect 34636 59220 34692 59948
rect 34188 59164 34356 59220
rect 34524 59164 34692 59220
rect 34188 58772 34244 59164
rect 34524 58996 34580 59164
rect 34188 58706 34244 58716
rect 34300 58940 34580 58996
rect 34300 58658 34356 58940
rect 34748 58884 34804 60284
rect 34972 60116 35028 60126
rect 35084 60116 35140 61516
rect 35308 61348 35364 61358
rect 35644 61348 35700 62190
rect 36092 62468 36148 62478
rect 36092 62242 36148 62412
rect 36092 62190 36094 62242
rect 36146 62190 36148 62242
rect 35308 61346 35700 61348
rect 35308 61294 35310 61346
rect 35362 61294 35700 61346
rect 35308 61292 35700 61294
rect 35756 61346 35812 61358
rect 35756 61294 35758 61346
rect 35810 61294 35812 61346
rect 35308 60564 35364 61292
rect 35756 61012 35812 61294
rect 35756 60956 36036 61012
rect 35420 60788 35476 60798
rect 35756 60788 35812 60798
rect 35420 60786 35588 60788
rect 35420 60734 35422 60786
rect 35474 60734 35588 60786
rect 35420 60732 35588 60734
rect 35420 60722 35476 60732
rect 35308 60498 35364 60508
rect 35196 60396 35460 60406
rect 35252 60340 35300 60396
rect 35356 60340 35404 60396
rect 35196 60330 35460 60340
rect 34972 60114 35140 60116
rect 34972 60062 34974 60114
rect 35026 60062 35140 60114
rect 34972 60060 35140 60062
rect 35420 60228 35476 60238
rect 34972 60050 35028 60060
rect 34860 59668 34916 59678
rect 34860 59218 34916 59612
rect 34860 59166 34862 59218
rect 34914 59166 34916 59218
rect 34860 58996 34916 59166
rect 34860 58930 34916 58940
rect 35084 59668 35140 59678
rect 34748 58818 34804 58828
rect 34300 58606 34302 58658
rect 34354 58606 34356 58658
rect 34300 58594 34356 58606
rect 34636 58772 34692 58782
rect 34076 58370 34132 58380
rect 34188 58548 34244 58558
rect 34188 58436 34244 58492
rect 34636 58436 34692 58716
rect 34188 58434 34580 58436
rect 34188 58382 34190 58434
rect 34242 58382 34580 58434
rect 34188 58380 34580 58382
rect 34188 58370 34244 58380
rect 34524 58324 34580 58380
rect 34300 58212 34356 58222
rect 33964 58156 34244 58212
rect 34076 57540 34132 57550
rect 33964 56980 34020 56990
rect 33964 56886 34020 56924
rect 33964 56084 34020 56094
rect 33964 55990 34020 56028
rect 33964 55412 34020 55422
rect 33964 55298 34020 55356
rect 33964 55246 33966 55298
rect 34018 55246 34020 55298
rect 33964 55234 34020 55246
rect 34076 55300 34132 57484
rect 34188 55412 34244 58156
rect 34300 58118 34356 58156
rect 34412 56866 34468 56878
rect 34412 56814 34414 56866
rect 34466 56814 34468 56866
rect 34412 56644 34468 56814
rect 34300 56196 34356 56206
rect 34300 56102 34356 56140
rect 34412 56084 34468 56588
rect 34412 56018 34468 56028
rect 34412 55412 34468 55422
rect 34188 55410 34468 55412
rect 34188 55358 34414 55410
rect 34466 55358 34468 55410
rect 34188 55356 34468 55358
rect 34412 55346 34468 55356
rect 34076 55244 34244 55300
rect 34076 54852 34132 54862
rect 34076 54740 34132 54796
rect 33628 53452 33908 53508
rect 33964 54738 34132 54740
rect 33964 54686 34078 54738
rect 34130 54686 34132 54738
rect 33964 54684 34132 54686
rect 33404 53060 33460 53070
rect 33404 52966 33460 53004
rect 33292 52780 33460 52836
rect 33292 52276 33348 52286
rect 33292 52182 33348 52220
rect 33180 51326 33182 51378
rect 33234 51326 33236 51378
rect 33180 51314 33236 51326
rect 33404 50596 33460 52780
rect 33404 50502 33460 50540
rect 33516 52276 33572 52286
rect 33516 52162 33572 52220
rect 33516 52110 33518 52162
rect 33570 52110 33572 52162
rect 32956 50372 33236 50428
rect 33068 48356 33124 48366
rect 33068 48262 33124 48300
rect 32844 47516 33124 47572
rect 32060 47458 32116 47470
rect 32060 47406 32062 47458
rect 32114 47406 32116 47458
rect 32060 47124 32116 47406
rect 32172 47460 32228 47470
rect 32508 47460 32564 47470
rect 32172 47458 32508 47460
rect 32172 47406 32174 47458
rect 32226 47406 32508 47458
rect 32172 47404 32508 47406
rect 32172 47394 32228 47404
rect 32508 47394 32564 47404
rect 32732 47460 32788 47470
rect 32732 47366 32788 47404
rect 32956 47346 33012 47358
rect 32956 47294 32958 47346
rect 33010 47294 33012 47346
rect 32508 47236 32564 47246
rect 32956 47236 33012 47294
rect 32508 47142 32564 47180
rect 32732 47180 33012 47236
rect 32060 47058 32116 47068
rect 32284 46900 32340 46910
rect 32284 46806 32340 46844
rect 32060 46676 32116 46686
rect 31948 46674 32116 46676
rect 31948 46622 32062 46674
rect 32114 46622 32116 46674
rect 31948 46620 32116 46622
rect 32060 46452 32116 46620
rect 32060 46386 32116 46396
rect 31948 45668 32004 45678
rect 31948 45106 32004 45612
rect 32396 45332 32452 45342
rect 32396 45218 32452 45276
rect 32620 45332 32676 45342
rect 32732 45332 32788 47180
rect 32620 45330 32788 45332
rect 32620 45278 32622 45330
rect 32674 45278 32788 45330
rect 32620 45276 32788 45278
rect 32844 47012 32900 47022
rect 32620 45266 32676 45276
rect 32396 45166 32398 45218
rect 32450 45166 32452 45218
rect 31948 45054 31950 45106
rect 32002 45054 32004 45106
rect 31948 45042 32004 45054
rect 32284 45108 32340 45118
rect 32284 45014 32340 45052
rect 32396 44212 32452 45166
rect 32396 44146 32452 44156
rect 32284 43764 32340 43774
rect 32284 43650 32340 43708
rect 32284 43598 32286 43650
rect 32338 43598 32340 43650
rect 32284 43586 32340 43598
rect 32620 43652 32676 43662
rect 32508 42868 32564 42878
rect 32508 42774 32564 42812
rect 31948 42642 32004 42654
rect 31948 42590 31950 42642
rect 32002 42590 32004 42642
rect 31948 41860 32004 42590
rect 31948 41794 32004 41804
rect 32508 41298 32564 41310
rect 32508 41246 32510 41298
rect 32562 41246 32564 41298
rect 32060 40404 32116 40414
rect 31836 39676 32004 39732
rect 30716 39566 30718 39618
rect 30770 39566 30772 39618
rect 30716 39554 30772 39566
rect 31052 39564 31220 39620
rect 31388 39620 31444 39630
rect 30268 38782 30270 38834
rect 30322 38782 30324 38834
rect 30268 38770 30324 38782
rect 30380 39396 30436 39406
rect 30044 38612 30324 38668
rect 30156 38164 30212 38174
rect 29932 37996 30100 38052
rect 29596 37828 29652 37838
rect 29932 37828 29988 37838
rect 29596 37826 29988 37828
rect 29596 37774 29598 37826
rect 29650 37774 29934 37826
rect 29986 37774 29988 37826
rect 29596 37772 29988 37774
rect 29596 37762 29652 37772
rect 29932 37762 29988 37772
rect 29820 37268 29876 37278
rect 29484 37266 29876 37268
rect 29484 37214 29822 37266
rect 29874 37214 29876 37266
rect 29484 37212 29876 37214
rect 29820 37202 29876 37212
rect 29372 36430 29374 36482
rect 29426 36430 29428 36482
rect 29372 36418 29428 36430
rect 29820 36484 29876 36494
rect 29820 36390 29876 36428
rect 29148 36260 29204 36270
rect 29148 36166 29204 36204
rect 29596 35700 29652 35710
rect 29372 35698 29652 35700
rect 29372 35646 29598 35698
rect 29650 35646 29652 35698
rect 29372 35644 29652 35646
rect 29260 34804 29316 34814
rect 29260 34690 29316 34748
rect 29260 34638 29262 34690
rect 29314 34638 29316 34690
rect 29260 33684 29316 34638
rect 29372 34020 29428 35644
rect 29596 35634 29652 35644
rect 30044 35308 30100 37996
rect 30156 37938 30212 38108
rect 30268 38050 30324 38612
rect 30268 37998 30270 38050
rect 30322 37998 30324 38050
rect 30268 37986 30324 37998
rect 30156 37886 30158 37938
rect 30210 37886 30212 37938
rect 30156 37492 30212 37886
rect 30380 37828 30436 39340
rect 30940 39394 30996 39406
rect 30940 39342 30942 39394
rect 30994 39342 30996 39394
rect 30716 39284 30772 39294
rect 30604 38612 30660 38622
rect 30604 38050 30660 38556
rect 30604 37998 30606 38050
rect 30658 37998 30660 38050
rect 30604 37986 30660 37998
rect 30716 37940 30772 39228
rect 30828 38722 30884 38734
rect 30828 38670 30830 38722
rect 30882 38670 30884 38722
rect 30828 38164 30884 38670
rect 30940 38668 30996 39342
rect 31052 38948 31108 39564
rect 31388 39526 31444 39564
rect 31836 39508 31892 39518
rect 31836 39414 31892 39452
rect 31164 39396 31220 39406
rect 31724 39396 31780 39406
rect 31164 39394 31780 39396
rect 31164 39342 31166 39394
rect 31218 39342 31726 39394
rect 31778 39342 31780 39394
rect 31164 39340 31780 39342
rect 31164 39330 31220 39340
rect 31724 39330 31780 39340
rect 31948 39284 32004 39676
rect 31836 39228 32004 39284
rect 31724 39060 31780 39070
rect 31724 38966 31780 39004
rect 31164 38948 31220 38958
rect 31052 38946 31220 38948
rect 31052 38894 31166 38946
rect 31218 38894 31220 38946
rect 31052 38892 31220 38894
rect 31164 38882 31220 38892
rect 31388 38834 31444 38846
rect 31388 38782 31390 38834
rect 31442 38782 31444 38834
rect 31388 38668 31444 38782
rect 31612 38834 31668 38846
rect 31612 38782 31614 38834
rect 31666 38782 31668 38834
rect 30940 38612 31108 38668
rect 30828 38098 30884 38108
rect 30716 37884 30996 37940
rect 30156 37426 30212 37436
rect 30268 37772 30436 37828
rect 30156 37268 30212 37278
rect 30268 37268 30324 37772
rect 30156 37266 30324 37268
rect 30156 37214 30158 37266
rect 30210 37214 30324 37266
rect 30156 37212 30324 37214
rect 30380 37378 30436 37390
rect 30380 37326 30382 37378
rect 30434 37326 30436 37378
rect 30156 37202 30212 37212
rect 30380 36708 30436 37326
rect 30492 37380 30548 37390
rect 30548 37324 30772 37380
rect 30492 37286 30548 37324
rect 30380 36652 30548 36708
rect 30156 36482 30212 36494
rect 30380 36484 30436 36494
rect 30156 36430 30158 36482
rect 30210 36430 30212 36482
rect 30156 36148 30212 36430
rect 30156 36082 30212 36092
rect 30268 36428 30380 36484
rect 30268 35812 30324 36428
rect 30380 36418 30436 36428
rect 30380 36260 30436 36270
rect 30380 36166 30436 36204
rect 30380 35812 30436 35822
rect 30268 35810 30436 35812
rect 30268 35758 30382 35810
rect 30434 35758 30436 35810
rect 30268 35756 30436 35758
rect 30380 35746 30436 35756
rect 29932 35252 30100 35308
rect 29596 34692 29652 34702
rect 29484 34244 29540 34254
rect 29484 34150 29540 34188
rect 29596 34130 29652 34636
rect 29596 34078 29598 34130
rect 29650 34078 29652 34130
rect 29596 34066 29652 34078
rect 29820 34356 29876 34366
rect 29820 34130 29876 34300
rect 29820 34078 29822 34130
rect 29874 34078 29876 34130
rect 29820 34066 29876 34078
rect 29708 34020 29764 34030
rect 29372 33964 29540 34020
rect 29260 33618 29316 33628
rect 29372 33236 29428 33246
rect 29372 33142 29428 33180
rect 29148 33124 29204 33134
rect 29148 33030 29204 33068
rect 29260 33122 29316 33134
rect 29260 33070 29262 33122
rect 29314 33070 29316 33122
rect 28924 32844 29092 32900
rect 28924 32452 28980 32844
rect 29036 32676 29092 32686
rect 29260 32676 29316 33070
rect 29484 33012 29540 33964
rect 29596 33124 29652 33134
rect 29596 33030 29652 33068
rect 29036 32674 29316 32676
rect 29036 32622 29038 32674
rect 29090 32622 29316 32674
rect 29036 32620 29316 32622
rect 29372 32956 29540 33012
rect 29036 32610 29092 32620
rect 28924 32396 29316 32452
rect 29148 31556 29204 31566
rect 28812 30716 29092 30772
rect 28700 30158 28702 30210
rect 28754 30158 28756 30210
rect 28700 30146 28756 30158
rect 28812 30548 28868 30558
rect 28588 28702 28590 28754
rect 28642 28702 28644 28754
rect 28588 28690 28644 28702
rect 27692 28418 27748 28430
rect 27692 28366 27694 28418
rect 27746 28366 27748 28418
rect 27692 28084 27748 28366
rect 28588 28420 28644 28430
rect 27916 28084 27972 28094
rect 27692 28028 27916 28084
rect 27916 27990 27972 28028
rect 27580 27748 27636 27758
rect 27244 27692 27580 27748
rect 27132 27186 27524 27188
rect 27132 27134 27134 27186
rect 27186 27134 27524 27186
rect 27132 27132 27524 27134
rect 27132 27122 27188 27132
rect 27468 27074 27524 27132
rect 27468 27022 27470 27074
rect 27522 27022 27524 27074
rect 27468 27010 27524 27022
rect 27580 26908 27636 27692
rect 28476 27748 28532 27758
rect 28588 27748 28644 28364
rect 28532 27692 28644 27748
rect 28476 27654 28532 27692
rect 27020 26852 27188 26908
rect 27132 26516 27188 26852
rect 27132 25506 27188 26460
rect 27356 26852 27636 26908
rect 27692 27076 27748 27086
rect 27244 26180 27300 26190
rect 27244 26086 27300 26124
rect 27132 25454 27134 25506
rect 27186 25454 27188 25506
rect 27132 25442 27188 25454
rect 27244 24612 27300 24622
rect 27356 24612 27412 26852
rect 27692 26628 27748 27020
rect 27244 24610 27412 24612
rect 27244 24558 27246 24610
rect 27298 24558 27412 24610
rect 27244 24556 27412 24558
rect 27468 26572 27748 26628
rect 28028 27074 28084 27086
rect 28028 27022 28030 27074
rect 28082 27022 28084 27074
rect 28028 26628 28084 27022
rect 27468 25394 27524 26572
rect 28028 26562 28084 26572
rect 28140 26964 28196 26974
rect 28812 26908 28868 30492
rect 29036 29876 29092 30716
rect 29148 30210 29204 31500
rect 29148 30158 29150 30210
rect 29202 30158 29204 30210
rect 29148 30146 29204 30158
rect 29036 29810 29092 29820
rect 29260 29652 29316 32396
rect 29372 32004 29428 32956
rect 29708 32676 29764 33964
rect 29372 31938 29428 31948
rect 29596 32620 29764 32676
rect 29932 32676 29988 35252
rect 30268 35028 30324 35038
rect 30044 33348 30100 33358
rect 30044 33254 30100 33292
rect 30156 33122 30212 33134
rect 30156 33070 30158 33122
rect 30210 33070 30212 33122
rect 30156 32788 30212 33070
rect 30156 32722 30212 32732
rect 29932 32620 30100 32676
rect 29484 31892 29540 31902
rect 29372 31780 29428 31790
rect 29372 31686 29428 31724
rect 29036 29596 29316 29652
rect 29372 31556 29428 31566
rect 29036 28308 29092 29596
rect 29260 29428 29316 29438
rect 29260 28866 29316 29372
rect 29260 28814 29262 28866
rect 29314 28814 29316 28866
rect 29260 28802 29316 28814
rect 29148 28532 29204 28542
rect 29148 28438 29204 28476
rect 29260 28420 29316 28430
rect 29260 28326 29316 28364
rect 29036 28252 29204 28308
rect 27468 25342 27470 25394
rect 27522 25342 27524 25394
rect 26908 23492 27076 23548
rect 26908 23044 26964 23054
rect 26908 22594 26964 22988
rect 27020 22820 27076 23492
rect 27132 23156 27188 23194
rect 27132 23090 27188 23100
rect 27244 23044 27300 24556
rect 27468 23492 27524 25342
rect 27468 23426 27524 23436
rect 27580 26404 27636 26414
rect 28140 26404 28196 26908
rect 27580 26180 27636 26348
rect 27916 26348 28196 26404
rect 28700 26852 28868 26908
rect 29036 27860 29092 27870
rect 27692 26180 27748 26190
rect 27580 26178 27748 26180
rect 27580 26126 27694 26178
rect 27746 26126 27748 26178
rect 27580 26124 27748 26126
rect 27356 23380 27412 23390
rect 27356 23268 27412 23324
rect 27468 23268 27524 23278
rect 27356 23266 27524 23268
rect 27356 23214 27470 23266
rect 27522 23214 27524 23266
rect 27356 23212 27524 23214
rect 27580 23268 27636 26124
rect 27692 26114 27748 26124
rect 27692 25508 27748 25518
rect 27692 24050 27748 25452
rect 27692 23998 27694 24050
rect 27746 23998 27748 24050
rect 27692 23986 27748 23998
rect 27692 23268 27748 23278
rect 27580 23212 27692 23268
rect 27468 23202 27524 23212
rect 27692 23202 27748 23212
rect 27804 23266 27860 23278
rect 27804 23214 27806 23266
rect 27858 23214 27860 23266
rect 27244 22978 27300 22988
rect 27804 23156 27860 23214
rect 27132 22820 27188 22830
rect 27020 22764 27132 22820
rect 27132 22754 27188 22764
rect 26908 22542 26910 22594
rect 26962 22542 26964 22594
rect 26908 22530 26964 22542
rect 26796 22418 26852 22428
rect 27692 22372 27748 22382
rect 26684 21410 26740 21420
rect 26908 22316 27188 22372
rect 26796 21364 26852 21374
rect 26908 21364 26964 22316
rect 27132 22258 27188 22316
rect 27692 22278 27748 22316
rect 27132 22206 27134 22258
rect 27186 22206 27188 22258
rect 27132 22194 27188 22206
rect 27020 22146 27076 22158
rect 27020 22094 27022 22146
rect 27074 22094 27076 22146
rect 27020 21700 27076 22094
rect 27020 21634 27076 21644
rect 27244 21924 27300 21934
rect 27244 21586 27300 21868
rect 27804 21924 27860 23100
rect 27804 21858 27860 21868
rect 27916 21700 27972 26348
rect 28588 26292 28644 26302
rect 28252 26290 28644 26292
rect 28252 26238 28590 26290
rect 28642 26238 28644 26290
rect 28252 26236 28644 26238
rect 28140 26178 28196 26190
rect 28140 26126 28142 26178
rect 28194 26126 28196 26178
rect 28140 25844 28196 26126
rect 28140 25778 28196 25788
rect 28140 25508 28196 25518
rect 28252 25508 28308 26236
rect 28588 26226 28644 26236
rect 28196 25452 28308 25508
rect 28140 25414 28196 25452
rect 28364 25396 28420 25406
rect 28420 25340 28644 25396
rect 28364 25302 28420 25340
rect 28252 24052 28308 24062
rect 28252 23958 28308 23996
rect 28588 24050 28644 25340
rect 28588 23998 28590 24050
rect 28642 23998 28644 24050
rect 28588 23828 28644 23998
rect 28588 23548 28644 23772
rect 28252 23492 28308 23502
rect 28140 22484 28196 22494
rect 28140 22390 28196 22428
rect 27244 21534 27246 21586
rect 27298 21534 27300 21586
rect 26796 21362 26964 21364
rect 26796 21310 26798 21362
rect 26850 21310 26964 21362
rect 26796 21308 26964 21310
rect 27020 21476 27076 21486
rect 26236 21196 26740 21252
rect 25788 19852 25956 19908
rect 26460 20690 26516 20702
rect 26460 20638 26462 20690
rect 26514 20638 26516 20690
rect 25340 19292 25508 19348
rect 25676 19348 25732 19358
rect 25340 18676 25396 19292
rect 25564 19236 25620 19246
rect 25676 19236 25732 19292
rect 25564 19234 25732 19236
rect 25564 19182 25566 19234
rect 25618 19182 25732 19234
rect 25564 19180 25732 19182
rect 25564 19170 25620 19180
rect 25452 19124 25508 19134
rect 25452 19030 25508 19068
rect 25676 19012 25732 19022
rect 25676 18918 25732 18956
rect 25340 18620 25508 18676
rect 24668 18562 24948 18564
rect 24668 18510 24670 18562
rect 24722 18510 24948 18562
rect 24668 18508 24948 18510
rect 24668 18498 24724 18508
rect 23996 17948 24500 18004
rect 23884 17714 23940 17724
rect 23548 17388 23716 17444
rect 23548 17220 23604 17230
rect 23548 16994 23604 17164
rect 23548 16942 23550 16994
rect 23602 16942 23604 16994
rect 23548 16930 23604 16942
rect 23660 16772 23716 17388
rect 24108 17220 24164 17948
rect 24108 17154 24164 17164
rect 24220 17778 24276 17790
rect 24220 17726 24222 17778
rect 24274 17726 24276 17778
rect 24220 17668 24276 17726
rect 24780 17668 24836 17678
rect 24220 17666 24836 17668
rect 24220 17614 24782 17666
rect 24834 17614 24836 17666
rect 24220 17612 24836 17614
rect 23884 16884 23940 16894
rect 24220 16884 24276 17612
rect 24780 17602 24836 17612
rect 24556 17444 24612 17454
rect 24892 17444 24948 18508
rect 24332 17442 24948 17444
rect 24332 17390 24558 17442
rect 24610 17390 24948 17442
rect 24332 17388 24948 17390
rect 25004 18228 25060 18238
rect 24332 17106 24388 17388
rect 24556 17378 24612 17388
rect 24332 17054 24334 17106
rect 24386 17054 24388 17106
rect 24332 17042 24388 17054
rect 24444 17220 24500 17230
rect 24444 16994 24500 17164
rect 24444 16942 24446 16994
rect 24498 16942 24500 16994
rect 24444 16930 24500 16942
rect 23884 16882 24276 16884
rect 23884 16830 23886 16882
rect 23938 16830 24276 16882
rect 23884 16828 24276 16830
rect 23884 16818 23940 16828
rect 23660 16706 23716 16716
rect 23884 16658 23940 16670
rect 23884 16606 23886 16658
rect 23938 16606 23940 16658
rect 23660 16098 23716 16110
rect 23660 16046 23662 16098
rect 23714 16046 23716 16098
rect 23660 15540 23716 16046
rect 23884 16098 23940 16606
rect 24332 16660 24388 16670
rect 24780 16660 24836 16670
rect 24332 16658 24612 16660
rect 24332 16606 24334 16658
rect 24386 16606 24612 16658
rect 24332 16604 24612 16606
rect 24332 16594 24388 16604
rect 23884 16046 23886 16098
rect 23938 16046 23940 16098
rect 23884 16034 23940 16046
rect 24556 16098 24612 16604
rect 24556 16046 24558 16098
rect 24610 16046 24612 16098
rect 24556 16034 24612 16046
rect 23660 15474 23716 15484
rect 23772 15986 23828 15998
rect 23772 15934 23774 15986
rect 23826 15934 23828 15986
rect 23324 15250 23380 15260
rect 23772 15314 23828 15934
rect 23772 15262 23774 15314
rect 23826 15262 23828 15314
rect 23548 15202 23604 15214
rect 23548 15150 23550 15202
rect 23602 15150 23604 15202
rect 23212 15092 23268 15102
rect 23212 14998 23268 15036
rect 23548 14756 23604 15150
rect 23772 14980 23828 15262
rect 23772 14914 23828 14924
rect 23884 15540 23940 15550
rect 23548 14690 23604 14700
rect 23100 14590 23102 14642
rect 23154 14590 23156 14642
rect 22988 12964 23044 12974
rect 22988 12870 23044 12908
rect 23100 12292 23156 14590
rect 23884 14642 23940 15484
rect 24668 15540 24724 15550
rect 24108 15314 24164 15326
rect 24108 15262 24110 15314
rect 24162 15262 24164 15314
rect 24108 14756 24164 15262
rect 24332 15316 24388 15326
rect 24332 15314 24500 15316
rect 24332 15262 24334 15314
rect 24386 15262 24500 15314
rect 24332 15260 24500 15262
rect 24332 15250 24388 15260
rect 24108 14690 24164 14700
rect 24220 15202 24276 15214
rect 24220 15150 24222 15202
rect 24274 15150 24276 15202
rect 23884 14590 23886 14642
rect 23938 14590 23940 14642
rect 23884 14578 23940 14590
rect 24108 14532 24164 14542
rect 24220 14532 24276 15150
rect 24108 14530 24276 14532
rect 24108 14478 24110 14530
rect 24162 14478 24276 14530
rect 24108 14476 24276 14478
rect 24332 15092 24388 15102
rect 24332 14530 24388 15036
rect 24332 14478 24334 14530
rect 24386 14478 24388 14530
rect 24108 14466 24164 14476
rect 24332 14466 24388 14478
rect 24444 14980 24500 15260
rect 24668 15314 24724 15484
rect 24668 15262 24670 15314
rect 24722 15262 24724 15314
rect 24668 15250 24724 15262
rect 24444 14420 24500 14924
rect 24780 14530 24836 16604
rect 25004 15148 25060 18172
rect 25228 17108 25284 18620
rect 25340 18338 25396 18350
rect 25340 18286 25342 18338
rect 25394 18286 25396 18338
rect 25340 18228 25396 18286
rect 25340 18162 25396 18172
rect 25340 17780 25396 17790
rect 25340 17686 25396 17724
rect 25340 17108 25396 17118
rect 25228 17106 25396 17108
rect 25228 17054 25342 17106
rect 25394 17054 25396 17106
rect 25228 17052 25396 17054
rect 25228 15540 25284 17052
rect 25340 17042 25396 17052
rect 25452 16994 25508 18620
rect 25788 18450 25844 19852
rect 26012 19460 26068 19470
rect 26012 19234 26068 19404
rect 26460 19348 26516 20638
rect 26460 19282 26516 19292
rect 26012 19182 26014 19234
rect 26066 19182 26068 19234
rect 26012 19170 26068 19182
rect 26124 19012 26180 19022
rect 26124 18918 26180 18956
rect 26236 19010 26292 19022
rect 26236 18958 26238 19010
rect 26290 18958 26292 19010
rect 25788 18398 25790 18450
rect 25842 18398 25844 18450
rect 25788 18228 25844 18398
rect 25788 18162 25844 18172
rect 25900 18676 25956 18686
rect 25900 18004 25956 18620
rect 26236 18564 26292 18958
rect 26460 19012 26516 19022
rect 26460 18918 26516 18956
rect 26236 18498 26292 18508
rect 25452 16942 25454 16994
rect 25506 16942 25508 16994
rect 25340 16660 25396 16670
rect 25340 16566 25396 16604
rect 25340 16212 25396 16222
rect 25452 16212 25508 16942
rect 25788 17948 25956 18004
rect 25340 16210 25732 16212
rect 25340 16158 25342 16210
rect 25394 16158 25732 16210
rect 25340 16156 25732 16158
rect 25340 16146 25396 16156
rect 25452 15988 25508 15998
rect 25340 15540 25396 15550
rect 25228 15538 25396 15540
rect 25228 15486 25342 15538
rect 25394 15486 25396 15538
rect 25228 15484 25396 15486
rect 25340 15474 25396 15484
rect 25228 15316 25284 15326
rect 25228 15222 25284 15260
rect 24780 14478 24782 14530
rect 24834 14478 24836 14530
rect 24780 14466 24836 14478
rect 24892 15092 25060 15148
rect 24444 14354 24500 14364
rect 24220 14308 24276 14318
rect 24220 14214 24276 14252
rect 24668 13748 24724 13758
rect 24668 13636 24724 13692
rect 24668 13634 24836 13636
rect 24668 13582 24670 13634
rect 24722 13582 24836 13634
rect 24668 13580 24836 13582
rect 24668 13570 24724 13580
rect 24444 13186 24500 13198
rect 24444 13134 24446 13186
rect 24498 13134 24500 13186
rect 23660 12962 23716 12974
rect 23660 12910 23662 12962
rect 23714 12910 23716 12962
rect 23100 12226 23156 12236
rect 23436 12852 23492 12862
rect 22652 11506 22932 11508
rect 22652 11454 22654 11506
rect 22706 11454 22932 11506
rect 22652 11452 22932 11454
rect 22652 11442 22708 11452
rect 22876 11396 22932 11452
rect 23324 11396 23380 11406
rect 22876 11394 23380 11396
rect 22876 11342 23326 11394
rect 23378 11342 23380 11394
rect 22876 11340 23380 11342
rect 23324 11330 23380 11340
rect 22428 11228 23156 11284
rect 21868 10612 21924 11228
rect 23100 11170 23156 11228
rect 23100 11118 23102 11170
rect 23154 11118 23156 11170
rect 23100 11106 23156 11118
rect 21868 10610 22260 10612
rect 21868 10558 21870 10610
rect 21922 10558 22260 10610
rect 21868 10556 22260 10558
rect 21868 10546 21924 10556
rect 22204 9826 22260 10556
rect 22540 10500 22596 10510
rect 22540 10498 22932 10500
rect 22540 10446 22542 10498
rect 22594 10446 22932 10498
rect 22540 10444 22932 10446
rect 22540 10434 22596 10444
rect 22204 9774 22206 9826
rect 22258 9774 22260 9826
rect 22204 9762 22260 9774
rect 21644 9604 21700 9614
rect 21420 9548 21644 9604
rect 21644 9510 21700 9548
rect 22876 9266 22932 10444
rect 22988 9716 23044 9726
rect 22988 9622 23044 9660
rect 22876 9214 22878 9266
rect 22930 9214 22932 9266
rect 22876 9202 22932 9214
rect 22988 9156 23044 9166
rect 22988 9062 23044 9100
rect 23436 9042 23492 12796
rect 23436 8990 23438 9042
rect 23490 8990 23492 9042
rect 22988 8932 23044 8942
rect 21420 3444 21476 3454
rect 21308 3442 21476 3444
rect 21308 3390 21422 3442
rect 21474 3390 21476 3442
rect 21308 3388 21476 3390
rect 20860 800 20916 3388
rect 21084 3378 21140 3388
rect 21420 3378 21476 3388
rect 21868 3444 21924 3454
rect 21868 3350 21924 3388
rect 22988 3442 23044 8876
rect 23436 8932 23492 8990
rect 23436 8866 23492 8876
rect 23548 4226 23604 4238
rect 23548 4174 23550 4226
rect 23602 4174 23604 4226
rect 22988 3390 22990 3442
rect 23042 3390 23044 3442
rect 22988 3378 23044 3390
rect 23212 3556 23268 3566
rect 23548 3556 23604 4174
rect 23212 3554 23604 3556
rect 23212 3502 23214 3554
rect 23266 3502 23604 3554
rect 23212 3500 23604 3502
rect 23212 2548 23268 3500
rect 23660 3442 23716 12910
rect 23996 12964 24052 12974
rect 23772 12292 23828 12302
rect 23772 12178 23828 12236
rect 23996 12290 24052 12908
rect 23996 12238 23998 12290
rect 24050 12238 24052 12290
rect 23996 12226 24052 12238
rect 24108 12962 24164 12974
rect 24108 12910 24110 12962
rect 24162 12910 24164 12962
rect 23772 12126 23774 12178
rect 23826 12126 23828 12178
rect 23772 12114 23828 12126
rect 24108 11844 24164 12910
rect 24108 11778 24164 11788
rect 24444 11060 24500 13134
rect 24668 12962 24724 12974
rect 24668 12910 24670 12962
rect 24722 12910 24724 12962
rect 24668 12180 24724 12910
rect 24780 12402 24836 13580
rect 24780 12350 24782 12402
rect 24834 12350 24836 12402
rect 24780 12338 24836 12350
rect 24668 11508 24724 12124
rect 24444 11004 24612 11060
rect 24444 9716 24500 9726
rect 24444 9266 24500 9660
rect 24444 9214 24446 9266
rect 24498 9214 24500 9266
rect 24444 9202 24500 9214
rect 24556 9154 24612 11004
rect 24668 10498 24724 11452
rect 24668 10446 24670 10498
rect 24722 10446 24724 10498
rect 24668 10434 24724 10446
rect 24556 9102 24558 9154
rect 24610 9102 24612 9154
rect 24556 9090 24612 9102
rect 23884 9044 23940 9054
rect 23884 8950 23940 8988
rect 24220 8932 24276 8942
rect 24220 8370 24276 8876
rect 24220 8318 24222 8370
rect 24274 8318 24276 8370
rect 24220 8306 24276 8318
rect 24332 4226 24388 4238
rect 24332 4174 24334 4226
rect 24386 4174 24388 4226
rect 24220 4114 24276 4126
rect 24220 4062 24222 4114
rect 24274 4062 24276 4114
rect 23660 3390 23662 3442
rect 23714 3390 23716 3442
rect 23660 3378 23716 3390
rect 23884 3556 23940 3566
rect 24220 3556 24276 4062
rect 23884 3554 24276 3556
rect 23884 3502 23886 3554
rect 23938 3502 24276 3554
rect 23884 3500 24276 3502
rect 23884 2548 23940 3500
rect 24332 3444 24388 4174
rect 24668 4226 24724 4238
rect 24668 4174 24670 4226
rect 24722 4174 24724 4226
rect 24668 4114 24724 4174
rect 24668 4062 24670 4114
rect 24722 4062 24724 4114
rect 24668 4050 24724 4062
rect 24556 3444 24612 3454
rect 24332 3442 24612 3444
rect 24332 3390 24558 3442
rect 24610 3390 24612 3442
rect 24332 3388 24612 3390
rect 24556 2548 24612 3388
rect 24892 3442 24948 15092
rect 25228 14756 25284 14766
rect 25228 14530 25284 14700
rect 25452 14642 25508 15932
rect 25676 15876 25732 16156
rect 25788 16098 25844 17948
rect 26460 16772 26516 16782
rect 25900 16660 25956 16670
rect 26236 16660 26292 16670
rect 25900 16658 26068 16660
rect 25900 16606 25902 16658
rect 25954 16606 26068 16658
rect 25900 16604 26068 16606
rect 25900 16594 25956 16604
rect 25788 16046 25790 16098
rect 25842 16046 25844 16098
rect 25788 16034 25844 16046
rect 25676 15820 25956 15876
rect 25564 15316 25620 15326
rect 25788 15316 25844 15326
rect 25564 15314 25844 15316
rect 25564 15262 25566 15314
rect 25618 15262 25790 15314
rect 25842 15262 25844 15314
rect 25564 15260 25844 15262
rect 25564 15250 25620 15260
rect 25788 15250 25844 15260
rect 25676 15092 25732 15102
rect 25452 14590 25454 14642
rect 25506 14590 25508 14642
rect 25452 14578 25508 14590
rect 25564 15036 25676 15092
rect 25228 14478 25230 14530
rect 25282 14478 25284 14530
rect 25116 14420 25172 14430
rect 25116 14326 25172 14364
rect 25228 13858 25284 14478
rect 25564 14084 25620 15036
rect 25676 15026 25732 15036
rect 25788 14420 25844 14430
rect 25228 13806 25230 13858
rect 25282 13806 25284 13858
rect 25228 13794 25284 13806
rect 25452 14028 25620 14084
rect 25676 14364 25788 14420
rect 25340 13748 25396 13758
rect 25340 13636 25396 13692
rect 25228 13580 25396 13636
rect 25004 12962 25060 12974
rect 25004 12910 25006 12962
rect 25058 12910 25060 12962
rect 25004 12292 25060 12910
rect 25228 12402 25284 13580
rect 25340 12964 25396 12974
rect 25340 12870 25396 12908
rect 25452 12962 25508 14028
rect 25452 12910 25454 12962
rect 25506 12910 25508 12962
rect 25452 12404 25508 12910
rect 25228 12350 25230 12402
rect 25282 12350 25284 12402
rect 25228 12338 25284 12350
rect 25340 12348 25508 12404
rect 25004 11172 25060 12236
rect 25004 9044 25060 11116
rect 25228 11844 25284 11854
rect 25116 10052 25172 10062
rect 25116 9938 25172 9996
rect 25116 9886 25118 9938
rect 25170 9886 25172 9938
rect 25116 9874 25172 9886
rect 25228 9156 25284 11788
rect 25340 11508 25396 12348
rect 25452 12180 25508 12190
rect 25452 12086 25508 12124
rect 25564 12068 25620 12078
rect 25676 12068 25732 14364
rect 25788 14354 25844 14364
rect 25900 13748 25956 15820
rect 26012 15764 26068 16604
rect 26236 16566 26292 16604
rect 26460 16212 26516 16716
rect 26236 16156 26516 16212
rect 26236 15988 26292 16156
rect 26460 15988 26516 15998
rect 26236 15922 26292 15932
rect 26348 15986 26516 15988
rect 26348 15934 26462 15986
rect 26514 15934 26516 15986
rect 26348 15932 26516 15934
rect 26012 15708 26292 15764
rect 26236 15538 26292 15708
rect 26236 15486 26238 15538
rect 26290 15486 26292 15538
rect 26236 15474 26292 15486
rect 26348 15538 26404 15932
rect 26460 15922 26516 15932
rect 26572 15988 26628 15998
rect 26348 15486 26350 15538
rect 26402 15486 26404 15538
rect 26348 15474 26404 15486
rect 26460 15540 26516 15550
rect 26572 15540 26628 15932
rect 26460 15538 26628 15540
rect 26460 15486 26462 15538
rect 26514 15486 26628 15538
rect 26460 15484 26628 15486
rect 26460 15474 26516 15484
rect 26124 14532 26180 14542
rect 26460 14532 26516 14542
rect 26124 14530 26516 14532
rect 26124 14478 26126 14530
rect 26178 14478 26462 14530
rect 26514 14478 26516 14530
rect 26124 14476 26516 14478
rect 26124 14466 26180 14476
rect 26460 14466 26516 14476
rect 26572 14420 26628 14430
rect 26572 14326 26628 14364
rect 25900 13654 25956 13692
rect 26348 13748 26404 13758
rect 26012 13634 26068 13646
rect 26012 13582 26014 13634
rect 26066 13582 26068 13634
rect 26012 13300 26068 13582
rect 26012 13244 26292 13300
rect 26236 12962 26292 13244
rect 26236 12910 26238 12962
rect 26290 12910 26292 12962
rect 26236 12898 26292 12910
rect 25564 12066 25732 12068
rect 25564 12014 25566 12066
rect 25618 12014 25732 12066
rect 25564 12012 25732 12014
rect 25788 12178 25844 12190
rect 25788 12126 25790 12178
rect 25842 12126 25844 12178
rect 25788 12068 25844 12126
rect 26124 12068 26180 12078
rect 25788 12012 26124 12068
rect 25564 12002 25620 12012
rect 26124 11974 26180 12012
rect 26348 11956 26404 13692
rect 26684 13300 26740 21196
rect 26796 20468 26852 21308
rect 26796 20402 26852 20412
rect 27020 19460 27076 21420
rect 27244 20802 27300 21534
rect 27244 20750 27246 20802
rect 27298 20750 27300 20802
rect 27244 19908 27300 20750
rect 27804 21644 27972 21700
rect 27804 20804 27860 21644
rect 27916 21476 27972 21486
rect 27916 21474 28196 21476
rect 27916 21422 27918 21474
rect 27970 21422 28196 21474
rect 27916 21420 28196 21422
rect 27916 21410 27972 21420
rect 28140 20914 28196 21420
rect 28252 21028 28308 23436
rect 28476 23492 28644 23548
rect 28364 23268 28420 23278
rect 28364 23174 28420 23212
rect 28252 20972 28420 21028
rect 28140 20862 28142 20914
rect 28194 20862 28196 20914
rect 28140 20850 28196 20862
rect 28252 20804 28308 20814
rect 27804 20748 27972 20804
rect 27804 20580 27860 20590
rect 27804 20486 27860 20524
rect 27692 19908 27748 19918
rect 27300 19852 27412 19908
rect 27244 19842 27300 19852
rect 27244 19460 27300 19470
rect 27020 19404 27244 19460
rect 27244 19366 27300 19404
rect 26908 19124 26964 19134
rect 26908 19030 26964 19068
rect 27356 18676 27412 19852
rect 27692 19814 27748 19852
rect 27692 19460 27748 19470
rect 27356 18610 27412 18620
rect 27468 19236 27524 19246
rect 26908 18564 26964 18574
rect 26908 17106 26964 18508
rect 27468 18564 27524 19180
rect 27692 19234 27748 19404
rect 27692 19182 27694 19234
rect 27746 19182 27748 19234
rect 27692 19170 27748 19182
rect 27804 19012 27860 19022
rect 27804 18676 27860 18956
rect 27916 18788 27972 20748
rect 28252 20710 28308 20748
rect 28028 20578 28084 20590
rect 28028 20526 28030 20578
rect 28082 20526 28084 20578
rect 28028 19010 28084 20526
rect 28252 20468 28308 20478
rect 28140 19236 28196 19246
rect 28140 19142 28196 19180
rect 28252 19234 28308 20412
rect 28252 19182 28254 19234
rect 28306 19182 28308 19234
rect 28252 19170 28308 19182
rect 28028 18958 28030 19010
rect 28082 18958 28084 19010
rect 28028 18946 28084 18958
rect 27916 18732 28308 18788
rect 27804 18610 27860 18620
rect 27468 18498 27524 18508
rect 28140 18564 28196 18574
rect 26908 17054 26910 17106
rect 26962 17054 26964 17106
rect 26908 17042 26964 17054
rect 27468 17052 28084 17108
rect 26796 16882 26852 16894
rect 26796 16830 26798 16882
rect 26850 16830 26852 16882
rect 26796 16660 26852 16830
rect 27020 16882 27076 16894
rect 27020 16830 27022 16882
rect 27074 16830 27076 16882
rect 27020 16772 27076 16830
rect 27468 16882 27524 17052
rect 27468 16830 27470 16882
rect 27522 16830 27524 16882
rect 27468 16818 27524 16830
rect 27692 16882 27748 16894
rect 27692 16830 27694 16882
rect 27746 16830 27748 16882
rect 27020 16706 27076 16716
rect 26796 15426 26852 16604
rect 27692 16660 27748 16830
rect 27916 16882 27972 16894
rect 27916 16830 27918 16882
rect 27970 16830 27972 16882
rect 27692 16594 27748 16604
rect 27804 16770 27860 16782
rect 27804 16718 27806 16770
rect 27858 16718 27860 16770
rect 27804 15988 27860 16718
rect 27916 16772 27972 16830
rect 27916 16706 27972 16716
rect 27804 15922 27860 15932
rect 26796 15374 26798 15426
rect 26850 15374 26852 15426
rect 26796 15362 26852 15374
rect 27692 15876 27748 15886
rect 27244 15316 27300 15326
rect 27132 14644 27188 14654
rect 27244 14644 27300 15260
rect 27692 15314 27748 15820
rect 28028 15538 28084 17052
rect 28140 17106 28196 18508
rect 28252 17890 28308 18732
rect 28252 17838 28254 17890
rect 28306 17838 28308 17890
rect 28252 17778 28308 17838
rect 28252 17726 28254 17778
rect 28306 17726 28308 17778
rect 28252 17714 28308 17726
rect 28364 17780 28420 20972
rect 28364 17714 28420 17724
rect 28476 17556 28532 23492
rect 28588 22146 28644 22158
rect 28588 22094 28590 22146
rect 28642 22094 28644 22146
rect 28588 21812 28644 22094
rect 28588 20804 28644 21756
rect 28700 21588 28756 26852
rect 28924 26516 28980 26526
rect 29036 26516 29092 27804
rect 29148 26908 29204 28252
rect 29372 28196 29428 31500
rect 29484 30322 29540 31836
rect 29484 30270 29486 30322
rect 29538 30270 29540 30322
rect 29484 30258 29540 30270
rect 29484 29540 29540 29550
rect 29484 29314 29540 29484
rect 29484 29262 29486 29314
rect 29538 29262 29540 29314
rect 29484 29250 29540 29262
rect 29260 28140 29428 28196
rect 29260 27074 29316 28140
rect 29484 28084 29540 28094
rect 29372 28028 29484 28084
rect 29372 27970 29428 28028
rect 29484 28018 29540 28028
rect 29372 27918 29374 27970
rect 29426 27918 29428 27970
rect 29372 27906 29428 27918
rect 29260 27022 29262 27074
rect 29314 27022 29316 27074
rect 29260 27010 29316 27022
rect 29596 26908 29652 32620
rect 29820 32564 29876 32574
rect 29820 32562 29988 32564
rect 29820 32510 29822 32562
rect 29874 32510 29988 32562
rect 29820 32508 29988 32510
rect 29820 32498 29876 32508
rect 29932 32004 29988 32508
rect 29932 31666 29988 31948
rect 29932 31614 29934 31666
rect 29986 31614 29988 31666
rect 29932 31556 29988 31614
rect 29932 31490 29988 31500
rect 29820 30322 29876 30334
rect 29820 30270 29822 30322
rect 29874 30270 29876 30322
rect 29820 29988 29876 30270
rect 29820 29538 29876 29932
rect 30044 29652 30100 32620
rect 30268 31780 30324 34972
rect 30380 33124 30436 33134
rect 30380 33030 30436 33068
rect 30268 31714 30324 31724
rect 30380 32564 30436 32574
rect 30268 30212 30324 30222
rect 30268 30118 30324 30156
rect 30044 29596 30324 29652
rect 29820 29486 29822 29538
rect 29874 29486 29876 29538
rect 29820 29474 29876 29486
rect 30044 29428 30100 29438
rect 30044 29334 30100 29372
rect 29932 29316 29988 29326
rect 29820 28756 29876 28766
rect 29820 28196 29876 28700
rect 29932 28530 29988 29260
rect 29932 28478 29934 28530
rect 29986 28478 29988 28530
rect 29932 28466 29988 28478
rect 30044 28418 30100 28430
rect 30044 28366 30046 28418
rect 30098 28366 30100 28418
rect 29820 28140 29988 28196
rect 29708 28084 29764 28094
rect 29708 27970 29764 28028
rect 29708 27918 29710 27970
rect 29762 27918 29764 27970
rect 29708 27906 29764 27918
rect 29820 27972 29876 27982
rect 29820 27878 29876 27916
rect 29820 27636 29876 27646
rect 29932 27636 29988 28140
rect 29820 27634 29988 27636
rect 29820 27582 29822 27634
rect 29874 27582 29988 27634
rect 29820 27580 29988 27582
rect 29820 27570 29876 27580
rect 29932 27188 29988 27198
rect 30044 27188 30100 28366
rect 30156 28420 30212 28430
rect 30156 28326 30212 28364
rect 30268 28082 30324 29596
rect 30268 28030 30270 28082
rect 30322 28030 30324 28082
rect 29932 27186 30100 27188
rect 29932 27134 29934 27186
rect 29986 27134 30100 27186
rect 29932 27132 30100 27134
rect 30156 27972 30212 27982
rect 29932 27122 29988 27132
rect 29148 26852 29316 26908
rect 29596 26852 29764 26908
rect 28924 26514 29092 26516
rect 28924 26462 28926 26514
rect 28978 26462 29092 26514
rect 28924 26460 29092 26462
rect 28924 26450 28980 26460
rect 29260 26404 29316 26852
rect 29260 26338 29316 26348
rect 29036 24612 29092 24622
rect 29484 24612 29540 24622
rect 28924 23044 28980 23054
rect 28924 22950 28980 22988
rect 29036 21812 29092 24556
rect 29260 24610 29540 24612
rect 29260 24558 29486 24610
rect 29538 24558 29540 24610
rect 29260 24556 29540 24558
rect 29260 24162 29316 24556
rect 29484 24546 29540 24556
rect 29260 24110 29262 24162
rect 29314 24110 29316 24162
rect 29260 24098 29316 24110
rect 29148 23826 29204 23838
rect 29148 23774 29150 23826
rect 29202 23774 29204 23826
rect 29148 22036 29204 23774
rect 29596 23828 29652 23838
rect 29596 23734 29652 23772
rect 29148 21970 29204 21980
rect 29036 21756 29204 21812
rect 28700 21532 28868 21588
rect 28588 20738 28644 20748
rect 28700 21364 28756 21374
rect 28700 20802 28756 21308
rect 28700 20750 28702 20802
rect 28754 20750 28756 20802
rect 28700 20738 28756 20750
rect 28812 18788 28868 21532
rect 28812 18722 28868 18732
rect 28924 20692 28980 20702
rect 28588 18338 28644 18350
rect 28588 18286 28590 18338
rect 28642 18286 28644 18338
rect 28588 18228 28644 18286
rect 28588 18162 28644 18172
rect 28140 17054 28142 17106
rect 28194 17054 28196 17106
rect 28140 17042 28196 17054
rect 28252 17500 28532 17556
rect 28588 17890 28644 17902
rect 28588 17838 28590 17890
rect 28642 17838 28644 17890
rect 28028 15486 28030 15538
rect 28082 15486 28084 15538
rect 28028 15474 28084 15486
rect 27692 15262 27694 15314
rect 27746 15262 27748 15314
rect 27692 15250 27748 15262
rect 28140 15426 28196 15438
rect 28140 15374 28142 15426
rect 28194 15374 28196 15426
rect 28140 15092 28196 15374
rect 27804 15036 28140 15092
rect 27804 14644 27860 15036
rect 28140 14998 28196 15036
rect 27132 14642 27860 14644
rect 27132 14590 27134 14642
rect 27186 14590 27806 14642
rect 27858 14590 27860 14642
rect 27132 14588 27860 14590
rect 27132 14578 27188 14588
rect 27804 14578 27860 14588
rect 27916 14754 27972 14766
rect 27916 14702 27918 14754
rect 27970 14702 27972 14754
rect 27916 14084 27972 14702
rect 28140 14644 28196 14654
rect 28140 14550 28196 14588
rect 27580 14028 27972 14084
rect 27580 13970 27636 14028
rect 28252 13972 28308 17500
rect 28588 17106 28644 17838
rect 28588 17054 28590 17106
rect 28642 17054 28644 17106
rect 28588 16548 28644 17054
rect 28924 17106 28980 20636
rect 28924 17054 28926 17106
rect 28978 17054 28980 17106
rect 28476 16492 28644 16548
rect 28700 16772 28756 16782
rect 28364 15316 28420 15354
rect 28364 15250 28420 15260
rect 28476 14754 28532 16492
rect 28476 14702 28478 14754
rect 28530 14702 28532 14754
rect 28476 14690 28532 14702
rect 28588 16210 28644 16222
rect 28588 16158 28590 16210
rect 28642 16158 28644 16210
rect 28588 15092 28644 16158
rect 28588 14642 28644 15036
rect 28588 14590 28590 14642
rect 28642 14590 28644 14642
rect 28588 14578 28644 14590
rect 28700 15314 28756 16716
rect 28700 15262 28702 15314
rect 28754 15262 28756 15314
rect 28700 14644 28756 15262
rect 28924 16100 28980 17054
rect 29036 18450 29092 18462
rect 29036 18398 29038 18450
rect 29090 18398 29092 18450
rect 29036 16212 29092 18398
rect 29036 16146 29092 16156
rect 28924 15316 28980 16044
rect 29036 15876 29092 15886
rect 29036 15782 29092 15820
rect 29148 15540 29204 21756
rect 29596 20804 29652 20814
rect 29484 20802 29652 20804
rect 29484 20750 29598 20802
rect 29650 20750 29652 20802
rect 29484 20748 29652 20750
rect 29260 19234 29316 19246
rect 29260 19182 29262 19234
rect 29314 19182 29316 19234
rect 29260 18228 29316 19182
rect 29260 18162 29316 18172
rect 29260 16100 29316 16110
rect 29316 16044 29428 16100
rect 29260 16034 29316 16044
rect 29372 15986 29428 16044
rect 29372 15934 29374 15986
rect 29426 15934 29428 15986
rect 29372 15922 29428 15934
rect 29148 15474 29204 15484
rect 29260 15874 29316 15886
rect 29260 15822 29262 15874
rect 29314 15822 29316 15874
rect 29148 15316 29204 15326
rect 28924 15314 29204 15316
rect 28924 15262 29150 15314
rect 29202 15262 29204 15314
rect 28924 15260 29204 15262
rect 29148 15250 29204 15260
rect 29260 15316 29316 15822
rect 29260 15250 29316 15260
rect 29372 15540 29428 15550
rect 29372 14754 29428 15484
rect 29372 14702 29374 14754
rect 29426 14702 29428 14754
rect 29372 14690 29428 14702
rect 28700 14578 28756 14588
rect 27580 13918 27582 13970
rect 27634 13918 27636 13970
rect 26908 13860 26964 13870
rect 27244 13860 27300 13870
rect 27580 13860 27636 13918
rect 26908 13858 27076 13860
rect 26908 13806 26910 13858
rect 26962 13806 27076 13858
rect 26908 13804 27076 13806
rect 26908 13794 26964 13804
rect 26684 13234 26740 13244
rect 26908 13412 26964 13422
rect 26908 13076 26964 13356
rect 26572 13020 26964 13076
rect 26572 12962 26628 13020
rect 27020 12964 27076 13804
rect 27244 13858 27636 13860
rect 27244 13806 27246 13858
rect 27298 13806 27636 13858
rect 27244 13804 27636 13806
rect 27244 13794 27300 13804
rect 27356 13636 27412 13646
rect 26572 12910 26574 12962
rect 26626 12910 26628 12962
rect 26572 12898 26628 12910
rect 26908 12908 27076 12964
rect 27132 13412 27188 13422
rect 26460 12738 26516 12750
rect 26460 12686 26462 12738
rect 26514 12686 26516 12738
rect 26460 12180 26516 12686
rect 26460 12114 26516 12124
rect 26572 12066 26628 12078
rect 26572 12014 26574 12066
rect 26626 12014 26628 12066
rect 26572 11956 26628 12014
rect 26908 12068 26964 12908
rect 27020 12740 27076 12750
rect 27132 12740 27188 13356
rect 27020 12738 27188 12740
rect 27020 12686 27022 12738
rect 27074 12686 27188 12738
rect 27020 12684 27188 12686
rect 27020 12674 27076 12684
rect 26908 12002 26964 12012
rect 26348 11900 26628 11956
rect 25340 11452 25620 11508
rect 25340 11284 25396 11294
rect 25396 11228 25508 11284
rect 25340 11190 25396 11228
rect 25452 10612 25508 11228
rect 25452 9826 25508 10556
rect 25564 10052 25620 11452
rect 27020 10612 27076 10622
rect 27020 10518 27076 10556
rect 25564 9986 25620 9996
rect 26572 10052 26628 10062
rect 25452 9774 25454 9826
rect 25506 9774 25508 9826
rect 25452 9762 25508 9774
rect 26236 9716 26292 9726
rect 26236 9714 26516 9716
rect 26236 9662 26238 9714
rect 26290 9662 26516 9714
rect 26236 9660 26516 9662
rect 26236 9650 26292 9660
rect 25340 9156 25396 9166
rect 25228 9154 25396 9156
rect 25228 9102 25342 9154
rect 25394 9102 25396 9154
rect 25228 9100 25396 9102
rect 25340 9090 25396 9100
rect 25004 8978 25060 8988
rect 25788 9042 25844 9054
rect 25788 8990 25790 9042
rect 25842 8990 25844 9042
rect 24892 3390 24894 3442
rect 24946 3390 24948 3442
rect 24892 3378 24948 3390
rect 25564 3442 25620 3454
rect 25564 3390 25566 3442
rect 25618 3390 25620 3442
rect 22876 2492 23268 2548
rect 23548 2492 23940 2548
rect 24220 2492 24612 2548
rect 25564 3220 25620 3390
rect 25788 3442 25844 8990
rect 26236 9044 26292 9054
rect 26236 8930 26292 8988
rect 26236 8878 26238 8930
rect 26290 8878 26292 8930
rect 26236 8866 26292 8878
rect 26460 8482 26516 9660
rect 26572 9042 26628 9996
rect 26572 8990 26574 9042
rect 26626 8990 26628 9042
rect 26572 8978 26628 8990
rect 26460 8430 26462 8482
rect 26514 8430 26516 8482
rect 26460 8418 26516 8430
rect 26572 8818 26628 8830
rect 26572 8766 26574 8818
rect 26626 8766 26628 8818
rect 26572 8370 26628 8766
rect 26572 8318 26574 8370
rect 26626 8318 26628 8370
rect 26572 8306 26628 8318
rect 26908 4564 26964 4574
rect 27356 4564 27412 13580
rect 27580 13074 27636 13804
rect 27916 13970 28308 13972
rect 27916 13918 28254 13970
rect 28306 13918 28308 13970
rect 27916 13916 28308 13918
rect 27916 13858 27972 13916
rect 27916 13806 27918 13858
rect 27970 13806 27972 13858
rect 27916 13794 27972 13806
rect 27580 13022 27582 13074
rect 27634 13022 27636 13074
rect 27580 13010 27636 13022
rect 28252 13076 28308 13916
rect 28588 13858 28644 13870
rect 28588 13806 28590 13858
rect 28642 13806 28644 13858
rect 28588 13524 28644 13806
rect 29036 13636 29092 13646
rect 29036 13542 29092 13580
rect 28588 13458 28644 13468
rect 28252 12982 28308 13020
rect 28700 13300 28756 13310
rect 26908 4562 27412 4564
rect 26908 4510 26910 4562
rect 26962 4510 27412 4562
rect 26908 4508 27412 4510
rect 26908 4498 26964 4508
rect 27244 4340 27300 4350
rect 27132 4116 27188 4126
rect 26236 3668 26292 3678
rect 25788 3390 25790 3442
rect 25842 3390 25844 3442
rect 25788 3378 25844 3390
rect 26012 3554 26068 3566
rect 26012 3502 26014 3554
rect 26066 3502 26068 3554
rect 26012 3220 26068 3502
rect 25564 3164 26068 3220
rect 22876 800 22932 2492
rect 23548 800 23604 2492
rect 24220 800 24276 2492
rect 25564 800 25620 3164
rect 26236 800 26292 3612
rect 26796 3444 26852 3454
rect 27132 3388 27188 4060
rect 27244 3556 27300 4284
rect 27356 4338 27412 4508
rect 27356 4286 27358 4338
rect 27410 4286 27412 4338
rect 27356 4274 27412 4286
rect 27692 12178 27748 12190
rect 27692 12126 27694 12178
rect 27746 12126 27748 12178
rect 27244 3462 27300 3500
rect 27580 3554 27636 3566
rect 27580 3502 27582 3554
rect 27634 3502 27636 3554
rect 26796 3350 26852 3388
rect 26908 3332 27188 3388
rect 27580 3444 27636 3502
rect 27692 3444 27748 12126
rect 28028 12178 28084 12190
rect 28700 12180 28756 13244
rect 29372 13076 29428 13086
rect 29372 12982 29428 13020
rect 28028 12126 28030 12178
rect 28082 12126 28084 12178
rect 28028 11396 28084 12126
rect 28364 12178 28756 12180
rect 28364 12126 28702 12178
rect 28754 12126 28756 12178
rect 28364 12124 28756 12126
rect 28140 12068 28196 12078
rect 28140 11974 28196 12012
rect 28028 11330 28084 11340
rect 27804 10500 27860 10510
rect 27804 10498 28084 10500
rect 27804 10446 27806 10498
rect 27858 10446 28084 10498
rect 27804 10444 28084 10446
rect 27804 10434 27860 10444
rect 27916 9940 27972 9950
rect 27804 9044 27860 9054
rect 27804 8950 27860 8988
rect 27916 8930 27972 9884
rect 27916 8878 27918 8930
rect 27970 8878 27972 8930
rect 27916 8866 27972 8878
rect 28028 8370 28084 10444
rect 28028 8318 28030 8370
rect 28082 8318 28084 8370
rect 28028 8306 28084 8318
rect 28140 10052 28196 10062
rect 28140 8370 28196 9996
rect 28364 9938 28420 12124
rect 28700 12114 28756 12124
rect 29260 12178 29316 12190
rect 29260 12126 29262 12178
rect 29314 12126 29316 12178
rect 28812 11954 28868 11966
rect 28812 11902 28814 11954
rect 28866 11902 28868 11954
rect 28812 10052 28868 11902
rect 28812 9986 28868 9996
rect 29260 11284 29316 12126
rect 29372 11396 29428 11406
rect 29372 11302 29428 11340
rect 28364 9886 28366 9938
rect 28418 9886 28420 9938
rect 28364 9044 28420 9886
rect 29260 9940 29316 11228
rect 29260 9874 29316 9884
rect 28364 8978 28420 8988
rect 28700 9828 28756 9838
rect 28700 8930 28756 9772
rect 28700 8878 28702 8930
rect 28754 8878 28756 8930
rect 28700 8866 28756 8878
rect 28140 8318 28142 8370
rect 28194 8318 28196 8370
rect 28140 8306 28196 8318
rect 28700 5124 28756 5134
rect 29148 5124 29204 5134
rect 28700 5122 29204 5124
rect 28700 5070 28702 5122
rect 28754 5070 29150 5122
rect 29202 5070 29204 5122
rect 28700 5068 29204 5070
rect 28140 4116 28196 4126
rect 28140 4022 28196 4060
rect 28364 3556 28420 3566
rect 28364 3462 28420 3500
rect 27804 3444 27860 3454
rect 27692 3442 27860 3444
rect 27692 3390 27806 3442
rect 27858 3390 27860 3442
rect 27692 3388 27860 3390
rect 26908 800 26964 3332
rect 27580 800 27636 3388
rect 27804 3378 27860 3388
rect 28700 3388 28756 5068
rect 29148 5058 29204 5068
rect 29484 5010 29540 20748
rect 29596 20738 29652 20748
rect 29708 20244 29764 26852
rect 29932 23716 29988 23726
rect 29932 23622 29988 23660
rect 30156 23044 30212 27916
rect 30268 27860 30324 28030
rect 30268 27794 30324 27804
rect 30380 26908 30436 32508
rect 30492 31332 30548 36652
rect 30716 36482 30772 37324
rect 30940 37378 30996 37884
rect 30940 37326 30942 37378
rect 30994 37326 30996 37378
rect 30940 37314 30996 37326
rect 30716 36430 30718 36482
rect 30770 36430 30772 36482
rect 30716 36260 30772 36430
rect 30828 37042 30884 37054
rect 30828 36990 30830 37042
rect 30882 36990 30884 37042
rect 30828 36484 30884 36990
rect 30828 36418 30884 36428
rect 31052 36482 31108 38612
rect 31276 38612 31444 38668
rect 31500 38722 31556 38734
rect 31500 38670 31502 38722
rect 31554 38670 31556 38722
rect 31164 37604 31220 37614
rect 31164 37044 31220 37548
rect 31276 37044 31332 38612
rect 31388 38164 31444 38174
rect 31500 38164 31556 38670
rect 31612 38276 31668 38782
rect 31836 38668 31892 39228
rect 31612 38210 31668 38220
rect 31724 38612 31892 38668
rect 31388 38162 31556 38164
rect 31388 38110 31390 38162
rect 31442 38110 31556 38162
rect 31388 38108 31556 38110
rect 31388 38098 31444 38108
rect 31388 37380 31444 37390
rect 31388 37286 31444 37324
rect 31500 37380 31556 37390
rect 31500 37378 31668 37380
rect 31500 37326 31502 37378
rect 31554 37326 31668 37378
rect 31500 37324 31668 37326
rect 31500 37314 31556 37324
rect 31500 37044 31556 37054
rect 31276 37042 31556 37044
rect 31276 36990 31502 37042
rect 31554 36990 31556 37042
rect 31276 36988 31556 36990
rect 31164 36932 31220 36988
rect 31500 36978 31556 36988
rect 31164 36876 31444 36932
rect 31052 36430 31054 36482
rect 31106 36430 31108 36482
rect 31052 36418 31108 36430
rect 30716 36194 30772 36204
rect 30828 36260 30884 36270
rect 30828 36258 31108 36260
rect 30828 36206 30830 36258
rect 30882 36206 31108 36258
rect 30828 36204 31108 36206
rect 30828 36194 30884 36204
rect 30604 35028 30660 35038
rect 30660 34972 30996 35028
rect 30604 34934 30660 34972
rect 30940 34354 30996 34972
rect 30940 34302 30942 34354
rect 30994 34302 30996 34354
rect 30940 34290 30996 34302
rect 30940 33572 30996 33582
rect 30828 33122 30884 33134
rect 30828 33070 30830 33122
rect 30882 33070 30884 33122
rect 30828 32676 30884 33070
rect 30940 32786 30996 33516
rect 30940 32734 30942 32786
rect 30994 32734 30996 32786
rect 30940 32722 30996 32734
rect 30828 32610 30884 32620
rect 30716 32452 30772 32462
rect 30716 32358 30772 32396
rect 30492 31108 30548 31276
rect 30828 31108 30884 31118
rect 30492 31106 30884 31108
rect 30492 31054 30830 31106
rect 30882 31054 30884 31106
rect 30492 31052 30884 31054
rect 30492 29540 30548 31052
rect 30828 31042 30884 31052
rect 30940 31108 30996 31118
rect 30940 29652 30996 31052
rect 30940 29586 30996 29596
rect 30492 29426 30548 29484
rect 30492 29374 30494 29426
rect 30546 29374 30548 29426
rect 30492 29362 30548 29374
rect 31052 29428 31108 36204
rect 31164 35364 31220 35374
rect 31164 33348 31220 35308
rect 31276 35252 31332 35262
rect 31276 34914 31332 35196
rect 31276 34862 31278 34914
rect 31330 34862 31332 34914
rect 31276 34850 31332 34862
rect 31276 34242 31332 34254
rect 31276 34190 31278 34242
rect 31330 34190 31332 34242
rect 31276 33460 31332 34190
rect 31276 33394 31332 33404
rect 31164 33282 31220 33292
rect 31164 33122 31220 33134
rect 31164 33070 31166 33122
rect 31218 33070 31220 33122
rect 31164 32900 31220 33070
rect 31164 32834 31220 32844
rect 31276 32788 31332 32798
rect 31276 32674 31332 32732
rect 31276 32622 31278 32674
rect 31330 32622 31332 32674
rect 31276 31108 31332 32622
rect 31388 32452 31444 36876
rect 31612 35028 31668 37324
rect 31500 34972 31668 35028
rect 31500 33684 31556 34972
rect 31612 34804 31668 34814
rect 31612 34710 31668 34748
rect 31724 34356 31780 38612
rect 32060 35138 32116 40348
rect 32396 39844 32452 39854
rect 32508 39844 32564 41246
rect 32452 39788 32564 39844
rect 32396 39730 32452 39788
rect 32396 39678 32398 39730
rect 32450 39678 32452 39730
rect 32172 39620 32228 39630
rect 32172 39060 32228 39564
rect 32396 39508 32452 39678
rect 32396 39442 32452 39452
rect 32172 38966 32228 39004
rect 32508 39284 32564 39294
rect 32508 39058 32564 39228
rect 32508 39006 32510 39058
rect 32562 39006 32564 39058
rect 32508 38994 32564 39006
rect 32172 38612 32228 38622
rect 32172 36482 32228 38556
rect 32620 37044 32676 43596
rect 32732 42754 32788 42766
rect 32732 42702 32734 42754
rect 32786 42702 32788 42754
rect 32732 42644 32788 42702
rect 32732 42578 32788 42588
rect 32844 38668 32900 46956
rect 33068 47012 33124 47516
rect 33068 46946 33124 46956
rect 33180 46788 33236 50372
rect 33404 49028 33460 49066
rect 33404 48962 33460 48972
rect 33292 48244 33348 48254
rect 33292 48150 33348 48188
rect 33516 47908 33572 52110
rect 33516 47124 33572 47852
rect 33516 47058 33572 47068
rect 33180 46732 33348 46788
rect 33180 46562 33236 46574
rect 33180 46510 33182 46562
rect 33234 46510 33236 46562
rect 33180 46452 33236 46510
rect 33180 46386 33236 46396
rect 33180 43316 33236 43326
rect 33180 42868 33236 43260
rect 33180 42754 33236 42812
rect 33180 42702 33182 42754
rect 33234 42702 33236 42754
rect 33180 42690 33236 42702
rect 32620 36978 32676 36988
rect 32732 38612 32900 38668
rect 32956 42530 33012 42542
rect 32956 42478 32958 42530
rect 33010 42478 33012 42530
rect 32956 38668 33012 42478
rect 33292 41972 33348 46732
rect 33516 46452 33572 46462
rect 33404 46450 33572 46452
rect 33404 46398 33518 46450
rect 33570 46398 33572 46450
rect 33404 46396 33572 46398
rect 33404 45780 33460 46396
rect 33516 46386 33572 46396
rect 33628 45892 33684 53452
rect 33964 53396 34020 54684
rect 34076 54674 34132 54684
rect 33852 53340 34020 53396
rect 34076 53508 34132 53518
rect 33852 52050 33908 53340
rect 33852 51998 33854 52050
rect 33906 51998 33908 52050
rect 33852 51986 33908 51998
rect 33964 51828 34020 51838
rect 33964 51490 34020 51772
rect 33964 51438 33966 51490
rect 34018 51438 34020 51490
rect 33964 51426 34020 51438
rect 34076 51716 34132 53452
rect 33852 50820 33908 50830
rect 33852 50706 33908 50764
rect 33852 50654 33854 50706
rect 33906 50654 33908 50706
rect 33852 50642 33908 50654
rect 33740 48916 33796 48926
rect 33740 48466 33796 48860
rect 33740 48414 33742 48466
rect 33794 48414 33796 48466
rect 33740 48402 33796 48414
rect 33852 47908 33908 47918
rect 33740 47458 33796 47470
rect 33740 47406 33742 47458
rect 33794 47406 33796 47458
rect 33740 46564 33796 47406
rect 33740 46004 33796 46508
rect 33740 45938 33796 45948
rect 33628 45826 33684 45836
rect 33404 45330 33460 45724
rect 33404 45278 33406 45330
rect 33458 45278 33460 45330
rect 33404 45266 33460 45278
rect 33516 45556 33572 45566
rect 33516 45330 33572 45500
rect 33740 45332 33796 45342
rect 33516 45278 33518 45330
rect 33570 45278 33572 45330
rect 33516 45266 33572 45278
rect 33628 45276 33740 45332
rect 33628 45218 33684 45276
rect 33740 45266 33796 45276
rect 33628 45166 33630 45218
rect 33682 45166 33684 45218
rect 33628 45154 33684 45166
rect 33404 44436 33460 44446
rect 33404 44342 33460 44380
rect 33740 43540 33796 43550
rect 33740 43446 33796 43484
rect 33628 42756 33684 42766
rect 33852 42756 33908 47852
rect 33964 47012 34020 47022
rect 33964 46786 34020 46956
rect 33964 46734 33966 46786
rect 34018 46734 34020 46786
rect 33964 45444 34020 46734
rect 34076 46788 34132 51660
rect 34188 47012 34244 55244
rect 34412 55188 34468 55198
rect 34412 54852 34468 55132
rect 34412 54738 34468 54796
rect 34412 54686 34414 54738
rect 34466 54686 34468 54738
rect 34412 54674 34468 54686
rect 34524 54516 34580 58268
rect 34636 57540 34692 58380
rect 34636 57474 34692 57484
rect 34860 58210 34916 58222
rect 34860 58158 34862 58210
rect 34914 58158 34916 58210
rect 34860 58100 34916 58158
rect 34860 56868 34916 58044
rect 34860 56802 34916 56812
rect 35084 56756 35140 59612
rect 35420 59108 35476 60172
rect 35532 60004 35588 60732
rect 35756 60786 35924 60788
rect 35756 60734 35758 60786
rect 35810 60734 35924 60786
rect 35756 60732 35924 60734
rect 35756 60722 35812 60732
rect 35532 59938 35588 59948
rect 35532 59780 35588 59790
rect 35532 59686 35588 59724
rect 35644 59778 35700 59790
rect 35644 59726 35646 59778
rect 35698 59726 35700 59778
rect 35532 59332 35588 59342
rect 35644 59332 35700 59726
rect 35532 59330 35700 59332
rect 35532 59278 35534 59330
rect 35586 59278 35700 59330
rect 35532 59276 35700 59278
rect 35756 59778 35812 59790
rect 35756 59726 35758 59778
rect 35810 59726 35812 59778
rect 35532 59266 35588 59276
rect 35756 59108 35812 59726
rect 35420 59052 35588 59108
rect 35196 58828 35460 58838
rect 35252 58772 35300 58828
rect 35356 58772 35404 58828
rect 35196 58762 35460 58772
rect 35196 58548 35252 58558
rect 35196 58322 35252 58492
rect 35196 58270 35198 58322
rect 35250 58270 35252 58322
rect 35196 58212 35252 58270
rect 35532 58324 35588 59052
rect 35756 59042 35812 59052
rect 35868 58996 35924 60732
rect 35980 60340 36036 60956
rect 35980 60114 36036 60284
rect 35980 60062 35982 60114
rect 36034 60062 36036 60114
rect 35980 60050 36036 60062
rect 36092 60228 36148 62190
rect 36764 62188 36820 65660
rect 37436 65604 37492 66220
rect 37324 65548 37492 65604
rect 37660 66274 37716 66286
rect 37660 66222 37662 66274
rect 37714 66222 37716 66274
rect 37660 66052 37716 66222
rect 37324 65492 37380 65548
rect 37212 64708 37268 64718
rect 37212 64594 37268 64652
rect 37212 64542 37214 64594
rect 37266 64542 37268 64594
rect 37100 63812 37156 63822
rect 37212 63812 37268 64542
rect 37324 64148 37380 65436
rect 37324 64082 37380 64092
rect 37436 65378 37492 65390
rect 37436 65326 37438 65378
rect 37490 65326 37492 65378
rect 37436 64706 37492 65326
rect 37436 64654 37438 64706
rect 37490 64654 37492 64706
rect 37436 63922 37492 64654
rect 37660 64148 37716 65996
rect 37772 64148 37828 64158
rect 37660 64146 37828 64148
rect 37660 64094 37774 64146
rect 37826 64094 37828 64146
rect 37660 64092 37828 64094
rect 37772 64082 37828 64092
rect 37996 64148 38052 64158
rect 37996 64054 38052 64092
rect 37436 63870 37438 63922
rect 37490 63870 37492 63922
rect 37436 63858 37492 63870
rect 36988 63756 37100 63812
rect 37156 63756 37268 63812
rect 36876 62916 36932 62926
rect 36876 62822 36932 62860
rect 36988 62188 37044 63756
rect 37100 63746 37156 63756
rect 37100 63476 37156 63486
rect 37100 63026 37156 63420
rect 37212 63140 37268 63756
rect 37884 63810 37940 63822
rect 37884 63758 37886 63810
rect 37938 63758 37940 63810
rect 37884 63364 37940 63758
rect 38108 63700 38164 66556
rect 38668 66274 38724 66286
rect 38668 66222 38670 66274
rect 38722 66222 38724 66274
rect 38668 65604 38724 66222
rect 38444 65548 38724 65604
rect 38444 65492 38500 65548
rect 38892 65492 38948 65502
rect 38220 65436 38500 65492
rect 38556 65436 38892 65492
rect 38220 64820 38276 65436
rect 38332 65268 38388 65278
rect 38388 65212 38500 65268
rect 38332 65202 38388 65212
rect 38220 64764 38388 64820
rect 38220 64594 38276 64606
rect 38220 64542 38222 64594
rect 38274 64542 38276 64594
rect 38220 63812 38276 64542
rect 38332 64260 38388 64764
rect 38332 63922 38388 64204
rect 38332 63870 38334 63922
rect 38386 63870 38388 63922
rect 38332 63858 38388 63870
rect 38220 63746 38276 63756
rect 37884 63298 37940 63308
rect 37996 63644 38164 63700
rect 37884 63140 37940 63150
rect 37212 63046 37268 63084
rect 37660 63084 37884 63140
rect 37100 62974 37102 63026
rect 37154 62974 37156 63026
rect 37100 62962 37156 62974
rect 36316 62132 36820 62188
rect 36876 62132 37044 62188
rect 37100 62692 37156 62702
rect 37100 62188 37156 62636
rect 37660 62578 37716 63084
rect 37884 63046 37940 63084
rect 37660 62526 37662 62578
rect 37714 62526 37716 62578
rect 37660 62514 37716 62526
rect 37324 62242 37380 62254
rect 37324 62190 37326 62242
rect 37378 62190 37380 62242
rect 37100 62132 37268 62188
rect 36204 61348 36260 61358
rect 36204 61254 36260 61292
rect 36092 59668 36148 60172
rect 36204 60228 36260 60238
rect 36316 60228 36372 62132
rect 36428 60676 36484 60686
rect 36428 60582 36484 60620
rect 36204 60226 36372 60228
rect 36204 60174 36206 60226
rect 36258 60174 36372 60226
rect 36204 60172 36372 60174
rect 36204 60162 36260 60172
rect 36092 59602 36148 59612
rect 36876 59220 36932 62132
rect 36988 60452 37044 60462
rect 36988 59332 37044 60396
rect 36988 59266 37044 59276
rect 37100 60002 37156 60014
rect 37100 59950 37102 60002
rect 37154 59950 37156 60002
rect 37100 59780 37156 59950
rect 35868 58930 35924 58940
rect 36652 59164 36932 59220
rect 36316 58884 36372 58894
rect 35532 58258 35588 58268
rect 36092 58324 36148 58334
rect 36092 58230 36148 58268
rect 35196 58146 35252 58156
rect 35644 58210 35700 58222
rect 35644 58158 35646 58210
rect 35698 58158 35700 58210
rect 35644 58100 35700 58158
rect 35644 58034 35700 58044
rect 35196 57260 35460 57270
rect 35252 57204 35300 57260
rect 35356 57204 35404 57260
rect 35196 57194 35460 57204
rect 36316 57090 36372 58828
rect 36316 57038 36318 57090
rect 36370 57038 36372 57090
rect 36316 57026 36372 57038
rect 36428 58660 36484 58670
rect 36428 56866 36484 58604
rect 36428 56814 36430 56866
rect 36482 56814 36484 56866
rect 36428 56802 36484 56814
rect 35196 56756 35252 56766
rect 35084 56754 35252 56756
rect 35084 56702 35198 56754
rect 35250 56702 35252 56754
rect 35084 56700 35252 56702
rect 35196 56690 35252 56700
rect 34860 56644 34916 56654
rect 34860 56550 34916 56588
rect 34972 56082 35028 56094
rect 34972 56030 34974 56082
rect 35026 56030 35028 56082
rect 34972 55410 35028 56030
rect 35196 55692 35460 55702
rect 35252 55636 35300 55692
rect 35356 55636 35404 55692
rect 35196 55626 35460 55636
rect 34972 55358 34974 55410
rect 35026 55358 35028 55410
rect 34972 55300 35028 55358
rect 36316 55524 36372 55534
rect 36204 55300 36260 55310
rect 34972 55234 35028 55244
rect 35756 55298 36260 55300
rect 35756 55246 36206 55298
rect 36258 55246 36260 55298
rect 35756 55244 36260 55246
rect 35644 55186 35700 55198
rect 35644 55134 35646 55186
rect 35698 55134 35700 55186
rect 35308 55074 35364 55086
rect 35308 55022 35310 55074
rect 35362 55022 35364 55074
rect 34860 54740 34916 54750
rect 34748 54626 34804 54638
rect 34748 54574 34750 54626
rect 34802 54574 34804 54626
rect 34300 54460 34580 54516
rect 34636 54516 34692 54526
rect 34300 50428 34356 54460
rect 34412 53730 34468 53742
rect 34412 53678 34414 53730
rect 34466 53678 34468 53730
rect 34412 53620 34468 53678
rect 34412 53554 34468 53564
rect 34524 53060 34580 53070
rect 34412 53058 34580 53060
rect 34412 53006 34526 53058
rect 34578 53006 34580 53058
rect 34412 53004 34580 53006
rect 34412 51940 34468 53004
rect 34524 52994 34580 53004
rect 34636 53058 34692 54460
rect 34748 54292 34804 54574
rect 34748 54226 34804 54236
rect 34860 54628 34916 54684
rect 35084 54628 35140 54638
rect 34860 54626 35140 54628
rect 34860 54574 35086 54626
rect 35138 54574 35140 54626
rect 34860 54572 35140 54574
rect 34860 53956 34916 54572
rect 35084 54562 35140 54572
rect 35308 54516 35364 55022
rect 35644 55076 35700 55134
rect 35644 55010 35700 55020
rect 35756 54852 35812 55244
rect 36204 55234 36260 55244
rect 35868 55076 35924 55086
rect 35868 54982 35924 55020
rect 35980 55076 36036 55086
rect 35980 55074 36148 55076
rect 35980 55022 35982 55074
rect 36034 55022 36148 55074
rect 35980 55020 36148 55022
rect 35980 55010 36036 55020
rect 35532 54796 35812 54852
rect 35532 54516 35588 54796
rect 35308 54514 35588 54516
rect 35308 54462 35310 54514
rect 35362 54462 35588 54514
rect 35308 54460 35588 54462
rect 35308 54450 35364 54460
rect 34748 53900 34916 53956
rect 34972 54404 35028 54414
rect 34748 53284 34804 53900
rect 34972 53842 35028 54348
rect 34972 53790 34974 53842
rect 35026 53790 35028 53842
rect 34972 53778 35028 53790
rect 35084 54292 35140 54302
rect 35084 53844 35140 54236
rect 35420 54292 35476 54330
rect 35420 54226 35476 54236
rect 35196 54124 35460 54134
rect 35252 54068 35300 54124
rect 35356 54068 35404 54124
rect 35196 54058 35460 54068
rect 35532 53956 35588 54460
rect 35084 53730 35140 53788
rect 35084 53678 35086 53730
rect 35138 53678 35140 53730
rect 35084 53666 35140 53678
rect 35308 53900 35588 53956
rect 35644 54514 35700 54526
rect 35644 54462 35646 54514
rect 35698 54462 35700 54514
rect 34860 53508 34916 53518
rect 34860 53414 34916 53452
rect 34748 53218 34804 53228
rect 35196 53172 35252 53182
rect 35308 53172 35364 53900
rect 35532 53730 35588 53742
rect 35532 53678 35534 53730
rect 35586 53678 35588 53730
rect 35252 53116 35364 53172
rect 35420 53284 35476 53294
rect 35420 53170 35476 53228
rect 35420 53118 35422 53170
rect 35474 53118 35476 53170
rect 35196 53078 35252 53116
rect 35420 53106 35476 53118
rect 35532 53170 35588 53678
rect 35532 53118 35534 53170
rect 35586 53118 35588 53170
rect 35532 53106 35588 53118
rect 34636 53006 34638 53058
rect 34690 53006 34692 53058
rect 34636 52994 34692 53006
rect 34860 52946 34916 52958
rect 34860 52894 34862 52946
rect 34914 52894 34916 52946
rect 34524 52724 34580 52734
rect 34860 52724 34916 52894
rect 35644 52948 35700 54462
rect 35756 54514 35812 54526
rect 35756 54462 35758 54514
rect 35810 54462 35812 54514
rect 35756 54292 35812 54462
rect 35756 54226 35812 54236
rect 35756 53956 35812 53966
rect 35756 53730 35812 53900
rect 35756 53678 35758 53730
rect 35810 53678 35812 53730
rect 35756 53666 35812 53678
rect 35980 53844 36036 53854
rect 35980 53730 36036 53788
rect 35980 53678 35982 53730
rect 36034 53678 36036 53730
rect 35980 53666 36036 53678
rect 35644 52882 35700 52892
rect 35868 53506 35924 53518
rect 35868 53454 35870 53506
rect 35922 53454 35924 53506
rect 34524 52722 34916 52724
rect 34524 52670 34526 52722
rect 34578 52670 34916 52722
rect 34524 52668 34916 52670
rect 34972 52836 35028 52846
rect 34524 52658 34580 52668
rect 34860 52276 34916 52286
rect 34972 52276 35028 52780
rect 35868 52836 35924 53454
rect 36092 53060 36148 55020
rect 36316 54738 36372 55468
rect 36316 54686 36318 54738
rect 36370 54686 36372 54738
rect 36316 54674 36372 54686
rect 36540 55298 36596 55310
rect 36540 55246 36542 55298
rect 36594 55246 36596 55298
rect 36204 54514 36260 54526
rect 36204 54462 36206 54514
rect 36258 54462 36260 54514
rect 36204 53844 36260 54462
rect 36428 54516 36484 54526
rect 36428 54422 36484 54460
rect 36428 53956 36484 53966
rect 36204 53508 36260 53788
rect 36204 53442 36260 53452
rect 36316 53900 36428 53956
rect 36092 52836 36148 53004
rect 36204 52836 36260 52846
rect 36092 52780 36204 52836
rect 35868 52770 35924 52780
rect 36204 52770 36260 52780
rect 35196 52556 35460 52566
rect 35252 52500 35300 52556
rect 35356 52500 35404 52556
rect 35196 52490 35460 52500
rect 34860 52274 35028 52276
rect 34860 52222 34862 52274
rect 34914 52222 35028 52274
rect 34860 52220 35028 52222
rect 34860 52210 34916 52220
rect 34412 51874 34468 51884
rect 34748 51938 34804 51950
rect 34748 51886 34750 51938
rect 34802 51886 34804 51938
rect 34748 51828 34804 51886
rect 34748 51762 34804 51772
rect 36316 51604 36372 53900
rect 36428 53890 36484 53900
rect 36428 53730 36484 53742
rect 36428 53678 36430 53730
rect 36482 53678 36484 53730
rect 36428 53170 36484 53678
rect 36540 53732 36596 55246
rect 36540 53666 36596 53676
rect 36428 53118 36430 53170
rect 36482 53118 36484 53170
rect 36428 53106 36484 53118
rect 36540 53058 36596 53070
rect 36540 53006 36542 53058
rect 36594 53006 36596 53058
rect 36540 52836 36596 53006
rect 36540 52770 36596 52780
rect 36428 51604 36484 51614
rect 36204 51602 36484 51604
rect 36204 51550 36430 51602
rect 36482 51550 36484 51602
rect 36204 51548 36484 51550
rect 35644 51492 35700 51502
rect 35196 50988 35460 50998
rect 35252 50932 35300 50988
rect 35356 50932 35404 50988
rect 35196 50922 35460 50932
rect 35644 50708 35700 51436
rect 36092 51268 36148 51278
rect 36092 51174 36148 51212
rect 35644 50706 35924 50708
rect 35644 50654 35646 50706
rect 35698 50654 35924 50706
rect 35644 50652 35924 50654
rect 35644 50642 35700 50652
rect 35868 50594 35924 50652
rect 36204 50596 36260 51548
rect 36428 51538 36484 51548
rect 36652 50932 36708 59164
rect 36876 58996 36932 59006
rect 36876 57538 36932 58940
rect 37100 58884 37156 59724
rect 37100 58434 37156 58828
rect 37100 58382 37102 58434
rect 37154 58382 37156 58434
rect 37100 58370 37156 58382
rect 36876 57486 36878 57538
rect 36930 57486 36932 57538
rect 36876 55300 36932 57486
rect 36988 56754 37044 56766
rect 36988 56702 36990 56754
rect 37042 56702 37044 56754
rect 36988 55524 37044 56702
rect 37100 56644 37156 56654
rect 37100 56550 37156 56588
rect 36988 55458 37044 55468
rect 36988 55300 37044 55310
rect 36876 55298 37044 55300
rect 36876 55246 36990 55298
rect 37042 55246 37044 55298
rect 36876 55244 37044 55246
rect 36764 54516 36820 54526
rect 36988 54516 37044 55244
rect 36764 54514 37044 54516
rect 36764 54462 36766 54514
rect 36818 54462 37044 54514
rect 36764 54460 37044 54462
rect 37100 55076 37156 55086
rect 36764 53620 36820 54460
rect 36764 53554 36820 53564
rect 37100 53618 37156 55020
rect 37100 53566 37102 53618
rect 37154 53566 37156 53618
rect 37100 53554 37156 53566
rect 37212 53284 37268 62132
rect 37324 61572 37380 62190
rect 37548 61572 37604 61582
rect 37324 61570 37604 61572
rect 37324 61518 37550 61570
rect 37602 61518 37604 61570
rect 37324 61516 37604 61518
rect 37324 61346 37380 61358
rect 37324 61294 37326 61346
rect 37378 61294 37380 61346
rect 37324 60452 37380 61294
rect 37548 61348 37604 61516
rect 37996 61458 38052 63644
rect 38108 63252 38164 63262
rect 38108 63138 38164 63196
rect 38332 63252 38388 63262
rect 38444 63252 38500 65212
rect 38332 63250 38500 63252
rect 38332 63198 38334 63250
rect 38386 63198 38500 63250
rect 38332 63196 38500 63198
rect 38332 63186 38388 63196
rect 38108 63086 38110 63138
rect 38162 63086 38164 63138
rect 38108 63074 38164 63086
rect 38220 63140 38276 63150
rect 38108 62580 38164 62590
rect 38220 62580 38276 63084
rect 38444 63026 38500 63038
rect 38444 62974 38446 63026
rect 38498 62974 38500 63026
rect 38444 62692 38500 62974
rect 38444 62626 38500 62636
rect 38108 62578 38276 62580
rect 38108 62526 38110 62578
rect 38162 62526 38276 62578
rect 38108 62524 38276 62526
rect 38556 62580 38612 65436
rect 38892 65426 38948 65436
rect 38892 65156 38948 65166
rect 38668 65100 38892 65156
rect 38668 64146 38724 65100
rect 38892 65090 38948 65100
rect 38668 64094 38670 64146
rect 38722 64094 38724 64146
rect 38668 64082 38724 64094
rect 38892 64148 38948 64158
rect 38892 64054 38948 64092
rect 38780 63812 38836 63822
rect 38780 63718 38836 63756
rect 38892 63700 38948 63710
rect 38892 63250 38948 63644
rect 38892 63198 38894 63250
rect 38946 63198 38948 63250
rect 38892 62916 38948 63198
rect 38892 62850 38948 62860
rect 38108 62514 38164 62524
rect 38556 62188 38612 62524
rect 38332 62132 38612 62188
rect 37996 61406 37998 61458
rect 38050 61406 38052 61458
rect 37996 61394 38052 61406
rect 38108 61682 38164 61694
rect 38108 61630 38110 61682
rect 38162 61630 38164 61682
rect 37548 61282 37604 61292
rect 37324 60386 37380 60396
rect 37436 60788 37492 60798
rect 37324 60002 37380 60014
rect 37324 59950 37326 60002
rect 37378 59950 37380 60002
rect 37324 59556 37380 59950
rect 37436 59778 37492 60732
rect 38108 60116 38164 61630
rect 37548 60114 38164 60116
rect 37548 60062 38110 60114
rect 38162 60062 38164 60114
rect 37548 60060 38164 60062
rect 37548 60002 37604 60060
rect 37548 59950 37550 60002
rect 37602 59950 37604 60002
rect 37548 59938 37604 59950
rect 37436 59726 37438 59778
rect 37490 59726 37492 59778
rect 37436 59714 37492 59726
rect 37324 59500 38052 59556
rect 37548 58434 37604 59500
rect 37996 59442 38052 59500
rect 37996 59390 37998 59442
rect 38050 59390 38052 59442
rect 37996 59378 38052 59390
rect 38108 59220 38164 60060
rect 38220 60002 38276 60014
rect 38220 59950 38222 60002
rect 38274 59950 38276 60002
rect 38220 59780 38276 59950
rect 38220 59714 38276 59724
rect 37772 59164 38164 59220
rect 37660 59106 37716 59118
rect 37660 59054 37662 59106
rect 37714 59054 37716 59106
rect 37660 58660 37716 59054
rect 37660 58594 37716 58604
rect 37548 58382 37550 58434
rect 37602 58382 37604 58434
rect 37548 58370 37604 58382
rect 37660 58210 37716 58222
rect 37660 58158 37662 58210
rect 37714 58158 37716 58210
rect 37660 57988 37716 58158
rect 37772 58210 37828 59164
rect 38220 58436 38276 58446
rect 37772 58158 37774 58210
rect 37826 58158 37828 58210
rect 37772 58146 37828 58158
rect 38108 58322 38164 58334
rect 38108 58270 38110 58322
rect 38162 58270 38164 58322
rect 38108 57988 38164 58270
rect 37660 57932 38164 57988
rect 38220 58322 38276 58380
rect 38220 58270 38222 58322
rect 38274 58270 38276 58322
rect 38220 57988 38276 58270
rect 38220 57922 38276 57932
rect 38332 57652 38388 62132
rect 38668 61570 38724 61582
rect 38668 61518 38670 61570
rect 38722 61518 38724 61570
rect 38668 61348 38724 61518
rect 39004 61572 39060 67788
rect 39116 66836 39172 68572
rect 39452 68628 39508 68638
rect 39788 68628 39844 68638
rect 39452 68626 39844 68628
rect 39452 68574 39454 68626
rect 39506 68574 39790 68626
rect 39842 68574 39844 68626
rect 39452 68572 39844 68574
rect 39452 68562 39508 68572
rect 39788 68562 39844 68572
rect 39900 68516 39956 69244
rect 40124 69188 40180 70142
rect 40348 70196 40404 70206
rect 40348 70102 40404 70140
rect 40908 70194 40964 70252
rect 41692 70306 41748 71484
rect 41692 70254 41694 70306
rect 41746 70254 41748 70306
rect 41692 70242 41748 70254
rect 41916 70978 41972 70990
rect 41916 70926 41918 70978
rect 41970 70926 41972 70978
rect 41916 70756 41972 70926
rect 41244 70196 41300 70206
rect 40908 70142 40910 70194
rect 40962 70142 40964 70194
rect 40460 69300 40516 69310
rect 40460 69206 40516 69244
rect 40124 68964 40180 69132
rect 40908 68964 40964 70142
rect 40124 68908 40516 68964
rect 40348 68738 40404 68750
rect 40348 68686 40350 68738
rect 40402 68686 40404 68738
rect 40124 68626 40180 68638
rect 40124 68574 40126 68626
rect 40178 68574 40180 68626
rect 40012 68516 40068 68526
rect 39900 68514 40068 68516
rect 39900 68462 40014 68514
rect 40066 68462 40068 68514
rect 39900 68460 40068 68462
rect 40012 68450 40068 68460
rect 40124 68516 40180 68574
rect 40124 68450 40180 68460
rect 39676 67620 39732 67630
rect 40236 67620 40292 67630
rect 39676 67284 39732 67564
rect 39676 67190 39732 67228
rect 40124 67564 40236 67620
rect 40348 67620 40404 68686
rect 40460 68740 40516 68908
rect 40908 68898 40964 68908
rect 41132 70140 41244 70196
rect 40460 68674 40516 68684
rect 40908 68626 40964 68638
rect 40908 68574 40910 68626
rect 40962 68574 40964 68626
rect 40796 68516 40852 68526
rect 40796 67842 40852 68460
rect 40908 68066 40964 68574
rect 40908 68014 40910 68066
rect 40962 68014 40964 68066
rect 40908 68002 40964 68014
rect 40796 67790 40798 67842
rect 40850 67790 40852 67842
rect 40796 67778 40852 67790
rect 41020 67730 41076 67742
rect 41020 67678 41022 67730
rect 41074 67678 41076 67730
rect 40572 67620 40628 67630
rect 40348 67618 40628 67620
rect 40348 67566 40574 67618
rect 40626 67566 40628 67618
rect 40348 67564 40628 67566
rect 39116 66770 39172 66780
rect 39900 66162 39956 66174
rect 39900 66110 39902 66162
rect 39954 66110 39956 66162
rect 39116 66050 39172 66062
rect 39116 65998 39118 66050
rect 39170 65998 39172 66050
rect 39116 65268 39172 65998
rect 39116 65202 39172 65212
rect 39228 66050 39284 66062
rect 39228 65998 39230 66050
rect 39282 65998 39284 66050
rect 39228 65156 39284 65998
rect 39340 66050 39396 66062
rect 39340 65998 39342 66050
rect 39394 65998 39396 66050
rect 39340 65380 39396 65998
rect 39564 66052 39620 66062
rect 39564 66050 39732 66052
rect 39564 65998 39566 66050
rect 39618 65998 39732 66050
rect 39564 65996 39732 65998
rect 39564 65986 39620 65996
rect 39340 65314 39396 65324
rect 39228 65090 39284 65100
rect 39340 64148 39396 64158
rect 39564 64148 39620 64158
rect 39396 64146 39620 64148
rect 39396 64094 39566 64146
rect 39618 64094 39620 64146
rect 39396 64092 39620 64094
rect 39340 64082 39396 64092
rect 39564 64082 39620 64092
rect 39340 63924 39396 63934
rect 39676 63924 39732 65996
rect 39340 63922 39732 63924
rect 39340 63870 39342 63922
rect 39394 63870 39732 63922
rect 39340 63868 39732 63870
rect 39788 66050 39844 66062
rect 39788 65998 39790 66050
rect 39842 65998 39844 66050
rect 39340 63858 39396 63868
rect 39788 63476 39844 65998
rect 39900 66052 39956 66110
rect 39900 65986 39956 65996
rect 40124 65492 40180 67564
rect 40236 67526 40292 67564
rect 40236 66946 40292 66958
rect 40236 66894 40238 66946
rect 40290 66894 40292 66946
rect 40236 66052 40292 66894
rect 40572 66836 40628 67564
rect 40572 66770 40628 66780
rect 41020 66500 41076 67678
rect 41132 67228 41188 70140
rect 41244 70130 41300 70140
rect 41468 69524 41524 69534
rect 41356 68852 41412 68862
rect 41356 68758 41412 68796
rect 41468 68852 41524 69468
rect 41468 68850 41636 68852
rect 41468 68798 41470 68850
rect 41522 68798 41636 68850
rect 41468 68796 41636 68798
rect 41468 68786 41524 68796
rect 41244 68740 41300 68750
rect 41244 68646 41300 68684
rect 41356 67954 41412 67966
rect 41356 67902 41358 67954
rect 41410 67902 41412 67954
rect 41132 67172 41300 67228
rect 41132 67058 41188 67070
rect 41132 67006 41134 67058
rect 41186 67006 41188 67058
rect 41132 66948 41188 67006
rect 41132 66882 41188 66892
rect 41132 66500 41188 66510
rect 41020 66498 41188 66500
rect 41020 66446 41134 66498
rect 41186 66446 41188 66498
rect 41020 66444 41188 66446
rect 41132 66434 41188 66444
rect 41244 66276 41300 67172
rect 41356 67172 41412 67902
rect 41356 67106 41412 67116
rect 41468 67170 41524 67182
rect 41468 67118 41470 67170
rect 41522 67118 41524 67170
rect 41468 66836 41524 67118
rect 41468 66770 41524 66780
rect 41580 66276 41636 68796
rect 41916 67620 41972 70700
rect 42700 70756 42756 70766
rect 42700 70662 42756 70700
rect 50556 70588 50820 70598
rect 50612 70532 50660 70588
rect 50716 70532 50764 70588
rect 50556 70522 50820 70532
rect 43820 70196 43876 70206
rect 43820 70082 43876 70140
rect 43820 70030 43822 70082
rect 43874 70030 43876 70082
rect 43820 70018 43876 70030
rect 42588 69524 42644 69534
rect 42588 69430 42644 69468
rect 43708 69298 43764 69310
rect 43708 69246 43710 69298
rect 43762 69246 43764 69298
rect 42924 69188 42980 69198
rect 42924 69094 42980 69132
rect 43260 69186 43316 69198
rect 43260 69134 43262 69186
rect 43314 69134 43316 69186
rect 42364 68964 42420 68974
rect 42364 68738 42420 68908
rect 42364 68686 42366 68738
rect 42418 68686 42420 68738
rect 42364 68674 42420 68686
rect 41916 67554 41972 67564
rect 43260 67396 43316 69134
rect 43596 69186 43652 69198
rect 43596 69134 43598 69186
rect 43650 69134 43652 69186
rect 43484 67956 43540 67966
rect 43596 67956 43652 69134
rect 43484 67954 43652 67956
rect 43484 67902 43486 67954
rect 43538 67902 43652 67954
rect 43484 67900 43652 67902
rect 43484 67890 43540 67900
rect 43260 67340 43540 67396
rect 42028 67284 42084 67294
rect 41804 67172 41860 67182
rect 41244 66182 41300 66220
rect 41356 66274 41636 66276
rect 41356 66222 41582 66274
rect 41634 66222 41636 66274
rect 41356 66220 41636 66222
rect 40348 66052 40404 66062
rect 41132 66052 41188 66062
rect 40236 65996 40348 66052
rect 40404 65996 40516 66052
rect 40348 65958 40404 65996
rect 40236 65492 40292 65502
rect 40124 65436 40236 65492
rect 40236 65398 40292 65436
rect 39900 65380 39956 65390
rect 39900 63810 39956 65324
rect 40124 65268 40180 65278
rect 40124 64596 40180 65212
rect 40124 63924 40180 64540
rect 39900 63758 39902 63810
rect 39954 63758 39956 63810
rect 39900 63746 39956 63758
rect 40012 63922 40180 63924
rect 40012 63870 40126 63922
rect 40178 63870 40180 63922
rect 40012 63868 40180 63870
rect 40460 64484 40516 65996
rect 41132 65958 41188 65996
rect 41356 65716 41412 66220
rect 41580 66210 41636 66220
rect 41692 67170 41860 67172
rect 41692 67118 41806 67170
rect 41858 67118 41860 67170
rect 41692 67116 41860 67118
rect 41132 65660 41412 65716
rect 41692 66052 41748 67116
rect 41804 67106 41860 67116
rect 42028 67058 42084 67228
rect 42028 67006 42030 67058
rect 42082 67006 42084 67058
rect 41916 66164 41972 66174
rect 41916 66070 41972 66108
rect 41692 65716 41748 65996
rect 41020 65380 41076 65390
rect 41020 65286 41076 65324
rect 40460 63924 40516 64428
rect 40908 65266 40964 65278
rect 40908 65214 40910 65266
rect 40962 65214 40964 65266
rect 40908 64148 40964 65214
rect 41132 64706 41188 65660
rect 41692 65650 41748 65660
rect 41244 65490 41300 65502
rect 41244 65438 41246 65490
rect 41298 65438 41300 65490
rect 41244 64932 41300 65438
rect 41804 65378 41860 65390
rect 41804 65326 41806 65378
rect 41858 65326 41860 65378
rect 41244 64866 41300 64876
rect 41468 65266 41524 65278
rect 41468 65214 41470 65266
rect 41522 65214 41524 65266
rect 41132 64654 41134 64706
rect 41186 64654 41188 64706
rect 41020 64594 41076 64606
rect 41020 64542 41022 64594
rect 41074 64542 41076 64594
rect 41020 64484 41076 64542
rect 41020 64418 41076 64428
rect 41020 64148 41076 64158
rect 40908 64146 41076 64148
rect 40908 64094 41022 64146
rect 41074 64094 41076 64146
rect 40908 64092 41076 64094
rect 41020 64082 41076 64092
rect 40684 63924 40740 63934
rect 40460 63868 40684 63924
rect 39788 63410 39844 63420
rect 40012 63364 40068 63868
rect 40124 63858 40180 63868
rect 39900 63308 40068 63364
rect 40348 63700 40404 63710
rect 39116 63252 39172 63262
rect 39116 62578 39172 63196
rect 39452 63252 39508 63262
rect 39900 63252 39956 63308
rect 39452 63250 39956 63252
rect 39452 63198 39454 63250
rect 39506 63198 39956 63250
rect 39452 63196 39956 63198
rect 40236 63252 40292 63262
rect 39452 63186 39508 63196
rect 40236 63158 40292 63196
rect 40012 63140 40068 63150
rect 40012 63138 40180 63140
rect 40012 63086 40014 63138
rect 40066 63086 40180 63138
rect 40012 63084 40180 63086
rect 40012 63074 40068 63084
rect 39340 62914 39396 62926
rect 39340 62862 39342 62914
rect 39394 62862 39396 62914
rect 39340 62692 39396 62862
rect 39564 62916 39620 62926
rect 39564 62914 39732 62916
rect 39564 62862 39566 62914
rect 39618 62862 39732 62914
rect 39564 62860 39732 62862
rect 39564 62850 39620 62860
rect 39340 62636 39620 62692
rect 39116 62526 39118 62578
rect 39170 62526 39172 62578
rect 39116 62514 39172 62526
rect 39452 62468 39508 62478
rect 39452 62374 39508 62412
rect 39564 62356 39620 62636
rect 39676 62580 39732 62860
rect 40124 62692 40180 63084
rect 40348 62916 40404 63644
rect 40012 62580 40068 62590
rect 39676 62524 40012 62580
rect 39676 62356 39732 62366
rect 39788 62356 39844 62366
rect 39564 62354 39788 62356
rect 39564 62302 39678 62354
rect 39730 62302 39788 62354
rect 39564 62300 39788 62302
rect 39676 62290 39732 62300
rect 39788 61572 39844 62300
rect 40012 62354 40068 62524
rect 40012 62302 40014 62354
rect 40066 62302 40068 62354
rect 40012 62290 40068 62302
rect 39900 62244 39956 62282
rect 39900 62178 39956 62188
rect 40012 62132 40068 62142
rect 39900 61572 39956 61582
rect 39004 61516 39284 61572
rect 39788 61570 39956 61572
rect 39788 61518 39902 61570
rect 39954 61518 39956 61570
rect 39788 61516 39956 61518
rect 39004 61348 39060 61358
rect 38668 61346 39060 61348
rect 38668 61294 39006 61346
rect 39058 61294 39060 61346
rect 38668 61292 39060 61294
rect 38556 60676 38612 60686
rect 38668 60676 38724 61292
rect 39004 61282 39060 61292
rect 38892 60788 38948 60798
rect 38556 60674 38724 60676
rect 38556 60622 38558 60674
rect 38610 60622 38724 60674
rect 38556 60620 38724 60622
rect 38780 60786 38948 60788
rect 38780 60734 38894 60786
rect 38946 60734 38948 60786
rect 38780 60732 38948 60734
rect 38556 60610 38612 60620
rect 38444 60004 38500 60014
rect 38444 59668 38500 59948
rect 38556 59892 38612 59902
rect 38556 59798 38612 59836
rect 38444 59612 38612 59668
rect 38444 59332 38500 59342
rect 38444 59238 38500 59276
rect 38556 59330 38612 59612
rect 38556 59278 38558 59330
rect 38610 59278 38612 59330
rect 38556 59266 38612 59278
rect 38668 59220 38724 59230
rect 38668 59126 38724 59164
rect 38780 58996 38836 60732
rect 38892 60722 38948 60732
rect 39116 60788 39172 60798
rect 39116 60694 39172 60732
rect 39004 60676 39060 60686
rect 39004 60582 39060 60620
rect 39228 60564 39284 61516
rect 39900 61506 39956 61516
rect 39340 61346 39396 61358
rect 39340 61294 39342 61346
rect 39394 61294 39396 61346
rect 39340 60676 39396 61294
rect 40012 60900 40068 62076
rect 40124 61458 40180 62636
rect 40236 62860 40404 62916
rect 40236 61570 40292 62860
rect 40460 62804 40516 62814
rect 40348 62748 40460 62804
rect 40348 62466 40404 62748
rect 40460 62738 40516 62748
rect 40348 62414 40350 62466
rect 40402 62414 40404 62466
rect 40348 62402 40404 62414
rect 40572 61684 40628 61694
rect 40572 61590 40628 61628
rect 40236 61518 40238 61570
rect 40290 61518 40292 61570
rect 40236 61506 40292 61518
rect 40124 61406 40126 61458
rect 40178 61406 40180 61458
rect 40124 61394 40180 61406
rect 39900 60844 40068 60900
rect 39564 60788 39620 60798
rect 39564 60786 39732 60788
rect 39564 60734 39566 60786
rect 39618 60734 39732 60786
rect 39564 60732 39732 60734
rect 39564 60722 39620 60732
rect 39340 60610 39396 60620
rect 39116 60508 39284 60564
rect 39004 60004 39060 60014
rect 39116 60004 39172 60508
rect 39564 60116 39620 60126
rect 39060 59948 39172 60004
rect 39340 60114 39620 60116
rect 39340 60062 39566 60114
rect 39618 60062 39620 60114
rect 39340 60060 39620 60062
rect 39340 60002 39396 60060
rect 39564 60050 39620 60060
rect 39340 59950 39342 60002
rect 39394 59950 39396 60002
rect 39004 59938 39060 59948
rect 39340 59938 39396 59950
rect 39564 59780 39620 59790
rect 39564 59686 39620 59724
rect 39452 59668 39508 59678
rect 39340 59444 39396 59454
rect 38444 58940 38836 58996
rect 38892 59388 39340 59444
rect 38444 58434 38500 58940
rect 38444 58382 38446 58434
rect 38498 58382 38500 58434
rect 38444 58370 38500 58382
rect 38780 58210 38836 58222
rect 38780 58158 38782 58210
rect 38834 58158 38836 58210
rect 38780 57988 38836 58158
rect 38780 57922 38836 57932
rect 38556 57652 38612 57662
rect 38332 57650 38836 57652
rect 38332 57598 38558 57650
rect 38610 57598 38836 57650
rect 38332 57596 38836 57598
rect 37436 56754 37492 56766
rect 37436 56702 37438 56754
rect 37490 56702 37492 56754
rect 37436 53842 37492 56702
rect 37548 56642 37604 56654
rect 37548 56590 37550 56642
rect 37602 56590 37604 56642
rect 37548 54626 37604 56590
rect 37660 56644 37716 56654
rect 37716 56588 37828 56644
rect 37660 56578 37716 56588
rect 37772 55410 37828 56588
rect 37996 56642 38052 56654
rect 37996 56590 37998 56642
rect 38050 56590 38052 56642
rect 37996 56532 38052 56590
rect 38332 56644 38388 56654
rect 38332 56550 38388 56588
rect 37996 56466 38052 56476
rect 38556 56194 38612 57596
rect 38780 57540 38836 57596
rect 38780 57474 38836 57484
rect 38556 56142 38558 56194
rect 38610 56142 38612 56194
rect 38556 56130 38612 56142
rect 38668 56754 38724 56766
rect 38668 56702 38670 56754
rect 38722 56702 38724 56754
rect 37772 55358 37774 55410
rect 37826 55358 37828 55410
rect 37772 55346 37828 55358
rect 38668 55412 38724 56702
rect 38668 55346 38724 55356
rect 37548 54574 37550 54626
rect 37602 54574 37604 54626
rect 37548 54562 37604 54574
rect 37436 53790 37438 53842
rect 37490 53790 37492 53842
rect 37436 53778 37492 53790
rect 37884 53956 37940 53966
rect 37884 53730 37940 53900
rect 37884 53678 37886 53730
rect 37938 53678 37940 53730
rect 37884 53666 37940 53678
rect 38220 53732 38276 53742
rect 38220 53638 38276 53676
rect 37324 53508 37380 53518
rect 37324 53414 37380 53452
rect 37548 53506 37604 53518
rect 37548 53454 37550 53506
rect 37602 53454 37604 53506
rect 37212 53228 37380 53284
rect 36764 53172 36820 53182
rect 36764 53078 36820 53116
rect 37100 53060 37156 53070
rect 37100 52946 37156 53004
rect 37100 52894 37102 52946
rect 37154 52894 37156 52946
rect 37100 52882 37156 52894
rect 37212 52948 37268 52958
rect 37212 52854 37268 52892
rect 36764 51378 36820 51390
rect 36764 51326 36766 51378
rect 36818 51326 36820 51378
rect 36764 51268 36820 51326
rect 36764 51044 36820 51212
rect 37212 51266 37268 51278
rect 37212 51214 37214 51266
rect 37266 51214 37268 51266
rect 36764 50988 37156 51044
rect 36652 50876 36932 50932
rect 36540 50820 36596 50830
rect 36540 50818 36820 50820
rect 36540 50766 36542 50818
rect 36594 50766 36820 50818
rect 36540 50764 36820 50766
rect 36540 50754 36596 50764
rect 35868 50542 35870 50594
rect 35922 50542 35924 50594
rect 35868 50530 35924 50542
rect 36092 50540 36260 50596
rect 34300 50372 34580 50428
rect 36092 50372 36148 50540
rect 36204 50372 36260 50382
rect 34300 48916 34356 48926
rect 34300 48356 34356 48860
rect 34412 48802 34468 48814
rect 34412 48750 34414 48802
rect 34466 48750 34468 48802
rect 34412 48580 34468 48750
rect 34524 48692 34580 50372
rect 35980 50370 36260 50372
rect 35980 50318 36206 50370
rect 36258 50318 36260 50370
rect 35980 50316 36260 50318
rect 35196 49924 35252 49934
rect 35084 49922 35252 49924
rect 35084 49870 35198 49922
rect 35250 49870 35252 49922
rect 35084 49868 35252 49870
rect 34748 49700 34804 49710
rect 35084 49700 35140 49868
rect 35196 49858 35252 49868
rect 35308 49812 35364 49822
rect 35308 49718 35364 49756
rect 34748 49698 35140 49700
rect 34748 49646 34750 49698
rect 34802 49646 35140 49698
rect 34748 49644 35140 49646
rect 35868 49698 35924 49710
rect 35868 49646 35870 49698
rect 35922 49646 35924 49698
rect 34636 49028 34692 49038
rect 34636 48934 34692 48972
rect 34748 48804 34804 49644
rect 35196 49588 35252 49598
rect 35868 49588 35924 49646
rect 35084 49586 35252 49588
rect 35084 49534 35198 49586
rect 35250 49534 35252 49586
rect 35084 49532 35252 49534
rect 34748 48738 34804 48748
rect 34972 48802 35028 48814
rect 34972 48750 34974 48802
rect 35026 48750 35028 48802
rect 34524 48636 34692 48692
rect 34636 48580 34692 48636
rect 34636 48524 34804 48580
rect 34412 48514 34468 48524
rect 34748 48356 34804 48524
rect 34300 48300 34468 48356
rect 34300 48130 34356 48142
rect 34300 48078 34302 48130
rect 34354 48078 34356 48130
rect 34300 47684 34356 48078
rect 34300 47618 34356 47628
rect 34300 47460 34356 47470
rect 34412 47460 34468 48300
rect 34300 47458 34468 47460
rect 34300 47406 34302 47458
rect 34354 47406 34468 47458
rect 34300 47404 34468 47406
rect 34524 48300 34804 48356
rect 34300 47394 34356 47404
rect 34188 46946 34244 46956
rect 34412 47236 34468 47246
rect 34076 46694 34132 46732
rect 34188 46676 34244 46686
rect 34188 46582 34244 46620
rect 34076 45892 34132 45902
rect 34132 45836 34244 45892
rect 34076 45826 34132 45836
rect 33964 45378 34020 45388
rect 33964 45220 34020 45230
rect 33964 45126 34020 45164
rect 34076 45106 34132 45118
rect 34076 45054 34078 45106
rect 34130 45054 34132 45106
rect 34076 44436 34132 45054
rect 34188 44772 34244 45836
rect 34188 44706 34244 44716
rect 34412 44548 34468 47180
rect 34412 44482 34468 44492
rect 34076 44370 34132 44380
rect 34524 44436 34580 48300
rect 34636 48230 34692 48242
rect 34636 48178 34638 48230
rect 34690 48178 34692 48230
rect 34636 47124 34692 48178
rect 34748 48020 34804 48030
rect 34748 47346 34804 47964
rect 34972 47460 35028 48750
rect 35084 47460 35140 49532
rect 35196 49522 35252 49532
rect 35644 49532 35924 49588
rect 35196 49420 35460 49430
rect 35252 49364 35300 49420
rect 35356 49364 35404 49420
rect 35196 49354 35460 49364
rect 35644 48804 35700 49532
rect 35980 49476 36036 50316
rect 36204 50306 36260 50316
rect 36428 50370 36484 50382
rect 36428 50318 36430 50370
rect 36482 50318 36484 50370
rect 35868 49420 36036 49476
rect 36204 49924 36260 49934
rect 36428 49924 36484 50318
rect 36540 50036 36596 50046
rect 36540 49942 36596 49980
rect 36204 49922 36484 49924
rect 36204 49870 36206 49922
rect 36258 49870 36484 49922
rect 36204 49868 36484 49870
rect 35756 49028 35812 49038
rect 35756 48934 35812 48972
rect 35868 49026 35924 49420
rect 35868 48974 35870 49026
rect 35922 48974 35924 49026
rect 35868 48962 35924 48974
rect 36204 49028 36260 49868
rect 36764 49810 36820 50764
rect 36764 49758 36766 49810
rect 36818 49758 36820 49810
rect 36764 49746 36820 49758
rect 36876 49588 36932 50876
rect 36988 50820 37044 50830
rect 36988 50594 37044 50764
rect 36988 50542 36990 50594
rect 37042 50542 37044 50594
rect 36988 50530 37044 50542
rect 37100 50482 37156 50988
rect 37212 50820 37268 51214
rect 37212 50754 37268 50764
rect 37100 50430 37102 50482
rect 37154 50430 37156 50482
rect 37100 50418 37156 50430
rect 36204 48962 36260 48972
rect 36316 49532 36932 49588
rect 37100 49812 37156 49822
rect 35980 48914 36036 48926
rect 35980 48862 35982 48914
rect 36034 48862 36036 48914
rect 35980 48804 36036 48862
rect 35644 48748 36036 48804
rect 35420 48132 35476 48142
rect 35756 48132 35812 48142
rect 35420 48130 35588 48132
rect 35420 48078 35422 48130
rect 35474 48078 35588 48130
rect 35420 48076 35588 48078
rect 35420 48066 35476 48076
rect 35196 47852 35460 47862
rect 35252 47796 35300 47852
rect 35356 47796 35404 47852
rect 35196 47786 35460 47796
rect 35196 47460 35252 47470
rect 35532 47460 35588 48076
rect 35084 47458 35252 47460
rect 35084 47406 35198 47458
rect 35250 47406 35252 47458
rect 35084 47404 35252 47406
rect 34972 47394 35028 47404
rect 35196 47394 35252 47404
rect 35420 47404 35588 47460
rect 35756 47458 35812 48076
rect 35980 47684 36036 48748
rect 35980 47618 36036 47628
rect 36204 48580 36260 48590
rect 35756 47406 35758 47458
rect 35810 47406 35812 47458
rect 34748 47294 34750 47346
rect 34802 47294 34804 47346
rect 34748 47282 34804 47294
rect 34972 47236 35028 47246
rect 34972 47142 35028 47180
rect 35084 47236 35140 47246
rect 35420 47236 35476 47404
rect 35756 47394 35812 47406
rect 36204 47458 36260 48524
rect 36204 47406 36206 47458
rect 36258 47406 36260 47458
rect 35084 47234 35476 47236
rect 35084 47182 35086 47234
rect 35138 47182 35476 47234
rect 35084 47180 35476 47182
rect 35532 47234 35588 47246
rect 35532 47182 35534 47234
rect 35586 47182 35588 47234
rect 35084 47170 35140 47180
rect 34636 47068 34916 47124
rect 34636 46674 34692 46686
rect 34636 46622 34638 46674
rect 34690 46622 34692 46674
rect 34636 46564 34692 46622
rect 34636 46498 34692 46508
rect 34748 46562 34804 46574
rect 34748 46510 34750 46562
rect 34802 46510 34804 46562
rect 34636 45892 34692 45902
rect 34636 45798 34692 45836
rect 34636 45444 34692 45454
rect 34636 45330 34692 45388
rect 34636 45278 34638 45330
rect 34690 45278 34692 45330
rect 34636 45266 34692 45278
rect 34748 45332 34804 46510
rect 34748 45266 34804 45276
rect 34860 45220 34916 47068
rect 34972 46788 35028 46798
rect 34972 46694 35028 46732
rect 35196 46676 35252 46686
rect 35196 46582 35252 46620
rect 35196 46284 35460 46294
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35196 46218 35460 46228
rect 35420 46004 35476 46014
rect 35308 45948 35420 46004
rect 35308 45890 35364 45948
rect 35420 45938 35476 45948
rect 35308 45838 35310 45890
rect 35362 45838 35364 45890
rect 35308 45826 35364 45838
rect 34972 45780 35028 45790
rect 34972 45686 35028 45724
rect 35532 45778 35588 47182
rect 35644 47234 35700 47246
rect 35644 47182 35646 47234
rect 35698 47182 35700 47234
rect 35644 46900 35700 47182
rect 35756 46900 35812 46910
rect 35644 46898 35812 46900
rect 35644 46846 35758 46898
rect 35810 46846 35812 46898
rect 35644 46844 35812 46846
rect 35756 46834 35812 46844
rect 36204 46900 36260 47406
rect 35980 46674 36036 46686
rect 35980 46622 35982 46674
rect 36034 46622 36036 46674
rect 35868 46564 35924 46574
rect 35532 45726 35534 45778
rect 35586 45726 35588 45778
rect 35308 45668 35364 45678
rect 35308 45574 35364 45612
rect 35532 45556 35588 45726
rect 35532 45490 35588 45500
rect 35644 46562 35924 46564
rect 35644 46510 35870 46562
rect 35922 46510 35924 46562
rect 35644 46508 35924 46510
rect 34972 45220 35028 45230
rect 34860 45164 34972 45220
rect 34860 45106 34916 45164
rect 34972 45154 35028 45164
rect 35644 45218 35700 46508
rect 35868 46498 35924 46508
rect 35868 46116 35924 46126
rect 35980 46116 36036 46622
rect 36204 46340 36260 46844
rect 36204 46274 36260 46284
rect 35868 46114 36036 46116
rect 35868 46062 35870 46114
rect 35922 46062 36036 46114
rect 35868 46060 36036 46062
rect 35868 46050 35924 46060
rect 35644 45166 35646 45218
rect 35698 45166 35700 45218
rect 35644 45154 35700 45166
rect 35868 45892 35924 45902
rect 34860 45054 34862 45106
rect 34914 45054 34916 45106
rect 34860 45042 34916 45054
rect 35196 44716 35460 44726
rect 34524 44342 34580 44380
rect 34972 44660 35028 44670
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35196 44650 35460 44660
rect 34076 44100 34132 44110
rect 33964 44098 34132 44100
rect 33964 44046 34078 44098
rect 34130 44046 34132 44098
rect 33964 44044 34132 44046
rect 33964 43876 34020 44044
rect 34076 44034 34132 44044
rect 33964 43810 34020 43820
rect 33964 43650 34020 43662
rect 33964 43598 33966 43650
rect 34018 43598 34020 43650
rect 33964 43540 34020 43598
rect 34748 43540 34804 43550
rect 33964 43538 34804 43540
rect 33964 43486 34750 43538
rect 34802 43486 34804 43538
rect 33964 43484 34804 43486
rect 34412 43426 34468 43484
rect 34748 43474 34804 43484
rect 34412 43374 34414 43426
rect 34466 43374 34468 43426
rect 34076 43204 34132 43214
rect 33852 42700 34020 42756
rect 33628 42662 33684 42700
rect 33404 42644 33460 42654
rect 33404 42550 33460 42588
rect 33852 42530 33908 42542
rect 33852 42478 33854 42530
rect 33906 42478 33908 42530
rect 33292 41906 33348 41916
rect 33404 41970 33460 41982
rect 33404 41918 33406 41970
rect 33458 41918 33460 41970
rect 33404 41524 33460 41918
rect 33404 41188 33460 41468
rect 33404 41122 33460 41132
rect 33852 40402 33908 42478
rect 33964 41858 34020 42700
rect 34076 42754 34132 43148
rect 34076 42702 34078 42754
rect 34130 42702 34132 42754
rect 34076 42690 34132 42702
rect 34188 42754 34244 42766
rect 34188 42702 34190 42754
rect 34242 42702 34244 42754
rect 34188 42644 34244 42702
rect 34188 42578 34244 42588
rect 34412 42420 34468 43374
rect 34636 42756 34692 42766
rect 34636 42662 34692 42700
rect 34972 42754 35028 44604
rect 35868 44436 35924 45836
rect 36204 45890 36260 45902
rect 36204 45838 36206 45890
rect 36258 45838 36260 45890
rect 36204 45556 36260 45838
rect 36204 45490 36260 45500
rect 35868 44342 35924 44380
rect 35308 44324 35364 44334
rect 35084 44212 35140 44222
rect 35084 44118 35140 44156
rect 35308 43876 35364 44268
rect 35308 43810 35364 43820
rect 35980 43652 36036 43662
rect 35980 43558 36036 43596
rect 35756 43538 35812 43550
rect 35756 43486 35758 43538
rect 35810 43486 35812 43538
rect 35196 43428 35252 43438
rect 35196 43334 35252 43372
rect 35196 43148 35460 43158
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35196 43082 35460 43092
rect 35756 42868 35812 43486
rect 36204 43316 36260 43326
rect 36092 43314 36260 43316
rect 36092 43262 36206 43314
rect 36258 43262 36260 43314
rect 36092 43260 36260 43262
rect 36092 42868 36148 43260
rect 36204 43250 36260 43260
rect 35756 42812 36148 42868
rect 34972 42702 34974 42754
rect 35026 42702 35028 42754
rect 34748 42532 34804 42542
rect 33964 41806 33966 41858
rect 34018 41806 34020 41858
rect 33964 41524 34020 41806
rect 33964 41458 34020 41468
rect 34188 42364 34468 42420
rect 34524 42530 34804 42532
rect 34524 42478 34750 42530
rect 34802 42478 34804 42530
rect 34524 42476 34804 42478
rect 34188 41188 34244 42364
rect 34188 41122 34244 41132
rect 34300 41970 34356 41982
rect 34300 41918 34302 41970
rect 34354 41918 34356 41970
rect 34300 40964 34356 41918
rect 34412 41410 34468 41422
rect 34412 41358 34414 41410
rect 34466 41358 34468 41410
rect 34412 41298 34468 41358
rect 34524 41412 34580 42476
rect 34748 42466 34804 42476
rect 34860 41972 34916 41982
rect 34860 41878 34916 41916
rect 34524 41356 34916 41412
rect 34412 41246 34414 41298
rect 34466 41246 34468 41298
rect 34412 41234 34468 41246
rect 34300 40898 34356 40908
rect 34748 40964 34804 40974
rect 34748 40870 34804 40908
rect 34748 40628 34804 40638
rect 34188 40516 34244 40526
rect 34188 40422 34244 40460
rect 33852 40350 33854 40402
rect 33906 40350 33908 40402
rect 33852 40338 33908 40350
rect 33964 40404 34020 40414
rect 33964 40310 34020 40348
rect 34412 40404 34468 40414
rect 34412 40310 34468 40348
rect 34748 40404 34804 40572
rect 34076 40290 34132 40302
rect 34076 40238 34078 40290
rect 34130 40238 34132 40290
rect 33964 39732 34020 39742
rect 34076 39732 34132 40238
rect 33964 39730 34132 39732
rect 33964 39678 33966 39730
rect 34018 39678 34132 39730
rect 33964 39676 34132 39678
rect 33964 39666 34020 39676
rect 33292 39618 33348 39630
rect 33292 39566 33294 39618
rect 33346 39566 33348 39618
rect 33292 38722 33348 39566
rect 33292 38670 33294 38722
rect 33346 38670 33348 38722
rect 32956 38612 33236 38668
rect 32172 36430 32174 36482
rect 32226 36430 32228 36482
rect 32172 36418 32228 36430
rect 32060 35086 32062 35138
rect 32114 35086 32116 35138
rect 32060 35074 32116 35086
rect 32508 35586 32564 35598
rect 32508 35534 32510 35586
rect 32562 35534 32564 35586
rect 32508 35476 32564 35534
rect 32508 34914 32564 35420
rect 32508 34862 32510 34914
rect 32562 34862 32564 34914
rect 32508 34850 32564 34862
rect 31948 34804 32004 34814
rect 31948 34710 32004 34748
rect 32060 34690 32116 34702
rect 32060 34638 32062 34690
rect 32114 34638 32116 34690
rect 31724 34354 31892 34356
rect 31724 34302 31726 34354
rect 31778 34302 31892 34354
rect 31724 34300 31892 34302
rect 31724 34290 31780 34300
rect 31500 33628 31668 33684
rect 31500 33460 31556 33470
rect 31500 33346 31556 33404
rect 31500 33294 31502 33346
rect 31554 33294 31556 33346
rect 31500 33282 31556 33294
rect 31612 32788 31668 33628
rect 31836 33572 31892 34300
rect 32060 34020 32116 34638
rect 32620 34244 32676 34254
rect 32060 33954 32116 33964
rect 32396 34020 32452 34030
rect 32396 33926 32452 33964
rect 31892 33516 32228 33572
rect 31836 33478 31892 33516
rect 32172 33234 32228 33516
rect 32620 33460 32676 34188
rect 32620 33366 32676 33404
rect 32172 33182 32174 33234
rect 32226 33182 32228 33234
rect 31836 33122 31892 33134
rect 31836 33070 31838 33122
rect 31890 33070 31892 33122
rect 31388 32386 31444 32396
rect 31500 32732 31668 32788
rect 31724 32900 31780 32910
rect 31500 32004 31556 32732
rect 31612 32562 31668 32574
rect 31612 32510 31614 32562
rect 31666 32510 31668 32562
rect 31612 32452 31668 32510
rect 31612 32386 31668 32396
rect 31500 31948 31668 32004
rect 31500 31780 31556 31790
rect 31500 31220 31556 31724
rect 31500 31126 31556 31164
rect 31276 31042 31332 31052
rect 31164 30996 31220 31006
rect 31164 30902 31220 30940
rect 31164 30322 31220 30334
rect 31164 30270 31166 30322
rect 31218 30270 31220 30322
rect 31164 30212 31220 30270
rect 31164 30146 31220 30156
rect 31276 30210 31332 30222
rect 31276 30158 31278 30210
rect 31330 30158 31332 30210
rect 30604 28644 30660 28654
rect 30604 28550 30660 28588
rect 31052 28642 31108 29372
rect 31276 29650 31332 30158
rect 31276 29598 31278 29650
rect 31330 29598 31332 29650
rect 31276 28868 31332 29598
rect 31388 30098 31444 30110
rect 31388 30046 31390 30098
rect 31442 30046 31444 30098
rect 31388 29540 31444 30046
rect 31612 29764 31668 31948
rect 31612 29698 31668 29708
rect 31724 30100 31780 32844
rect 31836 32676 31892 33070
rect 32172 32788 32228 33182
rect 32172 32722 32228 32732
rect 32284 33348 32340 33358
rect 31892 32620 32116 32676
rect 31836 32610 31892 32620
rect 32060 32004 32116 32620
rect 32172 32564 32228 32574
rect 32284 32564 32340 33292
rect 32228 32508 32340 32564
rect 32172 32470 32228 32508
rect 32060 31220 32116 31948
rect 32172 31220 32228 31230
rect 32060 31218 32228 31220
rect 32060 31166 32174 31218
rect 32226 31166 32228 31218
rect 32060 31164 32228 31166
rect 32172 31154 32228 31164
rect 31836 31106 31892 31118
rect 31836 31054 31838 31106
rect 31890 31054 31892 31106
rect 31836 30324 31892 31054
rect 32508 31108 32564 31118
rect 32508 31106 32676 31108
rect 32508 31054 32510 31106
rect 32562 31054 32676 31106
rect 32508 31052 32676 31054
rect 32508 31042 32564 31052
rect 32620 30548 32676 31052
rect 31836 30258 31892 30268
rect 32396 30492 32676 30548
rect 31724 29652 31780 30044
rect 32060 30210 32116 30222
rect 32060 30158 32062 30210
rect 32114 30158 32116 30210
rect 31724 29596 31892 29652
rect 31500 29540 31556 29550
rect 31388 29484 31500 29540
rect 31556 29484 31780 29540
rect 31500 29446 31556 29484
rect 31388 29316 31444 29326
rect 31388 29222 31444 29260
rect 31388 28868 31444 28878
rect 31276 28866 31556 28868
rect 31276 28814 31390 28866
rect 31442 28814 31556 28866
rect 31276 28812 31556 28814
rect 31388 28802 31444 28812
rect 31164 28756 31220 28766
rect 31164 28662 31220 28700
rect 31052 28590 31054 28642
rect 31106 28590 31108 28642
rect 31052 28578 31108 28590
rect 30940 28532 30996 28542
rect 30604 28084 30660 28094
rect 30604 27990 30660 28028
rect 30940 26908 30996 28476
rect 31164 28420 31220 28430
rect 31164 28082 31220 28364
rect 31164 28030 31166 28082
rect 31218 28030 31220 28082
rect 31164 28018 31220 28030
rect 31500 27858 31556 28812
rect 31500 27806 31502 27858
rect 31554 27806 31556 27858
rect 31500 27794 31556 27806
rect 31724 27858 31780 29484
rect 31836 29426 31892 29596
rect 31836 29374 31838 29426
rect 31890 29374 31892 29426
rect 31836 29362 31892 29374
rect 31948 29428 32004 29438
rect 31948 28084 32004 29372
rect 32060 28868 32116 30158
rect 32284 29652 32340 29662
rect 32284 29558 32340 29596
rect 32172 29428 32228 29438
rect 32172 29334 32228 29372
rect 32284 29202 32340 29214
rect 32284 29150 32286 29202
rect 32338 29150 32340 29202
rect 32060 28812 32228 28868
rect 32172 28420 32228 28812
rect 32284 28644 32340 29150
rect 32396 28756 32452 30492
rect 32620 30436 32676 30492
rect 32620 30370 32676 30380
rect 32508 30324 32564 30334
rect 32508 30212 32564 30268
rect 32508 30210 32676 30212
rect 32508 30158 32510 30210
rect 32562 30158 32676 30210
rect 32508 30156 32676 30158
rect 32508 30146 32564 30156
rect 32396 28700 32564 28756
rect 32284 28578 32340 28588
rect 32396 28530 32452 28542
rect 32396 28478 32398 28530
rect 32450 28478 32452 28530
rect 32284 28420 32340 28430
rect 32172 28418 32340 28420
rect 32172 28366 32286 28418
rect 32338 28366 32340 28418
rect 32172 28364 32340 28366
rect 32284 28354 32340 28364
rect 32172 28196 32228 28206
rect 32060 28084 32116 28094
rect 31948 28082 32116 28084
rect 31948 28030 32062 28082
rect 32114 28030 32116 28082
rect 31948 28028 32116 28030
rect 31724 27806 31726 27858
rect 31778 27806 31780 27858
rect 31724 27794 31780 27806
rect 32060 27186 32116 28028
rect 32060 27134 32062 27186
rect 32114 27134 32116 27186
rect 32060 27122 32116 27134
rect 32172 26908 32228 28140
rect 32284 27972 32340 27982
rect 32284 27878 32340 27916
rect 32396 27746 32452 28478
rect 32508 28084 32564 28700
rect 32620 28308 32676 30156
rect 32732 29988 32788 38612
rect 32956 36372 33012 36382
rect 32956 36278 33012 36316
rect 33180 35810 33236 38612
rect 33292 38612 33348 38670
rect 33292 38546 33348 38556
rect 33852 38276 33908 38286
rect 33852 38182 33908 38220
rect 34636 38276 34692 38286
rect 33516 38164 33572 38174
rect 33964 38164 34020 38174
rect 33572 38108 33684 38164
rect 33516 38070 33572 38108
rect 33628 37490 33684 38108
rect 33964 38070 34020 38108
rect 33628 37438 33630 37490
rect 33682 37438 33684 37490
rect 33628 37426 33684 37438
rect 33852 38052 33908 38062
rect 33516 36372 33572 36382
rect 33516 35922 33572 36316
rect 33516 35870 33518 35922
rect 33570 35870 33572 35922
rect 33516 35858 33572 35870
rect 33628 36036 33684 36046
rect 33628 35922 33684 35980
rect 33628 35870 33630 35922
rect 33682 35870 33684 35922
rect 33628 35858 33684 35870
rect 33740 35924 33796 35934
rect 33740 35830 33796 35868
rect 33180 35758 33182 35810
rect 33234 35758 33236 35810
rect 33180 35746 33236 35758
rect 33404 35700 33460 35710
rect 33292 35698 33460 35700
rect 33292 35646 33406 35698
rect 33458 35646 33460 35698
rect 33292 35644 33460 35646
rect 33180 35476 33236 35486
rect 33068 35420 33180 35476
rect 32844 34690 32900 34702
rect 32844 34638 32846 34690
rect 32898 34638 32900 34690
rect 32844 33236 32900 34638
rect 33068 34132 33124 35420
rect 33180 35410 33236 35420
rect 33292 35138 33348 35644
rect 33404 35634 33460 35644
rect 33292 35086 33294 35138
rect 33346 35086 33348 35138
rect 33292 35074 33348 35086
rect 33852 34916 33908 37996
rect 33740 34860 33908 34916
rect 33964 37940 34020 37950
rect 33180 34804 33236 34814
rect 33180 34710 33236 34748
rect 33292 34692 33348 34702
rect 33292 34244 33348 34636
rect 33292 34188 33572 34244
rect 33068 34076 33348 34132
rect 33292 34018 33348 34076
rect 33292 33966 33294 34018
rect 33346 33966 33348 34018
rect 33292 33954 33348 33966
rect 32844 33170 32900 33180
rect 33180 32562 33236 32574
rect 33180 32510 33182 32562
rect 33234 32510 33236 32562
rect 33068 31556 33124 31566
rect 33068 30994 33124 31500
rect 33068 30942 33070 30994
rect 33122 30942 33124 30994
rect 33068 30930 33124 30942
rect 33068 30324 33124 30334
rect 33180 30324 33236 32510
rect 33124 30268 33236 30324
rect 33292 32004 33348 32014
rect 33068 30258 33124 30268
rect 32956 30210 33012 30222
rect 33292 30212 33348 31948
rect 32956 30158 32958 30210
rect 33010 30158 33012 30210
rect 32956 30100 33012 30158
rect 33180 30156 33348 30212
rect 33404 31220 33460 31230
rect 33404 30212 33460 31164
rect 32956 30044 33124 30100
rect 32732 29932 33012 29988
rect 32732 29764 32788 29774
rect 32732 28644 32788 29708
rect 32732 28530 32788 28588
rect 32732 28478 32734 28530
rect 32786 28478 32788 28530
rect 32732 28466 32788 28478
rect 32844 29652 32900 29662
rect 32844 28530 32900 29596
rect 32844 28478 32846 28530
rect 32898 28478 32900 28530
rect 32844 28466 32900 28478
rect 32620 28242 32676 28252
rect 32956 28196 33012 29932
rect 33068 29876 33124 30044
rect 33068 29810 33124 29820
rect 33180 29650 33236 30156
rect 33404 30118 33460 30156
rect 33180 29598 33182 29650
rect 33234 29598 33236 29650
rect 33180 29586 33236 29598
rect 33068 28420 33124 28430
rect 33068 28418 33460 28420
rect 33068 28366 33070 28418
rect 33122 28366 33460 28418
rect 33068 28364 33460 28366
rect 33068 28354 33124 28364
rect 32956 28140 33236 28196
rect 32508 28028 33012 28084
rect 32396 27694 32398 27746
rect 32450 27694 32452 27746
rect 32396 27682 32452 27694
rect 32508 27858 32564 27870
rect 32508 27806 32510 27858
rect 32562 27806 32564 27858
rect 32508 27188 32564 27806
rect 32508 27094 32564 27132
rect 32620 27860 32676 27870
rect 30380 26852 30772 26908
rect 30940 26852 31108 26908
rect 30492 25396 30548 25406
rect 30380 25340 30492 25396
rect 30268 24724 30324 24734
rect 30268 24630 30324 24668
rect 30156 22978 30212 22988
rect 30268 22372 30324 22382
rect 30380 22372 30436 25340
rect 30492 25330 30548 25340
rect 30716 23380 30772 26852
rect 31052 25282 31108 26852
rect 32060 26852 32228 26908
rect 31276 25508 31332 25518
rect 31052 25230 31054 25282
rect 31106 25230 31108 25282
rect 31052 25060 31108 25230
rect 31052 24994 31108 25004
rect 31164 25506 31332 25508
rect 31164 25454 31278 25506
rect 31330 25454 31332 25506
rect 31164 25452 31332 25454
rect 31164 24722 31220 25452
rect 31276 25442 31332 25452
rect 31724 25396 31780 25406
rect 31724 25302 31780 25340
rect 31724 25060 31780 25070
rect 31164 24670 31166 24722
rect 31218 24670 31220 24722
rect 31164 23716 31220 24670
rect 31500 24836 31556 24846
rect 31500 24612 31556 24780
rect 31500 24610 31668 24612
rect 31500 24558 31502 24610
rect 31554 24558 31668 24610
rect 31500 24556 31668 24558
rect 31500 24546 31556 24556
rect 31164 23650 31220 23660
rect 30268 22370 30436 22372
rect 30268 22318 30270 22370
rect 30322 22318 30436 22370
rect 30268 22316 30436 22318
rect 30268 22306 30324 22316
rect 30268 22036 30324 22046
rect 29708 20178 29764 20188
rect 30044 21476 30100 21486
rect 29708 19124 29764 19134
rect 29708 19122 29876 19124
rect 29708 19070 29710 19122
rect 29762 19070 29876 19122
rect 29708 19068 29876 19070
rect 29708 19058 29764 19068
rect 29596 19012 29652 19022
rect 29596 18918 29652 18956
rect 29708 18564 29764 18574
rect 29708 18450 29764 18508
rect 29708 18398 29710 18450
rect 29762 18398 29764 18450
rect 29708 18386 29764 18398
rect 29820 17556 29876 19068
rect 29932 19122 29988 19134
rect 29932 19070 29934 19122
rect 29986 19070 29988 19122
rect 29932 17780 29988 19070
rect 29932 17714 29988 17724
rect 30044 17778 30100 21420
rect 30268 21026 30324 21980
rect 30268 20974 30270 21026
rect 30322 20974 30324 21026
rect 30268 20962 30324 20974
rect 30380 21252 30436 22316
rect 30492 23324 30772 23380
rect 30492 21698 30548 23324
rect 30828 23044 30884 23054
rect 30492 21646 30494 21698
rect 30546 21646 30548 21698
rect 30492 21588 30548 21646
rect 30716 22484 30772 22494
rect 30716 22370 30772 22428
rect 30716 22318 30718 22370
rect 30770 22318 30772 22370
rect 30492 21522 30548 21532
rect 30604 21586 30660 21598
rect 30604 21534 30606 21586
rect 30658 21534 30660 21586
rect 30604 21476 30660 21534
rect 30604 21410 30660 21420
rect 30492 21364 30548 21374
rect 30492 21270 30548 21308
rect 30156 20804 30212 20814
rect 30380 20804 30436 21196
rect 30156 20802 30436 20804
rect 30156 20750 30158 20802
rect 30210 20750 30436 20802
rect 30156 20748 30436 20750
rect 30156 20738 30212 20748
rect 30716 20244 30772 22318
rect 30828 22372 30884 22988
rect 31052 23042 31108 23054
rect 31052 22990 31054 23042
rect 31106 22990 31108 23042
rect 30828 20802 30884 22316
rect 30940 22594 30996 22606
rect 30940 22542 30942 22594
rect 30994 22542 30996 22594
rect 30940 21698 30996 22542
rect 31052 21810 31108 22990
rect 31052 21758 31054 21810
rect 31106 21758 31108 21810
rect 31052 21746 31108 21758
rect 31164 22708 31220 22718
rect 31164 22482 31220 22652
rect 31164 22430 31166 22482
rect 31218 22430 31220 22482
rect 31164 21812 31220 22430
rect 30940 21646 30942 21698
rect 30994 21646 30996 21698
rect 30940 21634 30996 21646
rect 30828 20750 30830 20802
rect 30882 20750 30884 20802
rect 30828 20738 30884 20750
rect 31052 20804 31108 20814
rect 31164 20804 31220 21756
rect 31500 21588 31556 21598
rect 31612 21588 31668 24556
rect 31724 22370 31780 25004
rect 31948 24724 32004 24734
rect 31948 23940 32004 24668
rect 32060 24722 32116 26852
rect 32172 25506 32228 25518
rect 32172 25454 32174 25506
rect 32226 25454 32228 25506
rect 32172 25396 32228 25454
rect 32172 25330 32228 25340
rect 32060 24670 32062 24722
rect 32114 24670 32116 24722
rect 32060 24388 32116 24670
rect 32396 24612 32452 24622
rect 32396 24518 32452 24556
rect 32060 24332 32564 24388
rect 31724 22318 31726 22370
rect 31778 22318 31780 22370
rect 31724 22306 31780 22318
rect 31836 23938 32004 23940
rect 31836 23886 31950 23938
rect 32002 23886 32004 23938
rect 31836 23884 32004 23886
rect 31836 23268 31892 23884
rect 31948 23874 32004 23884
rect 31836 23154 31892 23212
rect 31836 23102 31838 23154
rect 31890 23102 31892 23154
rect 31836 22148 31892 23102
rect 31836 22082 31892 22092
rect 32284 23828 32340 23838
rect 32284 22370 32340 23772
rect 32284 22318 32286 22370
rect 32338 22318 32340 22370
rect 31612 21532 31892 21588
rect 31500 21474 31556 21532
rect 31500 21422 31502 21474
rect 31554 21422 31556 21474
rect 31500 21364 31556 21422
rect 31500 21308 31780 21364
rect 31052 20802 31220 20804
rect 31052 20750 31054 20802
rect 31106 20750 31220 20802
rect 31052 20748 31220 20750
rect 31500 20802 31556 20814
rect 31500 20750 31502 20802
rect 31554 20750 31556 20802
rect 31052 20738 31108 20748
rect 31500 20580 31556 20750
rect 31500 20514 31556 20524
rect 30604 20188 30772 20244
rect 31276 20244 31332 20254
rect 30380 20020 30436 20030
rect 30268 19964 30380 20020
rect 30268 19234 30324 19964
rect 30380 19954 30436 19964
rect 30604 19908 30660 20188
rect 31164 20020 31220 20030
rect 31164 19926 31220 19964
rect 30604 19852 30772 19908
rect 30268 19182 30270 19234
rect 30322 19182 30324 19234
rect 30268 19170 30324 19182
rect 30380 19010 30436 19022
rect 30380 18958 30382 19010
rect 30434 18958 30436 19010
rect 30380 18564 30436 18958
rect 30492 19012 30548 19022
rect 30492 18918 30548 18956
rect 30380 18498 30436 18508
rect 30044 17726 30046 17778
rect 30098 17726 30100 17778
rect 29820 17490 29876 17500
rect 30044 17444 30100 17726
rect 30268 18452 30324 18462
rect 30268 17666 30324 18396
rect 30268 17614 30270 17666
rect 30322 17614 30324 17666
rect 30268 17602 30324 17614
rect 30044 17388 30660 17444
rect 30268 17220 30324 17230
rect 30268 17106 30324 17164
rect 30268 17054 30270 17106
rect 30322 17054 30324 17106
rect 30268 17042 30324 17054
rect 30604 16884 30660 17388
rect 30604 16770 30660 16828
rect 30604 16718 30606 16770
rect 30658 16718 30660 16770
rect 30604 16706 30660 16718
rect 30044 16660 30100 16670
rect 30044 16210 30100 16604
rect 30044 16158 30046 16210
rect 30098 16158 30100 16210
rect 29596 15764 29652 15774
rect 29596 15538 29652 15708
rect 30044 15652 30100 16158
rect 30604 16212 30660 16222
rect 30604 16118 30660 16156
rect 29596 15486 29598 15538
rect 29650 15486 29652 15538
rect 29596 13636 29652 15486
rect 29820 15596 30044 15652
rect 29820 15426 29876 15596
rect 30044 15586 30100 15596
rect 29820 15374 29822 15426
rect 29874 15374 29876 15426
rect 29820 15362 29876 15374
rect 29932 15426 29988 15438
rect 29932 15374 29934 15426
rect 29986 15374 29988 15426
rect 29932 15148 29988 15374
rect 30156 15316 30212 15326
rect 30492 15316 30548 15326
rect 30156 15314 30548 15316
rect 30156 15262 30158 15314
rect 30210 15262 30494 15314
rect 30546 15262 30548 15314
rect 30156 15260 30548 15262
rect 30156 15250 30212 15260
rect 30492 15250 30548 15260
rect 30716 15148 30772 19852
rect 31276 19348 31332 20188
rect 31388 20130 31444 20142
rect 31388 20078 31390 20130
rect 31442 20078 31444 20130
rect 31388 19908 31444 20078
rect 31724 20132 31780 21308
rect 31500 20020 31556 20030
rect 31500 20018 31668 20020
rect 31500 19966 31502 20018
rect 31554 19966 31668 20018
rect 31500 19964 31668 19966
rect 31500 19954 31556 19964
rect 31388 19842 31444 19852
rect 31276 19292 31556 19348
rect 30940 19236 30996 19246
rect 31164 19236 31220 19246
rect 30940 19234 31220 19236
rect 30940 19182 30942 19234
rect 30994 19182 31166 19234
rect 31218 19182 31220 19234
rect 30940 19180 31220 19182
rect 30940 19170 30996 19180
rect 31164 19170 31220 19180
rect 31500 19234 31556 19292
rect 31500 19182 31502 19234
rect 31554 19182 31556 19234
rect 31388 19010 31444 19022
rect 31388 18958 31390 19010
rect 31442 18958 31444 19010
rect 30828 17780 30884 17790
rect 30884 17724 31108 17780
rect 30828 17686 30884 17724
rect 31052 17666 31108 17724
rect 31052 17614 31054 17666
rect 31106 17614 31108 17666
rect 31052 17602 31108 17614
rect 31388 17668 31444 18958
rect 31388 17602 31444 17612
rect 31500 18452 31556 19182
rect 31388 17444 31444 17454
rect 31388 17220 31444 17388
rect 31388 17154 31444 17164
rect 30828 17108 30884 17118
rect 30828 17014 30884 17052
rect 31500 17106 31556 18396
rect 31612 17778 31668 19964
rect 31724 19124 31780 20076
rect 31836 19348 31892 21532
rect 31948 21474 32004 21486
rect 31948 21422 31950 21474
rect 32002 21422 32004 21474
rect 31948 19908 32004 21422
rect 32060 20916 32116 20926
rect 32284 20916 32340 22318
rect 32396 22372 32452 22382
rect 32396 22278 32452 22316
rect 32060 20914 32340 20916
rect 32060 20862 32062 20914
rect 32114 20862 32340 20914
rect 32060 20860 32340 20862
rect 32396 22148 32452 22158
rect 32060 20850 32116 20860
rect 31948 19814 32004 19852
rect 31836 19292 32004 19348
rect 31836 19124 31892 19134
rect 31724 19068 31836 19124
rect 31836 19058 31892 19068
rect 31948 18900 32004 19292
rect 32172 19236 32228 19246
rect 32396 19236 32452 22092
rect 32508 21810 32564 24332
rect 32508 21758 32510 21810
rect 32562 21758 32564 21810
rect 32508 21746 32564 21758
rect 32172 19234 32452 19236
rect 32172 19182 32174 19234
rect 32226 19182 32452 19234
rect 32172 19180 32452 19182
rect 32172 19170 32228 19180
rect 31612 17726 31614 17778
rect 31666 17726 31668 17778
rect 31612 17714 31668 17726
rect 31724 18844 32004 18900
rect 31500 17054 31502 17106
rect 31554 17054 31556 17106
rect 31500 17042 31556 17054
rect 31612 17556 31668 17566
rect 30940 16658 30996 16670
rect 30940 16606 30942 16658
rect 30994 16606 30996 16658
rect 29932 15092 30212 15148
rect 29708 14530 29764 14542
rect 29708 14478 29710 14530
rect 29762 14478 29764 14530
rect 29708 14420 29764 14478
rect 29932 14532 29988 14542
rect 29932 14438 29988 14476
rect 29708 14354 29764 14364
rect 29596 13570 29652 13580
rect 30156 12404 30212 15092
rect 30492 15092 30772 15148
rect 30828 15428 30884 15438
rect 30268 14868 30324 14878
rect 30268 14530 30324 14812
rect 30268 14478 30270 14530
rect 30322 14478 30324 14530
rect 30268 14466 30324 14478
rect 30268 13524 30324 13534
rect 30268 13074 30324 13468
rect 30268 13022 30270 13074
rect 30322 13022 30324 13074
rect 30268 13010 30324 13022
rect 30268 12404 30324 12414
rect 29932 12402 30324 12404
rect 29932 12350 30270 12402
rect 30322 12350 30324 12402
rect 29932 12348 30324 12350
rect 30492 12404 30548 15092
rect 30828 14980 30884 15372
rect 30940 15314 30996 16606
rect 30940 15262 30942 15314
rect 30994 15262 30996 15314
rect 30940 15250 30996 15262
rect 31500 15204 31556 15214
rect 30604 14924 30884 14980
rect 31276 15090 31332 15102
rect 31276 15038 31278 15090
rect 31330 15038 31332 15090
rect 30604 14756 30660 14924
rect 30604 14700 30772 14756
rect 30716 14642 30772 14700
rect 30716 14590 30718 14642
rect 30770 14590 30772 14642
rect 30716 14578 30772 14590
rect 30604 14532 30660 14542
rect 30604 14438 30660 14476
rect 31164 14530 31220 14542
rect 31164 14478 31166 14530
rect 31218 14478 31220 14530
rect 30828 14420 30884 14430
rect 30828 13186 30884 14364
rect 31164 14420 31220 14478
rect 31164 14354 31220 14364
rect 31276 14532 31332 15038
rect 31276 14418 31332 14476
rect 31276 14366 31278 14418
rect 31330 14366 31332 14418
rect 31276 14354 31332 14366
rect 31388 15092 31556 15148
rect 31388 14196 31444 15092
rect 31164 14140 31444 14196
rect 31164 13858 31220 14140
rect 31164 13806 31166 13858
rect 31218 13806 31220 13858
rect 31164 13794 31220 13806
rect 30828 13134 30830 13186
rect 30882 13134 30884 13186
rect 30828 13122 30884 13134
rect 31388 13524 31444 13534
rect 31052 13074 31108 13086
rect 31052 13022 31054 13074
rect 31106 13022 31108 13074
rect 30492 12348 30996 12404
rect 29708 12180 29764 12190
rect 29708 12086 29764 12124
rect 29820 11394 29876 11406
rect 29820 11342 29822 11394
rect 29874 11342 29876 11394
rect 29708 9604 29764 9614
rect 29708 9510 29764 9548
rect 29484 4958 29486 5010
rect 29538 4958 29540 5010
rect 29484 4946 29540 4958
rect 29596 5794 29652 5806
rect 29596 5742 29598 5794
rect 29650 5742 29652 5794
rect 29596 4788 29652 5742
rect 29820 5010 29876 11342
rect 29932 10498 29988 12348
rect 30268 12338 30324 12348
rect 30828 12180 30884 12190
rect 30716 11396 30772 11406
rect 30716 10724 30772 11340
rect 30828 11394 30884 12124
rect 30828 11342 30830 11394
rect 30882 11342 30884 11394
rect 30828 11330 30884 11342
rect 29932 10446 29934 10498
rect 29986 10446 29988 10498
rect 29932 10434 29988 10446
rect 30380 10610 30436 10622
rect 30380 10558 30382 10610
rect 30434 10558 30436 10610
rect 30380 9604 30436 10558
rect 30716 10498 30772 10668
rect 30716 10446 30718 10498
rect 30770 10446 30772 10498
rect 30492 9828 30548 9838
rect 30492 9826 30660 9828
rect 30492 9774 30494 9826
rect 30546 9774 30660 9826
rect 30492 9772 30660 9774
rect 30492 9762 30548 9772
rect 30380 9538 30436 9548
rect 30044 5124 30100 5134
rect 29820 4958 29822 5010
rect 29874 4958 29876 5010
rect 29820 4946 29876 4958
rect 29932 5122 30100 5124
rect 29932 5070 30046 5122
rect 30098 5070 30100 5122
rect 29932 5068 30100 5070
rect 29932 4788 29988 5068
rect 30044 5058 30100 5068
rect 29596 4732 29988 4788
rect 29372 3668 29428 3678
rect 29372 3574 29428 3612
rect 29932 3388 29988 4732
rect 30492 4338 30548 4350
rect 30492 4286 30494 4338
rect 30546 4286 30548 4338
rect 28700 3332 28980 3388
rect 28924 800 28980 3332
rect 29596 3332 29988 3388
rect 30268 4228 30324 4238
rect 30492 4228 30548 4286
rect 30268 4226 30548 4228
rect 30268 4174 30270 4226
rect 30322 4174 30548 4226
rect 30268 4172 30548 4174
rect 29596 800 29652 3332
rect 30268 800 30324 4172
rect 30604 3444 30660 9772
rect 30716 9826 30772 10446
rect 30716 9774 30718 9826
rect 30770 9774 30772 9826
rect 30716 9762 30772 9774
rect 30828 10164 30884 10174
rect 30828 9154 30884 10108
rect 30828 9102 30830 9154
rect 30882 9102 30884 9154
rect 30828 9090 30884 9102
rect 30828 8932 30884 8942
rect 30828 8258 30884 8876
rect 30828 8206 30830 8258
rect 30882 8206 30884 8258
rect 30828 8194 30884 8206
rect 30828 4564 30884 4574
rect 30940 4564 30996 12348
rect 31052 12402 31108 13022
rect 31052 12350 31054 12402
rect 31106 12350 31108 12402
rect 31052 12338 31108 12350
rect 31276 12292 31332 12302
rect 31052 11396 31108 11406
rect 31276 11396 31332 12236
rect 31388 12290 31444 13468
rect 31500 12964 31556 12974
rect 31500 12870 31556 12908
rect 31388 12238 31390 12290
rect 31442 12238 31444 12290
rect 31388 12226 31444 12238
rect 31612 12180 31668 17500
rect 31724 16660 31780 18844
rect 32284 18452 32340 18462
rect 32340 18396 32452 18452
rect 32284 18358 32340 18396
rect 31836 18338 31892 18350
rect 31836 18286 31838 18338
rect 31890 18286 31892 18338
rect 31836 17444 31892 18286
rect 32396 17892 32452 18396
rect 32060 17836 32452 17892
rect 31948 17444 32004 17454
rect 31836 17442 32004 17444
rect 31836 17390 31950 17442
rect 32002 17390 32004 17442
rect 31836 17388 32004 17390
rect 31948 17108 32004 17388
rect 31948 17042 32004 17052
rect 32060 17220 32116 17836
rect 32396 17778 32452 17836
rect 32396 17726 32398 17778
rect 32450 17726 32452 17778
rect 32396 17714 32452 17726
rect 32060 17106 32116 17164
rect 32060 17054 32062 17106
rect 32114 17054 32116 17106
rect 32060 17042 32116 17054
rect 32284 17668 32340 17678
rect 31948 16884 32004 16894
rect 31948 16790 32004 16828
rect 32060 16660 32116 16670
rect 31724 15988 31780 16604
rect 31724 15922 31780 15932
rect 31836 16658 32116 16660
rect 31836 16606 32062 16658
rect 32114 16606 32116 16658
rect 31836 16604 32116 16606
rect 31836 15314 31892 16604
rect 32060 16594 32116 16604
rect 32172 15764 32228 15774
rect 31836 15262 31838 15314
rect 31890 15262 31892 15314
rect 31836 15250 31892 15262
rect 32060 15652 32116 15662
rect 32060 15148 32116 15596
rect 32172 15426 32228 15708
rect 32284 15538 32340 17612
rect 32620 17332 32676 27804
rect 32732 24052 32788 24062
rect 32732 23958 32788 23996
rect 32956 20356 33012 28028
rect 33068 27858 33124 27870
rect 33068 27806 33070 27858
rect 33122 27806 33124 27858
rect 33068 24724 33124 27806
rect 33068 24658 33124 24668
rect 33180 23268 33236 28140
rect 33292 27412 33348 27422
rect 33292 27076 33348 27356
rect 33292 26982 33348 27020
rect 33404 27074 33460 28364
rect 33516 27860 33572 34188
rect 33628 33348 33684 33358
rect 33628 32674 33684 33292
rect 33628 32622 33630 32674
rect 33682 32622 33684 32674
rect 33628 32610 33684 32622
rect 33740 31556 33796 34860
rect 33852 34692 33908 34702
rect 33852 34598 33908 34636
rect 33852 34468 33908 34478
rect 33852 34354 33908 34412
rect 33852 34302 33854 34354
rect 33906 34302 33908 34354
rect 33852 34290 33908 34302
rect 33740 31490 33796 31500
rect 33852 31108 33908 31118
rect 33852 31014 33908 31052
rect 33628 30324 33684 30334
rect 33628 30098 33684 30268
rect 33628 30046 33630 30098
rect 33682 30046 33684 30098
rect 33628 30034 33684 30046
rect 33628 29876 33684 29886
rect 33628 29650 33684 29820
rect 33628 29598 33630 29650
rect 33682 29598 33684 29650
rect 33628 29586 33684 29598
rect 33964 29204 34020 37884
rect 34524 37828 34580 37838
rect 34524 37734 34580 37772
rect 34300 37266 34356 37278
rect 34300 37214 34302 37266
rect 34354 37214 34356 37266
rect 34300 35700 34356 37214
rect 34412 36036 34468 36046
rect 34412 35922 34468 35980
rect 34412 35870 34414 35922
rect 34466 35870 34468 35922
rect 34412 35858 34468 35870
rect 34524 35812 34580 35822
rect 34524 35718 34580 35756
rect 34300 35634 34356 35644
rect 34636 35252 34692 38220
rect 34748 37828 34804 40348
rect 34860 40402 34916 41356
rect 34972 41410 35028 42702
rect 35084 42754 35140 42766
rect 35084 42702 35086 42754
rect 35138 42702 35140 42754
rect 35084 42644 35140 42702
rect 35868 42644 35924 42654
rect 35140 42642 35924 42644
rect 35140 42590 35870 42642
rect 35922 42590 35924 42642
rect 35140 42588 35924 42590
rect 35084 42578 35140 42588
rect 35420 42194 35476 42588
rect 35868 42578 35924 42588
rect 35420 42142 35422 42194
rect 35474 42142 35476 42194
rect 35420 42130 35476 42142
rect 35644 41970 35700 41982
rect 35644 41918 35646 41970
rect 35698 41918 35700 41970
rect 35644 41748 35700 41918
rect 35644 41682 35700 41692
rect 35196 41580 35460 41590
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35196 41514 35460 41524
rect 34972 41358 34974 41410
rect 35026 41358 35028 41410
rect 34972 41346 35028 41358
rect 35196 41188 35252 41198
rect 35196 41094 35252 41132
rect 35868 40964 35924 40974
rect 35980 40964 36036 42812
rect 36204 42756 36260 42766
rect 36316 42756 36372 49532
rect 37100 49138 37156 49756
rect 37100 49086 37102 49138
rect 37154 49086 37156 49138
rect 37100 49074 37156 49086
rect 36428 48804 36484 48814
rect 36428 48710 36484 48748
rect 36988 48804 37044 48814
rect 37212 48804 37268 48814
rect 36988 48802 37156 48804
rect 36988 48750 36990 48802
rect 37042 48750 37156 48802
rect 36988 48748 37156 48750
rect 36988 48738 37044 48748
rect 37100 48692 37156 48748
rect 36876 48132 36932 48142
rect 36428 46676 36484 46686
rect 36428 46674 36708 46676
rect 36428 46622 36430 46674
rect 36482 46622 36708 46674
rect 36428 46620 36708 46622
rect 36428 46610 36484 46620
rect 36540 46452 36596 46462
rect 36428 46450 36596 46452
rect 36428 46398 36542 46450
rect 36594 46398 36596 46450
rect 36428 46396 36596 46398
rect 36428 46004 36484 46396
rect 36540 46386 36596 46396
rect 36652 46228 36708 46620
rect 36764 46564 36820 46574
rect 36764 46470 36820 46508
rect 36876 46450 36932 48076
rect 36988 47460 37044 47470
rect 36988 47366 37044 47404
rect 37100 47236 37156 48636
rect 37212 47684 37268 48748
rect 37212 47618 37268 47628
rect 37324 47908 37380 53228
rect 37436 53172 37492 53182
rect 37436 53078 37492 53116
rect 37548 52948 37604 53454
rect 37996 53506 38052 53518
rect 37996 53454 37998 53506
rect 38050 53454 38052 53506
rect 37996 53172 38052 53454
rect 37996 53106 38052 53116
rect 37548 52854 37604 52892
rect 38892 52500 38948 59388
rect 39340 59350 39396 59388
rect 39116 59220 39172 59230
rect 39116 58212 39172 59164
rect 39228 59218 39284 59230
rect 39228 59166 39230 59218
rect 39282 59166 39284 59218
rect 39228 58436 39284 59166
rect 39452 58772 39508 59612
rect 39564 59444 39620 59454
rect 39564 59350 39620 59388
rect 39676 59442 39732 60732
rect 39788 60004 39844 60014
rect 39788 59910 39844 59948
rect 39676 59390 39678 59442
rect 39730 59390 39732 59442
rect 39676 59378 39732 59390
rect 39900 59442 39956 60844
rect 40012 60674 40068 60686
rect 40012 60622 40014 60674
rect 40066 60622 40068 60674
rect 40012 60452 40068 60622
rect 40012 60386 40068 60396
rect 40348 60676 40404 60686
rect 40012 60228 40068 60238
rect 40012 60002 40068 60172
rect 40348 60004 40404 60620
rect 40012 59950 40014 60002
rect 40066 59950 40068 60002
rect 40012 59938 40068 59950
rect 40124 59948 40404 60004
rect 39900 59390 39902 59442
rect 39954 59390 39956 59442
rect 39900 59108 39956 59390
rect 40012 59780 40068 59790
rect 40124 59780 40180 59948
rect 40572 59890 40628 59902
rect 40572 59838 40574 59890
rect 40626 59838 40628 59890
rect 40068 59724 40180 59780
rect 40236 59780 40292 59790
rect 40236 59778 40404 59780
rect 40236 59726 40238 59778
rect 40290 59726 40404 59778
rect 40236 59724 40404 59726
rect 40012 59220 40068 59724
rect 40236 59714 40292 59724
rect 40012 59126 40068 59164
rect 39900 59042 39956 59052
rect 39452 58716 40292 58772
rect 39228 58434 39396 58436
rect 39228 58382 39230 58434
rect 39282 58382 39396 58434
rect 39228 58380 39396 58382
rect 39228 58370 39284 58380
rect 39116 58156 39284 58212
rect 39004 57428 39060 57438
rect 39004 56642 39060 57372
rect 39004 56590 39006 56642
rect 39058 56590 39060 56642
rect 39004 56578 39060 56590
rect 39116 57204 39172 57214
rect 39116 56196 39172 57148
rect 39116 55300 39172 56140
rect 39004 55244 39172 55300
rect 39004 52946 39060 55244
rect 39228 55188 39284 58156
rect 39340 56980 39396 58380
rect 39452 58434 39508 58716
rect 39564 58548 39620 58558
rect 39564 58454 39620 58492
rect 39452 58382 39454 58434
rect 39506 58382 39508 58434
rect 39452 58370 39508 58382
rect 39788 58434 39844 58446
rect 39788 58382 39790 58434
rect 39842 58382 39844 58434
rect 39340 56886 39396 56924
rect 39452 57428 39508 57438
rect 39004 52894 39006 52946
rect 39058 52894 39060 52946
rect 39004 52882 39060 52894
rect 39116 55132 39284 55188
rect 38780 52444 38948 52500
rect 38668 52276 38724 52286
rect 38556 52220 38668 52276
rect 38108 52164 38164 52174
rect 37996 51492 38052 51502
rect 37996 51398 38052 51436
rect 37884 51380 37940 51390
rect 37884 51286 37940 51324
rect 37996 51156 38052 51166
rect 37996 51062 38052 51100
rect 37996 50594 38052 50606
rect 37996 50542 37998 50594
rect 38050 50542 38052 50594
rect 37884 50372 37940 50382
rect 37436 50370 37940 50372
rect 37436 50318 37886 50370
rect 37938 50318 37940 50370
rect 37436 50316 37940 50318
rect 37436 49698 37492 50316
rect 37884 50306 37940 50316
rect 37548 50036 37604 50046
rect 37996 50036 38052 50542
rect 38108 50484 38164 52108
rect 38220 52164 38276 52174
rect 38444 52164 38500 52174
rect 38220 52162 38444 52164
rect 38220 52110 38222 52162
rect 38274 52110 38444 52162
rect 38220 52108 38444 52110
rect 38220 52098 38276 52108
rect 38444 52070 38500 52108
rect 38556 51602 38612 52220
rect 38668 52210 38724 52220
rect 38556 51550 38558 51602
rect 38610 51550 38612 51602
rect 38556 51538 38612 51550
rect 38668 52050 38724 52062
rect 38668 51998 38670 52050
rect 38722 51998 38724 52050
rect 38668 51380 38724 51998
rect 38780 51716 38836 52444
rect 38892 52276 38948 52286
rect 38892 52182 38948 52220
rect 38780 51650 38836 51660
rect 39004 52050 39060 52062
rect 39004 51998 39006 52050
rect 39058 51998 39060 52050
rect 39004 51604 39060 51998
rect 39004 51510 39060 51548
rect 38780 51380 38836 51390
rect 38668 51378 38836 51380
rect 38668 51326 38782 51378
rect 38834 51326 38836 51378
rect 38668 51324 38836 51326
rect 38108 50418 38164 50428
rect 38556 50594 38612 50606
rect 38556 50542 38558 50594
rect 38610 50542 38612 50594
rect 37604 49980 37716 50036
rect 37548 49970 37604 49980
rect 37436 49646 37438 49698
rect 37490 49646 37492 49698
rect 37436 48692 37492 49646
rect 37436 48626 37492 48636
rect 37548 49810 37604 49822
rect 37548 49758 37550 49810
rect 37602 49758 37604 49810
rect 37548 49026 37604 49758
rect 37548 48974 37550 49026
rect 37602 48974 37604 49026
rect 37548 48468 37604 48974
rect 37548 48402 37604 48412
rect 37548 48132 37604 48142
rect 37660 48132 37716 49980
rect 37996 49970 38052 49980
rect 38220 49924 38276 49934
rect 38220 49830 38276 49868
rect 38108 49028 38164 49038
rect 38108 48934 38164 48972
rect 37548 48130 37716 48132
rect 37548 48078 37550 48130
rect 37602 48078 37716 48130
rect 37548 48076 37716 48078
rect 37772 48802 37828 48814
rect 37772 48750 37774 48802
rect 37826 48750 37828 48802
rect 37548 48066 37604 48076
rect 37772 48020 37828 48750
rect 37884 48804 37940 48814
rect 37884 48356 37940 48748
rect 37996 48804 38052 48814
rect 37996 48802 38164 48804
rect 37996 48750 37998 48802
rect 38050 48750 38164 48802
rect 37996 48748 38164 48750
rect 37996 48738 38052 48748
rect 37996 48356 38052 48366
rect 37884 48354 38052 48356
rect 37884 48302 37998 48354
rect 38050 48302 38052 48354
rect 37884 48300 38052 48302
rect 37996 48290 38052 48300
rect 37772 47954 37828 47964
rect 38108 47908 38164 48748
rect 38220 48692 38276 48702
rect 38220 48466 38276 48636
rect 38220 48414 38222 48466
rect 38274 48414 38276 48466
rect 38220 48402 38276 48414
rect 38332 48468 38388 48478
rect 38108 47852 38276 47908
rect 37324 47572 37380 47852
rect 38108 47684 38164 47694
rect 38108 47590 38164 47628
rect 37436 47572 37492 47582
rect 37324 47570 37492 47572
rect 37324 47518 37438 47570
rect 37490 47518 37492 47570
rect 37324 47516 37492 47518
rect 37436 47506 37492 47516
rect 37884 47458 37940 47470
rect 37884 47406 37886 47458
rect 37938 47406 37940 47458
rect 37884 47236 37940 47406
rect 37100 47180 37940 47236
rect 37996 47236 38052 47246
rect 37996 47142 38052 47180
rect 38220 46788 38276 47852
rect 38332 47458 38388 48412
rect 38444 48356 38500 48366
rect 38444 48262 38500 48300
rect 38332 47406 38334 47458
rect 38386 47406 38388 47458
rect 38332 47236 38388 47406
rect 38444 48130 38500 48142
rect 38444 48078 38446 48130
rect 38498 48078 38500 48130
rect 38444 47460 38500 48078
rect 38444 47394 38500 47404
rect 38332 47170 38388 47180
rect 38108 46732 38276 46788
rect 37212 46676 37268 46686
rect 36876 46398 36878 46450
rect 36930 46398 36932 46450
rect 36876 46386 36932 46398
rect 36988 46452 37044 46462
rect 36652 46172 36932 46228
rect 36428 45910 36484 45948
rect 36876 45890 36932 46172
rect 36876 45838 36878 45890
rect 36930 45838 36932 45890
rect 36876 45826 36932 45838
rect 36988 43988 37044 46396
rect 37212 45778 37268 46620
rect 37212 45726 37214 45778
rect 37266 45726 37268 45778
rect 37100 45666 37156 45678
rect 37100 45614 37102 45666
rect 37154 45614 37156 45666
rect 37100 45332 37156 45614
rect 37212 45444 37268 45726
rect 37212 45378 37268 45388
rect 37436 46674 37492 46686
rect 37436 46622 37438 46674
rect 37490 46622 37492 46674
rect 37436 45780 37492 46622
rect 37772 46004 37828 46014
rect 37772 45780 37828 45948
rect 37436 45778 37828 45780
rect 37436 45726 37774 45778
rect 37826 45726 37828 45778
rect 37436 45724 37828 45726
rect 37100 44212 37156 45276
rect 37100 44146 37156 44156
rect 37436 45220 37492 45724
rect 37772 45714 37828 45724
rect 36988 43932 37156 43988
rect 36428 43426 36484 43438
rect 36428 43374 36430 43426
rect 36482 43374 36484 43426
rect 36428 43314 36484 43374
rect 36428 43262 36430 43314
rect 36482 43262 36484 43314
rect 36428 43250 36484 43262
rect 36204 42754 36372 42756
rect 36204 42702 36206 42754
rect 36258 42702 36372 42754
rect 36204 42700 36372 42702
rect 36204 41860 36260 42700
rect 36428 42644 36484 42654
rect 36428 42550 36484 42588
rect 36316 42530 36372 42542
rect 36316 42478 36318 42530
rect 36370 42478 36372 42530
rect 36316 42084 36372 42478
rect 36988 42530 37044 42542
rect 36988 42478 36990 42530
rect 37042 42478 37044 42530
rect 36764 42420 36820 42430
rect 36988 42420 37044 42478
rect 36820 42364 37044 42420
rect 36316 42028 36484 42084
rect 36316 41860 36372 41870
rect 36204 41858 36372 41860
rect 36204 41806 36318 41858
rect 36370 41806 36372 41858
rect 36204 41804 36372 41806
rect 36316 41794 36372 41804
rect 35924 40908 36036 40964
rect 35868 40898 35924 40908
rect 35532 40852 35588 40862
rect 35308 40628 35364 40638
rect 35308 40534 35364 40572
rect 34860 40350 34862 40402
rect 34914 40350 34916 40402
rect 34860 40338 34916 40350
rect 34972 40402 35028 40414
rect 34972 40350 34974 40402
rect 35026 40350 35028 40402
rect 34860 37828 34916 37838
rect 34748 37826 34916 37828
rect 34748 37774 34862 37826
rect 34914 37774 34916 37826
rect 34748 37772 34916 37774
rect 34748 35924 34804 37772
rect 34860 37762 34916 37772
rect 34972 37604 35028 40350
rect 35196 40404 35252 40414
rect 35196 40310 35252 40348
rect 34748 35858 34804 35868
rect 34860 37548 35028 37604
rect 35084 40290 35140 40302
rect 35084 40238 35086 40290
rect 35138 40238 35140 40290
rect 34076 35196 34692 35252
rect 34748 35588 34804 35598
rect 34076 33348 34132 35196
rect 34300 34916 34356 34926
rect 34748 34916 34804 35532
rect 34188 34914 34356 34916
rect 34188 34862 34302 34914
rect 34354 34862 34356 34914
rect 34188 34860 34356 34862
rect 34188 34468 34244 34860
rect 34300 34850 34356 34860
rect 34412 34914 34804 34916
rect 34412 34862 34750 34914
rect 34802 34862 34804 34914
rect 34412 34860 34804 34862
rect 34860 34916 34916 37548
rect 34972 37380 35028 37390
rect 35084 37380 35140 40238
rect 35196 40012 35460 40022
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35196 39946 35460 39956
rect 35532 38612 35588 40796
rect 36316 40628 36372 40638
rect 35756 40516 35812 40526
rect 35756 40422 35812 40460
rect 36316 40514 36372 40572
rect 36316 40462 36318 40514
rect 36370 40462 36372 40514
rect 36316 40450 36372 40462
rect 36204 40404 36260 40414
rect 36204 40310 36260 40348
rect 35868 40290 35924 40302
rect 35868 40238 35870 40290
rect 35922 40238 35924 40290
rect 35868 39732 35924 40238
rect 36092 39732 36148 39742
rect 35868 39730 36148 39732
rect 35868 39678 36094 39730
rect 36146 39678 36148 39730
rect 35868 39676 36148 39678
rect 36092 39508 36148 39676
rect 36092 39442 36148 39452
rect 35532 38546 35588 38556
rect 35196 38444 35460 38454
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35196 38378 35460 38388
rect 35420 37828 35476 37838
rect 35420 37734 35476 37772
rect 34972 37378 35140 37380
rect 34972 37326 34974 37378
rect 35026 37326 35140 37378
rect 34972 37324 35140 37326
rect 34972 37314 35028 37324
rect 35196 36876 35460 36886
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35196 36810 35460 36820
rect 35084 36594 35140 36606
rect 35084 36542 35086 36594
rect 35138 36542 35140 36594
rect 35084 35812 35140 36542
rect 35644 36482 35700 36494
rect 35644 36430 35646 36482
rect 35698 36430 35700 36482
rect 35644 35924 35700 36430
rect 36316 36484 36372 36494
rect 36428 36484 36484 42028
rect 36764 41972 36820 42364
rect 37100 42196 37156 43932
rect 37324 42756 37380 42766
rect 37324 42642 37380 42700
rect 37324 42590 37326 42642
rect 37378 42590 37380 42642
rect 37324 42532 37380 42590
rect 37324 42466 37380 42476
rect 36764 41878 36820 41916
rect 36988 42140 37156 42196
rect 36876 40290 36932 40302
rect 36876 40238 36878 40290
rect 36930 40238 36932 40290
rect 36876 39508 36932 40238
rect 36876 39442 36932 39452
rect 36316 36482 36484 36484
rect 36316 36430 36318 36482
rect 36370 36430 36484 36482
rect 36316 36428 36484 36430
rect 36316 36418 36372 36428
rect 35644 35858 35700 35868
rect 35868 36258 35924 36270
rect 35868 36206 35870 36258
rect 35922 36206 35924 36258
rect 35084 35746 35140 35756
rect 35308 35700 35364 35710
rect 35532 35700 35588 35710
rect 35308 35698 35532 35700
rect 35308 35646 35310 35698
rect 35362 35646 35532 35698
rect 35308 35644 35532 35646
rect 35308 35634 35364 35644
rect 35196 35308 35460 35318
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35196 35242 35460 35252
rect 35084 34916 35140 34926
rect 34860 34914 35140 34916
rect 34860 34862 35086 34914
rect 35138 34862 35140 34914
rect 34860 34860 35140 34862
rect 34188 34132 34244 34412
rect 34300 34356 34356 34366
rect 34412 34356 34468 34860
rect 34748 34850 34804 34860
rect 35084 34850 35140 34860
rect 35420 34804 35476 34814
rect 35420 34710 35476 34748
rect 35308 34692 35364 34702
rect 35308 34598 35364 34636
rect 34300 34354 34412 34356
rect 34300 34302 34302 34354
rect 34354 34302 34412 34354
rect 34300 34300 34412 34302
rect 34300 34290 34356 34300
rect 34412 34290 34468 34300
rect 34412 34132 34468 34142
rect 34188 34130 34468 34132
rect 34188 34078 34414 34130
rect 34466 34078 34468 34130
rect 34188 34076 34468 34078
rect 34412 34066 34468 34076
rect 34748 34130 34804 34142
rect 34748 34078 34750 34130
rect 34802 34078 34804 34130
rect 34636 34018 34692 34030
rect 34636 33966 34638 34018
rect 34690 33966 34692 34018
rect 34636 33684 34692 33966
rect 34412 33628 34692 33684
rect 34412 33570 34468 33628
rect 34412 33518 34414 33570
rect 34466 33518 34468 33570
rect 34412 33506 34468 33518
rect 34076 33282 34132 33292
rect 34188 33124 34244 33134
rect 34188 33030 34244 33068
rect 34300 33122 34356 33134
rect 34748 33124 34804 34078
rect 35084 34130 35140 34142
rect 35084 34078 35086 34130
rect 35138 34078 35140 34130
rect 35084 34020 35140 34078
rect 34972 33964 35084 34020
rect 34972 33908 35028 33964
rect 35084 33954 35140 33964
rect 35532 34130 35588 35644
rect 35868 35140 35924 36206
rect 35980 36258 36036 36270
rect 35980 36206 35982 36258
rect 36034 36206 36036 36258
rect 35980 35810 36036 36206
rect 35980 35758 35982 35810
rect 36034 35758 36036 35810
rect 35980 35746 36036 35758
rect 36092 36258 36148 36270
rect 36092 36206 36094 36258
rect 36146 36206 36148 36258
rect 35868 35074 35924 35084
rect 36092 34914 36148 36206
rect 36540 35812 36596 35822
rect 36540 35026 36596 35756
rect 36540 34974 36542 35026
rect 36594 34974 36596 35026
rect 36540 34962 36596 34974
rect 36092 34862 36094 34914
rect 36146 34862 36148 34914
rect 36092 34850 36148 34862
rect 35756 34804 35812 34814
rect 35756 34710 35812 34748
rect 35532 34078 35534 34130
rect 35586 34078 35588 34130
rect 34860 33852 35028 33908
rect 34860 33346 34916 33852
rect 35196 33740 35460 33750
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35196 33674 35460 33684
rect 35532 33572 35588 34078
rect 35532 33506 35588 33516
rect 35868 34690 35924 34702
rect 35868 34638 35870 34690
rect 35922 34638 35924 34690
rect 35868 33460 35924 34638
rect 36428 34692 36484 34702
rect 36204 34020 36260 34030
rect 35868 33394 35924 33404
rect 35980 34018 36260 34020
rect 35980 33966 36206 34018
rect 36258 33966 36260 34018
rect 35980 33964 36260 33966
rect 35980 33458 36036 33964
rect 36204 33954 36260 33964
rect 35980 33406 35982 33458
rect 36034 33406 36036 33458
rect 35980 33394 36036 33406
rect 34860 33294 34862 33346
rect 34914 33294 34916 33346
rect 34860 33282 34916 33294
rect 35084 33348 35140 33358
rect 35084 33254 35140 33292
rect 34972 33234 35028 33246
rect 34972 33182 34974 33234
rect 35026 33182 35028 33234
rect 34972 33124 35028 33182
rect 34300 33070 34302 33122
rect 34354 33070 34356 33122
rect 34188 32788 34244 32798
rect 34188 32694 34244 32732
rect 34300 32564 34356 33070
rect 34524 33068 35028 33124
rect 35532 33124 35588 33134
rect 34412 32788 34468 32798
rect 34412 32694 34468 32732
rect 34300 32498 34356 32508
rect 34076 30212 34132 30222
rect 34076 30118 34132 30156
rect 34076 29876 34132 29886
rect 34132 29820 34244 29876
rect 34076 29810 34132 29820
rect 33516 27794 33572 27804
rect 33628 29148 34020 29204
rect 33404 27022 33406 27074
rect 33458 27022 33460 27074
rect 33404 27010 33460 27022
rect 33292 26292 33348 26302
rect 33292 25506 33348 26236
rect 33292 25454 33294 25506
rect 33346 25454 33348 25506
rect 33292 24836 33348 25454
rect 33404 26180 33460 26190
rect 33404 25506 33460 26124
rect 33404 25454 33406 25506
rect 33458 25454 33460 25506
rect 33404 25442 33460 25454
rect 33516 25730 33572 25742
rect 33516 25678 33518 25730
rect 33570 25678 33572 25730
rect 33292 24770 33348 24780
rect 33404 24836 33460 24846
rect 33516 24836 33572 25678
rect 33404 24834 33572 24836
rect 33404 24782 33406 24834
rect 33458 24782 33572 24834
rect 33404 24780 33572 24782
rect 33404 24770 33460 24780
rect 33292 24610 33348 24622
rect 33292 24558 33294 24610
rect 33346 24558 33348 24610
rect 33292 24052 33348 24558
rect 33292 23986 33348 23996
rect 33404 24612 33460 24622
rect 33180 23212 33348 23268
rect 33180 23042 33236 23054
rect 33180 22990 33182 23042
rect 33234 22990 33236 23042
rect 33180 22484 33236 22990
rect 33180 22418 33236 22428
rect 33068 21812 33124 21822
rect 33068 21718 33124 21756
rect 32956 20300 33236 20356
rect 33068 20130 33124 20142
rect 33068 20078 33070 20130
rect 33122 20078 33124 20130
rect 32844 19122 32900 19134
rect 32844 19070 32846 19122
rect 32898 19070 32900 19122
rect 32844 18452 32900 19070
rect 32844 18386 32900 18396
rect 33068 18676 33124 20078
rect 32844 17668 32900 17678
rect 32844 17554 32900 17612
rect 32844 17502 32846 17554
rect 32898 17502 32900 17554
rect 32844 17490 32900 17502
rect 32620 17276 32900 17332
rect 32284 15486 32286 15538
rect 32338 15486 32340 15538
rect 32284 15474 32340 15486
rect 32620 16212 32676 16222
rect 32172 15374 32174 15426
rect 32226 15374 32228 15426
rect 32172 15362 32228 15374
rect 32508 15316 32564 15326
rect 32508 15222 32564 15260
rect 31836 15092 32116 15148
rect 31836 14642 31892 15092
rect 32620 14756 32676 16156
rect 32844 15764 32900 17276
rect 33068 15876 33124 18620
rect 33180 17780 33236 20300
rect 33180 17666 33236 17724
rect 33180 17614 33182 17666
rect 33234 17614 33236 17666
rect 33180 17602 33236 17614
rect 33180 17220 33236 17230
rect 33180 17106 33236 17164
rect 33180 17054 33182 17106
rect 33234 17054 33236 17106
rect 33180 17042 33236 17054
rect 33068 15810 33124 15820
rect 33292 15764 33348 23212
rect 33404 22484 33460 24556
rect 33516 22484 33572 22494
rect 33404 22482 33572 22484
rect 33404 22430 33518 22482
rect 33570 22430 33572 22482
rect 33404 22428 33572 22430
rect 33516 22418 33572 22428
rect 33516 21474 33572 21486
rect 33516 21422 33518 21474
rect 33570 21422 33572 21474
rect 33516 20580 33572 21422
rect 33516 20514 33572 20524
rect 33628 20356 33684 29148
rect 33740 28868 33796 28878
rect 33740 28866 34132 28868
rect 33740 28814 33742 28866
rect 33794 28814 34132 28866
rect 33740 28812 34132 28814
rect 33740 28802 33796 28812
rect 33852 28530 33908 28542
rect 33852 28478 33854 28530
rect 33906 28478 33908 28530
rect 33740 28420 33796 28430
rect 33740 28326 33796 28364
rect 33852 27972 33908 28478
rect 33740 27916 33908 27972
rect 33740 27300 33796 27916
rect 33740 27234 33796 27244
rect 33852 27746 33908 27758
rect 33852 27694 33854 27746
rect 33906 27694 33908 27746
rect 33852 27188 33908 27694
rect 33964 27188 34020 27198
rect 33852 27186 34020 27188
rect 33852 27134 33966 27186
rect 34018 27134 34020 27186
rect 33852 27132 34020 27134
rect 33964 27122 34020 27132
rect 34076 27074 34132 28812
rect 34188 28420 34244 29820
rect 34412 29540 34468 29550
rect 34412 29446 34468 29484
rect 34524 28868 34580 33068
rect 35532 33030 35588 33068
rect 35868 33122 35924 33134
rect 35868 33070 35870 33122
rect 35922 33070 35924 33122
rect 35196 32900 35252 32910
rect 35868 32900 35924 33070
rect 35196 32786 35252 32844
rect 35196 32734 35198 32786
rect 35250 32734 35252 32786
rect 35196 32722 35252 32734
rect 35532 32844 35924 32900
rect 35980 33124 36036 33134
rect 35532 32786 35588 32844
rect 35532 32734 35534 32786
rect 35586 32734 35588 32786
rect 35532 32722 35588 32734
rect 34748 32674 34804 32686
rect 34748 32622 34750 32674
rect 34802 32622 34804 32674
rect 34748 32340 34804 32622
rect 35980 32674 36036 33068
rect 35980 32622 35982 32674
rect 36034 32622 36036 32674
rect 35980 32610 36036 32622
rect 36092 33122 36148 33134
rect 36092 33070 36094 33122
rect 36146 33070 36148 33122
rect 35420 32564 35476 32574
rect 35644 32564 35700 32574
rect 35420 32562 35588 32564
rect 35420 32510 35422 32562
rect 35474 32510 35588 32562
rect 35420 32508 35588 32510
rect 35420 32498 35476 32508
rect 34748 32274 34804 32284
rect 35196 32172 35460 32182
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35196 32106 35460 32116
rect 35420 32004 35476 32014
rect 35308 31948 35420 32004
rect 34972 31780 35028 31790
rect 34972 31778 35140 31780
rect 34972 31726 34974 31778
rect 35026 31726 35140 31778
rect 34972 31724 35140 31726
rect 34972 31714 35028 31724
rect 34748 30324 34804 30334
rect 34188 28354 34244 28364
rect 34300 28812 34580 28868
rect 34636 29314 34692 29326
rect 34636 29262 34638 29314
rect 34690 29262 34692 29314
rect 34076 27022 34078 27074
rect 34130 27022 34132 27074
rect 34076 27010 34132 27022
rect 34188 27076 34244 27086
rect 33852 26962 33908 26974
rect 33852 26910 33854 26962
rect 33906 26910 33908 26962
rect 33852 26908 33908 26910
rect 34188 26908 34244 27020
rect 33852 26852 34244 26908
rect 34300 26292 34356 28812
rect 34524 28644 34580 28654
rect 34524 28550 34580 28588
rect 34412 27412 34468 27422
rect 34412 27074 34468 27356
rect 34412 27022 34414 27074
rect 34466 27022 34468 27074
rect 34412 27010 34468 27022
rect 34524 27076 34580 27114
rect 34524 27010 34580 27020
rect 34636 26908 34692 29262
rect 34748 27412 34804 30268
rect 35084 30324 35140 31724
rect 35308 31778 35364 31948
rect 35420 31938 35476 31948
rect 35308 31726 35310 31778
rect 35362 31726 35364 31778
rect 35308 31714 35364 31726
rect 35532 31780 35588 32508
rect 35644 32470 35700 32508
rect 36092 32228 36148 33070
rect 36428 33124 36484 34636
rect 36988 34244 37044 42140
rect 37324 41972 37380 41982
rect 37324 41878 37380 41916
rect 37212 40628 37268 40638
rect 37100 40572 37212 40628
rect 37100 37154 37156 40572
rect 37212 40534 37268 40572
rect 37212 39620 37268 39630
rect 37436 39620 37492 45164
rect 37772 45444 37828 45454
rect 37772 44994 37828 45388
rect 38108 45332 38164 46732
rect 38220 46564 38276 46574
rect 38220 46562 38500 46564
rect 38220 46510 38222 46562
rect 38274 46510 38500 46562
rect 38220 46508 38500 46510
rect 38220 46498 38276 46508
rect 38444 45332 38500 46508
rect 38556 46004 38612 50542
rect 38668 49924 38724 51324
rect 38780 51314 38836 51324
rect 38892 51380 38948 51390
rect 38892 51286 38948 51324
rect 39116 51156 39172 55132
rect 39452 54516 39508 57372
rect 39788 57204 39844 58382
rect 40236 58434 40292 58716
rect 40348 58548 40404 59724
rect 40460 59778 40516 59790
rect 40460 59726 40462 59778
rect 40514 59726 40516 59778
rect 40460 59444 40516 59726
rect 40460 59378 40516 59388
rect 40348 58492 40516 58548
rect 40236 58382 40238 58434
rect 40290 58382 40292 58434
rect 40236 58370 40292 58382
rect 39788 57138 39844 57148
rect 40124 58322 40180 58334
rect 40124 58270 40126 58322
rect 40178 58270 40180 58322
rect 40124 56980 40180 58270
rect 40348 58322 40404 58334
rect 40348 58270 40350 58322
rect 40402 58270 40404 58322
rect 40348 57764 40404 58270
rect 40460 58212 40516 58492
rect 40460 58146 40516 58156
rect 40572 57876 40628 59838
rect 40572 57810 40628 57820
rect 40348 57708 40516 57764
rect 40348 57540 40404 57550
rect 40124 56914 40180 56924
rect 40236 57092 40292 57102
rect 40236 56644 40292 57036
rect 39340 54460 39508 54516
rect 39900 55410 39956 55422
rect 39900 55358 39902 55410
rect 39954 55358 39956 55410
rect 39900 54516 39956 55358
rect 39228 52834 39284 52846
rect 39228 52782 39230 52834
rect 39282 52782 39284 52834
rect 39228 52052 39284 52782
rect 39340 52164 39396 54460
rect 39900 54450 39956 54460
rect 39676 54404 39732 54414
rect 39452 54402 39732 54404
rect 39452 54350 39678 54402
rect 39730 54350 39732 54402
rect 39452 54348 39732 54350
rect 39452 53060 39508 54348
rect 39676 54338 39732 54348
rect 40124 53732 40180 53742
rect 40124 53638 40180 53676
rect 39452 53058 39620 53060
rect 39452 53006 39454 53058
rect 39506 53006 39620 53058
rect 39452 53004 39620 53006
rect 39452 52994 39508 53004
rect 39564 52948 39620 53004
rect 39564 52724 39620 52892
rect 39676 52948 39732 52958
rect 39676 52946 40068 52948
rect 39676 52894 39678 52946
rect 39730 52894 40068 52946
rect 39676 52892 40068 52894
rect 39676 52882 39732 52892
rect 39564 52668 39956 52724
rect 39788 52164 39844 52174
rect 39340 52162 39844 52164
rect 39340 52110 39790 52162
rect 39842 52110 39844 52162
rect 39340 52108 39844 52110
rect 39788 52098 39844 52108
rect 39900 52162 39956 52668
rect 39900 52110 39902 52162
rect 39954 52110 39956 52162
rect 39900 52098 39956 52110
rect 40012 52162 40068 52892
rect 40012 52110 40014 52162
rect 40066 52110 40068 52162
rect 39228 51986 39284 51996
rect 39340 51940 39396 51950
rect 39340 51938 39732 51940
rect 39340 51886 39342 51938
rect 39394 51886 39732 51938
rect 39340 51884 39732 51886
rect 39340 51874 39396 51884
rect 39564 51716 39620 51726
rect 39228 51604 39284 51614
rect 39284 51548 39396 51604
rect 39228 51538 39284 51548
rect 38668 49858 38724 49868
rect 38780 51100 39172 51156
rect 39340 51156 39396 51548
rect 39452 51380 39508 51418
rect 39452 51314 39508 51324
rect 39452 51156 39508 51166
rect 39340 51154 39508 51156
rect 39340 51102 39454 51154
rect 39506 51102 39508 51154
rect 39340 51100 39508 51102
rect 38668 49700 38724 49710
rect 38668 49138 38724 49644
rect 38668 49086 38670 49138
rect 38722 49086 38724 49138
rect 38668 48804 38724 49086
rect 38668 48738 38724 48748
rect 38668 48242 38724 48254
rect 38668 48190 38670 48242
rect 38722 48190 38724 48242
rect 38668 47460 38724 48190
rect 38668 47394 38724 47404
rect 38556 45938 38612 45948
rect 38556 45332 38612 45342
rect 38444 45330 38612 45332
rect 38444 45278 38558 45330
rect 38610 45278 38612 45330
rect 38444 45276 38612 45278
rect 38108 45266 38164 45276
rect 38556 45266 38612 45276
rect 37772 44942 37774 44994
rect 37826 44942 37828 44994
rect 37772 44884 37828 44942
rect 38780 44996 38836 51100
rect 39228 51044 39284 51054
rect 38892 50932 38948 50942
rect 38892 47908 38948 50876
rect 39228 50706 39284 50988
rect 39228 50654 39230 50706
rect 39282 50654 39284 50706
rect 39228 50642 39284 50654
rect 39340 50260 39396 50270
rect 39228 49924 39284 49934
rect 39228 49830 39284 49868
rect 39340 49700 39396 50204
rect 39452 49810 39508 51100
rect 39564 50932 39620 51660
rect 39676 51380 39732 51884
rect 39900 51380 39956 51390
rect 39676 51324 39900 51380
rect 39900 51286 39956 51324
rect 40012 51268 40068 52110
rect 40012 51202 40068 51212
rect 39564 50866 39620 50876
rect 39676 51156 39732 51166
rect 39452 49758 39454 49810
rect 39506 49758 39508 49810
rect 39452 49746 39508 49758
rect 39340 49634 39396 49644
rect 39564 49140 39620 49150
rect 39004 49028 39060 49038
rect 39452 49028 39508 49038
rect 39004 49026 39508 49028
rect 39004 48974 39006 49026
rect 39058 48974 39454 49026
rect 39506 48974 39508 49026
rect 39004 48972 39508 48974
rect 39004 48962 39060 48972
rect 39452 48962 39508 48972
rect 39116 48804 39172 48814
rect 39116 48710 39172 48748
rect 39340 48804 39396 48814
rect 39340 48802 39508 48804
rect 39340 48750 39342 48802
rect 39394 48750 39508 48802
rect 39340 48748 39508 48750
rect 39340 48738 39396 48748
rect 39116 48468 39172 48478
rect 39116 48374 39172 48412
rect 39340 48244 39396 48254
rect 39340 48150 39396 48188
rect 39228 48132 39284 48142
rect 39228 48038 39284 48076
rect 38892 47852 39396 47908
rect 38892 47572 38948 47582
rect 38892 47478 38948 47516
rect 39228 47234 39284 47246
rect 39228 47182 39230 47234
rect 39282 47182 39284 47234
rect 38892 45220 38948 45230
rect 39228 45220 39284 47182
rect 38892 45218 39284 45220
rect 38892 45166 38894 45218
rect 38946 45166 39284 45218
rect 38892 45164 39284 45166
rect 38892 45154 38948 45164
rect 38780 44940 38948 44996
rect 37772 44828 38164 44884
rect 37996 43650 38052 43662
rect 37996 43598 37998 43650
rect 38050 43598 38052 43650
rect 37772 43538 37828 43550
rect 37772 43486 37774 43538
rect 37826 43486 37828 43538
rect 37660 42756 37716 42766
rect 37660 42662 37716 42700
rect 37548 41972 37604 41982
rect 37548 41878 37604 41916
rect 37660 41748 37716 41758
rect 37772 41748 37828 43486
rect 37996 43204 38052 43598
rect 37996 43138 38052 43148
rect 37884 42868 37940 42878
rect 37884 42194 37940 42812
rect 38108 42754 38164 44828
rect 38668 44212 38724 44222
rect 38668 44118 38724 44156
rect 38332 44098 38388 44110
rect 38332 44046 38334 44098
rect 38386 44046 38388 44098
rect 38332 43540 38388 44046
rect 38332 43474 38388 43484
rect 38780 43650 38836 43662
rect 38780 43598 38782 43650
rect 38834 43598 38836 43650
rect 38780 43428 38836 43598
rect 38668 43204 38724 43214
rect 38108 42702 38110 42754
rect 38162 42702 38164 42754
rect 38108 42690 38164 42702
rect 38332 42756 38388 42766
rect 38332 42662 38388 42700
rect 38668 42754 38724 43148
rect 38668 42702 38670 42754
rect 38722 42702 38724 42754
rect 38668 42690 38724 42702
rect 38780 42644 38836 43372
rect 38892 43652 38948 44940
rect 39340 43708 39396 47852
rect 39452 47012 39508 48748
rect 39564 48244 39620 49084
rect 39676 48914 39732 51100
rect 40236 50260 40292 56588
rect 40348 55972 40404 57484
rect 40460 57428 40516 57708
rect 40572 57428 40628 57438
rect 40460 57372 40572 57428
rect 40572 57362 40628 57372
rect 40348 55878 40404 55916
rect 40460 53506 40516 53518
rect 40460 53454 40462 53506
rect 40514 53454 40516 53506
rect 40460 53172 40516 53454
rect 40460 53106 40516 53116
rect 40684 50428 40740 63868
rect 40796 63922 40852 63934
rect 40796 63870 40798 63922
rect 40850 63870 40852 63922
rect 40796 63812 40852 63870
rect 41132 63922 41188 64654
rect 41244 64594 41300 64606
rect 41244 64542 41246 64594
rect 41298 64542 41300 64594
rect 41244 64372 41300 64542
rect 41244 64306 41300 64316
rect 41132 63870 41134 63922
rect 41186 63870 41188 63922
rect 41132 63858 41188 63870
rect 41356 63924 41412 63934
rect 41356 63830 41412 63868
rect 40796 63746 40852 63756
rect 41468 63812 41524 65214
rect 41804 65266 41860 65326
rect 41804 65214 41806 65266
rect 41858 65214 41860 65266
rect 41804 65202 41860 65214
rect 42028 65156 42084 67006
rect 42476 67170 42532 67182
rect 42476 67118 42478 67170
rect 42530 67118 42532 67170
rect 42252 66948 42308 66958
rect 42252 66274 42308 66892
rect 42476 66836 42532 67118
rect 42476 66770 42532 66780
rect 42588 67172 42644 67182
rect 42252 66222 42254 66274
rect 42306 66222 42308 66274
rect 42252 66210 42308 66222
rect 42476 66276 42532 66286
rect 42476 66162 42532 66220
rect 42476 66110 42478 66162
rect 42530 66110 42532 66162
rect 42476 66098 42532 66110
rect 42588 65604 42644 67116
rect 43260 67172 43316 67182
rect 43260 67078 43316 67116
rect 43484 67172 43540 67340
rect 43708 67284 43764 69246
rect 45276 69298 45332 69310
rect 45276 69246 45278 69298
rect 45330 69246 45332 69298
rect 44156 69188 44212 69226
rect 44156 69122 44212 69132
rect 44156 68964 44212 68974
rect 44156 67842 44212 68908
rect 45164 68964 45220 68974
rect 44156 67790 44158 67842
rect 44210 67790 44212 67842
rect 44156 67778 44212 67790
rect 44828 67954 44884 67966
rect 44828 67902 44830 67954
rect 44882 67902 44884 67954
rect 43484 67078 43540 67116
rect 43596 67228 43764 67284
rect 42700 67058 42756 67070
rect 42700 67006 42702 67058
rect 42754 67006 42756 67058
rect 42700 66500 42756 67006
rect 42812 67060 42868 67070
rect 42812 66946 42868 67004
rect 43036 67060 43092 67070
rect 43036 67058 43204 67060
rect 43036 67006 43038 67058
rect 43090 67006 43204 67058
rect 43036 67004 43204 67006
rect 43036 66994 43092 67004
rect 42812 66894 42814 66946
rect 42866 66894 42868 66946
rect 42812 66882 42868 66894
rect 42700 66444 42868 66500
rect 42700 66274 42756 66286
rect 42700 66222 42702 66274
rect 42754 66222 42756 66274
rect 42700 66164 42756 66222
rect 42700 66098 42756 66108
rect 42812 66052 42868 66444
rect 42812 65986 42868 65996
rect 43036 66052 43092 66062
rect 43036 65958 43092 65996
rect 43148 65828 43204 67004
rect 43372 66948 43428 66958
rect 43596 66948 43652 67228
rect 44492 67172 44548 67182
rect 44492 67078 44548 67116
rect 43372 66946 43652 66948
rect 43372 66894 43374 66946
rect 43426 66894 43652 66946
rect 43372 66892 43652 66894
rect 43932 67058 43988 67070
rect 43932 67006 43934 67058
rect 43986 67006 43988 67058
rect 43372 66882 43428 66892
rect 43260 66836 43316 66846
rect 43260 66162 43316 66780
rect 43372 66500 43428 66510
rect 43372 66406 43428 66444
rect 43932 66498 43988 67006
rect 43932 66446 43934 66498
rect 43986 66446 43988 66498
rect 43932 66434 43988 66446
rect 44044 67058 44100 67070
rect 44044 67006 44046 67058
rect 44098 67006 44100 67058
rect 44044 66500 44100 67006
rect 44716 67058 44772 67070
rect 44716 67006 44718 67058
rect 44770 67006 44772 67058
rect 44044 66434 44100 66444
rect 44604 66946 44660 66958
rect 44604 66894 44606 66946
rect 44658 66894 44660 66946
rect 44492 66388 44548 66398
rect 44156 66274 44212 66286
rect 44156 66222 44158 66274
rect 44210 66222 44212 66274
rect 43260 66110 43262 66162
rect 43314 66110 43316 66162
rect 43260 66098 43316 66110
rect 43596 66164 43652 66174
rect 43596 66070 43652 66108
rect 43708 66052 43764 66062
rect 43820 66052 43876 66062
rect 43764 66050 43876 66052
rect 43764 65998 43822 66050
rect 43874 65998 43876 66050
rect 43764 65996 43876 65998
rect 43148 65772 43652 65828
rect 43596 65714 43652 65772
rect 43596 65662 43598 65714
rect 43650 65662 43652 65714
rect 43596 65650 43652 65662
rect 42588 65538 42644 65548
rect 43372 65604 43428 65614
rect 43036 65492 43092 65502
rect 42028 65090 42084 65100
rect 42140 65378 42196 65390
rect 42140 65326 42142 65378
rect 42194 65326 42196 65378
rect 41692 64932 41748 64942
rect 41748 64876 42084 64932
rect 41692 64838 41748 64876
rect 42028 64706 42084 64876
rect 42028 64654 42030 64706
rect 42082 64654 42084 64706
rect 42028 64642 42084 64654
rect 42140 64484 42196 65326
rect 42588 65378 42644 65390
rect 42588 65326 42590 65378
rect 42642 65326 42644 65378
rect 42364 65266 42420 65278
rect 42364 65214 42366 65266
rect 42418 65214 42420 65266
rect 42252 64596 42308 64606
rect 42252 64502 42308 64540
rect 42140 64418 42196 64428
rect 42252 64260 42308 64270
rect 42364 64260 42420 65214
rect 42588 65266 42644 65326
rect 42588 65214 42590 65266
rect 42642 65214 42644 65266
rect 42588 65202 42644 65214
rect 42700 65380 42756 65390
rect 42700 64706 42756 65324
rect 43036 65378 43092 65436
rect 43036 65326 43038 65378
rect 43090 65326 43092 65378
rect 43036 64930 43092 65326
rect 43036 64878 43038 64930
rect 43090 64878 43092 64930
rect 43036 64866 43092 64878
rect 43260 65156 43316 65166
rect 42700 64654 42702 64706
rect 42754 64654 42756 64706
rect 42700 64642 42756 64654
rect 43036 64596 43092 64606
rect 43036 64502 43092 64540
rect 42476 64484 42532 64494
rect 42476 64482 42756 64484
rect 42476 64430 42478 64482
rect 42530 64430 42756 64482
rect 42476 64428 42756 64430
rect 42476 64418 42532 64428
rect 42308 64204 42420 64260
rect 42588 64260 42644 64270
rect 42252 64194 42308 64204
rect 42476 64148 42532 64158
rect 42364 64092 42476 64148
rect 41916 64036 41972 64046
rect 41468 63746 41524 63756
rect 41804 64034 41972 64036
rect 41804 63982 41918 64034
rect 41970 63982 41972 64034
rect 41804 63980 41972 63982
rect 41692 63252 41748 63262
rect 41692 63028 41748 63196
rect 41804 63140 41860 63980
rect 41916 63970 41972 63980
rect 42028 63924 42084 63934
rect 42252 63924 42308 63934
rect 42028 63922 42308 63924
rect 42028 63870 42030 63922
rect 42082 63870 42254 63922
rect 42306 63870 42308 63922
rect 42028 63868 42308 63870
rect 42028 63858 42084 63868
rect 42252 63858 42308 63868
rect 41916 63700 41972 63710
rect 42364 63700 42420 64092
rect 42476 64054 42532 64092
rect 42588 64034 42644 64204
rect 42588 63982 42590 64034
rect 42642 63982 42644 64034
rect 42588 63970 42644 63982
rect 41916 63606 41972 63644
rect 42028 63644 42420 63700
rect 41804 63084 41972 63140
rect 41692 62972 41860 63028
rect 41020 62804 41076 62814
rect 41020 62578 41076 62748
rect 41692 62692 41748 62702
rect 41020 62526 41022 62578
rect 41074 62526 41076 62578
rect 41020 62514 41076 62526
rect 41132 62580 41188 62590
rect 40908 62356 40964 62366
rect 40908 62262 40964 62300
rect 40796 62244 40852 62254
rect 41132 62188 41188 62524
rect 41692 62578 41748 62636
rect 41692 62526 41694 62578
rect 41746 62526 41748 62578
rect 41692 62514 41748 62526
rect 41356 62468 41412 62478
rect 41356 62374 41412 62412
rect 41804 62466 41860 62972
rect 41804 62414 41806 62466
rect 41858 62414 41860 62466
rect 40796 61794 40852 62188
rect 41020 62132 41188 62188
rect 41244 62356 41300 62366
rect 40796 61742 40798 61794
rect 40850 61742 40852 61794
rect 40796 61730 40852 61742
rect 40908 62020 40964 62030
rect 40908 61236 40964 61964
rect 41020 61460 41076 62132
rect 41132 61796 41188 61806
rect 41244 61796 41300 62300
rect 41804 62020 41860 62414
rect 41692 61964 41860 62020
rect 41132 61794 41300 61796
rect 41132 61742 41134 61794
rect 41186 61742 41300 61794
rect 41132 61740 41300 61742
rect 41468 61794 41524 61806
rect 41468 61742 41470 61794
rect 41522 61742 41524 61794
rect 41132 61730 41188 61740
rect 41356 61684 41412 61694
rect 41468 61684 41524 61742
rect 41412 61628 41524 61684
rect 41692 61684 41748 61964
rect 41804 61796 41860 61806
rect 41916 61796 41972 63084
rect 42028 62578 42084 63644
rect 42700 63364 42756 64428
rect 42700 63298 42756 63308
rect 43148 63922 43204 63934
rect 43148 63870 43150 63922
rect 43202 63870 43204 63922
rect 43148 63138 43204 63870
rect 43148 63086 43150 63138
rect 43202 63086 43204 63138
rect 42364 63028 42420 63038
rect 43148 63028 43204 63086
rect 42364 63026 42644 63028
rect 42364 62974 42366 63026
rect 42418 62974 42644 63026
rect 42364 62972 42644 62974
rect 42364 62962 42420 62972
rect 42028 62526 42030 62578
rect 42082 62526 42084 62578
rect 42028 62514 42084 62526
rect 42588 62578 42644 62972
rect 43148 62962 43204 62972
rect 42588 62526 42590 62578
rect 42642 62526 42644 62578
rect 42588 62514 42644 62526
rect 42924 62916 42980 62926
rect 42364 62354 42420 62366
rect 42364 62302 42366 62354
rect 42418 62302 42420 62354
rect 41804 61794 41916 61796
rect 41804 61742 41806 61794
rect 41858 61742 41916 61794
rect 41804 61740 41916 61742
rect 41804 61730 41860 61740
rect 41916 61702 41972 61740
rect 42140 61796 42196 61806
rect 42140 61702 42196 61740
rect 42364 61796 42420 62302
rect 42812 62356 42868 62366
rect 42812 62262 42868 62300
rect 42924 62188 42980 62860
rect 43260 62580 43316 65100
rect 43260 62486 43316 62524
rect 43372 62468 43428 65548
rect 43596 64930 43652 64942
rect 43596 64878 43598 64930
rect 43650 64878 43652 64930
rect 43596 64482 43652 64878
rect 43596 64430 43598 64482
rect 43650 64430 43652 64482
rect 43372 62188 43428 62412
rect 41356 61618 41412 61628
rect 41692 61618 41748 61628
rect 42252 61684 42308 61694
rect 41804 61460 41860 61470
rect 41020 61404 41188 61460
rect 40908 61170 40964 61180
rect 41020 60674 41076 60686
rect 41020 60622 41022 60674
rect 41074 60622 41076 60674
rect 41020 60564 41076 60622
rect 41020 60228 41076 60508
rect 41020 60162 41076 60172
rect 41020 59780 41076 59790
rect 41020 59686 41076 59724
rect 41132 59442 41188 61404
rect 41580 61346 41636 61358
rect 41580 61294 41582 61346
rect 41634 61294 41636 61346
rect 41580 61236 41636 61294
rect 41804 61236 41860 61404
rect 42252 61458 42308 61628
rect 42252 61406 42254 61458
rect 42306 61406 42308 61458
rect 42252 61236 42308 61406
rect 41636 61180 41972 61236
rect 41580 61170 41636 61180
rect 41692 61010 41748 61180
rect 41692 60958 41694 61010
rect 41746 60958 41748 61010
rect 41692 60946 41748 60958
rect 41916 61012 41972 61180
rect 42252 61170 42308 61180
rect 42140 61124 42196 61134
rect 41916 60956 42084 61012
rect 42028 60002 42084 60956
rect 42028 59950 42030 60002
rect 42082 59950 42084 60002
rect 42028 59938 42084 59950
rect 41580 59892 41636 59902
rect 41468 59780 41524 59790
rect 41468 59686 41524 59724
rect 41132 59390 41134 59442
rect 41186 59390 41188 59442
rect 41132 59378 41188 59390
rect 41580 59330 41636 59836
rect 41580 59278 41582 59330
rect 41634 59278 41636 59330
rect 41132 59218 41188 59230
rect 41132 59166 41134 59218
rect 41186 59166 41188 59218
rect 41132 58996 41188 59166
rect 41132 58940 41412 58996
rect 40796 58660 40852 58670
rect 41132 58660 41188 58940
rect 40796 58658 41188 58660
rect 40796 58606 40798 58658
rect 40850 58606 41188 58658
rect 40796 58604 41188 58606
rect 41244 58828 41300 58838
rect 40796 58594 40852 58604
rect 41244 58436 41300 58772
rect 40796 58380 41300 58436
rect 41356 58434 41412 58940
rect 41468 58548 41524 58558
rect 41468 58454 41524 58492
rect 41356 58382 41358 58434
rect 41410 58382 41412 58434
rect 40796 53732 40852 58380
rect 41356 58370 41412 58382
rect 41244 58212 41300 58222
rect 41300 58156 41524 58212
rect 41244 58146 41300 58156
rect 41132 58100 41188 58110
rect 41132 57762 41188 58044
rect 41132 57710 41134 57762
rect 41186 57710 41188 57762
rect 41132 57698 41188 57710
rect 41020 57650 41076 57662
rect 41020 57598 41022 57650
rect 41074 57598 41076 57650
rect 41020 56644 41076 57598
rect 41356 57652 41412 57662
rect 41356 57558 41412 57596
rect 41468 56978 41524 58156
rect 41580 58100 41636 59278
rect 41580 58034 41636 58044
rect 41804 59218 41860 59230
rect 41804 59166 41806 59218
rect 41858 59166 41860 59218
rect 41804 58658 41860 59166
rect 41804 58606 41806 58658
rect 41858 58606 41860 58658
rect 41804 57876 41860 58606
rect 42028 58100 42084 58110
rect 41580 57874 41860 57876
rect 41580 57822 41806 57874
rect 41858 57822 41860 57874
rect 41580 57820 41860 57822
rect 41580 57650 41636 57820
rect 41804 57810 41860 57820
rect 41916 57876 41972 57886
rect 41916 57782 41972 57820
rect 42028 57874 42084 58044
rect 42028 57822 42030 57874
rect 42082 57822 42084 57874
rect 42028 57810 42084 57822
rect 41580 57598 41582 57650
rect 41634 57598 41636 57650
rect 41580 57586 41636 57598
rect 41468 56926 41470 56978
rect 41522 56926 41524 56978
rect 41468 56914 41524 56926
rect 42140 56644 42196 61068
rect 42364 60676 42420 61740
rect 42812 62132 42980 62188
rect 43036 62132 43428 62188
rect 43484 64260 43540 64270
rect 42700 61460 42756 61470
rect 42700 61366 42756 61404
rect 42364 60674 42532 60676
rect 42364 60622 42366 60674
rect 42418 60622 42532 60674
rect 42364 60620 42532 60622
rect 42364 60610 42420 60620
rect 42252 60452 42308 60462
rect 42252 60116 42308 60396
rect 42252 60060 42420 60116
rect 42364 60002 42420 60060
rect 42364 59950 42366 60002
rect 42418 59950 42420 60002
rect 42364 59938 42420 59950
rect 42476 60004 42532 60620
rect 42588 60004 42644 60014
rect 42476 60002 42644 60004
rect 42476 59950 42590 60002
rect 42642 59950 42644 60002
rect 42476 59948 42644 59950
rect 42252 59890 42308 59902
rect 42252 59838 42254 59890
rect 42306 59838 42308 59890
rect 42252 59780 42308 59838
rect 42588 59892 42644 59948
rect 42588 59826 42644 59836
rect 42252 59714 42308 59724
rect 42364 59668 42420 59678
rect 42252 57762 42308 57774
rect 42252 57710 42254 57762
rect 42306 57710 42308 57762
rect 42252 57652 42308 57710
rect 42252 57586 42308 57596
rect 42252 57092 42308 57102
rect 42364 57092 42420 59612
rect 42588 59444 42644 59454
rect 42812 59444 42868 62132
rect 43036 60900 43092 62132
rect 43148 61346 43204 61358
rect 43148 61294 43150 61346
rect 43202 61294 43204 61346
rect 43148 61236 43204 61294
rect 43148 61170 43204 61180
rect 42588 59350 42644 59388
rect 42700 59388 42868 59444
rect 42924 60844 43092 60900
rect 42924 60002 42980 60844
rect 43036 60676 43092 60686
rect 43260 60676 43316 60686
rect 43036 60674 43316 60676
rect 43036 60622 43038 60674
rect 43090 60622 43262 60674
rect 43314 60622 43316 60674
rect 43036 60620 43316 60622
rect 43036 60610 43092 60620
rect 42924 59950 42926 60002
rect 42978 59950 42980 60002
rect 42924 59444 42980 59950
rect 43148 59778 43204 60620
rect 43260 60610 43316 60620
rect 43484 60340 43540 64204
rect 43596 63924 43652 64430
rect 43596 63858 43652 63868
rect 43596 62916 43652 62926
rect 43708 62916 43764 65996
rect 43820 65986 43876 65996
rect 43820 65716 43876 65726
rect 43820 65622 43876 65660
rect 44156 65714 44212 66222
rect 44156 65662 44158 65714
rect 44210 65662 44212 65714
rect 44156 65650 44212 65662
rect 44268 66164 44324 66174
rect 43932 65602 43988 65614
rect 43932 65550 43934 65602
rect 43986 65550 43988 65602
rect 43932 65492 43988 65550
rect 43932 65426 43988 65436
rect 44044 64594 44100 64606
rect 44044 64542 44046 64594
rect 44098 64542 44100 64594
rect 43932 64484 43988 64494
rect 43820 64482 43988 64484
rect 43820 64430 43934 64482
rect 43986 64430 43988 64482
rect 43820 64428 43988 64430
rect 43820 64034 43876 64428
rect 43932 64418 43988 64428
rect 44044 64484 44100 64542
rect 44044 64418 44100 64428
rect 43820 63982 43822 64034
rect 43874 63982 43876 64034
rect 43820 63970 43876 63982
rect 43652 62860 43764 62916
rect 43820 63026 43876 63038
rect 43820 62974 43822 63026
rect 43874 62974 43876 63026
rect 43596 62850 43652 62860
rect 43820 62578 43876 62974
rect 44044 62916 44100 62926
rect 44044 62822 44100 62860
rect 44268 62916 44324 66108
rect 44380 65716 44436 65726
rect 44380 65622 44436 65660
rect 44492 65604 44548 66332
rect 44604 66052 44660 66894
rect 44604 65986 44660 65996
rect 44716 65716 44772 67006
rect 44828 66388 44884 67902
rect 45052 67172 45108 67182
rect 44940 67060 44996 67070
rect 44940 66966 44996 67004
rect 44828 66322 44884 66332
rect 44716 65660 44996 65716
rect 44492 65602 44884 65604
rect 44492 65550 44494 65602
rect 44546 65550 44884 65602
rect 44492 65548 44884 65550
rect 44492 65538 44548 65548
rect 44716 64708 44772 64718
rect 44380 64706 44772 64708
rect 44380 64654 44718 64706
rect 44770 64654 44772 64706
rect 44380 64652 44772 64654
rect 44380 63362 44436 64652
rect 44716 64642 44772 64652
rect 44380 63310 44382 63362
rect 44434 63310 44436 63362
rect 44380 63298 44436 63310
rect 44716 64372 44772 64382
rect 44268 62822 44324 62860
rect 43820 62526 43822 62578
rect 43874 62526 43876 62578
rect 43820 62514 43876 62526
rect 44604 62580 44660 62590
rect 44604 62486 44660 62524
rect 43596 62466 43652 62478
rect 43596 62414 43598 62466
rect 43650 62414 43652 62466
rect 43596 62356 43652 62414
rect 44044 62466 44100 62478
rect 44044 62414 44046 62466
rect 44098 62414 44100 62466
rect 44044 62356 44100 62414
rect 44156 62468 44212 62478
rect 44156 62374 44212 62412
rect 43596 62300 44100 62356
rect 43596 61796 43652 61806
rect 43596 61682 43652 61740
rect 43596 61630 43598 61682
rect 43650 61630 43652 61682
rect 43596 61618 43652 61630
rect 44044 61236 44100 62300
rect 44380 61348 44436 61358
rect 44380 61254 44436 61292
rect 43820 61180 44100 61236
rect 43372 60284 43540 60340
rect 43596 60452 43652 60462
rect 43148 59726 43150 59778
rect 43202 59726 43204 59778
rect 43148 59668 43204 59726
rect 43148 59602 43204 59612
rect 43260 59778 43316 59790
rect 43260 59726 43262 59778
rect 43314 59726 43316 59778
rect 42476 59218 42532 59230
rect 42476 59166 42478 59218
rect 42530 59166 42532 59218
rect 42476 59108 42532 59166
rect 42588 59108 42644 59118
rect 42476 59052 42588 59108
rect 42588 59042 42644 59052
rect 42700 58996 42756 59388
rect 42924 59378 42980 59388
rect 42812 59220 42868 59230
rect 43260 59220 43316 59726
rect 42812 59218 43092 59220
rect 42812 59166 42814 59218
rect 42866 59166 43092 59218
rect 42812 59164 43092 59166
rect 42812 59154 42868 59164
rect 42700 58940 42980 58996
rect 42588 58884 42644 58894
rect 42588 58772 42868 58828
rect 42308 57036 42420 57092
rect 42588 58210 42644 58222
rect 42588 58158 42590 58210
rect 42642 58158 42644 58210
rect 42252 57026 42308 57036
rect 42252 56866 42308 56878
rect 42252 56814 42254 56866
rect 42306 56814 42308 56866
rect 42252 56756 42308 56814
rect 42252 56700 42532 56756
rect 42140 56588 42420 56644
rect 41020 55972 41076 56588
rect 40796 53638 40852 53676
rect 40908 55970 41076 55972
rect 40908 55918 41022 55970
rect 41074 55918 41076 55970
rect 40908 55916 41076 55918
rect 40908 52164 40964 55916
rect 41020 55906 41076 55916
rect 42364 56306 42420 56588
rect 42364 56254 42366 56306
rect 42418 56254 42420 56306
rect 42364 55412 42420 56254
rect 42364 55346 42420 55356
rect 42476 55972 42532 56700
rect 41580 55300 41636 55310
rect 41580 55206 41636 55244
rect 41020 55188 41076 55198
rect 41020 55094 41076 55132
rect 42252 55188 42308 55198
rect 42252 55094 42308 55132
rect 41132 55076 41188 55086
rect 41804 55076 41860 55086
rect 41132 55074 41412 55076
rect 41132 55022 41134 55074
rect 41186 55022 41412 55074
rect 41132 55020 41412 55022
rect 41132 55010 41188 55020
rect 41356 54740 41412 55020
rect 41804 54982 41860 55020
rect 42140 55074 42196 55086
rect 42140 55022 42142 55074
rect 42194 55022 42196 55074
rect 41356 54684 41748 54740
rect 41692 54626 41748 54684
rect 41692 54574 41694 54626
rect 41746 54574 41748 54626
rect 41692 54562 41748 54574
rect 41020 54516 41076 54526
rect 41020 54422 41076 54460
rect 42140 54404 42196 55022
rect 42140 53844 42196 54348
rect 41692 53788 42196 53844
rect 42364 55076 42420 55086
rect 42476 55076 42532 55916
rect 42588 55300 42644 58158
rect 42700 56196 42756 56206
rect 42700 56102 42756 56140
rect 42588 55234 42644 55244
rect 42700 55970 42756 55982
rect 42700 55918 42702 55970
rect 42754 55918 42756 55970
rect 42700 55298 42756 55918
rect 42700 55246 42702 55298
rect 42754 55246 42756 55298
rect 42700 55234 42756 55246
rect 42476 55020 42644 55076
rect 41356 53618 41412 53630
rect 41692 53620 41748 53788
rect 42364 53732 42420 55020
rect 42476 53732 42532 53742
rect 42364 53730 42532 53732
rect 42364 53678 42478 53730
rect 42530 53678 42532 53730
rect 42364 53676 42532 53678
rect 42476 53666 42532 53676
rect 41356 53566 41358 53618
rect 41410 53566 41412 53618
rect 41020 53506 41076 53518
rect 41020 53454 41022 53506
rect 41074 53454 41076 53506
rect 41020 53060 41076 53454
rect 41244 53506 41300 53518
rect 41244 53454 41246 53506
rect 41298 53454 41300 53506
rect 41244 53172 41300 53454
rect 41244 53106 41300 53116
rect 41356 53508 41412 53566
rect 41020 52994 41076 53004
rect 40908 52098 40964 52108
rect 41356 51492 41412 53452
rect 41244 51436 41412 51492
rect 41580 53618 41748 53620
rect 41580 53566 41694 53618
rect 41746 53566 41748 53618
rect 41580 53564 41748 53566
rect 41244 51266 41300 51436
rect 41244 51214 41246 51266
rect 41298 51214 41300 51266
rect 40236 50194 40292 50204
rect 40572 50372 40740 50428
rect 41132 50484 41188 50494
rect 41244 50484 41300 51214
rect 41356 51268 41412 51278
rect 41356 50708 41412 51212
rect 41356 50614 41412 50652
rect 41244 50428 41412 50484
rect 40124 50034 40180 50046
rect 40124 49982 40126 50034
rect 40178 49982 40180 50034
rect 40012 49812 40068 49822
rect 40012 49718 40068 49756
rect 39900 49028 39956 49038
rect 39676 48862 39678 48914
rect 39730 48862 39732 48914
rect 39676 48692 39732 48862
rect 39788 48916 39844 48926
rect 39788 48822 39844 48860
rect 39676 48626 39732 48636
rect 39676 48244 39732 48254
rect 39564 48242 39732 48244
rect 39564 48190 39678 48242
rect 39730 48190 39732 48242
rect 39564 48188 39732 48190
rect 39564 47572 39620 47582
rect 39564 47478 39620 47516
rect 39452 46946 39508 46956
rect 38892 42754 38948 43596
rect 38892 42702 38894 42754
rect 38946 42702 38948 42754
rect 38892 42690 38948 42702
rect 39004 43652 39396 43708
rect 39676 43708 39732 48188
rect 39788 47348 39844 47358
rect 39788 47254 39844 47292
rect 39564 43652 39620 43662
rect 39676 43652 39844 43708
rect 38780 42578 38836 42588
rect 37884 42142 37886 42194
rect 37938 42142 37940 42194
rect 37884 42130 37940 42142
rect 37996 42530 38052 42542
rect 37996 42478 37998 42530
rect 38050 42478 38052 42530
rect 37716 41692 37828 41748
rect 37660 41682 37716 41692
rect 37996 41524 38052 42478
rect 38556 41970 38612 41982
rect 38556 41918 38558 41970
rect 38610 41918 38612 41970
rect 37996 41468 38500 41524
rect 38108 41300 38164 41310
rect 38108 41206 38164 41244
rect 38444 40514 38500 41468
rect 38556 41300 38612 41918
rect 39004 41970 39060 43652
rect 39564 43558 39620 43596
rect 39116 43538 39172 43550
rect 39116 43486 39118 43538
rect 39170 43486 39172 43538
rect 39116 42868 39172 43486
rect 39116 42802 39172 42812
rect 39676 42756 39732 42766
rect 39340 42700 39676 42756
rect 39228 42644 39284 42654
rect 39228 42550 39284 42588
rect 39004 41918 39006 41970
rect 39058 41918 39060 41970
rect 39004 41906 39060 41918
rect 39116 42530 39172 42542
rect 39116 42478 39118 42530
rect 39170 42478 39172 42530
rect 38556 41234 38612 41244
rect 38444 40462 38446 40514
rect 38498 40462 38500 40514
rect 38444 40450 38500 40462
rect 38668 40404 38724 40414
rect 38556 40402 38724 40404
rect 38556 40350 38670 40402
rect 38722 40350 38724 40402
rect 38556 40348 38724 40350
rect 37884 40292 37940 40302
rect 37884 39730 37940 40236
rect 37884 39678 37886 39730
rect 37938 39678 37940 39730
rect 37884 39666 37940 39678
rect 37212 39618 37492 39620
rect 37212 39566 37214 39618
rect 37266 39566 37492 39618
rect 37212 39564 37492 39566
rect 37212 39554 37268 39564
rect 38220 39060 38276 39070
rect 38220 38162 38276 39004
rect 38332 38834 38388 38846
rect 38332 38782 38334 38834
rect 38386 38782 38388 38834
rect 38332 38724 38388 38782
rect 38332 38658 38388 38668
rect 38220 38110 38222 38162
rect 38274 38110 38276 38162
rect 38220 38098 38276 38110
rect 37100 37102 37102 37154
rect 37154 37102 37156 37154
rect 37100 37090 37156 37102
rect 37436 38050 37492 38062
rect 37436 37998 37438 38050
rect 37490 37998 37492 38050
rect 37436 37266 37492 37998
rect 37436 37214 37438 37266
rect 37490 37214 37492 37266
rect 37212 36372 37268 36382
rect 37436 36372 37492 37214
rect 37212 36370 37492 36372
rect 37212 36318 37214 36370
rect 37266 36318 37492 36370
rect 37212 36316 37492 36318
rect 38220 37154 38276 37166
rect 38220 37102 38222 37154
rect 38274 37102 38276 37154
rect 37212 35700 37268 36316
rect 38220 35924 38276 37102
rect 38220 35858 38276 35868
rect 38444 36372 38500 36382
rect 38444 36148 38500 36316
rect 38444 35810 38500 36092
rect 38444 35758 38446 35810
rect 38498 35758 38500 35810
rect 38444 35746 38500 35758
rect 37212 35634 37268 35644
rect 38108 35586 38164 35598
rect 38108 35534 38110 35586
rect 38162 35534 38164 35586
rect 37100 35140 37156 35150
rect 37436 35140 37492 35150
rect 37100 35046 37156 35084
rect 37212 35138 37492 35140
rect 37212 35086 37438 35138
rect 37490 35086 37492 35138
rect 37212 35084 37492 35086
rect 37212 35026 37268 35084
rect 37436 35074 37492 35084
rect 38108 35138 38164 35534
rect 38108 35086 38110 35138
rect 38162 35086 38164 35138
rect 37212 34974 37214 35026
rect 37266 34974 37268 35026
rect 37212 34962 37268 34974
rect 37660 34692 37716 34702
rect 36988 34178 37044 34188
rect 37548 34690 37716 34692
rect 37548 34638 37662 34690
rect 37714 34638 37716 34690
rect 37548 34636 37716 34638
rect 37212 34020 37268 34030
rect 36540 33348 36596 33358
rect 36876 33348 36932 33358
rect 36540 33346 36932 33348
rect 36540 33294 36542 33346
rect 36594 33294 36878 33346
rect 36930 33294 36932 33346
rect 36540 33292 36932 33294
rect 36540 33282 36596 33292
rect 36876 33282 36932 33292
rect 37212 33346 37268 33964
rect 37212 33294 37214 33346
rect 37266 33294 37268 33346
rect 37212 33282 37268 33294
rect 37436 33572 37492 33582
rect 36428 33068 36708 33124
rect 36092 32162 36148 32172
rect 36316 32562 36372 32574
rect 36316 32510 36318 32562
rect 36370 32510 36372 32562
rect 35644 31780 35700 31790
rect 35532 31724 35644 31780
rect 35644 31714 35700 31724
rect 36316 31780 36372 32510
rect 36540 32562 36596 32574
rect 36540 32510 36542 32562
rect 36594 32510 36596 32562
rect 36428 32450 36484 32462
rect 36428 32398 36430 32450
rect 36482 32398 36484 32450
rect 36428 32004 36484 32398
rect 36540 32452 36596 32510
rect 36540 32386 36596 32396
rect 36428 31938 36484 31948
rect 36316 31714 36372 31724
rect 36652 31668 36708 33068
rect 37100 33122 37156 33134
rect 37100 33070 37102 33122
rect 37154 33070 37156 33122
rect 37100 32340 37156 33070
rect 37436 32562 37492 33516
rect 37548 33460 37604 34636
rect 37660 34626 37716 34636
rect 37548 33394 37604 33404
rect 37660 33348 37716 33358
rect 37660 33254 37716 33292
rect 38108 33122 38164 35086
rect 38444 34916 38500 34926
rect 38556 34916 38612 40348
rect 38668 40338 38724 40348
rect 38892 40402 38948 40414
rect 38892 40350 38894 40402
rect 38946 40350 38948 40402
rect 38780 40292 38836 40302
rect 38780 40198 38836 40236
rect 38892 39508 38948 40350
rect 39004 40404 39060 40414
rect 39004 40310 39060 40348
rect 39116 39732 39172 42478
rect 39340 42194 39396 42700
rect 39676 42662 39732 42700
rect 39340 42142 39342 42194
rect 39394 42142 39396 42194
rect 39340 42130 39396 42142
rect 39676 41972 39732 41982
rect 39676 41300 39732 41916
rect 39676 41234 39732 41244
rect 39788 40852 39844 43652
rect 39900 42754 39956 48972
rect 40012 48468 40068 48478
rect 40124 48468 40180 49982
rect 40236 50036 40292 50046
rect 40236 49140 40292 49980
rect 40236 49046 40292 49084
rect 40068 48412 40404 48468
rect 40012 48374 40068 48412
rect 40236 48244 40292 48254
rect 40236 48150 40292 48188
rect 40124 48130 40180 48142
rect 40124 48078 40126 48130
rect 40178 48078 40180 48130
rect 40124 47458 40180 48078
rect 40124 47406 40126 47458
rect 40178 47406 40180 47458
rect 40124 47394 40180 47406
rect 40348 47458 40404 48412
rect 40348 47406 40350 47458
rect 40402 47406 40404 47458
rect 40348 47394 40404 47406
rect 40460 48356 40516 48366
rect 40460 48132 40516 48300
rect 40348 46564 40404 46574
rect 40460 46564 40516 48076
rect 40572 47796 40628 50372
rect 41132 49138 41188 50428
rect 41132 49086 41134 49138
rect 41186 49086 41188 49138
rect 41132 49028 41188 49086
rect 41188 48972 41300 49028
rect 41132 48962 41188 48972
rect 41020 48804 41076 48814
rect 41020 48466 41076 48748
rect 41020 48414 41022 48466
rect 41074 48414 41076 48466
rect 40796 48244 40852 48254
rect 40572 47740 40740 47796
rect 40572 47572 40628 47582
rect 40572 47478 40628 47516
rect 40348 46562 40516 46564
rect 40348 46510 40350 46562
rect 40402 46510 40516 46562
rect 40348 46508 40516 46510
rect 40348 43708 40404 46508
rect 40684 44212 40740 47740
rect 40796 47458 40852 48188
rect 40908 48132 40964 48142
rect 40908 48038 40964 48076
rect 41020 47682 41076 48414
rect 41020 47630 41022 47682
rect 41074 47630 41076 47682
rect 41020 47618 41076 47630
rect 40796 47406 40798 47458
rect 40850 47406 40852 47458
rect 40796 46898 40852 47406
rect 40796 46846 40798 46898
rect 40850 46846 40852 46898
rect 40796 46834 40852 46846
rect 41020 47460 41076 47470
rect 41020 46898 41076 47404
rect 41132 47348 41188 47358
rect 41132 47254 41188 47292
rect 41244 47346 41300 48972
rect 41244 47294 41246 47346
rect 41298 47294 41300 47346
rect 41244 47282 41300 47294
rect 41020 46846 41022 46898
rect 41074 46846 41076 46898
rect 41020 46834 41076 46846
rect 41132 47012 41188 47022
rect 41132 46786 41188 46956
rect 41356 46900 41412 50428
rect 41468 48916 41524 48926
rect 41468 48822 41524 48860
rect 41580 48804 41636 53564
rect 41692 53554 41748 53564
rect 41804 53506 41860 53518
rect 41804 53454 41806 53506
rect 41858 53454 41860 53506
rect 41804 53172 41860 53454
rect 42028 53508 42084 53518
rect 42252 53508 42308 53518
rect 42028 53506 42196 53508
rect 42028 53454 42030 53506
rect 42082 53454 42196 53506
rect 42028 53452 42196 53454
rect 42028 53442 42084 53452
rect 41804 53106 41860 53116
rect 42140 52948 42196 53452
rect 42252 53414 42308 53452
rect 42364 53506 42420 53518
rect 42364 53454 42366 53506
rect 42418 53454 42420 53506
rect 42364 53172 42420 53454
rect 42364 53106 42420 53116
rect 42476 53508 42532 53518
rect 42252 52948 42308 52958
rect 42140 52946 42308 52948
rect 42140 52894 42254 52946
rect 42306 52894 42308 52946
rect 42140 52892 42308 52894
rect 42252 52882 42308 52892
rect 42476 52834 42532 53452
rect 42588 53396 42644 55020
rect 42700 53620 42756 53630
rect 42700 53526 42756 53564
rect 42588 53340 42756 53396
rect 42588 53060 42644 53070
rect 42588 52966 42644 53004
rect 42476 52782 42478 52834
rect 42530 52782 42532 52834
rect 42476 52770 42532 52782
rect 42588 52164 42644 52174
rect 42700 52164 42756 53340
rect 42812 53172 42868 58772
rect 42924 58322 42980 58940
rect 42924 58270 42926 58322
rect 42978 58270 42980 58322
rect 42924 58258 42980 58270
rect 43036 58212 43092 59164
rect 43260 59154 43316 59164
rect 43148 59108 43204 59118
rect 43148 58996 43204 59052
rect 43372 58996 43428 60284
rect 43484 59890 43540 59902
rect 43484 59838 43486 59890
rect 43538 59838 43540 59890
rect 43484 59780 43540 59838
rect 43484 59714 43540 59724
rect 43596 59892 43652 60396
rect 43484 59218 43540 59230
rect 43484 59166 43486 59218
rect 43538 59166 43540 59218
rect 43484 59108 43540 59166
rect 43484 59042 43540 59052
rect 43148 58940 43428 58996
rect 43596 58828 43652 59836
rect 43708 60002 43764 60014
rect 43708 59950 43710 60002
rect 43762 59950 43764 60002
rect 43708 59442 43764 59950
rect 43708 59390 43710 59442
rect 43762 59390 43764 59442
rect 43708 59378 43764 59390
rect 43820 59444 43876 61180
rect 44716 60116 44772 64316
rect 44828 60228 44884 65548
rect 44940 65492 44996 65660
rect 44940 65426 44996 65436
rect 45052 64708 45108 67116
rect 45164 66274 45220 68908
rect 45276 67228 45332 69246
rect 45388 69188 45444 69198
rect 45388 69186 47012 69188
rect 45388 69134 45390 69186
rect 45442 69134 47012 69186
rect 45388 69132 47012 69134
rect 45388 69122 45444 69132
rect 45836 68626 45892 68638
rect 45836 68574 45838 68626
rect 45890 68574 45892 68626
rect 45836 67620 45892 68574
rect 46956 67954 47012 69132
rect 50556 69020 50820 69030
rect 50612 68964 50660 69020
rect 50716 68964 50764 69020
rect 50556 68954 50820 68964
rect 46956 67902 46958 67954
rect 47010 67902 47012 67954
rect 46956 67890 47012 67902
rect 47628 67844 47684 67854
rect 45836 67554 45892 67564
rect 47404 67842 47684 67844
rect 47404 67790 47630 67842
rect 47682 67790 47684 67842
rect 47404 67788 47684 67790
rect 45276 67172 45556 67228
rect 45500 67170 45556 67172
rect 45500 67118 45502 67170
rect 45554 67118 45556 67170
rect 45500 67106 45556 67118
rect 45388 67060 45444 67070
rect 45388 66966 45444 67004
rect 45612 67058 45668 67070
rect 45612 67006 45614 67058
rect 45666 67006 45668 67058
rect 45612 66388 45668 67006
rect 45612 66322 45668 66332
rect 45164 66222 45166 66274
rect 45218 66222 45220 66274
rect 45164 66210 45220 66222
rect 45948 66164 46004 66174
rect 45388 66162 46004 66164
rect 45388 66110 45950 66162
rect 46002 66110 46004 66162
rect 45388 66108 46004 66110
rect 45164 66052 45220 66062
rect 45220 65996 45332 66052
rect 45164 65986 45220 65996
rect 45276 65602 45332 65996
rect 45388 65714 45444 66108
rect 45948 66098 46004 66108
rect 45388 65662 45390 65714
rect 45442 65662 45444 65714
rect 45388 65650 45444 65662
rect 45276 65550 45278 65602
rect 45330 65550 45332 65602
rect 45276 65538 45332 65550
rect 45164 64708 45220 64718
rect 45052 64706 45220 64708
rect 45052 64654 45166 64706
rect 45218 64654 45220 64706
rect 45052 64652 45220 64654
rect 45164 64642 45220 64652
rect 45276 64484 45332 64494
rect 45276 64390 45332 64428
rect 45388 64484 45444 64494
rect 45948 64484 46004 64494
rect 45388 64482 46004 64484
rect 45388 64430 45390 64482
rect 45442 64430 45950 64482
rect 46002 64430 46004 64482
rect 45388 64428 46004 64430
rect 45388 64418 45444 64428
rect 45500 64148 45556 64158
rect 45276 64036 45332 64046
rect 45276 61682 45332 63980
rect 45388 63028 45444 63038
rect 45388 62354 45444 62972
rect 45388 62302 45390 62354
rect 45442 62302 45444 62354
rect 45388 62290 45444 62302
rect 45276 61630 45278 61682
rect 45330 61630 45332 61682
rect 45276 61618 45332 61630
rect 44940 61572 44996 61582
rect 44940 61458 44996 61516
rect 44940 61406 44942 61458
rect 44994 61406 44996 61458
rect 44940 61394 44996 61406
rect 45164 61348 45220 61358
rect 45052 61346 45220 61348
rect 45052 61294 45166 61346
rect 45218 61294 45220 61346
rect 45052 61292 45220 61294
rect 45052 60452 45108 61292
rect 45164 61282 45220 61292
rect 45388 61348 45444 61358
rect 45388 61254 45444 61292
rect 45388 60676 45444 60686
rect 45052 60386 45108 60396
rect 45164 60674 45444 60676
rect 45164 60622 45390 60674
rect 45442 60622 45444 60674
rect 45164 60620 45444 60622
rect 44828 60172 45108 60228
rect 44716 60060 44996 60116
rect 44828 59890 44884 59902
rect 44828 59838 44830 59890
rect 44882 59838 44884 59890
rect 44044 59780 44100 59790
rect 44828 59780 44884 59838
rect 44044 59778 44884 59780
rect 44044 59726 44046 59778
rect 44098 59726 44884 59778
rect 44044 59724 44884 59726
rect 44044 59714 44100 59724
rect 43820 59388 44212 59444
rect 43484 58772 43652 58828
rect 43708 59220 43764 59230
rect 43484 58548 43540 58772
rect 43708 58548 43764 59164
rect 43820 59218 43876 59230
rect 43820 59166 43822 59218
rect 43874 59166 43876 59218
rect 43820 58772 43876 59166
rect 44044 59218 44100 59230
rect 44044 59166 44046 59218
rect 44098 59166 44100 59218
rect 43820 58706 43876 58716
rect 43932 58996 43988 59006
rect 43708 58492 43876 58548
rect 43484 58482 43540 58492
rect 43708 58324 43764 58334
rect 43596 58266 43652 58278
rect 43596 58214 43598 58266
rect 43650 58214 43652 58266
rect 43596 58212 43652 58214
rect 43036 58156 43652 58212
rect 43708 58266 43764 58268
rect 43708 58214 43710 58266
rect 43762 58214 43764 58266
rect 43708 58202 43764 58214
rect 43820 58100 43876 58492
rect 43932 58436 43988 58940
rect 44044 58660 44100 59166
rect 44156 58828 44212 59388
rect 44940 59332 44996 60060
rect 44716 59276 44996 59332
rect 44268 59220 44324 59230
rect 44268 59126 44324 59164
rect 44156 58772 44324 58828
rect 44044 58594 44100 58604
rect 43932 58380 44212 58436
rect 43708 58044 43876 58100
rect 43932 58210 43988 58222
rect 43932 58158 43934 58210
rect 43986 58158 43988 58210
rect 43484 57876 43540 57886
rect 43484 57782 43540 57820
rect 43708 57874 43764 58044
rect 43708 57822 43710 57874
rect 43762 57822 43764 57874
rect 43708 57810 43764 57822
rect 43820 57764 43876 57774
rect 43932 57764 43988 58158
rect 43820 57762 43988 57764
rect 43820 57710 43822 57762
rect 43874 57710 43988 57762
rect 43820 57708 43988 57710
rect 43820 57698 43876 57708
rect 44044 56754 44100 56766
rect 44044 56702 44046 56754
rect 44098 56702 44100 56754
rect 43708 56642 43764 56654
rect 43932 56644 43988 56654
rect 43708 56590 43710 56642
rect 43762 56590 43764 56642
rect 43708 56194 43764 56590
rect 43708 56142 43710 56194
rect 43762 56142 43764 56194
rect 43708 56130 43764 56142
rect 43820 56642 43988 56644
rect 43820 56590 43934 56642
rect 43986 56590 43988 56642
rect 43820 56588 43988 56590
rect 43820 56308 43876 56588
rect 43932 56578 43988 56588
rect 42924 56084 42980 56094
rect 42924 54964 42980 56028
rect 43260 56082 43316 56094
rect 43260 56030 43262 56082
rect 43314 56030 43316 56082
rect 43036 55076 43092 55086
rect 43036 54982 43092 55020
rect 42924 54898 42980 54908
rect 43260 54740 43316 56030
rect 43820 55972 43876 56252
rect 44044 56196 44100 56702
rect 44156 56308 44212 58380
rect 44268 56532 44324 58772
rect 44380 58324 44436 58334
rect 44716 58324 44772 59276
rect 45052 59220 45108 60172
rect 45164 59890 45220 60620
rect 45388 60610 45444 60620
rect 45500 60116 45556 64092
rect 45948 63812 46004 64428
rect 46844 64482 46900 64494
rect 46844 64430 46846 64482
rect 46898 64430 46900 64482
rect 46844 64148 46900 64430
rect 46844 64082 46900 64092
rect 47180 64148 47236 64158
rect 47180 64054 47236 64092
rect 47068 64036 47124 64046
rect 47068 63922 47124 63980
rect 47292 64036 47348 64046
rect 47292 63924 47348 63980
rect 47068 63870 47070 63922
rect 47122 63870 47124 63922
rect 47068 63858 47124 63870
rect 47180 63868 47348 63924
rect 46396 63812 46452 63822
rect 45836 63810 46004 63812
rect 45836 63758 45950 63810
rect 46002 63758 46004 63810
rect 45836 63756 46004 63758
rect 45724 63364 45780 63374
rect 45724 61794 45780 63308
rect 45724 61742 45726 61794
rect 45778 61742 45780 61794
rect 45724 61730 45780 61742
rect 45500 60060 45780 60116
rect 45164 59838 45166 59890
rect 45218 59838 45220 59890
rect 45164 59826 45220 59838
rect 45500 59892 45556 59902
rect 45500 59798 45556 59836
rect 45612 59890 45668 59902
rect 45612 59838 45614 59890
rect 45666 59838 45668 59890
rect 45612 59668 45668 59838
rect 45612 59602 45668 59612
rect 44380 58322 44548 58324
rect 44380 58270 44382 58322
rect 44434 58270 44548 58322
rect 44380 58268 44548 58270
rect 44380 58258 44436 58268
rect 44492 58212 44548 58268
rect 44492 58146 44548 58156
rect 44604 58268 44772 58324
rect 44828 59164 45108 59220
rect 45164 59218 45220 59230
rect 45164 59166 45166 59218
rect 45218 59166 45220 59218
rect 44268 56466 44324 56476
rect 44492 56308 44548 56318
rect 44156 56306 44548 56308
rect 44156 56254 44158 56306
rect 44210 56254 44494 56306
rect 44546 56254 44548 56306
rect 44156 56252 44548 56254
rect 44156 56242 44212 56252
rect 44492 56242 44548 56252
rect 43932 56084 43988 56094
rect 43932 55990 43988 56028
rect 43596 55916 43876 55972
rect 43372 55412 43428 55422
rect 43372 55298 43428 55356
rect 43372 55246 43374 55298
rect 43426 55246 43428 55298
rect 43372 55234 43428 55246
rect 43036 54684 43316 54740
rect 43036 53730 43092 54684
rect 43596 54628 43652 55916
rect 44044 55860 44100 56140
rect 43708 55804 44100 55860
rect 44268 55858 44324 55870
rect 44268 55806 44270 55858
rect 44322 55806 44324 55858
rect 43708 55298 43764 55804
rect 43820 55524 43876 55534
rect 43820 55410 43876 55468
rect 43820 55358 43822 55410
rect 43874 55358 43876 55410
rect 43820 55346 43876 55358
rect 43708 55246 43710 55298
rect 43762 55246 43764 55298
rect 43708 55234 43764 55246
rect 43036 53678 43038 53730
rect 43090 53678 43092 53730
rect 43036 53666 43092 53678
rect 43260 54572 43652 54628
rect 43932 55076 43988 55086
rect 43260 53618 43316 54572
rect 43820 54404 43876 54414
rect 43820 54310 43876 54348
rect 43932 53730 43988 55020
rect 44156 54516 44212 54526
rect 44156 54422 44212 54460
rect 43932 53678 43934 53730
rect 43986 53678 43988 53730
rect 43932 53666 43988 53678
rect 44268 53730 44324 55806
rect 44380 55858 44436 55870
rect 44380 55806 44382 55858
rect 44434 55806 44436 55858
rect 44380 55298 44436 55806
rect 44380 55246 44382 55298
rect 44434 55246 44436 55298
rect 44380 55234 44436 55246
rect 44268 53678 44270 53730
rect 44322 53678 44324 53730
rect 44268 53666 44324 53678
rect 43260 53566 43262 53618
rect 43314 53566 43316 53618
rect 43260 53554 43316 53566
rect 43372 53618 43428 53630
rect 43372 53566 43374 53618
rect 43426 53566 43428 53618
rect 43372 53284 43428 53566
rect 43820 53620 43876 53630
rect 43820 53526 43876 53564
rect 43372 53218 43428 53228
rect 43708 53506 43764 53518
rect 43708 53454 43710 53506
rect 43762 53454 43764 53506
rect 43708 53284 43764 53454
rect 43708 53218 43764 53228
rect 43148 53172 43204 53182
rect 42812 53116 42980 53172
rect 42812 53002 42868 53014
rect 42812 52950 42814 53002
rect 42866 52950 42868 53002
rect 42812 52948 42868 52950
rect 42812 52882 42868 52892
rect 42644 52108 42756 52164
rect 41804 51492 41860 51502
rect 41804 50818 41860 51436
rect 41804 50766 41806 50818
rect 41858 50766 41860 50818
rect 41804 50754 41860 50766
rect 41916 50932 41972 50942
rect 41580 48710 41636 48748
rect 41692 50708 41748 50718
rect 41692 50594 41748 50652
rect 41692 50542 41694 50594
rect 41746 50542 41748 50594
rect 41468 48244 41524 48254
rect 41468 48150 41524 48188
rect 41692 47908 41748 50542
rect 41916 50708 41972 50876
rect 42364 50708 42420 50718
rect 41916 50652 42364 50708
rect 41804 50484 41860 50494
rect 41916 50484 41972 50652
rect 42364 50614 42420 50652
rect 41804 50482 41972 50484
rect 41804 50430 41806 50482
rect 41858 50430 41972 50482
rect 41804 50428 41972 50430
rect 41804 50418 41860 50428
rect 42252 49924 42308 49934
rect 42252 49922 42420 49924
rect 42252 49870 42254 49922
rect 42306 49870 42420 49922
rect 42252 49868 42420 49870
rect 42252 49858 42308 49868
rect 42140 49812 42196 49822
rect 41804 49810 42196 49812
rect 41804 49758 42142 49810
rect 42194 49758 42196 49810
rect 41804 49756 42196 49758
rect 41804 49026 41860 49756
rect 42140 49746 42196 49756
rect 42140 49588 42196 49598
rect 41804 48974 41806 49026
rect 41858 48974 41860 49026
rect 41804 48962 41860 48974
rect 42028 49028 42084 49038
rect 41356 46834 41412 46844
rect 41468 47852 41748 47908
rect 41804 48580 41860 48590
rect 41132 46734 41134 46786
rect 41186 46734 41188 46786
rect 41132 46722 41188 46734
rect 40908 46004 40964 46014
rect 40908 45106 40964 45948
rect 40908 45054 40910 45106
rect 40962 45054 40964 45106
rect 40908 45042 40964 45054
rect 40684 44146 40740 44156
rect 41356 44548 41412 44558
rect 40348 43652 40740 43708
rect 39900 42702 39902 42754
rect 39954 42702 39956 42754
rect 39900 42690 39956 42702
rect 40236 42754 40292 42766
rect 40236 42702 40238 42754
rect 40290 42702 40292 42754
rect 40236 42644 40292 42702
rect 40572 42756 40628 42766
rect 40572 42662 40628 42700
rect 40684 42754 40740 43652
rect 41356 43650 41412 44492
rect 41356 43598 41358 43650
rect 41410 43598 41412 43650
rect 41356 43586 41412 43598
rect 40908 43538 40964 43550
rect 40908 43486 40910 43538
rect 40962 43486 40964 43538
rect 40908 43428 40964 43486
rect 40684 42702 40686 42754
rect 40738 42702 40740 42754
rect 40684 42690 40740 42702
rect 40796 43372 40908 43428
rect 40236 42578 40292 42588
rect 39788 40786 39844 40796
rect 40012 42530 40068 42542
rect 40012 42478 40014 42530
rect 40066 42478 40068 42530
rect 39564 40404 39620 40414
rect 39564 40310 39620 40348
rect 39676 40402 39732 40414
rect 39676 40350 39678 40402
rect 39730 40350 39732 40402
rect 39116 39676 39620 39732
rect 38892 39452 39396 39508
rect 39340 39058 39396 39452
rect 39340 39006 39342 39058
rect 39394 39006 39396 39058
rect 39340 38994 39396 39006
rect 39452 38948 39508 38958
rect 39452 38854 39508 38892
rect 38892 38724 38948 38734
rect 39564 38724 39620 39676
rect 39676 38836 39732 40350
rect 39900 40402 39956 40414
rect 39900 40350 39902 40402
rect 39954 40350 39956 40402
rect 39788 40290 39844 40302
rect 39788 40238 39790 40290
rect 39842 40238 39844 40290
rect 39788 39060 39844 40238
rect 39788 38994 39844 39004
rect 39676 38770 39732 38780
rect 38892 38630 38948 38668
rect 39452 38668 39620 38724
rect 39900 38668 39956 40350
rect 40012 40402 40068 42478
rect 40796 42532 40852 43372
rect 40908 43362 40964 43372
rect 41132 43426 41188 43438
rect 41132 43374 41134 43426
rect 41186 43374 41188 43426
rect 41020 42644 41076 42654
rect 41020 42550 41076 42588
rect 40796 42466 40852 42476
rect 40908 42530 40964 42542
rect 40908 42478 40910 42530
rect 40962 42478 40964 42530
rect 40908 42084 40964 42478
rect 41020 42084 41076 42094
rect 40908 42082 41076 42084
rect 40908 42030 41022 42082
rect 41074 42030 41076 42082
rect 40908 42028 41076 42030
rect 41020 42018 41076 42028
rect 41020 41860 41076 41870
rect 40012 40350 40014 40402
rect 40066 40350 40068 40402
rect 40012 40338 40068 40350
rect 40908 41804 41020 41860
rect 40908 40404 40964 41804
rect 41020 41794 41076 41804
rect 41132 41636 41188 43374
rect 41356 42756 41412 42766
rect 41468 42756 41524 47852
rect 41580 47236 41636 47246
rect 41580 46898 41636 47180
rect 41580 46846 41582 46898
rect 41634 46846 41636 46898
rect 41580 46834 41636 46846
rect 41804 47234 41860 48524
rect 41804 47182 41806 47234
rect 41858 47182 41860 47234
rect 41804 46674 41860 47182
rect 41916 48244 41972 48254
rect 41916 47124 41972 48188
rect 42028 47682 42084 48972
rect 42028 47630 42030 47682
rect 42082 47630 42084 47682
rect 42028 47618 42084 47630
rect 41916 47012 42084 47068
rect 41804 46622 41806 46674
rect 41858 46622 41860 46674
rect 41692 46562 41748 46574
rect 41692 46510 41694 46562
rect 41746 46510 41748 46562
rect 41692 45218 41748 46510
rect 41804 45444 41860 46622
rect 42028 46674 42084 47012
rect 42028 46622 42030 46674
rect 42082 46622 42084 46674
rect 42028 46610 42084 46622
rect 42140 46340 42196 49532
rect 42252 48916 42308 48926
rect 42252 48822 42308 48860
rect 42364 48914 42420 49868
rect 42364 48862 42366 48914
rect 42418 48862 42420 48914
rect 42364 48468 42420 48862
rect 42364 48402 42420 48412
rect 42476 49810 42532 49822
rect 42476 49758 42478 49810
rect 42530 49758 42532 49810
rect 42476 48356 42532 49758
rect 42476 48290 42532 48300
rect 42476 48130 42532 48142
rect 42476 48078 42478 48130
rect 42530 48078 42532 48130
rect 42476 48018 42532 48078
rect 42476 47966 42478 48018
rect 42530 47966 42532 48018
rect 42476 47954 42532 47966
rect 42252 47682 42308 47694
rect 42252 47630 42254 47682
rect 42306 47630 42308 47682
rect 42252 47570 42308 47630
rect 42252 47518 42254 47570
rect 42306 47518 42308 47570
rect 42252 47506 42308 47518
rect 42588 47348 42644 52108
rect 42700 50260 42756 50270
rect 42700 49026 42756 50204
rect 42924 49588 42980 53116
rect 43148 53058 43204 53116
rect 43148 53006 43150 53058
rect 43202 53006 43204 53058
rect 43148 52994 43204 53006
rect 43260 52722 43316 52734
rect 43260 52670 43262 52722
rect 43314 52670 43316 52722
rect 43260 51492 43316 52670
rect 44268 52164 44324 52174
rect 44268 52070 44324 52108
rect 44156 52052 44212 52062
rect 43372 51492 43428 51502
rect 43260 51490 43428 51492
rect 43260 51438 43374 51490
rect 43426 51438 43428 51490
rect 43260 51436 43428 51438
rect 43372 51426 43428 51436
rect 44156 51378 44212 51996
rect 44156 51326 44158 51378
rect 44210 51326 44212 51378
rect 44156 51314 44212 51326
rect 43820 51268 43876 51278
rect 43148 50596 43204 50606
rect 43484 50596 43540 50606
rect 43148 50594 43484 50596
rect 43148 50542 43150 50594
rect 43202 50542 43484 50594
rect 43148 50540 43484 50542
rect 43148 50036 43204 50540
rect 43484 50502 43540 50540
rect 43820 50594 43876 51212
rect 43820 50542 43822 50594
rect 43874 50542 43876 50594
rect 43148 49970 43204 49980
rect 43820 50036 43876 50542
rect 43932 50540 44436 50596
rect 43932 50482 43988 50540
rect 43932 50430 43934 50482
rect 43986 50430 43988 50482
rect 43932 50418 43988 50430
rect 43820 49970 43876 49980
rect 44044 50370 44100 50382
rect 44044 50318 44046 50370
rect 44098 50318 44100 50370
rect 42924 49522 42980 49532
rect 43148 49810 43204 49822
rect 43148 49758 43150 49810
rect 43202 49758 43204 49810
rect 43148 49140 43204 49758
rect 43484 49812 43540 49822
rect 43484 49718 43540 49756
rect 43708 49812 43764 49822
rect 43932 49812 43988 49822
rect 44044 49812 44100 50318
rect 43708 49810 44100 49812
rect 43708 49758 43710 49810
rect 43762 49758 43934 49810
rect 43986 49758 44100 49810
rect 43708 49756 44100 49758
rect 44268 49812 44324 49822
rect 44380 49812 44436 50540
rect 44492 49812 44548 49822
rect 44380 49810 44548 49812
rect 44380 49758 44494 49810
rect 44546 49758 44548 49810
rect 44380 49756 44548 49758
rect 43596 49698 43652 49710
rect 43596 49646 43598 49698
rect 43650 49646 43652 49698
rect 43596 49252 43652 49646
rect 43484 49196 43652 49252
rect 43148 49138 43428 49140
rect 43148 49086 43150 49138
rect 43202 49086 43428 49138
rect 43148 49084 43428 49086
rect 43148 49074 43204 49084
rect 42700 48974 42702 49026
rect 42754 48974 42756 49026
rect 42700 48018 42756 48974
rect 42924 48804 42980 48814
rect 42924 48710 42980 48748
rect 43148 48804 43204 48814
rect 43148 48710 43204 48748
rect 43372 48466 43428 49084
rect 43372 48414 43374 48466
rect 43426 48414 43428 48466
rect 43372 48402 43428 48414
rect 43260 48356 43316 48366
rect 43260 48262 43316 48300
rect 42700 47966 42702 48018
rect 42754 47966 42756 48018
rect 42700 47954 42756 47966
rect 42924 48130 42980 48142
rect 42924 48078 42926 48130
rect 42978 48078 42980 48130
rect 42924 47908 42980 48078
rect 42924 47842 42980 47852
rect 42476 47292 42644 47348
rect 42924 47348 42980 47358
rect 42476 47068 42532 47292
rect 42924 47254 42980 47292
rect 43372 47346 43428 47358
rect 43372 47294 43374 47346
rect 43426 47294 43428 47346
rect 42700 47234 42756 47246
rect 42700 47182 42702 47234
rect 42754 47182 42756 47234
rect 42364 47012 42420 47022
rect 42476 47012 42644 47068
rect 42364 46676 42420 46956
rect 42588 46788 42644 47012
rect 42700 46900 42756 47182
rect 42812 47234 42868 47246
rect 42812 47182 42814 47234
rect 42866 47182 42868 47234
rect 42812 47068 42868 47182
rect 43260 47236 43316 47246
rect 43260 47142 43316 47180
rect 42812 47012 43316 47068
rect 43260 46946 43316 46956
rect 42700 46844 43092 46900
rect 42588 46722 42644 46732
rect 42476 46676 42532 46686
rect 42364 46674 42532 46676
rect 42364 46622 42478 46674
rect 42530 46622 42532 46674
rect 42364 46620 42532 46622
rect 42476 46610 42532 46620
rect 42924 46676 42980 46686
rect 42924 46582 42980 46620
rect 43036 46676 43092 46844
rect 43036 46674 43316 46676
rect 43036 46622 43038 46674
rect 43090 46622 43316 46674
rect 43036 46620 43316 46622
rect 43036 46610 43092 46620
rect 42252 46562 42308 46574
rect 42252 46510 42254 46562
rect 42306 46510 42308 46562
rect 42252 46452 42308 46510
rect 42700 46562 42756 46574
rect 42700 46510 42702 46562
rect 42754 46510 42756 46562
rect 42700 46452 42756 46510
rect 42252 46396 42756 46452
rect 42812 46564 42868 46574
rect 42140 46284 42308 46340
rect 41804 45378 41860 45388
rect 41692 45166 41694 45218
rect 41746 45166 41748 45218
rect 41692 45154 41748 45166
rect 41580 44212 41636 44222
rect 41580 44118 41636 44156
rect 42140 44212 42196 44222
rect 42140 43650 42196 44156
rect 42252 43708 42308 46284
rect 42812 45890 42868 46508
rect 43260 46114 43316 46620
rect 43260 46062 43262 46114
rect 43314 46062 43316 46114
rect 43260 46050 43316 46062
rect 42812 45838 42814 45890
rect 42866 45838 42868 45890
rect 42812 44546 42868 45838
rect 42812 44494 42814 44546
rect 42866 44494 42868 44546
rect 42812 44436 42868 44494
rect 42812 44370 42868 44380
rect 42924 45220 42980 45230
rect 42924 44434 42980 45164
rect 43372 44996 43428 47294
rect 43484 46676 43540 49196
rect 43596 48916 43652 48926
rect 43596 48822 43652 48860
rect 43708 48692 43764 49756
rect 43932 49746 43988 49756
rect 44268 49718 44324 49756
rect 44492 49746 44548 49756
rect 44156 49698 44212 49710
rect 44156 49646 44158 49698
rect 44210 49646 44212 49698
rect 44156 49364 44212 49646
rect 43820 49308 44212 49364
rect 43820 49250 43876 49308
rect 43820 49198 43822 49250
rect 43874 49198 43876 49250
rect 43820 49186 43876 49198
rect 44604 49140 44660 58268
rect 44716 58100 44772 58110
rect 44716 56308 44772 58044
rect 44828 57764 44884 59164
rect 44940 58884 44996 58894
rect 44940 58436 44996 58828
rect 45164 58772 45220 59166
rect 45500 59108 45556 59118
rect 45276 58996 45332 59006
rect 45276 58902 45332 58940
rect 45500 58828 45556 59052
rect 45724 59108 45780 60060
rect 45724 59042 45780 59052
rect 45836 58828 45892 63756
rect 45948 63746 46004 63756
rect 46060 63810 46452 63812
rect 46060 63758 46398 63810
rect 46450 63758 46452 63810
rect 46060 63756 46452 63758
rect 46060 63028 46116 63756
rect 46396 63746 46452 63756
rect 47180 63698 47236 63868
rect 47180 63646 47182 63698
rect 47234 63646 47236 63698
rect 47180 63634 47236 63646
rect 44940 58380 45108 58436
rect 44940 58212 44996 58222
rect 44940 58118 44996 58156
rect 45052 57876 45108 58380
rect 45164 58212 45220 58716
rect 45388 58772 45556 58828
rect 45612 58772 45892 58828
rect 45948 62972 46116 63028
rect 45948 61570 46004 62972
rect 46060 62242 46116 62254
rect 46060 62190 46062 62242
rect 46114 62190 46116 62242
rect 46060 62188 46116 62190
rect 47404 62244 47460 67788
rect 47628 67778 47684 67788
rect 50556 67452 50820 67462
rect 50612 67396 50660 67452
rect 50716 67396 50764 67452
rect 50556 67386 50820 67396
rect 48076 66386 48132 66398
rect 48076 66334 48078 66386
rect 48130 66334 48132 66386
rect 46060 62132 46340 62188
rect 46284 61682 46340 62132
rect 46284 61630 46286 61682
rect 46338 61630 46340 61682
rect 46284 61618 46340 61630
rect 47292 62132 47460 62188
rect 47516 65602 47572 65614
rect 47516 65550 47518 65602
rect 47570 65550 47572 65602
rect 47516 65492 47572 65550
rect 47516 62188 47572 65436
rect 47852 65492 47908 65502
rect 48076 65492 48132 66334
rect 50556 65884 50820 65894
rect 50612 65828 50660 65884
rect 50716 65828 50764 65884
rect 50556 65818 50820 65828
rect 47852 65490 48132 65492
rect 47852 65438 47854 65490
rect 47906 65438 48132 65490
rect 47852 65436 48132 65438
rect 47852 65426 47908 65436
rect 47628 64036 47684 64046
rect 47628 63942 47684 63980
rect 47852 63922 47908 63934
rect 47852 63870 47854 63922
rect 47906 63870 47908 63922
rect 47740 63810 47796 63822
rect 47740 63758 47742 63810
rect 47794 63758 47796 63810
rect 47740 62188 47796 63758
rect 47852 63028 47908 63870
rect 47964 63476 48020 65436
rect 50556 64316 50820 64326
rect 50612 64260 50660 64316
rect 50716 64260 50764 64316
rect 50556 64250 50820 64260
rect 48188 64036 48244 64046
rect 48076 63476 48132 63486
rect 47964 63420 48076 63476
rect 48076 63410 48132 63420
rect 47852 62962 47908 62972
rect 48188 62242 48244 63980
rect 48972 64036 49028 64046
rect 48972 63942 49028 63980
rect 48188 62190 48190 62242
rect 48242 62190 48244 62242
rect 47516 62132 47684 62188
rect 47740 62132 48132 62188
rect 48188 62178 48244 62190
rect 48300 63922 48356 63934
rect 48300 63870 48302 63922
rect 48354 63870 48356 63922
rect 48300 62188 48356 63870
rect 48748 63924 48804 63934
rect 48748 63138 48804 63868
rect 49420 63924 49476 63934
rect 49420 63830 49476 63868
rect 48860 63700 48916 63710
rect 48860 63698 49140 63700
rect 48860 63646 48862 63698
rect 48914 63646 49140 63698
rect 48860 63644 49140 63646
rect 48860 63634 48916 63644
rect 48748 63086 48750 63138
rect 48802 63086 48804 63138
rect 48748 62354 48804 63086
rect 48748 62302 48750 62354
rect 48802 62302 48804 62354
rect 48748 62290 48804 62302
rect 48860 63476 48916 63486
rect 48300 62132 48804 62188
rect 45948 61518 45950 61570
rect 46002 61518 46004 61570
rect 45948 60340 46004 61518
rect 46396 61572 46452 61582
rect 47292 61572 47348 62132
rect 46396 61478 46452 61516
rect 47180 61570 47348 61572
rect 47180 61518 47294 61570
rect 47346 61518 47348 61570
rect 47180 61516 47348 61518
rect 46172 61460 46228 61470
rect 46172 61366 46228 61404
rect 46956 61348 47012 61358
rect 46844 61346 47012 61348
rect 46844 61294 46958 61346
rect 47010 61294 47012 61346
rect 46844 61292 47012 61294
rect 46172 60788 46228 60798
rect 46172 60694 46228 60732
rect 45276 58660 45332 58670
rect 45276 58546 45332 58604
rect 45276 58494 45278 58546
rect 45330 58494 45332 58546
rect 45276 58482 45332 58494
rect 45388 58212 45444 58772
rect 45164 58118 45220 58156
rect 45276 58210 45444 58212
rect 45276 58158 45390 58210
rect 45442 58158 45444 58210
rect 45276 58156 45444 58158
rect 45276 58100 45332 58156
rect 45388 58146 45444 58156
rect 45276 58034 45332 58044
rect 45388 57988 45444 57998
rect 45164 57876 45220 57886
rect 45052 57874 45220 57876
rect 45052 57822 45166 57874
rect 45218 57822 45220 57874
rect 45052 57820 45220 57822
rect 45164 57810 45220 57820
rect 44828 57698 44884 57708
rect 45276 57764 45332 57774
rect 44940 57650 44996 57662
rect 44940 57598 44942 57650
rect 44994 57598 44996 57650
rect 44940 57204 44996 57598
rect 45276 57650 45332 57708
rect 45276 57598 45278 57650
rect 45330 57598 45332 57650
rect 45276 57586 45332 57598
rect 44716 56252 44884 56308
rect 44716 56084 44772 56094
rect 44716 55990 44772 56028
rect 44828 53844 44884 56252
rect 44940 55300 44996 57148
rect 45388 56532 45444 57932
rect 45612 57876 45668 58772
rect 45948 58660 46004 60284
rect 46396 60564 46452 60574
rect 46396 60002 46452 60508
rect 46844 60564 46900 61292
rect 46956 61282 47012 61292
rect 46396 59950 46398 60002
rect 46450 59950 46452 60002
rect 46396 59938 46452 59950
rect 46732 60004 46788 60014
rect 46732 59910 46788 59948
rect 46060 59778 46116 59790
rect 46060 59726 46062 59778
rect 46114 59726 46116 59778
rect 46060 59668 46116 59726
rect 46060 59444 46116 59612
rect 46844 59444 46900 60508
rect 46956 60786 47012 60798
rect 46956 60734 46958 60786
rect 47010 60734 47012 60786
rect 46956 60114 47012 60734
rect 46956 60062 46958 60114
rect 47010 60062 47012 60114
rect 46956 60050 47012 60062
rect 47180 60788 47236 61516
rect 47292 61506 47348 61516
rect 47516 61572 47572 61582
rect 46956 59892 47012 59902
rect 46956 59798 47012 59836
rect 46060 59388 46676 59444
rect 46844 59388 47124 59444
rect 46172 59218 46228 59230
rect 46172 59166 46174 59218
rect 46226 59166 46228 59218
rect 45948 58594 46004 58604
rect 46060 59108 46116 59118
rect 45948 58434 46004 58446
rect 45948 58382 45950 58434
rect 46002 58382 46004 58434
rect 45836 58212 45892 58222
rect 45836 58118 45892 58156
rect 45276 56476 45444 56532
rect 45500 57820 45668 57876
rect 45948 57876 46004 58382
rect 46060 58100 46116 59052
rect 46172 58884 46228 59166
rect 46172 58818 46228 58828
rect 46508 59218 46564 59230
rect 46508 59166 46510 59218
rect 46562 59166 46564 59218
rect 46060 58034 46116 58044
rect 46508 57876 46564 59166
rect 46620 58100 46676 59388
rect 46956 59220 47012 59230
rect 46844 59164 46956 59220
rect 46844 58436 46900 59164
rect 46956 59126 47012 59164
rect 46844 58434 47012 58436
rect 46844 58382 46846 58434
rect 46898 58382 47012 58434
rect 46844 58380 47012 58382
rect 46844 58370 46900 58380
rect 46732 58324 46788 58334
rect 46732 58230 46788 58268
rect 46620 58044 46900 58100
rect 46732 57876 46788 57886
rect 45948 57874 46788 57876
rect 45948 57822 46734 57874
rect 46786 57822 46788 57874
rect 45948 57820 46788 57822
rect 45164 56196 45220 56206
rect 45052 56194 45220 56196
rect 45052 56142 45166 56194
rect 45218 56142 45220 56194
rect 45052 56140 45220 56142
rect 45052 56082 45108 56140
rect 45164 56130 45220 56140
rect 45052 56030 45054 56082
rect 45106 56030 45108 56082
rect 45052 56018 45108 56030
rect 45276 56084 45332 56476
rect 45500 56420 45556 57820
rect 46732 57810 46788 57820
rect 45612 57650 45668 57662
rect 45612 57598 45614 57650
rect 45666 57598 45668 57650
rect 45612 57540 45668 57598
rect 46060 57650 46116 57662
rect 46060 57598 46062 57650
rect 46114 57598 46116 57650
rect 46060 57540 46116 57598
rect 46172 57652 46228 57662
rect 46172 57558 46228 57596
rect 46284 57652 46340 57662
rect 46284 57650 46564 57652
rect 46284 57598 46286 57650
rect 46338 57598 46564 57650
rect 46284 57596 46564 57598
rect 46284 57586 46340 57596
rect 45612 57474 45668 57484
rect 45836 57484 46060 57540
rect 45836 56978 45892 57484
rect 46060 57474 46116 57484
rect 45836 56926 45838 56978
rect 45890 56926 45892 56978
rect 45836 56914 45892 56926
rect 46508 57428 46564 57596
rect 45388 56308 45444 56318
rect 45388 56214 45444 56252
rect 45500 56194 45556 56364
rect 46396 56420 46452 56430
rect 46396 56306 46452 56364
rect 46396 56254 46398 56306
rect 46450 56254 46452 56306
rect 46396 56242 46452 56254
rect 45500 56142 45502 56194
rect 45554 56142 45556 56194
rect 45500 56130 45556 56142
rect 45276 56028 45444 56084
rect 44940 55244 45108 55300
rect 44940 54402 44996 54414
rect 44940 54350 44942 54402
rect 44994 54350 44996 54402
rect 44940 53954 44996 54350
rect 44940 53902 44942 53954
rect 44994 53902 44996 53954
rect 44940 53890 44996 53902
rect 44716 53788 44884 53844
rect 44716 50596 44772 53788
rect 45052 53732 45108 55244
rect 45164 55298 45220 55310
rect 45164 55246 45166 55298
rect 45218 55246 45220 55298
rect 45164 54516 45220 55246
rect 45164 54450 45220 54460
rect 44940 53676 45108 53732
rect 44828 53620 44884 53630
rect 44828 53526 44884 53564
rect 44828 51492 44884 51502
rect 44940 51492 44996 53676
rect 45052 53284 45108 53294
rect 45108 53228 45220 53284
rect 45052 53218 45108 53228
rect 45052 52836 45108 52846
rect 45052 51602 45108 52780
rect 45052 51550 45054 51602
rect 45106 51550 45108 51602
rect 45052 51538 45108 51550
rect 44828 51490 44996 51492
rect 44828 51438 44830 51490
rect 44882 51438 44996 51490
rect 44828 51436 44996 51438
rect 45164 51490 45220 53228
rect 45388 53060 45444 56028
rect 45836 55970 45892 55982
rect 46508 55972 46564 57372
rect 46732 57092 46788 57102
rect 46732 56644 46788 57036
rect 46732 56550 46788 56588
rect 45836 55918 45838 55970
rect 45890 55918 45892 55970
rect 45836 55524 45892 55918
rect 46396 55916 46564 55972
rect 45836 55458 45892 55468
rect 45948 55858 46004 55870
rect 45948 55806 45950 55858
rect 46002 55806 46004 55858
rect 45948 55410 46004 55806
rect 45948 55358 45950 55410
rect 46002 55358 46004 55410
rect 45948 55346 46004 55358
rect 45388 52966 45444 53004
rect 45500 54516 45556 54526
rect 45500 52274 45556 54460
rect 45948 53284 46004 53294
rect 45948 53058 46004 53228
rect 45948 53006 45950 53058
rect 46002 53006 46004 53058
rect 45948 52994 46004 53006
rect 46060 53060 46116 53070
rect 46396 53060 46452 55916
rect 46732 53844 46788 53854
rect 46732 53730 46788 53788
rect 46732 53678 46734 53730
rect 46786 53678 46788 53730
rect 46508 53506 46564 53518
rect 46508 53454 46510 53506
rect 46562 53454 46564 53506
rect 46508 53172 46564 53454
rect 46620 53508 46676 53518
rect 46620 53414 46676 53452
rect 46508 53106 46564 53116
rect 46060 53058 46452 53060
rect 46060 53006 46062 53058
rect 46114 53006 46452 53058
rect 46060 53004 46452 53006
rect 46060 52994 46116 53004
rect 45500 52222 45502 52274
rect 45554 52222 45556 52274
rect 45500 52052 45556 52222
rect 45164 51438 45166 51490
rect 45218 51438 45220 51490
rect 44828 51426 44884 51436
rect 45164 51426 45220 51438
rect 45388 51492 45444 51502
rect 45388 51398 45444 51436
rect 44716 50530 44772 50540
rect 45388 49698 45444 49710
rect 45388 49646 45390 49698
rect 45442 49646 45444 49698
rect 44940 49140 44996 49150
rect 44268 49138 45220 49140
rect 44268 49086 44942 49138
rect 44994 49086 45220 49138
rect 44268 49084 45220 49086
rect 43596 48636 43764 48692
rect 43932 48804 43988 48814
rect 43596 48466 43652 48636
rect 43596 48414 43598 48466
rect 43650 48414 43652 48466
rect 43596 48402 43652 48414
rect 43820 48468 43876 48478
rect 43820 48374 43876 48412
rect 43932 48132 43988 48748
rect 44156 48804 44212 48814
rect 44156 48710 44212 48748
rect 43932 48038 43988 48076
rect 43596 48020 43652 48030
rect 43596 47458 43652 47964
rect 43596 47406 43598 47458
rect 43650 47406 43652 47458
rect 43596 47394 43652 47406
rect 44044 47572 44100 47582
rect 44268 47572 44324 49084
rect 44940 49074 44996 49084
rect 44828 48468 44884 48478
rect 45164 48468 45220 49084
rect 45276 48914 45332 48926
rect 45276 48862 45278 48914
rect 45330 48862 45332 48914
rect 45276 48804 45332 48862
rect 45276 48738 45332 48748
rect 45388 48580 45444 49646
rect 45388 48514 45444 48524
rect 44884 48412 45108 48468
rect 45164 48412 45332 48468
rect 44828 48374 44884 48412
rect 45052 48356 45108 48412
rect 45052 48300 45220 48356
rect 44044 47458 44100 47516
rect 44044 47406 44046 47458
rect 44098 47406 44100 47458
rect 44044 47394 44100 47406
rect 44156 47516 44324 47572
rect 44380 48130 44436 48142
rect 44380 48078 44382 48130
rect 44434 48078 44436 48130
rect 44380 48020 44436 48078
rect 43932 47236 43988 47246
rect 43932 47142 43988 47180
rect 43484 45892 43540 46620
rect 43708 47012 43764 47022
rect 43708 46452 43764 46956
rect 43708 46358 43764 46396
rect 43820 46900 43876 46910
rect 43484 45826 43540 45836
rect 43820 45890 43876 46844
rect 44156 46676 44212 47516
rect 44268 47346 44324 47358
rect 44268 47294 44270 47346
rect 44322 47294 44324 47346
rect 44268 47012 44324 47294
rect 44268 46946 44324 46956
rect 44380 46786 44436 47964
rect 45164 47572 45220 48300
rect 45164 47458 45220 47516
rect 45164 47406 45166 47458
rect 45218 47406 45220 47458
rect 45164 47394 45220 47406
rect 45276 47458 45332 48412
rect 45388 48244 45444 48254
rect 45500 48244 45556 51996
rect 45724 52946 45780 52958
rect 45724 52894 45726 52946
rect 45778 52894 45780 52946
rect 45724 51492 45780 52894
rect 46508 52948 46564 52958
rect 46508 52722 46564 52892
rect 46508 52670 46510 52722
rect 46562 52670 46564 52722
rect 46508 52388 46564 52670
rect 45724 51426 45780 51436
rect 46284 52332 46564 52388
rect 46172 51380 46228 51390
rect 46284 51380 46340 52332
rect 46732 51492 46788 53678
rect 46732 51398 46788 51436
rect 46172 51378 46340 51380
rect 46172 51326 46174 51378
rect 46226 51326 46340 51378
rect 46172 51324 46340 51326
rect 46172 51314 46228 51324
rect 46396 51268 46452 51278
rect 46396 51174 46452 51212
rect 46732 50708 46788 50718
rect 46732 50614 46788 50652
rect 45948 50036 46004 50046
rect 45836 49980 45948 50036
rect 45836 49922 45892 49980
rect 45948 49970 46004 49980
rect 45836 49870 45838 49922
rect 45890 49870 45892 49922
rect 45836 49028 45892 49870
rect 45948 49252 46004 49262
rect 45948 49250 46340 49252
rect 45948 49198 45950 49250
rect 46002 49198 46340 49250
rect 45948 49196 46340 49198
rect 45948 49186 46004 49196
rect 46172 49028 46228 49038
rect 45836 49026 46228 49028
rect 45836 48974 46174 49026
rect 46226 48974 46228 49026
rect 45836 48972 46228 48974
rect 45612 48804 45668 48814
rect 45612 48802 46116 48804
rect 45612 48750 45614 48802
rect 45666 48750 46116 48802
rect 45612 48748 46116 48750
rect 45612 48738 45668 48748
rect 46060 48354 46116 48748
rect 46060 48302 46062 48354
rect 46114 48302 46116 48354
rect 46060 48290 46116 48302
rect 45388 48242 45556 48244
rect 45388 48190 45390 48242
rect 45442 48190 45556 48242
rect 45388 48188 45556 48190
rect 46172 48244 46228 48972
rect 45388 48178 45444 48188
rect 46172 48178 46228 48188
rect 45276 47406 45278 47458
rect 45330 47406 45332 47458
rect 45276 47394 45332 47406
rect 45724 47460 45780 47470
rect 45724 47366 45780 47404
rect 44492 47348 44548 47358
rect 44492 46898 44548 47292
rect 45052 47346 45108 47358
rect 45948 47348 46004 47358
rect 45052 47294 45054 47346
rect 45106 47294 45108 47346
rect 45052 47012 45108 47294
rect 44492 46846 44494 46898
rect 44546 46846 44548 46898
rect 44492 46834 44548 46846
rect 44604 46900 44660 46910
rect 44380 46734 44382 46786
rect 44434 46734 44436 46786
rect 44380 46722 44436 46734
rect 43820 45838 43822 45890
rect 43874 45838 43876 45890
rect 43820 45826 43876 45838
rect 43932 46620 44212 46676
rect 44604 46674 44660 46844
rect 45052 46788 45108 46956
rect 45836 47292 45948 47348
rect 45052 46732 45332 46788
rect 44604 46622 44606 46674
rect 44658 46622 44660 46674
rect 43708 45778 43764 45790
rect 43708 45726 43710 45778
rect 43762 45726 43764 45778
rect 43708 45668 43764 45726
rect 43932 45668 43988 46620
rect 44604 46610 44660 46622
rect 44940 46676 44996 46686
rect 44940 46674 45220 46676
rect 44940 46622 44942 46674
rect 44994 46622 45220 46674
rect 44940 46620 45220 46622
rect 44940 46610 44996 46620
rect 44044 46452 44100 46462
rect 44828 46452 44884 46462
rect 44044 46450 44436 46452
rect 44044 46398 44046 46450
rect 44098 46398 44436 46450
rect 44044 46396 44436 46398
rect 44044 46386 44100 46396
rect 43708 45612 43988 45668
rect 44044 45890 44100 45902
rect 44044 45838 44046 45890
rect 44098 45838 44100 45890
rect 43708 45220 43764 45612
rect 43708 45154 43764 45164
rect 44044 45220 44100 45838
rect 44156 45332 44212 45342
rect 44156 45238 44212 45276
rect 44380 45330 44436 46396
rect 44828 45890 44884 46396
rect 44828 45838 44830 45890
rect 44882 45838 44884 45890
rect 44828 45826 44884 45838
rect 45052 45892 45108 45902
rect 45052 45798 45108 45836
rect 44380 45278 44382 45330
rect 44434 45278 44436 45330
rect 44380 45266 44436 45278
rect 44940 45666 44996 45678
rect 44940 45614 44942 45666
rect 44994 45614 44996 45666
rect 44940 45332 44996 45614
rect 44940 45266 44996 45276
rect 45164 45332 45220 46620
rect 45276 45892 45332 46732
rect 45500 46674 45556 46686
rect 45500 46622 45502 46674
rect 45554 46622 45556 46674
rect 45276 45826 45332 45836
rect 45388 46340 45444 46350
rect 45500 46340 45556 46622
rect 45444 46284 45556 46340
rect 45388 45892 45444 46284
rect 45836 46116 45892 47292
rect 45948 47282 46004 47292
rect 46060 47348 46116 47358
rect 46060 47346 46228 47348
rect 46060 47294 46062 47346
rect 46114 47294 46228 47346
rect 46060 47292 46228 47294
rect 46060 47282 46116 47292
rect 45948 47124 46004 47134
rect 45948 46898 46004 47068
rect 45948 46846 45950 46898
rect 46002 46846 46004 46898
rect 45948 46834 46004 46846
rect 46172 46788 46228 47292
rect 46284 47234 46340 49196
rect 46508 48916 46564 48926
rect 46508 48822 46564 48860
rect 46396 48802 46452 48814
rect 46396 48750 46398 48802
rect 46450 48750 46452 48802
rect 46396 48580 46452 48750
rect 46620 48804 46676 48814
rect 46620 48710 46676 48748
rect 46396 48514 46452 48524
rect 46284 47182 46286 47234
rect 46338 47182 46340 47234
rect 46284 47170 46340 47182
rect 46396 48356 46452 48366
rect 46396 47458 46452 48300
rect 46396 47406 46398 47458
rect 46450 47406 46452 47458
rect 46396 47124 46452 47406
rect 46620 47460 46676 47470
rect 46620 47366 46676 47404
rect 46844 47236 46900 58044
rect 46956 57650 47012 58380
rect 46956 57598 46958 57650
rect 47010 57598 47012 57650
rect 46956 57586 47012 57598
rect 47068 57428 47124 59388
rect 47180 58434 47236 60732
rect 47404 61348 47460 61358
rect 47404 60676 47460 61292
rect 47516 60786 47572 61516
rect 47516 60734 47518 60786
rect 47570 60734 47572 60786
rect 47516 60722 47572 60734
rect 47404 60582 47460 60620
rect 47292 60562 47348 60574
rect 47628 60564 47684 62132
rect 48076 61682 48132 62132
rect 48076 61630 48078 61682
rect 48130 61630 48132 61682
rect 48076 61618 48132 61630
rect 48748 61012 48804 62132
rect 47292 60510 47294 60562
rect 47346 60510 47348 60562
rect 47292 59444 47348 60510
rect 47516 60508 47684 60564
rect 48636 60956 48804 61012
rect 47516 60004 47572 60508
rect 48076 60452 48132 60462
rect 48076 60226 48132 60396
rect 48076 60174 48078 60226
rect 48130 60174 48132 60226
rect 48076 60162 48132 60174
rect 47516 59910 47572 59948
rect 47404 59892 47460 59902
rect 47404 59668 47460 59836
rect 47628 59890 47684 59902
rect 47628 59838 47630 59890
rect 47682 59838 47684 59890
rect 47628 59780 47684 59838
rect 47628 59724 48020 59780
rect 47404 59612 47908 59668
rect 47516 59444 47572 59454
rect 47292 59442 47572 59444
rect 47292 59390 47518 59442
rect 47570 59390 47572 59442
rect 47292 59388 47572 59390
rect 47292 59220 47348 59230
rect 47292 59126 47348 59164
rect 47180 58382 47182 58434
rect 47234 58382 47236 58434
rect 47180 58370 47236 58382
rect 47404 59106 47460 59118
rect 47404 59054 47406 59106
rect 47458 59054 47460 59106
rect 47292 58212 47348 58222
rect 47180 58156 47292 58212
rect 47180 57874 47236 58156
rect 47292 58146 47348 58156
rect 47404 58100 47460 59054
rect 47516 58324 47572 59388
rect 47740 59332 47796 59342
rect 47516 58258 47572 58268
rect 47628 59330 47796 59332
rect 47628 59278 47742 59330
rect 47794 59278 47796 59330
rect 47628 59276 47796 59278
rect 47628 58212 47684 59276
rect 47740 59266 47796 59276
rect 47852 59220 47908 59612
rect 47964 59332 48020 59724
rect 48636 59442 48692 60956
rect 48860 60898 48916 63420
rect 48860 60846 48862 60898
rect 48914 60846 48916 60898
rect 48860 60834 48916 60846
rect 48972 63028 49028 63038
rect 48860 60676 48916 60686
rect 48860 60582 48916 60620
rect 48748 60228 48804 60238
rect 48972 60228 49028 62972
rect 49084 61572 49140 63644
rect 50556 62748 50820 62758
rect 50612 62692 50660 62748
rect 50716 62692 50764 62748
rect 50556 62682 50820 62692
rect 50764 62244 50820 62254
rect 50764 62150 50820 62188
rect 50204 61682 50260 61694
rect 50204 61630 50206 61682
rect 50258 61630 50260 61682
rect 50204 61572 50260 61630
rect 49140 61516 49364 61572
rect 49084 61506 49140 61516
rect 49196 61348 49252 61358
rect 49084 61292 49196 61348
rect 49084 60786 49140 61292
rect 49196 61282 49252 61292
rect 49084 60734 49086 60786
rect 49138 60734 49140 60786
rect 49084 60722 49140 60734
rect 49196 60676 49252 60686
rect 48748 60226 49028 60228
rect 48748 60174 48750 60226
rect 48802 60174 49028 60226
rect 48748 60172 49028 60174
rect 49084 60452 49140 60462
rect 49084 60226 49140 60396
rect 49084 60174 49086 60226
rect 49138 60174 49140 60226
rect 48748 60162 48804 60172
rect 49084 60162 49140 60174
rect 49196 60226 49252 60620
rect 49196 60174 49198 60226
rect 49250 60174 49252 60226
rect 49196 60162 49252 60174
rect 48860 60004 48916 60014
rect 49308 60004 49364 61516
rect 49868 60788 49924 60798
rect 50204 60788 50260 61516
rect 50876 61572 50932 61582
rect 50876 61478 50932 61516
rect 49868 60786 50260 60788
rect 49868 60734 49870 60786
rect 49922 60734 50260 60786
rect 49868 60732 50260 60734
rect 50316 61348 50372 61358
rect 50540 61348 50596 61358
rect 50316 61010 50372 61292
rect 50316 60958 50318 61010
rect 50370 60958 50372 61010
rect 49868 60722 49924 60732
rect 50316 60004 50372 60958
rect 48860 60002 49364 60004
rect 48860 59950 48862 60002
rect 48914 59950 49364 60002
rect 48860 59948 49364 59950
rect 49980 59948 50372 60004
rect 50428 61346 50596 61348
rect 50428 61294 50542 61346
rect 50594 61294 50596 61346
rect 50428 61292 50596 61294
rect 48860 59938 48916 59948
rect 49756 59778 49812 59790
rect 49756 59726 49758 59778
rect 49810 59726 49812 59778
rect 48636 59390 48638 59442
rect 48690 59390 48692 59442
rect 48636 59378 48692 59390
rect 48860 59444 48916 59454
rect 49420 59444 49476 59454
rect 48860 59442 49700 59444
rect 48860 59390 48862 59442
rect 48914 59390 49422 59442
rect 49474 59390 49700 59442
rect 48860 59388 49700 59390
rect 48860 59378 48916 59388
rect 49420 59378 49476 59388
rect 47964 59266 48020 59276
rect 48748 59332 48804 59342
rect 47852 59154 47908 59164
rect 47628 58146 47684 58156
rect 47740 58324 47796 58334
rect 47404 58034 47460 58044
rect 47180 57822 47182 57874
rect 47234 57822 47236 57874
rect 47180 57810 47236 57822
rect 47292 57876 47348 57886
rect 47740 57876 47796 58268
rect 46956 57372 47124 57428
rect 46956 56306 47012 57372
rect 47180 57316 47236 57326
rect 47180 56532 47236 57260
rect 47292 56866 47348 57820
rect 47516 57820 47796 57876
rect 47964 58322 48020 58334
rect 47964 58270 47966 58322
rect 48018 58270 48020 58322
rect 47404 57652 47460 57662
rect 47516 57652 47572 57820
rect 47404 57650 47572 57652
rect 47404 57598 47406 57650
rect 47458 57598 47572 57650
rect 47404 57596 47572 57598
rect 47628 57650 47684 57662
rect 47852 57652 47908 57662
rect 47628 57598 47630 57650
rect 47682 57598 47684 57650
rect 47404 57586 47460 57596
rect 47516 57204 47572 57214
rect 47628 57204 47684 57598
rect 47572 57148 47684 57204
rect 47740 57650 47908 57652
rect 47740 57598 47854 57650
rect 47906 57598 47908 57650
rect 47740 57596 47908 57598
rect 47516 57138 47572 57148
rect 47740 56980 47796 57596
rect 47852 57586 47908 57596
rect 47964 57092 48020 58270
rect 48076 57762 48132 57774
rect 48076 57710 48078 57762
rect 48130 57710 48132 57762
rect 48076 57316 48132 57710
rect 48076 57250 48132 57260
rect 48188 57650 48244 57662
rect 48188 57598 48190 57650
rect 48242 57598 48244 57650
rect 48188 57540 48244 57598
rect 47292 56814 47294 56866
rect 47346 56814 47348 56866
rect 47292 56802 47348 56814
rect 47404 56924 47796 56980
rect 47852 57036 48020 57092
rect 47404 56754 47460 56924
rect 47852 56868 47908 57036
rect 47404 56702 47406 56754
rect 47458 56702 47460 56754
rect 47404 56690 47460 56702
rect 47628 56812 47908 56868
rect 47628 56754 47684 56812
rect 47628 56702 47630 56754
rect 47682 56702 47684 56754
rect 47628 56690 47684 56702
rect 47964 56698 48020 56710
rect 47964 56646 47966 56698
rect 48018 56646 48020 56698
rect 47964 56644 48020 56646
rect 47852 56588 48020 56644
rect 47180 56476 47460 56532
rect 46956 56254 46958 56306
rect 47010 56254 47012 56306
rect 46956 56084 47012 56254
rect 47292 56308 47348 56318
rect 47292 56214 47348 56252
rect 46956 56018 47012 56028
rect 47068 54404 47124 54414
rect 47068 54402 47236 54404
rect 47068 54350 47070 54402
rect 47122 54350 47236 54402
rect 47068 54348 47236 54350
rect 47068 54338 47124 54348
rect 47068 53730 47124 53742
rect 47068 53678 47070 53730
rect 47122 53678 47124 53730
rect 46956 53172 47012 53182
rect 46956 52276 47012 53116
rect 46956 51378 47012 52220
rect 47068 51604 47124 53678
rect 47180 53284 47236 54348
rect 47404 53284 47460 56476
rect 47852 56196 47908 56588
rect 47852 56102 47908 56140
rect 48076 56194 48132 56206
rect 48076 56142 48078 56194
rect 48130 56142 48132 56194
rect 47628 56084 47684 56094
rect 47628 55990 47684 56028
rect 48076 56084 48132 56142
rect 48076 56018 48132 56028
rect 47740 55858 47796 55870
rect 48188 55860 48244 57484
rect 48748 56980 48804 59276
rect 48972 59220 49028 59230
rect 48972 59126 49028 59164
rect 48860 57540 48916 57550
rect 48860 57446 48916 57484
rect 49308 57540 49364 57550
rect 49308 57446 49364 57484
rect 49420 57092 49476 57102
rect 48748 56978 49140 56980
rect 48748 56926 48750 56978
rect 48802 56926 49140 56978
rect 48748 56924 49140 56926
rect 48748 56914 48804 56924
rect 47740 55806 47742 55858
rect 47794 55806 47796 55858
rect 47628 54514 47684 54526
rect 47628 54462 47630 54514
rect 47682 54462 47684 54514
rect 47628 53956 47684 54462
rect 47628 53890 47684 53900
rect 47740 53730 47796 55806
rect 47852 55804 48244 55860
rect 48300 56754 48356 56766
rect 48300 56702 48302 56754
rect 48354 56702 48356 56754
rect 47852 54516 47908 55804
rect 48076 55410 48132 55422
rect 48076 55358 48078 55410
rect 48130 55358 48132 55410
rect 48076 55076 48132 55358
rect 48300 55076 48356 56702
rect 48636 56308 48692 56318
rect 48692 56252 48804 56308
rect 48636 56242 48692 56252
rect 48636 55410 48692 55422
rect 48636 55358 48638 55410
rect 48690 55358 48692 55410
rect 48524 55186 48580 55198
rect 48524 55134 48526 55186
rect 48578 55134 48580 55186
rect 48524 55076 48580 55134
rect 48076 55020 48580 55076
rect 47964 54740 48020 54750
rect 48636 54740 48692 55358
rect 48748 55298 48804 56252
rect 48972 56196 49028 56206
rect 48972 56102 49028 56140
rect 49084 56194 49140 56924
rect 49084 56142 49086 56194
rect 49138 56142 49140 56194
rect 49084 56130 49140 56142
rect 48748 55246 48750 55298
rect 48802 55246 48804 55298
rect 48748 55234 48804 55246
rect 48860 56084 48916 56094
rect 47964 54646 48020 54684
rect 48188 54684 48692 54740
rect 48188 54626 48244 54684
rect 48188 54574 48190 54626
rect 48242 54574 48244 54626
rect 48188 54562 48244 54574
rect 48524 54516 48580 54526
rect 47852 54460 48020 54516
rect 47852 53844 47908 53854
rect 47852 53750 47908 53788
rect 47740 53678 47742 53730
rect 47794 53678 47796 53730
rect 47740 53666 47796 53678
rect 47964 53620 48020 54460
rect 48412 54460 48524 54516
rect 47852 53564 48020 53620
rect 48076 54402 48132 54414
rect 48076 54350 48078 54402
rect 48130 54350 48132 54402
rect 47516 53508 47572 53518
rect 47572 53452 47684 53508
rect 47516 53442 47572 53452
rect 47404 53228 47572 53284
rect 47180 53218 47236 53228
rect 47180 52948 47236 52958
rect 47180 52854 47236 52892
rect 47292 52836 47348 52846
rect 47292 52742 47348 52780
rect 47068 51538 47124 51548
rect 47516 51490 47572 53228
rect 47516 51438 47518 51490
rect 47570 51438 47572 51490
rect 46956 51326 46958 51378
rect 47010 51326 47012 51378
rect 46956 51314 47012 51326
rect 47068 51380 47124 51390
rect 47068 50708 47124 51324
rect 47404 51380 47460 51390
rect 47404 51286 47460 51324
rect 47516 50708 47572 51438
rect 47628 51380 47684 53452
rect 47852 52836 47908 53564
rect 48076 53508 48132 54350
rect 47964 53452 48132 53508
rect 47964 53058 48020 53452
rect 48300 53172 48356 53182
rect 48412 53172 48468 54460
rect 48524 54450 48580 54460
rect 48300 53170 48468 53172
rect 48300 53118 48302 53170
rect 48354 53118 48468 53170
rect 48300 53116 48468 53118
rect 48524 53956 48580 53966
rect 48524 53730 48580 53900
rect 48636 53844 48692 54684
rect 48636 53750 48692 53788
rect 48748 54404 48804 54414
rect 48524 53678 48526 53730
rect 48578 53678 48580 53730
rect 48300 53106 48356 53116
rect 47964 53006 47966 53058
rect 48018 53006 48020 53058
rect 47964 52994 48020 53006
rect 48076 53060 48132 53070
rect 48076 52966 48132 53004
rect 47852 52780 48244 52836
rect 47740 51604 47796 51614
rect 48076 51604 48132 51614
rect 47740 51602 48132 51604
rect 47740 51550 47742 51602
rect 47794 51550 48078 51602
rect 48130 51550 48132 51602
rect 47740 51548 48132 51550
rect 47740 51538 47796 51548
rect 48076 51538 48132 51548
rect 47964 51380 48020 51390
rect 47628 51378 48020 51380
rect 47628 51326 47966 51378
rect 48018 51326 48020 51378
rect 47628 51324 48020 51326
rect 47964 51314 48020 51324
rect 48076 51156 48132 51166
rect 48076 51062 48132 51100
rect 47068 50706 47348 50708
rect 47068 50654 47070 50706
rect 47122 50654 47348 50706
rect 47068 50652 47348 50654
rect 47068 50642 47124 50652
rect 47180 50372 47236 50382
rect 47180 49026 47236 50316
rect 47180 48974 47182 49026
rect 47234 48974 47236 49026
rect 47180 48962 47236 48974
rect 47180 47460 47236 47470
rect 46284 46900 46340 46910
rect 46284 46788 46340 46844
rect 46172 46786 46340 46788
rect 46172 46734 46174 46786
rect 46226 46734 46340 46786
rect 46172 46732 46340 46734
rect 46172 46722 46228 46732
rect 46060 46676 46116 46686
rect 46396 46676 46452 47068
rect 46620 47180 46900 47236
rect 46956 47346 47012 47358
rect 46956 47294 46958 47346
rect 47010 47294 47012 47346
rect 46956 47236 47012 47294
rect 47180 47346 47236 47404
rect 47180 47294 47182 47346
rect 47234 47294 47236 47346
rect 47180 47282 47236 47294
rect 46508 46676 46564 46686
rect 46396 46674 46564 46676
rect 46396 46622 46510 46674
rect 46562 46622 46564 46674
rect 46396 46620 46564 46622
rect 46060 46582 46116 46620
rect 46508 46610 46564 46620
rect 45836 46060 46004 46116
rect 45836 45892 45892 45902
rect 45388 45890 45892 45892
rect 45388 45838 45390 45890
rect 45442 45838 45838 45890
rect 45890 45838 45892 45890
rect 45388 45836 45892 45838
rect 45388 45556 45444 45836
rect 45836 45826 45892 45836
rect 45948 45556 46004 46060
rect 46396 46002 46452 46014
rect 46396 45950 46398 46002
rect 46450 45950 46452 46002
rect 46396 45892 46452 45950
rect 46396 45826 46452 45836
rect 45164 45266 45220 45276
rect 45276 45500 45444 45556
rect 45836 45500 46452 45556
rect 44044 45154 44100 45164
rect 44828 45108 44884 45118
rect 45052 45108 45108 45118
rect 44828 45014 44884 45052
rect 44940 45106 45108 45108
rect 44940 45054 45054 45106
rect 45106 45054 45108 45106
rect 44940 45052 45108 45054
rect 45276 45108 45332 45500
rect 45388 45332 45444 45342
rect 45836 45332 45892 45500
rect 45388 45330 45892 45332
rect 45388 45278 45390 45330
rect 45442 45278 45838 45330
rect 45890 45278 45892 45330
rect 45388 45276 45892 45278
rect 45388 45266 45444 45276
rect 45836 45266 45892 45276
rect 45948 45332 46004 45342
rect 45612 45108 45668 45118
rect 45276 45052 45556 45108
rect 43372 44930 43428 44940
rect 43820 44996 43876 45006
rect 43820 44902 43876 44940
rect 44268 44994 44324 45006
rect 44268 44942 44270 44994
rect 44322 44942 44324 44994
rect 42924 44382 42926 44434
rect 42978 44382 42980 44434
rect 42252 43652 42532 43708
rect 42140 43598 42142 43650
rect 42194 43598 42196 43650
rect 42140 43586 42196 43598
rect 41580 43540 41636 43550
rect 41916 43540 41972 43550
rect 41580 43538 41972 43540
rect 41580 43486 41582 43538
rect 41634 43486 41918 43538
rect 41970 43486 41972 43538
rect 41580 43484 41972 43486
rect 41580 43204 41636 43484
rect 41916 43474 41972 43484
rect 42364 43428 42420 43438
rect 41580 43138 41636 43148
rect 42028 43426 42420 43428
rect 42028 43374 42366 43426
rect 42418 43374 42420 43426
rect 42028 43372 42420 43374
rect 41580 42756 41636 42766
rect 41468 42754 41636 42756
rect 41468 42702 41582 42754
rect 41634 42702 41636 42754
rect 41468 42700 41636 42702
rect 41356 42662 41412 42700
rect 41580 42690 41636 42700
rect 41916 42644 41972 42654
rect 41916 42550 41972 42588
rect 41804 42530 41860 42542
rect 41804 42478 41806 42530
rect 41858 42478 41860 42530
rect 40012 39730 40068 39742
rect 40012 39678 40014 39730
rect 40066 39678 40068 39730
rect 40012 38948 40068 39678
rect 40684 39618 40740 39630
rect 40684 39566 40686 39618
rect 40738 39566 40740 39618
rect 40684 39284 40740 39566
rect 40908 39506 40964 40348
rect 40908 39454 40910 39506
rect 40962 39454 40964 39506
rect 40908 39396 40964 39454
rect 40908 39330 40964 39340
rect 41020 41580 41188 41636
rect 41244 41970 41300 41982
rect 41244 41918 41246 41970
rect 41298 41918 41300 41970
rect 40684 39218 40740 39228
rect 40012 38882 40068 38892
rect 40908 39060 40964 39070
rect 41020 39060 41076 41580
rect 41132 41412 41188 41422
rect 41132 41188 41188 41356
rect 41244 41300 41300 41918
rect 41468 41972 41524 41982
rect 41468 41878 41524 41916
rect 41580 41970 41636 41982
rect 41580 41918 41582 41970
rect 41634 41918 41636 41970
rect 41356 41858 41412 41870
rect 41356 41806 41358 41858
rect 41410 41806 41412 41858
rect 41356 41524 41412 41806
rect 41580 41860 41636 41918
rect 41580 41794 41636 41804
rect 41804 41636 41860 42478
rect 41804 41580 41972 41636
rect 41356 41468 41860 41524
rect 41244 41244 41412 41300
rect 41132 41186 41300 41188
rect 41132 41134 41134 41186
rect 41186 41134 41300 41186
rect 41132 41132 41300 41134
rect 41132 41122 41188 41132
rect 41244 40402 41300 41132
rect 41244 40350 41246 40402
rect 41298 40350 41300 40402
rect 41244 40338 41300 40350
rect 41356 39620 41412 41244
rect 41804 41298 41860 41468
rect 41804 41246 41806 41298
rect 41858 41246 41860 41298
rect 41804 41234 41860 41246
rect 41580 40404 41636 40414
rect 41244 39564 41412 39620
rect 41468 39732 41524 39742
rect 41468 39618 41524 39676
rect 41580 39730 41636 40348
rect 41580 39678 41582 39730
rect 41634 39678 41636 39730
rect 41580 39666 41636 39678
rect 41468 39566 41470 39618
rect 41522 39566 41524 39618
rect 41244 39172 41300 39564
rect 41468 39554 41524 39566
rect 41916 39618 41972 41580
rect 42028 40628 42084 43372
rect 42364 43362 42420 43372
rect 42476 42868 42532 43652
rect 42588 43538 42644 43550
rect 42588 43486 42590 43538
rect 42642 43486 42644 43538
rect 42588 43204 42644 43486
rect 42924 43540 42980 44382
rect 43372 44546 43428 44558
rect 43372 44494 43374 44546
rect 43426 44494 43428 44546
rect 43372 44098 43428 44494
rect 43372 44046 43374 44098
rect 43426 44046 43428 44098
rect 42924 43474 42980 43484
rect 43036 43538 43092 43550
rect 43036 43486 43038 43538
rect 43090 43486 43092 43538
rect 42588 43138 42644 43148
rect 42140 42812 42532 42868
rect 42140 42196 42196 42812
rect 42476 42754 42532 42812
rect 42476 42702 42478 42754
rect 42530 42702 42532 42754
rect 42476 42690 42532 42702
rect 42700 43092 42756 43102
rect 42700 42754 42756 43036
rect 42700 42702 42702 42754
rect 42754 42702 42756 42754
rect 42700 42690 42756 42702
rect 42252 42642 42308 42654
rect 42252 42590 42254 42642
rect 42306 42590 42308 42642
rect 42252 42532 42308 42590
rect 42252 42466 42308 42476
rect 42364 42530 42420 42542
rect 42364 42478 42366 42530
rect 42418 42478 42420 42530
rect 42252 42196 42308 42206
rect 42140 42194 42308 42196
rect 42140 42142 42254 42194
rect 42306 42142 42308 42194
rect 42140 42140 42308 42142
rect 42252 42130 42308 42140
rect 42028 40572 42196 40628
rect 42028 40404 42084 40414
rect 42028 40310 42084 40348
rect 41916 39566 41918 39618
rect 41970 39566 41972 39618
rect 41916 39554 41972 39566
rect 41356 39396 41412 39406
rect 41356 39302 41412 39340
rect 41692 39394 41748 39406
rect 41692 39342 41694 39394
rect 41746 39342 41748 39394
rect 41244 39116 41636 39172
rect 41020 39004 41412 39060
rect 40908 38836 40964 39004
rect 41020 38836 41076 38846
rect 38780 36372 38836 36382
rect 38836 36316 38948 36372
rect 38780 36306 38836 36316
rect 38780 35810 38836 35822
rect 38780 35758 38782 35810
rect 38834 35758 38836 35810
rect 38780 35028 38836 35758
rect 38780 34962 38836 34972
rect 38444 34914 38612 34916
rect 38444 34862 38446 34914
rect 38498 34862 38612 34914
rect 38444 34860 38612 34862
rect 38444 34850 38500 34860
rect 38780 34802 38836 34814
rect 38780 34750 38782 34802
rect 38834 34750 38836 34802
rect 38220 34692 38276 34702
rect 38668 34692 38724 34702
rect 38220 34598 38276 34636
rect 38332 34690 38724 34692
rect 38332 34638 38670 34690
rect 38722 34638 38724 34690
rect 38332 34636 38724 34638
rect 38332 34020 38388 34636
rect 38668 34626 38724 34636
rect 38780 34692 38836 34750
rect 38780 34626 38836 34636
rect 38780 34356 38836 34366
rect 38892 34356 38948 36316
rect 39452 35810 39508 38668
rect 39676 38612 39956 38668
rect 40348 38834 41076 38836
rect 40348 38782 41022 38834
rect 41074 38782 41076 38834
rect 40348 38780 41076 38782
rect 39676 36260 39732 38612
rect 40348 38162 40404 38780
rect 41020 38770 41076 38780
rect 41132 38836 41188 38846
rect 41132 38668 41188 38780
rect 41356 38668 41412 39004
rect 40908 38612 41188 38668
rect 41244 38612 41412 38668
rect 40908 38610 40964 38612
rect 40908 38558 40910 38610
rect 40962 38558 40964 38610
rect 40908 38546 40964 38558
rect 40348 38110 40350 38162
rect 40402 38110 40404 38162
rect 40348 38098 40404 38110
rect 40348 37154 40404 37166
rect 40348 37102 40350 37154
rect 40402 37102 40404 37154
rect 40348 36932 40404 37102
rect 40348 36866 40404 36876
rect 41132 37154 41188 37166
rect 41132 37102 41134 37154
rect 41186 37102 41188 37154
rect 41132 36932 41188 37102
rect 39452 35758 39454 35810
rect 39506 35758 39508 35810
rect 39452 35746 39508 35758
rect 39564 36204 39732 36260
rect 38780 34354 38948 34356
rect 38780 34302 38782 34354
rect 38834 34302 38948 34354
rect 38780 34300 38948 34302
rect 39340 34692 39396 34702
rect 38780 34290 38836 34300
rect 39340 34244 39396 34636
rect 39564 34356 39620 36204
rect 41020 36036 41076 36046
rect 41132 36036 41188 36876
rect 41076 35980 41188 36036
rect 39788 35924 39844 35934
rect 39788 35830 39844 35868
rect 40124 35924 40180 35934
rect 39676 35700 39732 35710
rect 39900 35700 39956 35710
rect 39676 35698 39844 35700
rect 39676 35646 39678 35698
rect 39730 35646 39844 35698
rect 39676 35644 39844 35646
rect 39676 35634 39732 35644
rect 39676 34804 39732 34814
rect 39676 34710 39732 34748
rect 39676 34356 39732 34366
rect 39564 34354 39732 34356
rect 39564 34302 39678 34354
rect 39730 34302 39732 34354
rect 39564 34300 39732 34302
rect 39676 34290 39732 34300
rect 39788 34354 39844 35644
rect 39900 35606 39956 35644
rect 40124 35698 40180 35868
rect 41020 35810 41076 35980
rect 41244 35924 41300 38612
rect 41468 37828 41524 37838
rect 41468 37492 41524 37772
rect 41468 37398 41524 37436
rect 41020 35758 41022 35810
rect 41074 35758 41076 35810
rect 41020 35746 41076 35758
rect 41132 35868 41300 35924
rect 41356 37268 41412 37278
rect 40124 35646 40126 35698
rect 40178 35646 40180 35698
rect 40124 35634 40180 35646
rect 40908 35700 40964 35710
rect 40908 35606 40964 35644
rect 41132 35588 41188 35868
rect 41356 35698 41412 37212
rect 41580 36484 41636 39116
rect 41692 37044 41748 39342
rect 42028 38724 42084 38734
rect 41916 37268 41972 37278
rect 41916 37174 41972 37212
rect 41692 36978 41748 36988
rect 41356 35646 41358 35698
rect 41410 35646 41412 35698
rect 41356 35634 41412 35646
rect 41468 36428 41636 36484
rect 42028 36484 42084 38668
rect 42140 36708 42196 40572
rect 42252 38052 42308 38062
rect 42364 38052 42420 42478
rect 42924 41972 42980 41982
rect 42924 39842 42980 41916
rect 43036 41412 43092 43486
rect 43036 40404 43092 41356
rect 43372 41188 43428 44046
rect 44268 43708 44324 44942
rect 44940 44324 44996 45052
rect 45052 45042 45108 45052
rect 45500 44434 45556 45052
rect 45612 45014 45668 45052
rect 45948 45106 46004 45276
rect 46396 45330 46452 45500
rect 46396 45278 46398 45330
rect 46450 45278 46452 45330
rect 46396 45266 46452 45278
rect 45948 45054 45950 45106
rect 46002 45054 46004 45106
rect 45500 44382 45502 44434
rect 45554 44382 45556 44434
rect 45500 44370 45556 44382
rect 44940 44230 44996 44268
rect 43820 43652 44324 43708
rect 43820 43650 43876 43652
rect 43820 43598 43822 43650
rect 43874 43598 43876 43650
rect 43820 43586 43876 43598
rect 45948 43426 46004 45054
rect 45948 43374 45950 43426
rect 46002 43374 46004 43426
rect 45612 43204 45668 43214
rect 45052 42980 45108 42990
rect 44828 42644 44884 42654
rect 44828 42550 44884 42588
rect 43372 41122 43428 41132
rect 43932 41298 43988 41310
rect 43932 41246 43934 41298
rect 43986 41246 43988 41298
rect 43036 40338 43092 40348
rect 42924 39790 42926 39842
rect 42978 39790 42980 39842
rect 42924 39778 42980 39790
rect 43484 40068 43540 40078
rect 43372 39732 43428 39742
rect 43372 39638 43428 39676
rect 43484 39730 43540 40012
rect 43484 39678 43486 39730
rect 43538 39678 43540 39730
rect 43484 39666 43540 39678
rect 43036 39620 43092 39630
rect 43036 39526 43092 39564
rect 43932 39620 43988 41246
rect 45052 40740 45108 42924
rect 45388 42754 45444 42766
rect 45388 42702 45390 42754
rect 45442 42702 45444 42754
rect 45388 42644 45444 42702
rect 45388 42578 45444 42588
rect 45164 42532 45220 42542
rect 45164 42438 45220 42476
rect 45612 42196 45668 43148
rect 45836 42756 45892 42766
rect 45948 42756 46004 43374
rect 45836 42754 46004 42756
rect 45836 42702 45838 42754
rect 45890 42702 46004 42754
rect 45836 42700 46004 42702
rect 46060 43764 46116 43774
rect 46060 42756 46116 43708
rect 46396 43428 46452 43438
rect 46620 43428 46676 47180
rect 46956 47170 47012 47180
rect 47068 47234 47124 47246
rect 47068 47182 47070 47234
rect 47122 47182 47124 47234
rect 47068 47068 47124 47182
rect 46732 47012 47124 47068
rect 46732 46900 46788 47012
rect 46732 46674 46788 46844
rect 47068 46788 47124 46798
rect 47068 46694 47124 46732
rect 46732 46622 46734 46674
rect 46786 46622 46788 46674
rect 46732 46610 46788 46622
rect 46844 44324 46900 44334
rect 46844 43764 46900 44268
rect 47292 43708 47348 50652
rect 47516 50642 47572 50652
rect 48188 50428 48244 52780
rect 47628 50372 48244 50428
rect 48524 50372 48580 53678
rect 48748 52948 48804 54348
rect 48860 53284 48916 56028
rect 49308 55298 49364 55310
rect 49308 55246 49310 55298
rect 49362 55246 49364 55298
rect 49308 54404 49364 55246
rect 49308 54338 49364 54348
rect 49420 54068 49476 57036
rect 49308 54012 49476 54068
rect 49532 55858 49588 55870
rect 49532 55806 49534 55858
rect 49586 55806 49588 55858
rect 49532 54740 49588 55806
rect 49084 53284 49140 53294
rect 48860 53228 49084 53284
rect 49084 53170 49140 53228
rect 49084 53118 49086 53170
rect 49138 53118 49140 53170
rect 49084 53106 49140 53118
rect 49308 53172 49364 54012
rect 49532 53954 49588 54684
rect 49532 53902 49534 53954
rect 49586 53902 49588 53954
rect 49532 53890 49588 53902
rect 49420 53844 49476 53854
rect 49420 53750 49476 53788
rect 49644 53620 49700 59388
rect 49756 59332 49812 59726
rect 49756 59266 49812 59276
rect 49868 59444 49924 59454
rect 49868 59220 49924 59388
rect 49868 59154 49924 59164
rect 49756 57538 49812 57550
rect 49756 57486 49758 57538
rect 49810 57486 49812 57538
rect 49756 57316 49812 57486
rect 49756 57250 49812 57260
rect 49980 56308 50036 59948
rect 50204 59780 50260 59790
rect 50428 59780 50484 61292
rect 50540 61282 50596 61292
rect 50556 61180 50820 61190
rect 50612 61124 50660 61180
rect 50716 61124 50764 61180
rect 50556 61114 50820 61124
rect 50204 59778 50484 59780
rect 50204 59726 50206 59778
rect 50258 59726 50484 59778
rect 50204 59724 50484 59726
rect 52108 59780 52164 59790
rect 50204 59714 50260 59724
rect 50316 59444 50372 59724
rect 50556 59612 50820 59622
rect 50612 59556 50660 59612
rect 50716 59556 50764 59612
rect 50556 59546 50820 59556
rect 50316 59106 50372 59388
rect 50316 59054 50318 59106
rect 50370 59054 50372 59106
rect 50092 58546 50148 58558
rect 50092 58494 50094 58546
rect 50146 58494 50148 58546
rect 50092 57540 50148 58494
rect 50092 57474 50148 57484
rect 49980 56242 50036 56252
rect 49868 55074 49924 55086
rect 49868 55022 49870 55074
rect 49922 55022 49924 55074
rect 49868 54516 49924 55022
rect 49980 55076 50036 55086
rect 49980 54982 50036 55020
rect 50092 55074 50148 55086
rect 50092 55022 50094 55074
rect 50146 55022 50148 55074
rect 49868 54450 49924 54460
rect 50092 54292 50148 55022
rect 49868 54236 50148 54292
rect 49756 53956 49812 53966
rect 49756 53862 49812 53900
rect 49868 53954 49924 54236
rect 50316 54180 50372 59054
rect 50556 58044 50820 58054
rect 50612 57988 50660 58044
rect 50716 57988 50764 58044
rect 50556 57978 50820 57988
rect 50556 56476 50820 56486
rect 50612 56420 50660 56476
rect 50716 56420 50764 56476
rect 50556 56410 50820 56420
rect 49868 53902 49870 53954
rect 49922 53902 49924 53954
rect 49868 53890 49924 53902
rect 49980 54124 50372 54180
rect 50428 55298 50484 55310
rect 50428 55246 50430 55298
rect 50482 55246 50484 55298
rect 49980 53732 50036 54124
rect 49308 53116 49476 53172
rect 49308 52948 49364 52958
rect 48748 52946 49364 52948
rect 48748 52894 49310 52946
rect 49362 52894 49364 52946
rect 48748 52892 49364 52894
rect 49308 52882 49364 52892
rect 49084 52724 49140 52734
rect 49420 52724 49476 53116
rect 48636 52276 48692 52286
rect 48692 52220 48804 52276
rect 48636 52210 48692 52220
rect 48748 51490 48804 52220
rect 48860 51604 48916 51614
rect 48860 51510 48916 51548
rect 48748 51438 48750 51490
rect 48802 51438 48804 51490
rect 48748 51426 48804 51438
rect 48972 51492 49028 51502
rect 48972 51378 49028 51436
rect 48972 51326 48974 51378
rect 49026 51326 49028 51378
rect 48972 51314 49028 51326
rect 47628 49588 47684 50372
rect 48524 50316 48804 50372
rect 47628 49532 48132 49588
rect 47852 48916 47908 48926
rect 47852 48822 47908 48860
rect 47740 47460 47796 47470
rect 47628 47346 47684 47358
rect 47628 47294 47630 47346
rect 47682 47294 47684 47346
rect 47628 47068 47684 47294
rect 47740 47346 47796 47404
rect 47740 47294 47742 47346
rect 47794 47294 47796 47346
rect 47740 47282 47796 47294
rect 47964 47234 48020 47246
rect 47964 47182 47966 47234
rect 48018 47182 48020 47234
rect 47628 47012 47796 47068
rect 47628 46788 47684 46798
rect 47628 46694 47684 46732
rect 47404 46676 47460 46686
rect 47404 46582 47460 46620
rect 47516 46564 47572 46574
rect 47516 46470 47572 46508
rect 47628 46340 47684 46350
rect 47740 46340 47796 47012
rect 47964 46674 48020 47182
rect 47964 46622 47966 46674
rect 48018 46622 48020 46674
rect 47964 46610 48020 46622
rect 47684 46284 47796 46340
rect 47628 46274 47684 46284
rect 47964 45892 48020 45902
rect 46844 43538 46900 43708
rect 46844 43486 46846 43538
rect 46898 43486 46900 43538
rect 46844 43474 46900 43486
rect 47068 43652 47348 43708
rect 47516 44212 47572 44222
rect 47068 43538 47124 43652
rect 47068 43486 47070 43538
rect 47122 43486 47124 43538
rect 47068 43474 47124 43486
rect 47404 43540 47460 43550
rect 47516 43540 47572 44156
rect 47964 43650 48020 45836
rect 47964 43598 47966 43650
rect 48018 43598 48020 43650
rect 47964 43586 48020 43598
rect 48076 43708 48132 49532
rect 48748 48804 48804 50316
rect 48748 48738 48804 48748
rect 48188 48132 48244 48142
rect 48188 45780 48244 48076
rect 48300 47572 48356 47582
rect 48300 47478 48356 47516
rect 48748 47572 48804 47582
rect 48748 47478 48804 47516
rect 48300 46564 48356 46574
rect 48356 46508 48580 46564
rect 48300 46498 48356 46508
rect 48524 46002 48580 46508
rect 48524 45950 48526 46002
rect 48578 45950 48580 46002
rect 48524 45938 48580 45950
rect 48188 45724 48580 45780
rect 48412 44324 48468 44334
rect 48412 44230 48468 44268
rect 48524 44322 48580 45724
rect 49084 45668 49140 52668
rect 49308 52668 49476 52724
rect 49308 51604 49364 52668
rect 49308 51490 49364 51548
rect 49308 51438 49310 51490
rect 49362 51438 49364 51490
rect 49308 51426 49364 51438
rect 49420 52164 49476 52174
rect 49196 51156 49252 51166
rect 49196 50706 49252 51100
rect 49196 50654 49198 50706
rect 49250 50654 49252 50706
rect 49196 50642 49252 50654
rect 49308 50372 49364 50382
rect 49308 50036 49364 50316
rect 49196 49980 49364 50036
rect 49196 45890 49252 49980
rect 49308 49812 49364 49822
rect 49420 49812 49476 52108
rect 49644 50036 49700 53564
rect 49868 53676 50036 53732
rect 50428 53732 50484 55246
rect 50876 55076 50932 55086
rect 50556 54908 50820 54918
rect 50612 54852 50660 54908
rect 50716 54852 50764 54908
rect 50556 54842 50820 54852
rect 50876 54626 50932 55020
rect 50876 54574 50878 54626
rect 50930 54574 50932 54626
rect 50876 54562 50932 54574
rect 51660 54514 51716 54526
rect 51660 54462 51662 54514
rect 51714 54462 51716 54514
rect 50540 53732 50596 53742
rect 50428 53730 50596 53732
rect 50428 53678 50542 53730
rect 50594 53678 50596 53730
rect 50428 53676 50596 53678
rect 49756 51604 49812 51614
rect 49756 51510 49812 51548
rect 49644 49980 49812 50036
rect 49644 49812 49700 49822
rect 49308 49810 49700 49812
rect 49308 49758 49310 49810
rect 49362 49758 49646 49810
rect 49698 49758 49700 49810
rect 49308 49756 49700 49758
rect 49308 49746 49364 49756
rect 49644 49746 49700 49756
rect 49756 47572 49812 49980
rect 49756 47506 49812 47516
rect 49196 45838 49198 45890
rect 49250 45838 49252 45890
rect 49196 45826 49252 45838
rect 49084 45612 49252 45668
rect 48524 44270 48526 44322
rect 48578 44270 48580 44322
rect 48524 44258 48580 44270
rect 49084 44322 49140 44334
rect 49084 44270 49086 44322
rect 49138 44270 49140 44322
rect 48860 44212 48916 44222
rect 49084 44212 49140 44270
rect 49196 44324 49252 45612
rect 49420 44324 49476 44334
rect 49196 44322 49476 44324
rect 49196 44270 49422 44322
rect 49474 44270 49476 44322
rect 49196 44268 49476 44270
rect 49420 44258 49476 44268
rect 49644 44324 49700 44334
rect 49644 44230 49700 44268
rect 48916 44156 49140 44212
rect 48860 44118 48916 44156
rect 48748 44098 48804 44110
rect 48748 44046 48750 44098
rect 48802 44046 48804 44098
rect 48748 43708 48804 44046
rect 49308 44098 49364 44110
rect 49308 44046 49310 44098
rect 49362 44046 49364 44098
rect 49308 43708 49364 44046
rect 48076 43652 48468 43708
rect 48748 43652 49140 43708
rect 49308 43652 49700 43708
rect 47404 43538 47572 43540
rect 47404 43486 47406 43538
rect 47458 43486 47518 43538
rect 47570 43486 47572 43538
rect 47404 43484 47572 43486
rect 47404 43474 47460 43484
rect 46396 43426 46676 43428
rect 46396 43374 46398 43426
rect 46450 43374 46676 43426
rect 46396 43372 46676 43374
rect 46396 43362 46452 43372
rect 46284 43204 46340 43214
rect 46340 43148 46452 43204
rect 46284 43138 46340 43148
rect 46060 42754 46340 42756
rect 46060 42702 46062 42754
rect 46114 42702 46340 42754
rect 46060 42700 46340 42702
rect 45836 42690 45892 42700
rect 46060 42690 46116 42700
rect 45724 42532 45780 42542
rect 46172 42532 46228 42542
rect 45724 42530 46004 42532
rect 45724 42478 45726 42530
rect 45778 42478 46004 42530
rect 45724 42476 46004 42478
rect 45724 42466 45780 42476
rect 45836 42196 45892 42206
rect 45612 42194 45892 42196
rect 45612 42142 45838 42194
rect 45890 42142 45892 42194
rect 45612 42140 45892 42142
rect 45836 42130 45892 42140
rect 45164 41188 45220 41198
rect 45164 41094 45220 41132
rect 45052 40674 45108 40684
rect 45276 40628 45332 40638
rect 44940 40404 44996 40414
rect 44940 40310 44996 40348
rect 44156 40290 44212 40302
rect 44156 40238 44158 40290
rect 44210 40238 44212 40290
rect 44156 40068 44212 40238
rect 44156 40002 44212 40012
rect 43932 39554 43988 39564
rect 45164 39508 45220 39518
rect 43260 38724 43316 38734
rect 43260 38162 43316 38668
rect 43260 38110 43262 38162
rect 43314 38110 43316 38162
rect 43260 38098 43316 38110
rect 42252 38050 42420 38052
rect 42252 37998 42254 38050
rect 42306 37998 42420 38050
rect 42252 37996 42420 37998
rect 45164 38052 45220 39452
rect 45276 39060 45332 40572
rect 45612 40292 45668 40302
rect 45612 40290 45892 40292
rect 45612 40238 45614 40290
rect 45666 40238 45892 40290
rect 45612 40236 45892 40238
rect 45612 40226 45668 40236
rect 45388 39618 45444 39630
rect 45388 39566 45390 39618
rect 45442 39566 45444 39618
rect 45388 39284 45444 39566
rect 45388 39218 45444 39228
rect 45612 39394 45668 39406
rect 45612 39342 45614 39394
rect 45666 39342 45668 39394
rect 45276 38994 45332 39004
rect 45612 39060 45668 39342
rect 45836 39396 45892 40236
rect 45948 39618 46004 42476
rect 46172 41970 46228 42476
rect 46284 42196 46340 42700
rect 46396 42754 46452 43148
rect 46396 42702 46398 42754
rect 46450 42702 46452 42754
rect 46396 42690 46452 42702
rect 46620 42754 46676 43372
rect 47180 43426 47236 43438
rect 47180 43374 47182 43426
rect 47234 43374 47236 43426
rect 46620 42702 46622 42754
rect 46674 42702 46676 42754
rect 46620 42690 46676 42702
rect 46956 42756 47012 42766
rect 46956 42662 47012 42700
rect 46620 42530 46676 42542
rect 47180 42532 47236 43374
rect 47292 43204 47348 43214
rect 47292 42754 47348 43148
rect 47292 42702 47294 42754
rect 47346 42702 47348 42754
rect 47292 42690 47348 42702
rect 46620 42478 46622 42530
rect 46674 42478 46676 42530
rect 46508 42196 46564 42206
rect 46284 42194 46564 42196
rect 46284 42142 46510 42194
rect 46562 42142 46564 42194
rect 46284 42140 46564 42142
rect 46508 42130 46564 42140
rect 46172 41918 46174 41970
rect 46226 41918 46228 41970
rect 46172 40180 46228 41918
rect 46172 40114 46228 40124
rect 46508 41972 46564 41982
rect 46284 39620 46340 39630
rect 45948 39566 45950 39618
rect 46002 39566 46004 39618
rect 45948 39554 46004 39566
rect 46060 39618 46340 39620
rect 46060 39566 46286 39618
rect 46338 39566 46340 39618
rect 46060 39564 46340 39566
rect 46508 39620 46564 41916
rect 46620 40404 46676 42478
rect 47068 42476 47236 42532
rect 47404 42530 47460 42542
rect 47404 42478 47406 42530
rect 47458 42478 47460 42530
rect 47068 42308 47124 42476
rect 47404 42420 47460 42478
rect 47068 42242 47124 42252
rect 47180 42364 47460 42420
rect 47180 42196 47236 42364
rect 47516 42308 47572 43484
rect 47740 43426 47796 43438
rect 47740 43374 47742 43426
rect 47794 43374 47796 43426
rect 47628 42868 47684 42878
rect 47628 42754 47684 42812
rect 47628 42702 47630 42754
rect 47682 42702 47684 42754
rect 47628 42690 47684 42702
rect 47180 42130 47236 42140
rect 47292 42252 47572 42308
rect 47628 42420 47684 42430
rect 46732 41972 46788 41982
rect 47180 41972 47236 41982
rect 46732 41970 47236 41972
rect 46732 41918 46734 41970
rect 46786 41918 47182 41970
rect 47234 41918 47236 41970
rect 46732 41916 47236 41918
rect 46732 41412 46788 41916
rect 47180 41906 47236 41916
rect 46732 41346 46788 41356
rect 46620 40348 47236 40404
rect 46956 40180 47012 40190
rect 46508 39564 46900 39620
rect 46060 39396 46116 39564
rect 46284 39554 46340 39564
rect 45836 39340 46116 39396
rect 46172 39394 46228 39406
rect 46172 39342 46174 39394
rect 46226 39342 46228 39394
rect 45612 38994 45668 39004
rect 46172 38668 46228 39342
rect 46396 39396 46452 39406
rect 46396 39302 46452 39340
rect 46508 39394 46564 39406
rect 46508 39342 46510 39394
rect 46562 39342 46564 39394
rect 46508 39060 46564 39342
rect 46620 39060 46676 39070
rect 46508 39004 46620 39060
rect 46620 38994 46676 39004
rect 42252 37986 42308 37996
rect 45164 37986 45220 37996
rect 46060 38612 46228 38668
rect 46844 38668 46900 39564
rect 46956 39618 47012 40124
rect 46956 39566 46958 39618
rect 47010 39566 47012 39618
rect 46956 39554 47012 39566
rect 46844 38612 47012 38668
rect 43820 37938 43876 37950
rect 43820 37886 43822 37938
rect 43874 37886 43876 37938
rect 42364 37826 42420 37838
rect 42364 37774 42366 37826
rect 42418 37774 42420 37826
rect 42364 36932 42420 37774
rect 42476 37826 42532 37838
rect 42476 37774 42478 37826
rect 42530 37774 42532 37826
rect 42476 37380 42532 37774
rect 42588 37828 42644 37838
rect 42588 37734 42644 37772
rect 42700 37826 42756 37838
rect 42700 37774 42702 37826
rect 42754 37774 42756 37826
rect 42588 37380 42644 37390
rect 42476 37378 42644 37380
rect 42476 37326 42590 37378
rect 42642 37326 42644 37378
rect 42476 37324 42644 37326
rect 42588 37314 42644 37324
rect 42364 36866 42420 36876
rect 42140 36652 42420 36708
rect 42252 36484 42308 36494
rect 42028 36482 42308 36484
rect 42028 36430 42254 36482
rect 42306 36430 42308 36482
rect 42028 36428 42308 36430
rect 41020 35532 41188 35588
rect 40460 34916 40516 34926
rect 40124 34804 40180 34814
rect 40460 34804 40516 34860
rect 40124 34690 40180 34748
rect 40124 34638 40126 34690
rect 40178 34638 40180 34690
rect 40124 34468 40180 34638
rect 40124 34402 40180 34412
rect 40236 34802 40516 34804
rect 40236 34750 40462 34802
rect 40514 34750 40516 34802
rect 40236 34748 40516 34750
rect 39788 34302 39790 34354
rect 39842 34302 39844 34354
rect 39788 34290 39844 34302
rect 39340 34150 39396 34188
rect 39452 34242 39508 34254
rect 39452 34190 39454 34242
rect 39506 34190 39508 34242
rect 38332 33926 38388 33964
rect 38108 33070 38110 33122
rect 38162 33070 38164 33122
rect 38108 32676 38164 33070
rect 38108 32610 38164 32620
rect 38444 33124 38500 33134
rect 37436 32510 37438 32562
rect 37490 32510 37492 32562
rect 37436 32498 37492 32510
rect 37100 32274 37156 32284
rect 37324 32452 37380 32462
rect 36988 32228 37044 32238
rect 36988 32002 37044 32172
rect 36988 31950 36990 32002
rect 37042 31950 37044 32002
rect 36988 31938 37044 31950
rect 37324 31890 37380 32396
rect 37324 31838 37326 31890
rect 37378 31838 37380 31890
rect 37324 31826 37380 31838
rect 38220 32450 38276 32462
rect 38220 32398 38222 32450
rect 38274 32398 38276 32450
rect 38220 31892 38276 32398
rect 38220 31826 38276 31836
rect 36540 31612 36708 31668
rect 37548 31780 37604 31790
rect 35420 31554 35476 31566
rect 35420 31502 35422 31554
rect 35474 31502 35476 31554
rect 35420 31108 35476 31502
rect 35532 31556 35588 31566
rect 35532 31462 35588 31500
rect 35756 31554 35812 31566
rect 35756 31502 35758 31554
rect 35810 31502 35812 31554
rect 35420 31042 35476 31052
rect 35756 30772 35812 31502
rect 36316 31556 36372 31566
rect 36316 31462 36372 31500
rect 36316 31108 36372 31118
rect 36092 31106 36372 31108
rect 36092 31054 36318 31106
rect 36370 31054 36372 31106
rect 36092 31052 36372 31054
rect 35756 30706 35812 30716
rect 35980 30884 36036 30894
rect 36092 30884 36148 31052
rect 36316 31042 36372 31052
rect 36428 31108 36484 31118
rect 36428 31014 36484 31052
rect 35980 30882 36148 30884
rect 35980 30830 35982 30882
rect 36034 30830 36148 30882
rect 35980 30828 36148 30830
rect 35196 30604 35460 30614
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35196 30538 35460 30548
rect 35756 30548 35812 30558
rect 35196 30324 35252 30334
rect 35084 30322 35252 30324
rect 35084 30270 35198 30322
rect 35250 30270 35252 30322
rect 35084 30268 35252 30270
rect 34972 29428 35028 29438
rect 34972 29334 35028 29372
rect 34972 28644 35028 28654
rect 34972 28550 35028 28588
rect 34972 28196 35028 28206
rect 34748 27346 34804 27356
rect 34860 28140 34972 28196
rect 34860 27076 34916 28140
rect 34972 28130 35028 28140
rect 34300 26198 34356 26236
rect 34524 26852 34692 26908
rect 34748 26964 34804 27002
rect 34860 26982 34916 27020
rect 34748 26852 34804 26908
rect 33740 26178 33796 26190
rect 33740 26126 33742 26178
rect 33794 26126 33796 26178
rect 33740 25506 33796 26126
rect 34524 25732 34580 26852
rect 34748 26796 34916 26852
rect 34748 26290 34804 26302
rect 34748 26238 34750 26290
rect 34802 26238 34804 26290
rect 34748 26180 34804 26238
rect 34748 26114 34804 26124
rect 34860 25956 34916 26796
rect 34188 25676 34580 25732
rect 34748 25900 34916 25956
rect 34972 26180 35028 26190
rect 33740 25454 33742 25506
rect 33794 25454 33796 25506
rect 33740 23828 33796 25454
rect 33964 25506 34020 25518
rect 33964 25454 33966 25506
rect 34018 25454 34020 25506
rect 33740 23762 33796 23772
rect 33852 25284 33908 25294
rect 33852 24834 33908 25228
rect 33964 25060 34020 25454
rect 33964 24994 34020 25004
rect 34076 24948 34132 24958
rect 33852 24782 33854 24834
rect 33906 24782 33908 24834
rect 33852 21588 33908 24782
rect 33964 24836 34020 24846
rect 33964 24742 34020 24780
rect 33964 21588 34020 21598
rect 33852 21586 34020 21588
rect 33852 21534 33966 21586
rect 34018 21534 34020 21586
rect 33852 21532 34020 21534
rect 33964 21522 34020 21532
rect 33628 20290 33684 20300
rect 33404 20132 33460 20142
rect 33964 20132 34020 20142
rect 34076 20132 34132 24892
rect 34188 24946 34244 25676
rect 34748 25060 34804 25900
rect 34748 24994 34804 25004
rect 34860 25506 34916 25518
rect 34860 25454 34862 25506
rect 34914 25454 34916 25506
rect 34188 24894 34190 24946
rect 34242 24894 34244 24946
rect 34188 24882 34244 24894
rect 34860 24836 34916 25454
rect 34636 24612 34692 24622
rect 34636 24518 34692 24556
rect 34636 24164 34692 24174
rect 34524 23716 34580 23726
rect 34412 21924 34468 21934
rect 34300 20692 34356 20702
rect 34300 20598 34356 20636
rect 34300 20244 34356 20254
rect 33404 20130 34076 20132
rect 33404 20078 33406 20130
rect 33458 20078 33966 20130
rect 34018 20078 34076 20130
rect 33404 20076 34076 20078
rect 33404 20066 33460 20076
rect 33964 20066 34020 20076
rect 34076 20038 34132 20076
rect 34188 20188 34300 20244
rect 34412 20244 34468 21868
rect 34524 21810 34580 23660
rect 34524 21758 34526 21810
rect 34578 21758 34580 21810
rect 34524 21746 34580 21758
rect 34636 23154 34692 24108
rect 34860 24050 34916 24780
rect 34860 23998 34862 24050
rect 34914 23998 34916 24050
rect 34860 23986 34916 23998
rect 34636 23102 34638 23154
rect 34690 23102 34692 23154
rect 34412 20188 34580 20244
rect 34188 20130 34244 20188
rect 34300 20178 34356 20188
rect 34188 20078 34190 20130
rect 34242 20078 34244 20130
rect 34188 20066 34244 20078
rect 34412 20018 34468 20030
rect 34412 19966 34414 20018
rect 34466 19966 34468 20018
rect 33516 19908 33572 19918
rect 33404 18338 33460 18350
rect 33404 18286 33406 18338
rect 33458 18286 33460 18338
rect 33404 18228 33460 18286
rect 33404 18162 33460 18172
rect 33516 17220 33572 19852
rect 34300 19906 34356 19918
rect 34300 19854 34302 19906
rect 34354 19854 34356 19906
rect 34300 19124 34356 19854
rect 33628 19068 34356 19124
rect 33628 18674 33684 19068
rect 34412 18900 34468 19966
rect 34412 18834 34468 18844
rect 34524 18788 34580 20188
rect 34524 18722 34580 18732
rect 33628 18622 33630 18674
rect 33682 18622 33684 18674
rect 33628 18610 33684 18622
rect 34076 18562 34132 18574
rect 34076 18510 34078 18562
rect 34130 18510 34132 18562
rect 33740 18452 33796 18462
rect 33740 18358 33796 18396
rect 33852 18450 33908 18462
rect 33852 18398 33854 18450
rect 33906 18398 33908 18450
rect 33852 18116 33908 18398
rect 33852 18050 33908 18060
rect 33964 18452 34020 18462
rect 33628 17780 33684 17790
rect 33628 17686 33684 17724
rect 33516 17154 33572 17164
rect 33964 17666 34020 18396
rect 34076 17890 34132 18510
rect 34524 18452 34580 18462
rect 34412 18450 34580 18452
rect 34412 18398 34526 18450
rect 34578 18398 34580 18450
rect 34412 18396 34580 18398
rect 34076 17838 34078 17890
rect 34130 17838 34132 17890
rect 34076 17826 34132 17838
rect 34188 18340 34244 18350
rect 33964 17614 33966 17666
rect 34018 17614 34020 17666
rect 33964 17106 34020 17614
rect 34076 17668 34132 17678
rect 34076 17554 34132 17612
rect 34076 17502 34078 17554
rect 34130 17502 34132 17554
rect 34076 17490 34132 17502
rect 33964 17054 33966 17106
rect 34018 17054 34020 17106
rect 33964 17042 34020 17054
rect 34188 17108 34244 18284
rect 34412 18116 34468 18396
rect 34524 18386 34580 18396
rect 34412 18050 34468 18060
rect 34524 18228 34580 18238
rect 34524 17556 34580 18172
rect 34524 17490 34580 17500
rect 34188 16772 34244 17052
rect 34188 16706 34244 16716
rect 34636 16100 34692 23102
rect 34972 21812 35028 26124
rect 35084 24164 35140 30268
rect 35196 30258 35252 30268
rect 35756 30324 35812 30492
rect 35756 30322 35924 30324
rect 35756 30270 35758 30322
rect 35810 30270 35924 30322
rect 35756 30268 35924 30270
rect 35756 30258 35812 30268
rect 35868 29540 35924 30268
rect 35980 29652 36036 30828
rect 36204 30772 36260 30782
rect 36428 30772 36484 30782
rect 36260 30770 36484 30772
rect 36260 30718 36430 30770
rect 36482 30718 36484 30770
rect 36260 30716 36484 30718
rect 36204 30706 36260 30716
rect 36428 30706 36484 30716
rect 35980 29596 36484 29652
rect 35868 29484 36148 29540
rect 35644 29428 35700 29438
rect 35196 29036 35460 29046
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35196 28970 35460 28980
rect 35644 28754 35700 29372
rect 35756 29428 35812 29438
rect 36092 29428 36148 29484
rect 35756 29426 36036 29428
rect 35756 29374 35758 29426
rect 35810 29374 36036 29426
rect 35756 29372 36036 29374
rect 35756 29362 35812 29372
rect 35644 28702 35646 28754
rect 35698 28702 35700 28754
rect 35644 28690 35700 28702
rect 35980 28756 36036 29372
rect 36092 29334 36148 29372
rect 36316 28868 36372 28878
rect 35980 28700 36148 28756
rect 35532 28644 35588 28654
rect 35532 28550 35588 28588
rect 35868 28644 35924 28654
rect 35924 28588 36036 28644
rect 35868 28550 35924 28588
rect 35196 28530 35252 28542
rect 35196 28478 35198 28530
rect 35250 28478 35252 28530
rect 35196 28196 35252 28478
rect 35196 28130 35252 28140
rect 35980 27746 36036 28588
rect 36092 28642 36148 28700
rect 36092 28590 36094 28642
rect 36146 28590 36148 28642
rect 36092 28578 36148 28590
rect 36316 28530 36372 28812
rect 36428 28756 36484 29596
rect 36428 28642 36484 28700
rect 36428 28590 36430 28642
rect 36482 28590 36484 28642
rect 36428 28578 36484 28590
rect 36316 28478 36318 28530
rect 36370 28478 36372 28530
rect 36316 28466 36372 28478
rect 35980 27694 35982 27746
rect 36034 27694 36036 27746
rect 35980 27682 36036 27694
rect 35196 27468 35460 27478
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35196 27402 35460 27412
rect 35196 27300 35252 27310
rect 35196 27206 35252 27244
rect 35756 27076 35812 27086
rect 35308 26964 35364 27002
rect 35308 26898 35364 26908
rect 35532 26964 35588 27002
rect 35756 26982 35812 27020
rect 35532 26898 35588 26908
rect 36316 26964 36372 27002
rect 35196 26404 35252 26414
rect 35196 26290 35252 26348
rect 35196 26238 35198 26290
rect 35250 26238 35252 26290
rect 35196 26226 35252 26238
rect 36092 26292 36148 26302
rect 36092 26198 36148 26236
rect 35868 26180 35924 26190
rect 35868 26066 35924 26124
rect 35868 26014 35870 26066
rect 35922 26014 35924 26066
rect 35868 26002 35924 26014
rect 35196 25900 35460 25910
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35196 25834 35460 25844
rect 35196 25618 35252 25630
rect 35196 25566 35198 25618
rect 35250 25566 35252 25618
rect 35196 25060 35252 25566
rect 36204 25508 36260 25518
rect 35868 25284 35924 25294
rect 35868 25190 35924 25228
rect 35196 24994 35252 25004
rect 36204 24722 36260 25452
rect 36204 24670 36206 24722
rect 36258 24670 36260 24722
rect 35196 24332 35460 24342
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35196 24266 35460 24276
rect 35084 24098 35140 24108
rect 36204 24050 36260 24670
rect 36204 23998 36206 24050
rect 36258 23998 36260 24050
rect 36204 23986 36260 23998
rect 35756 23938 35812 23950
rect 35756 23886 35758 23938
rect 35810 23886 35812 23938
rect 35196 23716 35252 23726
rect 35196 23622 35252 23660
rect 35756 23604 35812 23886
rect 35756 23538 35812 23548
rect 36316 23492 36372 26908
rect 36204 23436 36372 23492
rect 36428 26290 36484 26302
rect 36428 26238 36430 26290
rect 36482 26238 36484 26290
rect 35644 23268 35700 23278
rect 35532 23212 35644 23268
rect 35196 22764 35460 22774
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35196 22698 35460 22708
rect 35532 22596 35588 23212
rect 35644 23174 35700 23212
rect 34972 21746 35028 21756
rect 35420 22540 35588 22596
rect 35196 21588 35252 21598
rect 35196 21494 35252 21532
rect 35420 21364 35476 22540
rect 35644 22484 35700 22494
rect 35644 22390 35700 22428
rect 35868 21812 35924 21822
rect 35532 21698 35588 21710
rect 35532 21646 35534 21698
rect 35586 21646 35588 21698
rect 35532 21476 35588 21646
rect 35868 21698 35924 21756
rect 35868 21646 35870 21698
rect 35922 21646 35924 21698
rect 35868 21634 35924 21646
rect 35532 21420 35924 21476
rect 35420 21308 35588 21364
rect 35196 21196 35460 21206
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35196 21130 35460 21140
rect 35532 21028 35588 21308
rect 35420 20972 35588 21028
rect 34972 20690 35028 20702
rect 34972 20638 34974 20690
rect 35026 20638 35028 20690
rect 34748 20578 34804 20590
rect 34748 20526 34750 20578
rect 34802 20526 34804 20578
rect 34748 19796 34804 20526
rect 34860 20578 34916 20590
rect 34860 20526 34862 20578
rect 34914 20526 34916 20578
rect 34860 20244 34916 20526
rect 34860 20178 34916 20188
rect 34860 20020 34916 20030
rect 34860 19926 34916 19964
rect 34748 19730 34804 19740
rect 34972 19572 35028 20638
rect 34748 19516 35028 19572
rect 35084 20244 35140 20254
rect 34748 17780 34804 19516
rect 34972 19348 35028 19358
rect 34972 19254 35028 19292
rect 35084 19124 35140 20188
rect 35420 20018 35476 20972
rect 35420 19966 35422 20018
rect 35474 19966 35476 20018
rect 35420 19954 35476 19966
rect 35532 20578 35588 20590
rect 35532 20526 35534 20578
rect 35586 20526 35588 20578
rect 35196 19628 35460 19638
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35196 19562 35460 19572
rect 35308 19460 35364 19470
rect 35308 19366 35364 19404
rect 35420 19348 35476 19358
rect 34860 19068 35252 19124
rect 34860 18450 34916 19068
rect 34860 18398 34862 18450
rect 34914 18398 34916 18450
rect 34860 18386 34916 18398
rect 35084 18900 35140 18910
rect 35084 18340 35140 18844
rect 35196 18452 35252 19068
rect 35420 18564 35476 19292
rect 35308 18452 35364 18462
rect 35196 18450 35364 18452
rect 35196 18398 35310 18450
rect 35362 18398 35364 18450
rect 35196 18396 35364 18398
rect 35308 18386 35364 18396
rect 35084 18246 35140 18284
rect 34972 18228 35028 18238
rect 35420 18228 35476 18508
rect 35532 18450 35588 20526
rect 35644 20578 35700 20590
rect 35644 20526 35646 20578
rect 35698 20526 35700 20578
rect 35644 20356 35700 20526
rect 35756 20580 35812 20590
rect 35756 20486 35812 20524
rect 35868 20356 35924 21420
rect 36204 21028 36260 23436
rect 36316 23268 36372 23278
rect 36316 22372 36372 23212
rect 36428 22820 36484 26238
rect 36428 22754 36484 22764
rect 36316 22278 36372 22316
rect 36428 21700 36484 21710
rect 36428 21606 36484 21644
rect 36204 20972 36372 21028
rect 36204 20802 36260 20814
rect 36204 20750 36206 20802
rect 36258 20750 36260 20802
rect 35644 20290 35700 20300
rect 35756 20300 35924 20356
rect 36092 20356 36148 20366
rect 35644 19460 35700 19470
rect 35644 18900 35700 19404
rect 35756 19236 35812 20300
rect 36092 20130 36148 20300
rect 36092 20078 36094 20130
rect 36146 20078 36148 20130
rect 36092 20066 36148 20078
rect 36204 19460 36260 20750
rect 36204 19394 36260 19404
rect 35756 19142 35812 19180
rect 36092 19348 36148 19358
rect 36092 19234 36148 19292
rect 36092 19182 36094 19234
rect 36146 19182 36148 19234
rect 36092 19170 36148 19182
rect 35868 19124 35924 19134
rect 35868 19122 36036 19124
rect 35868 19070 35870 19122
rect 35922 19070 36036 19122
rect 35868 19068 36036 19070
rect 35868 19058 35924 19068
rect 35644 18844 35812 18900
rect 35756 18788 35812 18844
rect 35756 18732 35924 18788
rect 35532 18398 35534 18450
rect 35586 18398 35588 18450
rect 35532 18386 35588 18398
rect 35644 18676 35700 18686
rect 35420 18172 35588 18228
rect 34860 17780 34916 17790
rect 34748 17778 34916 17780
rect 34748 17726 34862 17778
rect 34914 17726 34916 17778
rect 34748 17724 34916 17726
rect 34860 17714 34916 17724
rect 34972 17666 35028 18172
rect 35196 18060 35460 18070
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35196 17994 35460 18004
rect 35532 17892 35588 18172
rect 35308 17836 35588 17892
rect 34972 17614 34974 17666
rect 35026 17614 35028 17666
rect 34972 17602 35028 17614
rect 35196 17668 35252 17678
rect 34748 17556 34804 17566
rect 34748 17462 34804 17500
rect 35196 17106 35252 17612
rect 35308 17666 35364 17836
rect 35308 17614 35310 17666
rect 35362 17614 35364 17666
rect 35308 17602 35364 17614
rect 35196 17054 35198 17106
rect 35250 17054 35252 17106
rect 35196 17042 35252 17054
rect 35644 17332 35700 18620
rect 35756 18450 35812 18462
rect 35756 18398 35758 18450
rect 35810 18398 35812 18450
rect 35756 18340 35812 18398
rect 35868 18450 35924 18732
rect 35868 18398 35870 18450
rect 35922 18398 35924 18450
rect 35868 18386 35924 18398
rect 35756 17444 35812 18284
rect 35980 18228 36036 19068
rect 36316 18788 36372 20972
rect 36540 19012 36596 31612
rect 37548 31220 37604 31724
rect 38220 31220 38276 31230
rect 37548 31218 38276 31220
rect 37548 31166 38222 31218
rect 38274 31166 38276 31218
rect 37548 31164 38276 31166
rect 38220 31154 38276 31164
rect 36988 31108 37044 31118
rect 36988 30882 37044 31052
rect 38108 30996 38164 31006
rect 38108 30902 38164 30940
rect 38332 30994 38388 31006
rect 38332 30942 38334 30994
rect 38386 30942 38388 30994
rect 36988 30830 36990 30882
rect 37042 30830 37044 30882
rect 36988 30772 37044 30830
rect 38332 30884 38388 30942
rect 38332 30818 38388 30828
rect 36988 30706 37044 30716
rect 37324 30212 37380 30222
rect 37884 30212 37940 30222
rect 37324 30210 37940 30212
rect 37324 30158 37326 30210
rect 37378 30158 37886 30210
rect 37938 30158 37940 30210
rect 37324 30156 37940 30158
rect 37324 30146 37380 30156
rect 37884 30146 37940 30156
rect 38332 30210 38388 30222
rect 38332 30158 38334 30210
rect 38386 30158 38388 30210
rect 36988 30098 37044 30110
rect 36988 30046 36990 30098
rect 37042 30046 37044 30098
rect 36652 29652 36708 29662
rect 36652 29314 36708 29596
rect 36652 29262 36654 29314
rect 36706 29262 36708 29314
rect 36652 28196 36708 29262
rect 36988 28868 37044 30046
rect 38332 30100 38388 30158
rect 38332 30034 38388 30044
rect 37100 29988 37156 29998
rect 37100 29894 37156 29932
rect 38444 29876 38500 33068
rect 39452 32004 39508 34190
rect 40012 34242 40068 34254
rect 40012 34190 40014 34242
rect 40066 34190 40068 34242
rect 39564 33124 39620 33134
rect 40012 33124 40068 34190
rect 40124 34244 40180 34254
rect 40236 34244 40292 34748
rect 40460 34738 40516 34748
rect 40796 34916 40852 34926
rect 41020 34916 41076 35532
rect 41244 34916 41300 34926
rect 41020 34914 41300 34916
rect 41020 34862 41246 34914
rect 41298 34862 41300 34914
rect 41020 34860 41300 34862
rect 40124 34242 40292 34244
rect 40124 34190 40126 34242
rect 40178 34190 40292 34242
rect 40124 34188 40292 34190
rect 40124 34178 40180 34188
rect 40684 34132 40740 34142
rect 39564 33122 40068 33124
rect 39564 33070 39566 33122
rect 39618 33070 40068 33122
rect 39564 33068 40068 33070
rect 40348 34076 40684 34132
rect 39564 32004 39620 33068
rect 40348 32452 40404 34076
rect 40684 34066 40740 34076
rect 40796 33348 40852 34860
rect 41244 34850 41300 34860
rect 40908 34804 40964 34814
rect 40908 34244 40964 34748
rect 41356 34690 41412 34702
rect 41356 34638 41358 34690
rect 41410 34638 41412 34690
rect 41132 34580 41188 34590
rect 41132 34356 41188 34524
rect 41244 34356 41300 34366
rect 41132 34354 41300 34356
rect 41132 34302 41246 34354
rect 41298 34302 41300 34354
rect 41132 34300 41300 34302
rect 41244 34290 41300 34300
rect 40908 34150 40964 34188
rect 41020 34242 41076 34254
rect 41020 34190 41022 34242
rect 41074 34190 41076 34242
rect 41020 34132 41076 34190
rect 41020 34066 41076 34076
rect 40908 33348 40964 33358
rect 40796 33346 40964 33348
rect 40796 33294 40910 33346
rect 40962 33294 40964 33346
rect 40796 33292 40964 33294
rect 40908 33282 40964 33292
rect 41244 33348 41300 33358
rect 41356 33348 41412 34638
rect 41468 34580 41524 36428
rect 41580 36260 41636 36270
rect 41580 34914 41636 36204
rect 42140 35586 42196 35598
rect 42140 35534 42142 35586
rect 42194 35534 42196 35586
rect 41692 35028 41748 35038
rect 41692 35026 42084 35028
rect 41692 34974 41694 35026
rect 41746 34974 42084 35026
rect 41692 34972 42084 34974
rect 41692 34962 41748 34972
rect 41580 34862 41582 34914
rect 41634 34862 41636 34914
rect 41580 34850 41636 34862
rect 41692 34692 41748 34702
rect 41692 34690 41860 34692
rect 41692 34638 41694 34690
rect 41746 34638 41860 34690
rect 41692 34636 41860 34638
rect 41692 34626 41748 34636
rect 41468 34514 41524 34524
rect 41804 34580 41860 34636
rect 41804 34514 41860 34524
rect 42028 34356 42084 34972
rect 42140 34468 42196 35534
rect 42252 35588 42308 36428
rect 42252 35522 42308 35532
rect 42252 34916 42308 34926
rect 42364 34916 42420 36652
rect 42588 36372 42644 36382
rect 42700 36372 42756 37774
rect 43708 37828 43764 37838
rect 43708 37734 43764 37772
rect 42812 37492 42868 37502
rect 42812 36484 42868 37436
rect 42812 36390 42868 36428
rect 43260 37044 43316 37054
rect 42588 36370 42756 36372
rect 42588 36318 42590 36370
rect 42642 36318 42756 36370
rect 42588 36316 42756 36318
rect 42588 36306 42644 36316
rect 42700 35924 42756 36316
rect 42252 34914 42420 34916
rect 42252 34862 42254 34914
rect 42306 34862 42420 34914
rect 42252 34860 42420 34862
rect 42588 35476 42644 35486
rect 42588 34914 42644 35420
rect 42588 34862 42590 34914
rect 42642 34862 42644 34914
rect 42252 34850 42308 34860
rect 42588 34850 42644 34862
rect 42700 34914 42756 35868
rect 43260 35138 43316 36988
rect 43820 37044 43876 37886
rect 45164 37268 45220 37278
rect 45220 37212 45444 37268
rect 45164 37174 45220 37212
rect 43820 36978 43876 36988
rect 44716 37154 44772 37166
rect 44716 37102 44718 37154
rect 44770 37102 44772 37154
rect 44716 37044 44772 37102
rect 44716 36978 44772 36988
rect 44940 36932 44996 36942
rect 43484 36596 43540 36606
rect 43484 36502 43540 36540
rect 44380 36596 44436 36606
rect 44268 36370 44324 36382
rect 44268 36318 44270 36370
rect 44322 36318 44324 36370
rect 43372 36260 43428 36270
rect 43372 36166 43428 36204
rect 44156 36258 44212 36270
rect 44156 36206 44158 36258
rect 44210 36206 44212 36258
rect 44156 35476 44212 36206
rect 44268 35700 44324 36318
rect 44268 35586 44324 35644
rect 44268 35534 44270 35586
rect 44322 35534 44324 35586
rect 44268 35522 44324 35534
rect 44156 35410 44212 35420
rect 43260 35086 43262 35138
rect 43314 35086 43316 35138
rect 43260 35074 43316 35086
rect 42700 34862 42702 34914
rect 42754 34862 42756 34914
rect 42364 34692 42420 34702
rect 42364 34598 42420 34636
rect 42476 34690 42532 34702
rect 42476 34638 42478 34690
rect 42530 34638 42532 34690
rect 42476 34468 42532 34638
rect 42700 34580 42756 34862
rect 43148 34804 43204 34814
rect 43148 34710 43204 34748
rect 43932 34804 43988 34814
rect 43932 34710 43988 34748
rect 42700 34514 42756 34524
rect 43260 34690 43316 34702
rect 43260 34638 43262 34690
rect 43314 34638 43316 34690
rect 42140 34412 42532 34468
rect 42028 34300 42308 34356
rect 42252 34242 42308 34300
rect 42252 34190 42254 34242
rect 42306 34190 42308 34242
rect 42252 34178 42308 34190
rect 41244 33346 41412 33348
rect 41244 33294 41246 33346
rect 41298 33294 41412 33346
rect 41244 33292 41412 33294
rect 41468 34130 41524 34142
rect 41468 34078 41470 34130
rect 41522 34078 41524 34130
rect 41244 33282 41300 33292
rect 40684 33124 40740 33134
rect 40684 33030 40740 33068
rect 41020 33124 41076 33134
rect 41020 33030 41076 33068
rect 40012 32450 40404 32452
rect 40012 32398 40350 32450
rect 40402 32398 40404 32450
rect 40012 32396 40404 32398
rect 39900 32340 39956 32350
rect 39564 31948 39844 32004
rect 39452 31938 39508 31948
rect 39004 31892 39060 31902
rect 39004 31798 39060 31836
rect 39452 31780 39508 31790
rect 39676 31780 39732 31790
rect 39452 31778 39732 31780
rect 39452 31726 39454 31778
rect 39506 31726 39678 31778
rect 39730 31726 39732 31778
rect 39452 31724 39732 31726
rect 39452 31714 39508 31724
rect 39676 31714 39732 31724
rect 38892 31556 38948 31566
rect 38892 31462 38948 31500
rect 39116 31554 39172 31566
rect 39116 31502 39118 31554
rect 39170 31502 39172 31554
rect 39004 31220 39060 31230
rect 39116 31220 39172 31502
rect 39004 31218 39172 31220
rect 39004 31166 39006 31218
rect 39058 31166 39172 31218
rect 39004 31164 39172 31166
rect 39004 31154 39060 31164
rect 38668 30994 38724 31006
rect 38668 30942 38670 30994
rect 38722 30942 38724 30994
rect 38220 29820 38500 29876
rect 38556 29988 38612 29998
rect 37436 29540 37492 29550
rect 37212 29428 37268 29438
rect 37212 29334 37268 29372
rect 36988 28812 37156 28868
rect 36988 28644 37044 28654
rect 36988 28550 37044 28588
rect 37100 28532 37156 28812
rect 37100 28466 37156 28476
rect 36652 28130 36708 28140
rect 36988 28196 37044 28206
rect 36652 27972 36708 27982
rect 36652 19348 36708 27916
rect 36876 26180 36932 26190
rect 36876 26086 36932 26124
rect 36764 26066 36820 26078
rect 36764 26014 36766 26066
rect 36818 26014 36820 26066
rect 36764 22484 36820 26014
rect 36988 25956 37044 28140
rect 37436 27860 37492 29484
rect 37548 29538 37604 29550
rect 37548 29486 37550 29538
rect 37602 29486 37604 29538
rect 37548 29428 37604 29486
rect 37548 29362 37604 29372
rect 38108 29316 38164 29326
rect 38108 29222 38164 29260
rect 37548 28868 37604 28878
rect 37548 28754 37604 28812
rect 37548 28702 37550 28754
rect 37602 28702 37604 28754
rect 37548 28690 37604 28702
rect 36764 22418 36820 22428
rect 36876 25900 37044 25956
rect 37100 27858 37492 27860
rect 37100 27806 37438 27858
rect 37490 27806 37492 27858
rect 37100 27804 37492 27806
rect 36876 21924 36932 25900
rect 37100 25506 37156 27804
rect 37436 27794 37492 27804
rect 37996 28530 38052 28542
rect 37996 28478 37998 28530
rect 38050 28478 38052 28530
rect 37996 27186 38052 28478
rect 38108 28420 38164 28430
rect 38108 28326 38164 28364
rect 38220 28196 38276 29820
rect 38332 29428 38388 29438
rect 38332 28756 38388 29372
rect 38332 28690 38388 28700
rect 38556 29426 38612 29932
rect 38556 29374 38558 29426
rect 38610 29374 38612 29426
rect 37996 27134 37998 27186
rect 38050 27134 38052 27186
rect 37996 27122 38052 27134
rect 38108 28140 38276 28196
rect 38332 28418 38388 28430
rect 38332 28366 38334 28418
rect 38386 28366 38388 28418
rect 37772 27076 37828 27086
rect 37324 26964 37380 27002
rect 37324 26898 37380 26908
rect 37548 26964 37604 27002
rect 37772 26982 37828 27020
rect 37548 26898 37604 26908
rect 37996 26852 38052 26862
rect 37996 26758 38052 26796
rect 37100 25454 37102 25506
rect 37154 25454 37156 25506
rect 37100 25442 37156 25454
rect 37212 26628 37268 26638
rect 37100 24610 37156 24622
rect 37100 24558 37102 24610
rect 37154 24558 37156 24610
rect 37100 24164 37156 24558
rect 37100 24098 37156 24108
rect 36988 23828 37044 23838
rect 36988 23734 37044 23772
rect 37212 23044 37268 26572
rect 37884 26292 37940 26302
rect 37884 26198 37940 26236
rect 37324 26178 37380 26190
rect 37324 26126 37326 26178
rect 37378 26126 37380 26178
rect 37324 23828 37380 26126
rect 37436 26068 37492 26078
rect 37436 26066 37828 26068
rect 37436 26014 37438 26066
rect 37490 26014 37828 26066
rect 37436 26012 37828 26014
rect 37436 26002 37492 26012
rect 37772 25618 37828 26012
rect 37772 25566 37774 25618
rect 37826 25566 37828 25618
rect 37772 25554 37828 25566
rect 37436 23940 37492 23950
rect 37436 23846 37492 23884
rect 37996 23940 38052 23950
rect 37996 23846 38052 23884
rect 37324 23762 37380 23772
rect 36876 21858 36932 21868
rect 36988 22988 37268 23044
rect 36988 19908 37044 22988
rect 37100 22820 37156 22830
rect 37100 21700 37156 22764
rect 37548 22372 37604 22382
rect 37548 22278 37604 22316
rect 37996 21812 38052 21822
rect 37100 21698 37268 21700
rect 37100 21646 37102 21698
rect 37154 21646 37268 21698
rect 37100 21644 37268 21646
rect 37100 21634 37156 21644
rect 37212 21364 37268 21644
rect 37548 21588 37604 21598
rect 37548 21586 37716 21588
rect 37548 21534 37550 21586
rect 37602 21534 37716 21586
rect 37548 21532 37716 21534
rect 37548 21522 37604 21532
rect 37212 21308 37604 21364
rect 37548 20802 37604 21308
rect 37548 20750 37550 20802
rect 37602 20750 37604 20802
rect 37548 20738 37604 20750
rect 37100 20580 37156 20590
rect 37660 20580 37716 21532
rect 37996 21474 38052 21756
rect 37996 21422 37998 21474
rect 38050 21422 38052 21474
rect 37996 21252 38052 21422
rect 38108 21476 38164 28140
rect 38220 27746 38276 27758
rect 38220 27694 38222 27746
rect 38274 27694 38276 27746
rect 38220 26908 38276 27694
rect 38332 27074 38388 28366
rect 38332 27022 38334 27074
rect 38386 27022 38388 27074
rect 38332 27010 38388 27022
rect 38556 27076 38612 29374
rect 38668 29314 38724 30942
rect 38780 30996 38836 31006
rect 38780 30324 38836 30940
rect 39340 30996 39396 31006
rect 39340 30902 39396 30940
rect 39452 30884 39508 30894
rect 39564 30884 39620 30894
rect 39508 30882 39620 30884
rect 39508 30830 39566 30882
rect 39618 30830 39620 30882
rect 39508 30828 39620 30830
rect 38780 30322 38948 30324
rect 38780 30270 38782 30322
rect 38834 30270 38948 30322
rect 38780 30268 38948 30270
rect 38780 30258 38836 30268
rect 38892 30100 38948 30268
rect 39228 30212 39284 30222
rect 39228 30118 39284 30156
rect 39116 30100 39172 30110
rect 38892 30098 39172 30100
rect 38892 30046 39118 30098
rect 39170 30046 39172 30098
rect 38892 30044 39172 30046
rect 39116 30034 39172 30044
rect 39340 29988 39396 30026
rect 39452 29988 39508 30828
rect 39564 30818 39620 30828
rect 39564 30660 39620 30670
rect 39564 30098 39620 30604
rect 39564 30046 39566 30098
rect 39618 30046 39620 30098
rect 39564 30034 39620 30046
rect 39396 29932 39508 29988
rect 39340 29922 39396 29932
rect 38780 29876 38836 29886
rect 39004 29876 39060 29886
rect 38780 29650 38836 29820
rect 38780 29598 38782 29650
rect 38834 29598 38836 29650
rect 38780 29586 38836 29598
rect 38892 29820 39004 29876
rect 38668 29262 38670 29314
rect 38722 29262 38724 29314
rect 38668 29250 38724 29262
rect 38668 28756 38724 28766
rect 38668 28662 38724 28700
rect 38556 27010 38612 27020
rect 38444 26962 38500 26974
rect 38444 26910 38446 26962
rect 38498 26910 38500 26962
rect 38444 26908 38500 26910
rect 38220 26852 38500 26908
rect 38556 26850 38612 26862
rect 38556 26798 38558 26850
rect 38610 26798 38612 26850
rect 38332 26628 38388 26638
rect 38556 26628 38612 26798
rect 38556 26572 38836 26628
rect 38332 26516 38388 26572
rect 38332 26514 38612 26516
rect 38332 26462 38334 26514
rect 38386 26462 38612 26514
rect 38332 26460 38612 26462
rect 38332 26450 38388 26460
rect 38556 26290 38612 26460
rect 38780 26514 38836 26572
rect 38780 26462 38782 26514
rect 38834 26462 38836 26514
rect 38780 26450 38836 26462
rect 38556 26238 38558 26290
rect 38610 26238 38612 26290
rect 38556 26226 38612 26238
rect 38780 24164 38836 24174
rect 38780 24050 38836 24108
rect 38780 23998 38782 24050
rect 38834 23998 38836 24050
rect 38780 23986 38836 23998
rect 38668 23828 38724 23838
rect 38332 22258 38388 22270
rect 38332 22206 38334 22258
rect 38386 22206 38388 22258
rect 38332 21812 38388 22206
rect 38332 21746 38388 21756
rect 38556 21588 38612 21598
rect 38556 21494 38612 21532
rect 38108 21410 38164 21420
rect 38668 21362 38724 23772
rect 38892 23548 38948 29820
rect 39004 29810 39060 29820
rect 39788 29876 39844 31948
rect 39788 29810 39844 29820
rect 39900 31666 39956 32284
rect 39900 31614 39902 31666
rect 39954 31614 39956 31666
rect 39900 31220 39956 31614
rect 39340 29708 39732 29764
rect 39340 29650 39396 29708
rect 39340 29598 39342 29650
rect 39394 29598 39396 29650
rect 39340 29586 39396 29598
rect 39676 29652 39732 29708
rect 39900 29652 39956 31164
rect 40012 31778 40068 32396
rect 40348 32386 40404 32396
rect 40012 31726 40014 31778
rect 40066 31726 40068 31778
rect 40012 30100 40068 31726
rect 41132 31780 41188 31790
rect 41468 31780 41524 34078
rect 43036 32788 43092 32798
rect 43036 32694 43092 32732
rect 43260 32676 43316 34638
rect 43596 34692 43652 34702
rect 43596 34598 43652 34636
rect 43820 34690 43876 34702
rect 43820 34638 43822 34690
rect 43874 34638 43876 34690
rect 43820 33684 43876 34638
rect 44380 34018 44436 36540
rect 44716 35588 44772 35598
rect 44716 35494 44772 35532
rect 44940 35138 44996 36876
rect 45164 36484 45220 36494
rect 45164 35924 45220 36428
rect 45164 35830 45220 35868
rect 45388 35476 45444 37212
rect 45836 37156 45892 37166
rect 45836 37062 45892 37100
rect 45500 35924 45556 35934
rect 45500 35830 45556 35868
rect 45836 35924 45892 35934
rect 45836 35830 45892 35868
rect 45388 35410 45444 35420
rect 44940 35086 44942 35138
rect 44994 35086 44996 35138
rect 44940 35074 44996 35086
rect 45724 34914 45780 34926
rect 45724 34862 45726 34914
rect 45778 34862 45780 34914
rect 44828 34804 44884 34814
rect 44828 34710 44884 34748
rect 44940 34690 44996 34702
rect 44940 34638 44942 34690
rect 44994 34638 44996 34690
rect 44828 34020 44884 34030
rect 44940 34020 44996 34638
rect 45724 34468 45780 34862
rect 45948 34692 46004 34702
rect 45948 34598 46004 34636
rect 45724 34356 45780 34412
rect 45948 34356 46004 34366
rect 45724 34354 46004 34356
rect 45724 34302 45950 34354
rect 46002 34302 46004 34354
rect 45724 34300 46004 34302
rect 45948 34290 46004 34300
rect 45612 34244 45668 34254
rect 45612 34150 45668 34188
rect 44380 33966 44382 34018
rect 44434 33966 44436 34018
rect 44380 33908 44436 33966
rect 44380 33842 44436 33852
rect 44716 34018 44996 34020
rect 44716 33966 44830 34018
rect 44882 33966 44996 34018
rect 44716 33964 44996 33966
rect 43596 33628 43876 33684
rect 43372 33124 43428 33134
rect 43596 33124 43652 33628
rect 43372 33122 43652 33124
rect 43372 33070 43374 33122
rect 43426 33070 43652 33122
rect 43372 33068 43652 33070
rect 44156 33124 44212 33134
rect 43372 33058 43428 33068
rect 43148 32620 43316 32676
rect 43148 31892 43204 32620
rect 42924 31836 43148 31892
rect 41132 31778 41524 31780
rect 41132 31726 41134 31778
rect 41186 31726 41524 31778
rect 41132 31724 41524 31726
rect 42812 31780 42868 31790
rect 40572 30212 40628 30222
rect 40572 30118 40628 30156
rect 40796 30100 40852 30110
rect 40012 30034 40068 30044
rect 40684 30044 40796 30100
rect 40460 29988 40516 29998
rect 40460 29894 40516 29932
rect 39676 29596 39956 29652
rect 40460 29652 40516 29662
rect 40684 29652 40740 30044
rect 40796 30034 40852 30044
rect 40460 29650 40740 29652
rect 40460 29598 40462 29650
rect 40514 29598 40740 29650
rect 40460 29596 40740 29598
rect 40460 29586 40516 29596
rect 40236 29538 40292 29550
rect 40236 29486 40238 29538
rect 40290 29486 40292 29538
rect 39116 29428 39172 29438
rect 39004 29426 39172 29428
rect 39004 29374 39118 29426
rect 39170 29374 39172 29426
rect 39004 29372 39172 29374
rect 39004 27074 39060 29372
rect 39116 29362 39172 29372
rect 39452 29426 39508 29438
rect 39452 29374 39454 29426
rect 39506 29374 39508 29426
rect 39452 29204 39508 29374
rect 40124 29426 40180 29438
rect 40124 29374 40126 29426
rect 40178 29374 40180 29426
rect 39452 29138 39508 29148
rect 40012 29204 40068 29214
rect 39788 28866 39844 28878
rect 39788 28814 39790 28866
rect 39842 28814 39844 28866
rect 39788 28642 39844 28814
rect 39788 28590 39790 28642
rect 39842 28590 39844 28642
rect 39116 28532 39172 28542
rect 39116 28438 39172 28476
rect 39788 27972 39844 28590
rect 39788 27906 39844 27916
rect 40012 28084 40068 29148
rect 40124 28866 40180 29374
rect 40124 28814 40126 28866
rect 40178 28814 40180 28866
rect 40124 28802 40180 28814
rect 40236 28644 40292 29486
rect 41132 29540 41188 31724
rect 41916 31668 41972 31678
rect 41916 31666 42196 31668
rect 41916 31614 41918 31666
rect 41970 31614 42196 31666
rect 41916 31612 42196 31614
rect 41916 31602 41972 31612
rect 41244 31220 41300 31230
rect 41244 31126 41300 31164
rect 42140 31218 42196 31612
rect 42140 31166 42142 31218
rect 42194 31166 42196 31218
rect 42140 31154 42196 31166
rect 42252 31220 42308 31230
rect 42700 31220 42756 31230
rect 42252 31218 42756 31220
rect 42252 31166 42254 31218
rect 42306 31166 42702 31218
rect 42754 31166 42756 31218
rect 42252 31164 42756 31166
rect 42252 31154 42308 31164
rect 42700 31154 42756 31164
rect 42812 31220 42868 31724
rect 42812 31154 42868 31164
rect 41356 30996 41412 31006
rect 41580 30996 41636 31006
rect 41356 30902 41412 30940
rect 41468 30994 41636 30996
rect 41468 30942 41582 30994
rect 41634 30942 41636 30994
rect 41468 30940 41636 30942
rect 41244 30772 41300 30782
rect 41468 30772 41524 30940
rect 41580 30930 41636 30940
rect 42028 30996 42084 31006
rect 42476 30996 42532 31006
rect 42028 30994 42420 30996
rect 42028 30942 42030 30994
rect 42082 30942 42420 30994
rect 42028 30940 42420 30942
rect 42028 30930 42084 30940
rect 41244 30770 41524 30772
rect 41244 30718 41246 30770
rect 41298 30718 41524 30770
rect 41244 30716 41524 30718
rect 42252 30772 42308 30782
rect 41244 30706 41300 30716
rect 42140 30322 42196 30334
rect 42140 30270 42142 30322
rect 42194 30270 42196 30322
rect 41468 30210 41524 30222
rect 41468 30158 41470 30210
rect 41522 30158 41524 30210
rect 41132 29446 41188 29484
rect 41356 30098 41412 30110
rect 41356 30046 41358 30098
rect 41410 30046 41412 30098
rect 41356 29876 41412 30046
rect 41468 29988 41524 30158
rect 42140 30100 42196 30270
rect 42252 30210 42308 30716
rect 42252 30158 42254 30210
rect 42306 30158 42308 30210
rect 42252 30146 42308 30158
rect 42140 30034 42196 30044
rect 41468 29922 41524 29932
rect 40460 29428 40516 29438
rect 40348 28756 40404 28766
rect 40460 28756 40516 29372
rect 41356 28866 41412 29820
rect 41356 28814 41358 28866
rect 41410 28814 41412 28866
rect 41356 28802 41412 28814
rect 42364 28866 42420 30940
rect 42364 28814 42366 28866
rect 42418 28814 42420 28866
rect 42364 28802 42420 28814
rect 40348 28754 40516 28756
rect 40348 28702 40350 28754
rect 40402 28702 40516 28754
rect 40348 28700 40516 28702
rect 40348 28690 40404 28700
rect 40236 28578 40292 28588
rect 39004 27022 39006 27074
rect 39058 27022 39060 27074
rect 39004 27010 39060 27022
rect 39116 27020 39508 27076
rect 39116 26964 39172 27020
rect 39452 26962 39508 27020
rect 38668 21310 38670 21362
rect 38722 21310 38724 21362
rect 38668 21298 38724 21310
rect 38780 23492 38948 23548
rect 39004 26852 39060 26862
rect 39004 26402 39060 26796
rect 39004 26350 39006 26402
rect 39058 26350 39060 26402
rect 37996 21196 38500 21252
rect 38444 20914 38500 21196
rect 38444 20862 38446 20914
rect 38498 20862 38500 20914
rect 38444 20850 38500 20862
rect 37156 20524 37268 20580
rect 37100 20486 37156 20524
rect 36876 19852 37044 19908
rect 36876 19572 36932 19852
rect 37212 19684 37268 20524
rect 37212 19618 37268 19628
rect 37548 20524 37660 20580
rect 36876 19516 37044 19572
rect 36708 19292 36932 19348
rect 36652 19282 36708 19292
rect 36540 18946 36596 18956
rect 36316 18722 36372 18732
rect 35980 18162 36036 18172
rect 36092 18564 36148 18574
rect 36316 18564 36372 18574
rect 35868 18116 35924 18126
rect 35868 17666 35924 18060
rect 36092 17892 36148 18508
rect 35980 17836 36148 17892
rect 36204 18562 36372 18564
rect 36204 18510 36318 18562
rect 36370 18510 36372 18562
rect 36204 18508 36372 18510
rect 35980 17778 36036 17836
rect 35980 17726 35982 17778
rect 36034 17726 36036 17778
rect 35980 17714 36036 17726
rect 35868 17614 35870 17666
rect 35922 17614 35924 17666
rect 35868 17602 35924 17614
rect 36204 17666 36260 18508
rect 36316 18498 36372 18508
rect 36540 18450 36596 18462
rect 36540 18398 36542 18450
rect 36594 18398 36596 18450
rect 36204 17614 36206 17666
rect 36258 17614 36260 17666
rect 36204 17444 36260 17614
rect 35756 17388 35924 17444
rect 34748 16884 34804 16894
rect 34972 16884 35028 16894
rect 34748 16790 34804 16828
rect 34860 16882 35028 16884
rect 34860 16830 34974 16882
rect 35026 16830 35028 16882
rect 34860 16828 35028 16830
rect 34748 16100 34804 16110
rect 34636 16044 34748 16100
rect 34748 16034 34804 16044
rect 34860 15876 34916 16828
rect 34972 16818 35028 16828
rect 35308 16882 35364 16894
rect 35308 16830 35310 16882
rect 35362 16830 35364 16882
rect 35308 16660 35364 16830
rect 35644 16884 35700 17276
rect 35756 17108 35812 17118
rect 35756 17014 35812 17052
rect 35644 16818 35700 16828
rect 35420 16660 35476 16670
rect 32844 15148 32900 15708
rect 33180 15708 33348 15764
rect 34636 15820 34916 15876
rect 35084 16604 35420 16660
rect 33180 15652 33236 15708
rect 31836 14590 31838 14642
rect 31890 14590 31892 14642
rect 31836 14578 31892 14590
rect 31948 14700 32676 14756
rect 31948 13746 32004 14700
rect 31948 13694 31950 13746
rect 32002 13694 32004 13746
rect 31948 13682 32004 13694
rect 32172 14530 32228 14542
rect 32172 14478 32174 14530
rect 32226 14478 32228 14530
rect 32172 13524 32228 14478
rect 32620 14530 32676 14700
rect 32620 14478 32622 14530
rect 32674 14478 32676 14530
rect 32620 14466 32676 14478
rect 32732 15092 32900 15148
rect 32956 15596 33236 15652
rect 33404 15652 33460 15662
rect 32396 13634 32452 13646
rect 32396 13582 32398 13634
rect 32450 13582 32452 13634
rect 32284 13524 32340 13534
rect 32172 13522 32340 13524
rect 32172 13470 32286 13522
rect 32338 13470 32340 13522
rect 32172 13468 32340 13470
rect 32284 13458 32340 13468
rect 32396 13074 32452 13582
rect 32396 13022 32398 13074
rect 32450 13022 32452 13074
rect 32396 13010 32452 13022
rect 31612 12114 31668 12124
rect 31948 12962 32004 12974
rect 31948 12910 31950 12962
rect 32002 12910 32004 12962
rect 31836 12068 31892 12078
rect 31948 12068 32004 12910
rect 32508 12964 32564 12974
rect 32732 12964 32788 15092
rect 32564 12908 32788 12964
rect 32508 12850 32564 12908
rect 32508 12798 32510 12850
rect 32562 12798 32564 12850
rect 32284 12738 32340 12750
rect 32284 12686 32286 12738
rect 32338 12686 32340 12738
rect 32284 12292 32340 12686
rect 32396 12404 32452 12414
rect 32508 12404 32564 12798
rect 32396 12402 32508 12404
rect 32396 12350 32398 12402
rect 32450 12350 32508 12402
rect 32396 12348 32508 12350
rect 32396 12338 32452 12348
rect 32508 12310 32564 12348
rect 32284 12226 32340 12236
rect 31836 12066 32004 12068
rect 31836 12014 31838 12066
rect 31890 12014 32004 12066
rect 31836 12012 32004 12014
rect 31836 12002 31892 12012
rect 31948 11732 32004 12012
rect 31948 11666 32004 11676
rect 32620 11956 32676 11966
rect 32060 11620 32116 11630
rect 32060 11618 32564 11620
rect 32060 11566 32062 11618
rect 32114 11566 32564 11618
rect 32060 11564 32564 11566
rect 32060 11554 32116 11564
rect 31948 11506 32004 11518
rect 31948 11454 31950 11506
rect 32002 11454 32004 11506
rect 31500 11396 31556 11406
rect 31276 11394 31556 11396
rect 31276 11342 31502 11394
rect 31554 11342 31556 11394
rect 31276 11340 31556 11342
rect 31052 9938 31108 11340
rect 31052 9886 31054 9938
rect 31106 9886 31108 9938
rect 31052 9874 31108 9886
rect 31276 9828 31332 9838
rect 31388 9828 31444 11340
rect 31500 11330 31556 11340
rect 31948 11284 32004 11454
rect 32508 11506 32564 11564
rect 32508 11454 32510 11506
rect 32562 11454 32564 11506
rect 32508 11442 32564 11454
rect 32620 11284 32676 11900
rect 32956 11396 33012 15596
rect 33292 15540 33348 15550
rect 33292 15446 33348 15484
rect 33068 15428 33124 15438
rect 33068 15314 33124 15372
rect 33404 15316 33460 15596
rect 33068 15262 33070 15314
rect 33122 15262 33124 15314
rect 33068 15250 33124 15262
rect 33292 15260 33460 15316
rect 33516 15426 33572 15438
rect 33516 15374 33518 15426
rect 33570 15374 33572 15426
rect 33516 15316 33572 15374
rect 33180 15204 33236 15242
rect 33180 15138 33236 15148
rect 33180 13076 33236 13086
rect 33292 13076 33348 15260
rect 33516 15250 33572 15260
rect 33964 15316 34020 15354
rect 33964 15250 34020 15260
rect 34188 15314 34244 15326
rect 34188 15262 34190 15314
rect 34242 15262 34244 15314
rect 34076 15202 34132 15214
rect 34076 15150 34078 15202
rect 34130 15150 34132 15202
rect 34076 15148 34132 15150
rect 33404 15092 34132 15148
rect 33404 14642 33460 15092
rect 33404 14590 33406 14642
rect 33458 14590 33460 14642
rect 33404 14578 33460 14590
rect 33628 14980 33684 14990
rect 33404 13860 33460 13870
rect 33404 13766 33460 13804
rect 33628 13636 33684 14924
rect 34188 13972 34244 15262
rect 34636 15314 34692 15820
rect 34636 15262 34638 15314
rect 34690 15262 34692 15314
rect 34636 15250 34692 15262
rect 34748 15314 34804 15326
rect 34748 15262 34750 15314
rect 34802 15262 34804 15314
rect 34748 14868 34804 15262
rect 34748 14802 34804 14812
rect 35084 14756 35140 16604
rect 35420 16594 35476 16604
rect 35196 16492 35460 16502
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35196 16426 35460 16436
rect 35644 16100 35700 16110
rect 35196 15652 35252 15662
rect 35196 15538 35252 15596
rect 35196 15486 35198 15538
rect 35250 15486 35252 15538
rect 35196 15474 35252 15486
rect 35308 15316 35364 15326
rect 35308 15222 35364 15260
rect 35420 15314 35476 15326
rect 35420 15262 35422 15314
rect 35474 15262 35476 15314
rect 35420 15092 35476 15262
rect 35420 15026 35476 15036
rect 35644 15204 35700 16044
rect 35868 15538 35924 17388
rect 36204 17378 36260 17388
rect 36316 18338 36372 18350
rect 36316 18286 36318 18338
rect 36370 18286 36372 18338
rect 36204 17108 36260 17118
rect 36204 16100 36260 17052
rect 36316 16996 36372 18286
rect 36540 17668 36596 18398
rect 36652 18452 36708 18462
rect 36652 17780 36708 18396
rect 36652 17714 36708 17724
rect 36764 18450 36820 18462
rect 36764 18398 36766 18450
rect 36818 18398 36820 18450
rect 36540 17602 36596 17612
rect 36428 17554 36484 17566
rect 36428 17502 36430 17554
rect 36482 17502 36484 17554
rect 36428 17444 36484 17502
rect 36764 17444 36820 18398
rect 36428 17388 36820 17444
rect 36540 17220 36596 17230
rect 36540 17106 36596 17164
rect 36540 17054 36542 17106
rect 36594 17054 36596 17106
rect 36540 17042 36596 17054
rect 36652 17108 36708 17388
rect 36652 17042 36708 17052
rect 36428 16996 36484 17006
rect 36316 16994 36484 16996
rect 36316 16942 36430 16994
rect 36482 16942 36484 16994
rect 36316 16940 36484 16942
rect 36428 16930 36484 16940
rect 36540 16884 36596 16894
rect 36540 16658 36596 16828
rect 36540 16606 36542 16658
rect 36594 16606 36596 16658
rect 36540 16594 36596 16606
rect 36204 16044 36820 16100
rect 35980 15876 36036 15886
rect 36204 15876 36260 15886
rect 36036 15874 36260 15876
rect 36036 15822 36206 15874
rect 36258 15822 36260 15874
rect 36036 15820 36260 15822
rect 35980 15810 36036 15820
rect 36204 15810 36260 15820
rect 36316 15876 36372 15886
rect 35868 15486 35870 15538
rect 35922 15486 35924 15538
rect 35868 15474 35924 15486
rect 35980 15652 36036 15662
rect 36316 15652 36372 15820
rect 35980 15538 36036 15596
rect 35980 15486 35982 15538
rect 36034 15486 36036 15538
rect 35980 15474 36036 15486
rect 36204 15596 36372 15652
rect 35196 14924 35460 14934
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35196 14858 35460 14868
rect 33516 13634 33684 13636
rect 33516 13582 33630 13634
rect 33682 13582 33684 13634
rect 33516 13580 33684 13582
rect 33404 13188 33460 13198
rect 33516 13188 33572 13580
rect 33628 13570 33684 13580
rect 33740 13916 34244 13972
rect 34972 14700 35084 14756
rect 35644 14756 35700 15148
rect 35756 15314 35812 15326
rect 35756 15262 35758 15314
rect 35810 15262 35812 15314
rect 35756 14980 35812 15262
rect 35980 15092 36036 15102
rect 35980 14980 36036 15036
rect 35756 14924 36036 14980
rect 35644 14700 35924 14756
rect 33404 13186 33572 13188
rect 33404 13134 33406 13186
rect 33458 13134 33572 13186
rect 33404 13132 33572 13134
rect 33740 13186 33796 13916
rect 34300 13860 34356 13870
rect 34300 13746 34356 13804
rect 34972 13860 35028 14700
rect 35084 14690 35140 14700
rect 35532 14644 35588 14654
rect 35532 14642 35812 14644
rect 35532 14590 35534 14642
rect 35586 14590 35812 14642
rect 35532 14588 35812 14590
rect 35532 14578 35588 14588
rect 35756 14532 35812 14588
rect 35756 14466 35812 14476
rect 35532 14420 35588 14430
rect 34300 13694 34302 13746
rect 34354 13694 34356 13746
rect 34300 13682 34356 13694
rect 34524 13748 34580 13758
rect 34860 13748 34916 13758
rect 34524 13746 34916 13748
rect 34524 13694 34526 13746
rect 34578 13694 34862 13746
rect 34914 13694 34916 13746
rect 34524 13692 34916 13694
rect 34524 13682 34580 13692
rect 34860 13682 34916 13692
rect 33740 13134 33742 13186
rect 33794 13134 33796 13186
rect 33404 13122 33460 13132
rect 33740 13122 33796 13134
rect 34076 13636 34132 13646
rect 33180 13074 33348 13076
rect 33180 13022 33182 13074
rect 33234 13022 33348 13074
rect 33180 13020 33348 13022
rect 33180 13010 33236 13020
rect 33964 12852 34020 12862
rect 33292 12404 33348 12414
rect 33292 12310 33348 12348
rect 33964 12178 34020 12796
rect 34076 12404 34132 13580
rect 34972 13524 35028 13804
rect 35084 14308 35140 14318
rect 35084 13970 35140 14252
rect 35084 13918 35086 13970
rect 35138 13918 35140 13970
rect 35084 13748 35140 13918
rect 35196 13860 35252 13870
rect 35196 13766 35252 13804
rect 35084 13682 35140 13692
rect 34972 13468 35140 13524
rect 35084 13188 35140 13468
rect 35196 13356 35460 13366
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35196 13290 35460 13300
rect 35084 13132 35364 13188
rect 35308 13074 35364 13132
rect 35308 13022 35310 13074
rect 35362 13022 35364 13074
rect 35308 13010 35364 13022
rect 34188 12852 34244 12862
rect 34188 12758 34244 12796
rect 34748 12852 34804 12862
rect 34748 12850 34916 12852
rect 34748 12798 34750 12850
rect 34802 12798 34916 12850
rect 34748 12796 34916 12798
rect 34748 12786 34804 12796
rect 34636 12740 34692 12750
rect 34300 12738 34692 12740
rect 34300 12686 34638 12738
rect 34690 12686 34692 12738
rect 34300 12684 34692 12686
rect 34076 12348 34244 12404
rect 33964 12126 33966 12178
rect 34018 12126 34020 12178
rect 33964 12114 34020 12126
rect 33628 12068 33684 12078
rect 33628 12066 33796 12068
rect 33628 12014 33630 12066
rect 33682 12014 33796 12066
rect 33628 12012 33796 12014
rect 33628 12002 33684 12012
rect 31948 10724 32004 11228
rect 32508 11228 32676 11284
rect 32844 11394 33012 11396
rect 32844 11342 32958 11394
rect 33010 11342 33012 11394
rect 32844 11340 33012 11342
rect 32396 11170 32452 11182
rect 32396 11118 32398 11170
rect 32450 11118 32452 11170
rect 31948 10722 32116 10724
rect 31948 10670 31950 10722
rect 32002 10670 32116 10722
rect 31948 10668 32116 10670
rect 31948 10658 32004 10668
rect 31612 10498 31668 10510
rect 31612 10446 31614 10498
rect 31666 10446 31668 10498
rect 31332 9772 31444 9828
rect 31500 10386 31556 10398
rect 31500 10334 31502 10386
rect 31554 10334 31556 10386
rect 31276 9734 31332 9772
rect 31500 8370 31556 10334
rect 31612 10050 31668 10446
rect 31612 9998 31614 10050
rect 31666 9998 31668 10050
rect 31612 9986 31668 9998
rect 32060 9826 32116 10668
rect 32396 10164 32452 11118
rect 32508 10834 32564 11228
rect 32844 10948 32900 11340
rect 32956 11330 33012 11340
rect 33180 11956 33236 11966
rect 33180 11282 33236 11900
rect 33180 11230 33182 11282
rect 33234 11230 33236 11282
rect 33180 11218 33236 11230
rect 33628 11394 33684 11406
rect 33628 11342 33630 11394
rect 33682 11342 33684 11394
rect 32508 10782 32510 10834
rect 32562 10782 32564 10834
rect 32508 10770 32564 10782
rect 32620 10892 32900 10948
rect 32396 10098 32452 10108
rect 32060 9774 32062 9826
rect 32114 9774 32116 9826
rect 32060 9762 32116 9774
rect 32508 9828 32564 9838
rect 32508 9734 32564 9772
rect 32620 9266 32676 10892
rect 33068 10724 33124 10734
rect 33068 10630 33124 10668
rect 33404 10610 33460 10622
rect 33404 10558 33406 10610
rect 33458 10558 33460 10610
rect 32620 9214 32622 9266
rect 32674 9214 32676 9266
rect 32620 9202 32676 9214
rect 33180 9940 33236 9950
rect 33180 9826 33236 9884
rect 33180 9774 33182 9826
rect 33234 9774 33236 9826
rect 31612 9042 31668 9054
rect 31612 8990 31614 9042
rect 31666 8990 31668 9042
rect 31612 8932 31668 8990
rect 31612 8866 31668 8876
rect 33180 8932 33236 9774
rect 33404 9716 33460 10558
rect 33628 10052 33684 11342
rect 33740 11396 33796 12012
rect 33740 10500 33796 11340
rect 33740 10434 33796 10444
rect 34188 10612 34244 12348
rect 34300 11506 34356 12684
rect 34636 12674 34692 12684
rect 34748 12178 34804 12190
rect 34748 12126 34750 12178
rect 34802 12126 34804 12178
rect 34748 11956 34804 12126
rect 34748 11890 34804 11900
rect 34300 11454 34302 11506
rect 34354 11454 34356 11506
rect 34300 11442 34356 11454
rect 34300 10612 34356 10622
rect 34188 10610 34356 10612
rect 34188 10558 34302 10610
rect 34354 10558 34356 10610
rect 34188 10556 34356 10558
rect 33516 9996 33684 10052
rect 34076 10386 34132 10398
rect 34076 10334 34078 10386
rect 34130 10334 34132 10386
rect 33516 9940 33572 9996
rect 33516 9874 33572 9884
rect 33628 9828 33684 9838
rect 33404 9660 33572 9716
rect 33180 8866 33236 8876
rect 31500 8318 31502 8370
rect 31554 8318 31556 8370
rect 31500 8306 31556 8318
rect 30828 4562 30996 4564
rect 30828 4510 30830 4562
rect 30882 4510 30996 4562
rect 30828 4508 30996 4510
rect 30828 4498 30884 4508
rect 31388 4228 31444 4238
rect 31388 4226 31556 4228
rect 31388 4174 31390 4226
rect 31442 4174 31556 4226
rect 31388 4172 31556 4174
rect 31388 4162 31444 4172
rect 31500 3554 31556 4172
rect 31500 3502 31502 3554
rect 31554 3502 31556 3554
rect 31276 3444 31332 3454
rect 30604 3442 31332 3444
rect 30604 3390 31278 3442
rect 31330 3390 31332 3442
rect 30604 3388 31332 3390
rect 31276 3378 31332 3388
rect 31500 2548 31556 3502
rect 30940 2492 31556 2548
rect 32956 3444 33012 3482
rect 33180 3444 33236 3454
rect 32956 3442 33236 3444
rect 32956 3390 32958 3442
rect 33010 3390 33182 3442
rect 33234 3390 33236 3442
rect 32956 3388 33236 3390
rect 30940 800 30996 2492
rect 32956 800 33012 3388
rect 33180 3378 33236 3388
rect 33516 3442 33572 9660
rect 33628 8370 33684 9772
rect 33852 9714 33908 9726
rect 33852 9662 33854 9714
rect 33906 9662 33908 9714
rect 33852 8484 33908 9662
rect 33964 8484 34020 8494
rect 33852 8482 34020 8484
rect 33852 8430 33966 8482
rect 34018 8430 34020 8482
rect 33852 8428 34020 8430
rect 33964 8418 34020 8428
rect 33628 8318 33630 8370
rect 33682 8318 33684 8370
rect 33628 8306 33684 8318
rect 34076 8370 34132 10334
rect 34188 9828 34244 10556
rect 34300 10546 34356 10556
rect 34748 10610 34804 10622
rect 34748 10558 34750 10610
rect 34802 10558 34804 10610
rect 34748 10500 34804 10558
rect 34748 10434 34804 10444
rect 34860 10388 34916 12796
rect 35308 12068 35364 12078
rect 35308 11974 35364 12012
rect 35196 11788 35460 11798
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35196 11722 35460 11732
rect 35532 10612 35588 14364
rect 35868 13636 35924 14700
rect 36204 14530 36260 15596
rect 36316 15316 36372 15326
rect 36316 14754 36372 15260
rect 36316 14702 36318 14754
rect 36370 14702 36372 14754
rect 36316 14690 36372 14702
rect 36428 15314 36484 15326
rect 36428 15262 36430 15314
rect 36482 15262 36484 15314
rect 36428 14756 36484 15262
rect 36764 15316 36820 16044
rect 36876 15538 36932 19292
rect 36988 18116 37044 19516
rect 37100 19460 37156 19470
rect 37436 19460 37492 19470
rect 37100 19366 37156 19404
rect 37212 19458 37492 19460
rect 37212 19406 37438 19458
rect 37490 19406 37492 19458
rect 37212 19404 37492 19406
rect 37212 19234 37268 19404
rect 37436 19394 37492 19404
rect 37212 19182 37214 19234
rect 37266 19182 37268 19234
rect 37212 19170 37268 19182
rect 37100 19124 37156 19134
rect 37100 19030 37156 19068
rect 37324 18564 37380 18574
rect 37324 18470 37380 18508
rect 36988 17556 37044 18060
rect 37100 18450 37156 18462
rect 37100 18398 37102 18450
rect 37154 18398 37156 18450
rect 37100 17892 37156 18398
rect 37212 18340 37268 18350
rect 37212 18246 37268 18284
rect 37548 18116 37604 20524
rect 37660 20486 37716 20524
rect 37996 20802 38052 20814
rect 37996 20750 37998 20802
rect 38050 20750 38052 20802
rect 37884 19458 37940 19470
rect 37884 19406 37886 19458
rect 37938 19406 37940 19458
rect 37660 19348 37716 19358
rect 37660 19254 37716 19292
rect 37884 18564 37940 19406
rect 37996 18676 38052 20750
rect 38108 20244 38164 20254
rect 38668 20244 38724 20254
rect 38780 20244 38836 23492
rect 39004 22484 39060 26350
rect 39116 26290 39172 26908
rect 39116 26238 39118 26290
rect 39170 26238 39172 26290
rect 39116 26226 39172 26238
rect 39340 26908 39396 26918
rect 39452 26910 39454 26962
rect 39506 26910 39508 26962
rect 39452 26898 39508 26910
rect 40012 27074 40068 28028
rect 40348 27860 40404 27870
rect 40348 27746 40404 27804
rect 40348 27694 40350 27746
rect 40402 27694 40404 27746
rect 40348 27682 40404 27694
rect 40012 27022 40014 27074
rect 40066 27022 40068 27074
rect 39340 26404 39396 26852
rect 40012 26852 40068 27022
rect 40348 27076 40404 27086
rect 40348 26982 40404 27020
rect 40012 26786 40068 26796
rect 39340 25060 39396 26348
rect 39900 25618 39956 25630
rect 39900 25566 39902 25618
rect 39954 25566 39956 25618
rect 39900 25060 39956 25566
rect 40236 25394 40292 25406
rect 40236 25342 40238 25394
rect 40290 25342 40292 25394
rect 40236 25284 40292 25342
rect 40236 25218 40292 25228
rect 40348 25282 40404 25294
rect 40348 25230 40350 25282
rect 40402 25230 40404 25282
rect 39340 25004 39956 25060
rect 39116 24052 39172 24062
rect 39116 23958 39172 23996
rect 39228 23940 39284 23950
rect 39228 23378 39284 23884
rect 39228 23326 39230 23378
rect 39282 23326 39284 23378
rect 39228 23314 39284 23326
rect 38108 19346 38164 20188
rect 38332 20242 38836 20244
rect 38332 20190 38670 20242
rect 38722 20190 38836 20242
rect 38332 20188 38836 20190
rect 38892 21476 38948 21486
rect 38220 19906 38276 19918
rect 38220 19854 38222 19906
rect 38274 19854 38276 19906
rect 38220 19458 38276 19854
rect 38220 19406 38222 19458
rect 38274 19406 38276 19458
rect 38220 19394 38276 19406
rect 38108 19294 38110 19346
rect 38162 19294 38164 19346
rect 38108 19236 38164 19294
rect 38108 19170 38164 19180
rect 37996 18620 38164 18676
rect 37884 18508 38052 18564
rect 37772 18452 37828 18462
rect 37772 18450 37940 18452
rect 37772 18398 37774 18450
rect 37826 18398 37940 18450
rect 37772 18396 37940 18398
rect 37772 18386 37828 18396
rect 37436 18060 37604 18116
rect 37660 18340 37716 18350
rect 37660 18116 37716 18284
rect 37660 18060 37828 18116
rect 37436 17892 37492 18060
rect 37100 17836 37268 17892
rect 37436 17836 37604 17892
rect 36988 17490 37044 17500
rect 37100 17666 37156 17678
rect 37100 17614 37102 17666
rect 37154 17614 37156 17666
rect 36988 17108 37044 17118
rect 36988 16994 37044 17052
rect 36988 16942 36990 16994
rect 37042 16942 37044 16994
rect 36988 16930 37044 16942
rect 37100 16884 37156 17614
rect 37212 16996 37268 17836
rect 37212 16930 37268 16940
rect 37324 17556 37380 17566
rect 37100 16818 37156 16828
rect 37100 16212 37156 16222
rect 37324 16212 37380 17500
rect 37100 16210 37380 16212
rect 37100 16158 37102 16210
rect 37154 16158 37380 16210
rect 37100 16156 37380 16158
rect 37100 16146 37156 16156
rect 36876 15486 36878 15538
rect 36930 15486 36932 15538
rect 36876 15474 36932 15486
rect 37324 15876 37380 15886
rect 36764 15260 36932 15316
rect 36876 15148 36932 15260
rect 36876 15092 37156 15148
rect 36876 14756 36932 14766
rect 36428 14754 36932 14756
rect 36428 14702 36878 14754
rect 36930 14702 36932 14754
rect 36428 14700 36932 14702
rect 36876 14690 36932 14700
rect 36204 14478 36206 14530
rect 36258 14478 36260 14530
rect 36204 13972 36260 14478
rect 36988 14420 37044 14430
rect 36988 14326 37044 14364
rect 36316 14308 36372 14318
rect 36316 14306 36484 14308
rect 36316 14254 36318 14306
rect 36370 14254 36484 14306
rect 36316 14252 36484 14254
rect 36316 14242 36372 14252
rect 36316 13972 36372 13982
rect 36204 13970 36372 13972
rect 36204 13918 36318 13970
rect 36370 13918 36372 13970
rect 36204 13916 36372 13918
rect 36316 13906 36372 13916
rect 35868 13634 36036 13636
rect 35868 13582 35870 13634
rect 35922 13582 36036 13634
rect 35868 13580 36036 13582
rect 35868 13570 35924 13580
rect 35868 13076 35924 13086
rect 35868 12982 35924 13020
rect 35980 12852 36036 13580
rect 36428 12962 36484 14252
rect 37100 14084 37156 15092
rect 37324 14420 37380 15820
rect 37324 14354 37380 14364
rect 37436 14418 37492 14430
rect 37436 14366 37438 14418
rect 37490 14366 37492 14418
rect 37212 14308 37268 14318
rect 37212 14214 37268 14252
rect 37436 14084 37492 14366
rect 37100 14028 37492 14084
rect 36764 13860 36820 13870
rect 36764 13766 36820 13804
rect 36428 12910 36430 12962
rect 36482 12910 36484 12962
rect 36316 12852 36372 12862
rect 35980 12796 36148 12852
rect 35756 12068 35812 12078
rect 35756 10724 35812 12012
rect 35756 10630 35812 10668
rect 35644 10612 35700 10622
rect 35532 10610 35644 10612
rect 35532 10558 35534 10610
rect 35586 10558 35644 10610
rect 35532 10556 35644 10558
rect 35532 10546 35588 10556
rect 34972 10388 35028 10398
rect 34860 10332 34972 10388
rect 34972 10322 35028 10332
rect 35196 10220 35460 10230
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35196 10154 35460 10164
rect 35644 10164 35700 10556
rect 35644 10108 36036 10164
rect 35980 9938 36036 10108
rect 35980 9886 35982 9938
rect 36034 9886 36036 9938
rect 35980 9874 36036 9886
rect 34188 9762 34244 9772
rect 36092 9268 36148 12796
rect 36204 12178 36260 12190
rect 36204 12126 36206 12178
rect 36258 12126 36260 12178
rect 36204 12068 36260 12126
rect 36204 12002 36260 12012
rect 36204 10388 36260 10398
rect 36204 10294 36260 10332
rect 36316 9940 36372 12796
rect 36428 11506 36484 12910
rect 36764 13076 36820 13086
rect 36764 12178 36820 13020
rect 36764 12126 36766 12178
rect 36818 12126 36820 12178
rect 36428 11454 36430 11506
rect 36482 11454 36484 11506
rect 36428 11442 36484 11454
rect 36540 11954 36596 11966
rect 36540 11902 36542 11954
rect 36594 11902 36596 11954
rect 36428 9940 36484 9950
rect 36316 9884 36428 9940
rect 36428 9846 36484 9884
rect 36204 9268 36260 9278
rect 36092 9212 36204 9268
rect 36204 9202 36260 9212
rect 36316 8932 36372 8942
rect 36316 8838 36372 8876
rect 36540 8708 36596 11902
rect 36764 11788 36820 12126
rect 36652 11732 36820 11788
rect 37100 12962 37156 12974
rect 37100 12910 37102 12962
rect 37154 12910 37156 12962
rect 37100 11732 37156 12910
rect 37212 12404 37268 14028
rect 37436 13858 37492 13870
rect 37436 13806 37438 13858
rect 37490 13806 37492 13858
rect 37324 13746 37380 13758
rect 37324 13694 37326 13746
rect 37378 13694 37380 13746
rect 37324 13524 37380 13694
rect 37436 13748 37492 13806
rect 37436 13682 37492 13692
rect 37324 12852 37380 13468
rect 37324 12786 37380 12796
rect 37436 13522 37492 13534
rect 37436 13470 37438 13522
rect 37490 13470 37492 13522
rect 37324 12404 37380 12414
rect 37212 12348 37324 12404
rect 37324 12338 37380 12348
rect 37436 12180 37492 13470
rect 37436 12114 37492 12124
rect 37324 12066 37380 12078
rect 37324 12014 37326 12066
rect 37378 12014 37380 12066
rect 37212 11732 37268 11742
rect 36652 10610 36708 11732
rect 37100 11676 37212 11732
rect 37212 11666 37268 11676
rect 37324 11508 37380 12014
rect 37212 11396 37268 11406
rect 37100 11394 37268 11396
rect 37100 11342 37214 11394
rect 37266 11342 37268 11394
rect 37100 11340 37268 11342
rect 36988 11284 37044 11294
rect 36652 10558 36654 10610
rect 36706 10558 36708 10610
rect 36652 10546 36708 10558
rect 36764 11282 37044 11284
rect 36764 11230 36990 11282
rect 37042 11230 37044 11282
rect 36764 11228 37044 11230
rect 36764 10724 36820 11228
rect 36988 11218 37044 11228
rect 36764 10610 36820 10668
rect 36764 10558 36766 10610
rect 36818 10558 36820 10610
rect 36764 10546 36820 10558
rect 37100 11172 37156 11340
rect 37212 11330 37268 11340
rect 36988 9940 37044 9950
rect 36988 9826 37044 9884
rect 36988 9774 36990 9826
rect 37042 9774 37044 9826
rect 36988 9762 37044 9774
rect 35196 8652 35460 8662
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35196 8586 35460 8596
rect 36316 8652 36596 8708
rect 36988 8932 37044 8942
rect 34076 8318 34078 8370
rect 34130 8318 34132 8370
rect 34076 8306 34132 8318
rect 36316 8370 36372 8652
rect 36316 8318 36318 8370
rect 36370 8318 36372 8370
rect 36316 8306 36372 8318
rect 36988 8258 37044 8876
rect 36988 8206 36990 8258
rect 37042 8206 37044 8258
rect 36988 8194 37044 8206
rect 36428 8148 36484 8158
rect 36428 8054 36484 8092
rect 37100 7364 37156 11116
rect 37212 10612 37268 10622
rect 37212 10518 37268 10556
rect 37324 9940 37380 11452
rect 37436 9940 37492 9950
rect 37324 9938 37492 9940
rect 37324 9886 37438 9938
rect 37490 9886 37492 9938
rect 37324 9884 37492 9886
rect 37436 9874 37492 9884
rect 37436 7364 37492 7374
rect 37100 7362 37492 7364
rect 37100 7310 37438 7362
rect 37490 7310 37492 7362
rect 37100 7308 37492 7310
rect 37436 7298 37492 7308
rect 35196 7084 35460 7094
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35196 7018 35460 7028
rect 35196 5516 35460 5526
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35196 5450 35460 5460
rect 34860 5012 34916 5022
rect 33516 3390 33518 3442
rect 33570 3390 33572 3442
rect 33516 3378 33572 3390
rect 33628 4226 33684 4238
rect 33628 4174 33630 4226
rect 33682 4174 33684 4226
rect 33628 3556 33684 4174
rect 34300 4226 34356 4238
rect 34300 4174 34302 4226
rect 34354 4174 34356 4226
rect 33852 3556 33908 3566
rect 33628 3554 33908 3556
rect 33628 3502 33854 3554
rect 33906 3502 33908 3554
rect 33628 3500 33908 3502
rect 33628 800 33684 3500
rect 33852 3490 33908 3500
rect 34300 3556 34356 4174
rect 34524 3556 34580 3566
rect 34300 3554 34580 3556
rect 34300 3502 34526 3554
rect 34578 3502 34580 3554
rect 34300 3500 34580 3502
rect 34188 3444 34244 3482
rect 34188 3378 34244 3388
rect 34300 800 34356 3500
rect 34524 3490 34580 3500
rect 34860 3442 34916 4956
rect 36428 4228 36484 4238
rect 37100 4228 37156 4238
rect 36428 4226 36708 4228
rect 36428 4174 36430 4226
rect 36482 4174 36708 4226
rect 36428 4172 36708 4174
rect 36428 4162 36484 4172
rect 35196 3948 35460 3958
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35196 3882 35460 3892
rect 36652 3554 36708 4172
rect 37100 4226 37380 4228
rect 37100 4174 37102 4226
rect 37154 4174 37380 4226
rect 37100 4172 37380 4174
rect 37100 4162 37156 4172
rect 36652 3502 36654 3554
rect 36706 3502 36708 3554
rect 34860 3390 34862 3442
rect 34914 3390 34916 3442
rect 34860 3378 34916 3390
rect 35532 3444 35588 3454
rect 35980 3444 36036 3454
rect 35532 3442 36036 3444
rect 35532 3390 35534 3442
rect 35586 3390 35982 3442
rect 36034 3390 36036 3442
rect 35532 3388 36036 3390
rect 35532 3378 35588 3388
rect 35644 800 35700 3388
rect 35980 3378 36036 3388
rect 36316 3444 36372 3482
rect 36316 3378 36372 3388
rect 36652 2548 36708 3502
rect 37324 3554 37380 4172
rect 37324 3502 37326 3554
rect 37378 3502 37380 3554
rect 36988 3444 37044 3454
rect 37212 3444 37268 3454
rect 36988 3442 37212 3444
rect 36988 3390 36990 3442
rect 37042 3390 37212 3442
rect 36988 3388 37212 3390
rect 36988 3378 37044 3388
rect 37212 3378 37268 3388
rect 37324 2548 37380 3502
rect 37548 3444 37604 17836
rect 37772 17778 37828 18060
rect 37884 18004 37940 18396
rect 37884 17938 37940 17948
rect 37772 17726 37774 17778
rect 37826 17726 37828 17778
rect 37772 17714 37828 17726
rect 37660 17108 37716 17118
rect 37660 16884 37716 17052
rect 37660 16882 37828 16884
rect 37660 16830 37662 16882
rect 37714 16830 37828 16882
rect 37660 16828 37828 16830
rect 37660 16818 37716 16828
rect 37772 15988 37828 16828
rect 37884 16772 37940 16782
rect 37996 16772 38052 18508
rect 38108 17892 38164 18620
rect 38332 18338 38388 20188
rect 38668 20178 38724 20188
rect 38556 19124 38612 19134
rect 38556 19030 38612 19068
rect 38332 18286 38334 18338
rect 38386 18286 38388 18338
rect 38332 18116 38388 18286
rect 38332 18050 38388 18060
rect 38668 18450 38724 18462
rect 38668 18398 38670 18450
rect 38722 18398 38724 18450
rect 38108 17836 38500 17892
rect 38332 16772 38388 16782
rect 37884 16770 38388 16772
rect 37884 16718 37886 16770
rect 37938 16718 38334 16770
rect 38386 16718 38388 16770
rect 37884 16716 38388 16718
rect 37884 16706 37940 16716
rect 37996 16098 38052 16716
rect 38332 16706 38388 16716
rect 38444 16548 38500 17836
rect 38668 17780 38724 18398
rect 38892 18228 38948 21420
rect 39004 20802 39060 22428
rect 39564 21586 39620 25004
rect 40348 24052 40404 25230
rect 40460 24164 40516 28700
rect 41132 28756 41188 28766
rect 40796 28642 40852 28654
rect 40796 28590 40798 28642
rect 40850 28590 40852 28642
rect 40796 26908 40852 28590
rect 41020 28644 41076 28654
rect 40908 28084 40964 28094
rect 40908 27990 40964 28028
rect 40572 26852 40852 26908
rect 40572 25506 40628 26852
rect 41020 25620 41076 28588
rect 40572 25454 40574 25506
rect 40626 25454 40628 25506
rect 40572 25442 40628 25454
rect 40684 25564 41076 25620
rect 40460 24098 40516 24108
rect 40348 23986 40404 23996
rect 40236 23940 40292 23950
rect 40236 23378 40292 23884
rect 40236 23326 40238 23378
rect 40290 23326 40292 23378
rect 40236 23314 40292 23326
rect 39788 23268 39844 23278
rect 39788 23154 39844 23212
rect 39788 23102 39790 23154
rect 39842 23102 39844 23154
rect 39788 21700 39844 23102
rect 40684 22932 40740 25564
rect 41132 25508 41188 28700
rect 41356 28642 41412 28654
rect 41356 28590 41358 28642
rect 41410 28590 41412 28642
rect 41244 27860 41300 27870
rect 41244 27766 41300 27804
rect 41356 27748 41412 28590
rect 41804 28642 41860 28654
rect 41804 28590 41806 28642
rect 41858 28590 41860 28642
rect 41692 27970 41748 27982
rect 41692 27918 41694 27970
rect 41746 27918 41748 27970
rect 41692 27860 41748 27918
rect 41692 27794 41748 27804
rect 41580 27748 41636 27758
rect 41356 27746 41636 27748
rect 41356 27694 41582 27746
rect 41634 27694 41636 27746
rect 41356 27692 41636 27694
rect 41580 27682 41636 27692
rect 40460 22876 40740 22932
rect 40796 25452 41188 25508
rect 41244 27636 41300 27646
rect 41244 25618 41300 27580
rect 41580 27188 41636 27198
rect 41580 27094 41636 27132
rect 41804 27074 41860 28590
rect 42476 28196 42532 30940
rect 42588 30994 42644 31006
rect 42588 30942 42590 30994
rect 42642 30942 42644 30994
rect 42588 30436 42644 30942
rect 42812 30994 42868 31006
rect 42812 30942 42814 30994
rect 42866 30942 42868 30994
rect 42700 30436 42756 30446
rect 42588 30434 42756 30436
rect 42588 30382 42702 30434
rect 42754 30382 42756 30434
rect 42588 30380 42756 30382
rect 42700 29988 42756 30380
rect 42700 28866 42756 29932
rect 42700 28814 42702 28866
rect 42754 28814 42756 28866
rect 42700 28802 42756 28814
rect 42812 29876 42868 30942
rect 42924 30772 42980 31836
rect 43148 31826 43204 31836
rect 43260 32450 43316 32462
rect 43260 32398 43262 32450
rect 43314 32398 43316 32450
rect 43260 31780 43316 32398
rect 43260 31714 43316 31724
rect 43484 31444 43540 33068
rect 43708 32788 43764 32798
rect 43708 32562 43764 32732
rect 43708 32510 43710 32562
rect 43762 32510 43764 32562
rect 43708 32498 43764 32510
rect 44156 32450 44212 33068
rect 44156 32398 44158 32450
rect 44210 32398 44212 32450
rect 44156 32386 44212 32398
rect 44044 31892 44100 31902
rect 44044 31798 44100 31836
rect 42924 30706 42980 30716
rect 43036 31388 43540 31444
rect 42812 28756 42868 29820
rect 42924 28756 42980 28766
rect 42812 28754 42980 28756
rect 42812 28702 42926 28754
rect 42978 28702 42980 28754
rect 42812 28700 42980 28702
rect 42924 28690 42980 28700
rect 42476 28130 42532 28140
rect 42700 28644 42756 28654
rect 42364 27746 42420 27758
rect 42364 27694 42366 27746
rect 42418 27694 42420 27746
rect 41804 27022 41806 27074
rect 41858 27022 41860 27074
rect 41804 27010 41860 27022
rect 41916 27634 41972 27646
rect 41916 27582 41918 27634
rect 41970 27582 41972 27634
rect 41916 27076 41972 27582
rect 42140 27076 42196 27086
rect 42364 27076 42420 27694
rect 41916 27020 42140 27076
rect 42196 27020 42420 27076
rect 42476 27188 42532 27198
rect 42476 27074 42532 27132
rect 42476 27022 42478 27074
rect 42530 27022 42532 27074
rect 42140 26982 42196 27020
rect 42476 27010 42532 27022
rect 42700 27074 42756 28588
rect 43036 28532 43092 31388
rect 43148 30996 43204 31006
rect 43148 30660 43204 30940
rect 43148 30594 43204 30604
rect 43260 30772 43316 30782
rect 43260 30436 43316 30716
rect 42700 27022 42702 27074
rect 42754 27022 42756 27074
rect 42700 27010 42756 27022
rect 42812 28476 43092 28532
rect 43148 30380 43316 30436
rect 42812 26908 42868 28476
rect 43148 28420 43204 30380
rect 43260 30212 43316 30222
rect 43260 30118 43316 30156
rect 42028 26852 42084 26862
rect 42028 26758 42084 26796
rect 42252 26852 42868 26908
rect 42924 28364 43204 28420
rect 43372 30098 43428 30110
rect 43372 30046 43374 30098
rect 43426 30046 43428 30098
rect 42924 26962 42980 28364
rect 43036 27300 43092 27310
rect 43372 27300 43428 30046
rect 44380 29986 44436 29998
rect 44380 29934 44382 29986
rect 44434 29934 44436 29986
rect 44380 29652 44436 29934
rect 44380 29586 44436 29596
rect 44268 29204 44324 29214
rect 43484 28642 43540 28654
rect 43484 28590 43486 28642
rect 43538 28590 43540 28642
rect 43484 28420 43540 28590
rect 43484 28354 43540 28364
rect 43596 28642 43652 28654
rect 43596 28590 43598 28642
rect 43650 28590 43652 28642
rect 43036 27298 43428 27300
rect 43036 27246 43038 27298
rect 43090 27246 43428 27298
rect 43036 27244 43428 27246
rect 43484 28196 43540 28206
rect 43484 27300 43540 28140
rect 43036 27234 43092 27244
rect 43484 27188 43540 27244
rect 43372 27132 43540 27188
rect 43260 27076 43316 27086
rect 43260 26982 43316 27020
rect 42924 26910 42926 26962
rect 42978 26910 42980 26962
rect 42924 26898 42980 26910
rect 43372 26962 43428 27132
rect 43596 27074 43652 28590
rect 44268 28530 44324 29148
rect 44268 28478 44270 28530
rect 44322 28478 44324 28530
rect 44268 28466 44324 28478
rect 44044 28420 44100 28430
rect 43932 27300 43988 27310
rect 43932 27186 43988 27244
rect 43932 27134 43934 27186
rect 43986 27134 43988 27186
rect 43932 27122 43988 27134
rect 43596 27022 43598 27074
rect 43650 27022 43652 27074
rect 43596 27010 43652 27022
rect 43372 26910 43374 26962
rect 43426 26910 43428 26962
rect 43372 26898 43428 26910
rect 41244 25566 41246 25618
rect 41298 25566 41300 25618
rect 40460 22482 40516 22876
rect 40796 22820 40852 25452
rect 41020 25284 41076 25294
rect 41076 25228 41188 25284
rect 41020 25190 41076 25228
rect 40908 23154 40964 23166
rect 40908 23102 40910 23154
rect 40962 23102 40964 23154
rect 40908 22932 40964 23102
rect 40908 22866 40964 22876
rect 40460 22430 40462 22482
rect 40514 22430 40516 22482
rect 40124 21812 40180 21822
rect 40124 21718 40180 21756
rect 39564 21534 39566 21586
rect 39618 21534 39620 21586
rect 39564 21522 39620 21534
rect 39676 21698 39844 21700
rect 39676 21646 39790 21698
rect 39842 21646 39844 21698
rect 39676 21644 39844 21646
rect 39676 21364 39732 21644
rect 39788 21634 39844 21644
rect 39004 20750 39006 20802
rect 39058 20750 39060 20802
rect 39004 20738 39060 20750
rect 39564 21308 39732 21364
rect 40012 21588 40068 21598
rect 39564 20802 39620 21308
rect 39564 20750 39566 20802
rect 39618 20750 39620 20802
rect 39564 20738 39620 20750
rect 40012 20802 40068 21532
rect 40460 21588 40516 22430
rect 40460 21522 40516 21532
rect 40572 22764 40852 22820
rect 40236 21474 40292 21486
rect 40236 21422 40238 21474
rect 40290 21422 40292 21474
rect 40236 21026 40292 21422
rect 40236 20974 40238 21026
rect 40290 20974 40292 21026
rect 40236 20962 40292 20974
rect 40012 20750 40014 20802
rect 40066 20750 40068 20802
rect 40012 20738 40068 20750
rect 40348 20804 40404 20814
rect 39452 20132 39508 20142
rect 39676 20132 39732 20142
rect 40012 20132 40068 20142
rect 39508 20130 39732 20132
rect 39508 20078 39678 20130
rect 39730 20078 39732 20130
rect 39508 20076 39732 20078
rect 39452 20038 39508 20076
rect 39676 20066 39732 20076
rect 39900 20130 40068 20132
rect 39900 20078 40014 20130
rect 40066 20078 40068 20130
rect 39900 20076 40068 20078
rect 39900 19796 39956 20076
rect 40012 20066 40068 20076
rect 39340 19234 39396 19246
rect 39340 19182 39342 19234
rect 39394 19182 39396 19234
rect 39004 19010 39060 19022
rect 39004 18958 39006 19010
rect 39058 18958 39060 19010
rect 39004 18452 39060 18958
rect 39116 18452 39172 18462
rect 39004 18396 39116 18452
rect 39116 18358 39172 18396
rect 39340 18452 39396 19182
rect 38892 18172 39060 18228
rect 37996 16046 37998 16098
rect 38050 16046 38052 16098
rect 37996 16034 38052 16046
rect 38220 16492 38500 16548
rect 38556 16884 38612 16894
rect 37884 15988 37940 15998
rect 37772 15986 37940 15988
rect 37772 15934 37886 15986
rect 37938 15934 37940 15986
rect 37772 15932 37940 15934
rect 37884 15922 37940 15932
rect 37660 15874 37716 15886
rect 37660 15822 37662 15874
rect 37714 15822 37716 15874
rect 37660 15314 37716 15822
rect 37660 15262 37662 15314
rect 37714 15262 37716 15314
rect 37660 15250 37716 15262
rect 37884 15316 37940 15326
rect 37884 15202 37940 15260
rect 37884 15150 37886 15202
rect 37938 15150 37940 15202
rect 37884 15138 37940 15150
rect 38220 15148 38276 16492
rect 38332 16322 38388 16334
rect 38332 16270 38334 16322
rect 38386 16270 38388 16322
rect 38332 15314 38388 16270
rect 38556 15988 38612 16828
rect 38668 16882 38724 17724
rect 38892 18004 38948 18014
rect 38892 17106 38948 17948
rect 38892 17054 38894 17106
rect 38946 17054 38948 17106
rect 38892 17042 38948 17054
rect 38668 16830 38670 16882
rect 38722 16830 38724 16882
rect 38668 16818 38724 16830
rect 38668 16658 38724 16670
rect 38668 16606 38670 16658
rect 38722 16606 38724 16658
rect 38668 16322 38724 16606
rect 38668 16270 38670 16322
rect 38722 16270 38724 16322
rect 38668 16258 38724 16270
rect 38444 15876 38500 15886
rect 38444 15782 38500 15820
rect 38332 15262 38334 15314
rect 38386 15262 38388 15314
rect 38332 15250 38388 15262
rect 38108 15090 38164 15102
rect 38220 15092 38500 15148
rect 38108 15038 38110 15090
rect 38162 15038 38164 15090
rect 37884 14980 37940 14990
rect 37884 14418 37940 14924
rect 38108 14532 38164 15038
rect 37884 14366 37886 14418
rect 37938 14366 37940 14418
rect 37884 14354 37940 14366
rect 37996 14530 38164 14532
rect 37996 14478 38110 14530
rect 38162 14478 38164 14530
rect 37996 14476 38164 14478
rect 37996 14420 38052 14476
rect 38108 14466 38164 14476
rect 38332 14532 38388 14542
rect 38332 14438 38388 14476
rect 37996 14196 38052 14364
rect 37884 14140 38052 14196
rect 38220 14306 38276 14318
rect 38444 14308 38500 15092
rect 38220 14254 38222 14306
rect 38274 14254 38276 14306
rect 37884 13746 37940 14140
rect 38220 13972 38276 14254
rect 38220 13906 38276 13916
rect 38332 14252 38500 14308
rect 38332 13748 38388 14252
rect 37884 13694 37886 13746
rect 37938 13694 37940 13746
rect 37884 13682 37940 13694
rect 38220 13692 38388 13748
rect 38444 13748 38500 13758
rect 37996 13636 38052 13646
rect 37660 13412 37716 13422
rect 37660 12068 37716 13356
rect 37884 13076 37940 13086
rect 37996 13076 38052 13580
rect 38108 13524 38164 13534
rect 38108 13430 38164 13468
rect 37884 13074 38052 13076
rect 37884 13022 37886 13074
rect 37938 13022 38052 13074
rect 37884 13020 38052 13022
rect 37884 13010 37940 13020
rect 37660 12002 37716 12012
rect 37772 12852 37828 12862
rect 37660 10500 37716 10510
rect 37660 10406 37716 10444
rect 37772 9492 37828 12796
rect 37772 9426 37828 9436
rect 37884 12178 37940 12190
rect 37884 12126 37886 12178
rect 37938 12126 37940 12178
rect 37772 8148 37828 8158
rect 37772 8054 37828 8092
rect 37772 4226 37828 4238
rect 37772 4174 37774 4226
rect 37826 4174 37828 4226
rect 37660 3444 37716 3454
rect 37548 3442 37716 3444
rect 37548 3390 37662 3442
rect 37714 3390 37716 3442
rect 37548 3388 37716 3390
rect 37660 3378 37716 3388
rect 37772 2548 37828 4174
rect 37884 3444 37940 12126
rect 38108 12068 38164 12078
rect 37996 11508 38052 11518
rect 37996 11394 38052 11452
rect 37996 11342 37998 11394
rect 38050 11342 38052 11394
rect 37996 11330 38052 11342
rect 38108 11394 38164 12012
rect 38108 11342 38110 11394
rect 38162 11342 38164 11394
rect 38108 11060 38164 11342
rect 38108 10994 38164 11004
rect 38220 9828 38276 13692
rect 38444 13654 38500 13692
rect 38332 12178 38388 12190
rect 38332 12126 38334 12178
rect 38386 12126 38388 12178
rect 38332 11284 38388 12126
rect 38556 11732 38612 15932
rect 39004 15426 39060 18172
rect 39228 18116 39284 18126
rect 39228 17108 39284 18060
rect 39116 16996 39172 17006
rect 39116 15538 39172 16940
rect 39228 16994 39284 17052
rect 39228 16942 39230 16994
rect 39282 16942 39284 16994
rect 39228 16930 39284 16942
rect 39340 16884 39396 18396
rect 39452 18562 39508 18574
rect 39452 18510 39454 18562
rect 39506 18510 39508 18562
rect 39452 16996 39508 18510
rect 39900 18562 39956 19740
rect 40236 19796 40292 19806
rect 40124 19124 40180 19134
rect 39900 18510 39902 18562
rect 39954 18510 39956 18562
rect 39900 18116 39956 18510
rect 40012 19122 40180 19124
rect 40012 19070 40126 19122
rect 40178 19070 40180 19122
rect 40012 19068 40180 19070
rect 40012 18340 40068 19068
rect 40124 19058 40180 19068
rect 40236 18788 40292 19740
rect 40124 18732 40236 18788
rect 40124 18674 40180 18732
rect 40236 18722 40292 18732
rect 40124 18622 40126 18674
rect 40178 18622 40180 18674
rect 40124 18610 40180 18622
rect 40348 18676 40404 20748
rect 40348 18582 40404 18620
rect 40236 18564 40292 18574
rect 40236 18450 40292 18508
rect 40236 18398 40238 18450
rect 40290 18398 40292 18450
rect 40236 18386 40292 18398
rect 40012 18274 40068 18284
rect 39900 18060 40068 18116
rect 39564 17780 39620 17790
rect 39900 17780 39956 17790
rect 39620 17778 39956 17780
rect 39620 17726 39902 17778
rect 39954 17726 39956 17778
rect 39620 17724 39956 17726
rect 39564 17714 39620 17724
rect 39900 17714 39956 17724
rect 40012 17556 40068 18060
rect 39900 17500 40068 17556
rect 40572 17556 40628 22764
rect 40796 22596 40852 22606
rect 40796 22372 40852 22540
rect 40796 22370 41076 22372
rect 40796 22318 40798 22370
rect 40850 22318 41076 22370
rect 40796 22316 41076 22318
rect 40796 22306 40852 22316
rect 40796 21924 40852 21934
rect 40684 20580 40740 20590
rect 40684 20486 40740 20524
rect 40796 19236 40852 21868
rect 41020 21924 41076 22316
rect 41020 21810 41076 21868
rect 41020 21758 41022 21810
rect 41074 21758 41076 21810
rect 41020 21746 41076 21758
rect 41132 20580 41188 25228
rect 41244 24724 41300 25566
rect 41468 24724 41524 24734
rect 41244 24722 41524 24724
rect 41244 24670 41470 24722
rect 41522 24670 41524 24722
rect 41244 24668 41524 24670
rect 41244 23828 41300 23838
rect 41244 23734 41300 23772
rect 41356 23154 41412 23166
rect 41356 23102 41358 23154
rect 41410 23102 41412 23154
rect 41244 22932 41300 22942
rect 41244 22482 41300 22876
rect 41244 22430 41246 22482
rect 41298 22430 41300 22482
rect 41244 22418 41300 22430
rect 41356 20916 41412 23102
rect 41468 23156 41524 24668
rect 41580 24722 41636 24734
rect 41580 24670 41582 24722
rect 41634 24670 41636 24722
rect 41580 23268 41636 24670
rect 41580 23202 41636 23212
rect 41692 24052 41748 24062
rect 41468 23090 41524 23100
rect 41692 22370 41748 23996
rect 42028 23938 42084 23950
rect 42028 23886 42030 23938
rect 42082 23886 42084 23938
rect 42028 23604 42084 23886
rect 42028 23538 42084 23548
rect 42140 23156 42196 23166
rect 42140 23062 42196 23100
rect 42140 22484 42196 22494
rect 42140 22390 42196 22428
rect 41692 22318 41694 22370
rect 41746 22318 41748 22370
rect 41692 22306 41748 22318
rect 41916 21924 41972 21934
rect 42252 21924 42308 26852
rect 42364 26292 42420 26302
rect 42364 24722 42420 26236
rect 43148 26292 43204 26302
rect 43148 26198 43204 26236
rect 43932 26290 43988 26302
rect 43932 26238 43934 26290
rect 43986 26238 43988 26290
rect 42364 24670 42366 24722
rect 42418 24670 42420 24722
rect 42364 24658 42420 24670
rect 42700 26180 42756 26190
rect 42700 24610 42756 26124
rect 42700 24558 42702 24610
rect 42754 24558 42756 24610
rect 42588 23716 42644 23726
rect 41468 21812 41524 21822
rect 41468 21718 41524 21756
rect 41916 21810 41972 21868
rect 41916 21758 41918 21810
rect 41970 21758 41972 21810
rect 41916 21746 41972 21758
rect 42140 21868 42308 21924
rect 42476 23714 42644 23716
rect 42476 23662 42590 23714
rect 42642 23662 42644 23714
rect 42476 23660 42644 23662
rect 42140 21812 42196 21868
rect 41132 20514 41188 20524
rect 41244 20692 41300 20702
rect 41244 20242 41300 20636
rect 41244 20190 41246 20242
rect 41298 20190 41300 20242
rect 41244 20178 41300 20190
rect 40796 19170 40852 19180
rect 40684 18788 40740 18798
rect 40684 17780 40740 18732
rect 40796 18676 40852 18686
rect 40796 17892 40852 18620
rect 40908 18564 40964 18574
rect 40908 18470 40964 18508
rect 41132 18450 41188 18462
rect 41132 18398 41134 18450
rect 41186 18398 41188 18450
rect 41020 18340 41076 18350
rect 41020 18246 41076 18284
rect 40908 17892 40964 17902
rect 40796 17890 40964 17892
rect 40796 17838 40910 17890
rect 40962 17838 40964 17890
rect 40796 17836 40964 17838
rect 41132 17892 41188 18398
rect 41244 17892 41300 17902
rect 41132 17890 41300 17892
rect 41132 17838 41246 17890
rect 41298 17838 41300 17890
rect 41132 17836 41300 17838
rect 40908 17826 40964 17836
rect 41244 17826 41300 17836
rect 40684 17778 40852 17780
rect 40684 17726 40686 17778
rect 40738 17726 40852 17778
rect 40684 17724 40852 17726
rect 40684 17714 40740 17724
rect 40796 17668 40852 17724
rect 41356 17668 41412 20860
rect 41580 20804 41636 20814
rect 41580 20710 41636 20748
rect 41468 20692 41524 20702
rect 41468 20598 41524 20636
rect 41692 20690 41748 20702
rect 41692 20638 41694 20690
rect 41746 20638 41748 20690
rect 41692 20188 41748 20638
rect 41580 20132 41748 20188
rect 41580 19348 41636 20132
rect 41692 20020 41748 20030
rect 41692 19926 41748 19964
rect 41804 20018 41860 20030
rect 41804 19966 41806 20018
rect 41858 19966 41860 20018
rect 41580 19282 41636 19292
rect 41804 19124 41860 19966
rect 42028 20020 42084 20030
rect 42140 20020 42196 21756
rect 42252 21700 42308 21710
rect 42476 21700 42532 23660
rect 42588 23650 42644 23660
rect 42588 23156 42644 23166
rect 42700 23156 42756 24558
rect 42924 26178 42980 26190
rect 42924 26126 42926 26178
rect 42978 26126 42980 26178
rect 42924 25956 42980 26126
rect 43932 26180 43988 26238
rect 43932 26114 43988 26124
rect 42644 23100 42756 23156
rect 42812 23716 42868 23726
rect 42588 23062 42644 23100
rect 42812 22930 42868 23660
rect 42924 23492 42980 25900
rect 43372 25396 43428 25406
rect 43372 25394 43540 25396
rect 43372 25342 43374 25394
rect 43426 25342 43540 25394
rect 43372 25340 43540 25342
rect 43372 25330 43428 25340
rect 43372 24948 43428 24958
rect 43372 24722 43428 24892
rect 43372 24670 43374 24722
rect 43426 24670 43428 24722
rect 43372 24658 43428 24670
rect 43036 24500 43092 24510
rect 43036 24406 43092 24444
rect 43484 24162 43540 25340
rect 43596 25284 43652 25294
rect 43596 24834 43652 25228
rect 44044 24948 44100 28364
rect 44156 28418 44212 28430
rect 44156 28366 44158 28418
rect 44210 28366 44212 28418
rect 44156 27972 44212 28366
rect 44492 27972 44548 27982
rect 44156 27970 44548 27972
rect 44156 27918 44494 27970
rect 44546 27918 44548 27970
rect 44156 27916 44548 27918
rect 44492 27906 44548 27916
rect 44492 27300 44548 27310
rect 44380 26290 44436 26302
rect 44380 26238 44382 26290
rect 44434 26238 44436 26290
rect 43596 24782 43598 24834
rect 43650 24782 43652 24834
rect 43596 24770 43652 24782
rect 43820 24892 44100 24948
rect 44156 25506 44212 25518
rect 44156 25454 44158 25506
rect 44210 25454 44212 25506
rect 43708 24612 43764 24622
rect 43484 24110 43486 24162
rect 43538 24110 43540 24162
rect 43484 24098 43540 24110
rect 43596 24500 43652 24510
rect 43596 24050 43652 24444
rect 43596 23998 43598 24050
rect 43650 23998 43652 24050
rect 43596 23986 43652 23998
rect 43148 23938 43204 23950
rect 43148 23886 43150 23938
rect 43202 23886 43204 23938
rect 42924 23436 43092 23492
rect 43036 23380 43092 23436
rect 43036 23314 43092 23324
rect 42924 23268 42980 23278
rect 42924 23154 42980 23212
rect 42924 23102 42926 23154
rect 42978 23102 42980 23154
rect 42924 23090 42980 23102
rect 43036 23154 43092 23166
rect 43036 23102 43038 23154
rect 43090 23102 43092 23154
rect 43036 22932 43092 23102
rect 43148 23156 43204 23886
rect 43372 23604 43428 23614
rect 43708 23604 43764 24556
rect 43148 23090 43204 23100
rect 43260 23492 43316 23502
rect 42812 22878 42814 22930
rect 42866 22878 42868 22930
rect 42812 22866 42868 22878
rect 42924 22876 43092 22932
rect 42812 22484 42868 22494
rect 42924 22484 42980 22876
rect 43148 22484 43204 22494
rect 43260 22484 43316 23436
rect 42868 22428 42980 22484
rect 43036 22482 43316 22484
rect 43036 22430 43150 22482
rect 43202 22430 43316 22482
rect 43036 22428 43316 22430
rect 42812 22418 42868 22428
rect 42588 22146 42644 22158
rect 42588 22094 42590 22146
rect 42642 22094 42644 22146
rect 42588 21924 42644 22094
rect 42588 21858 42644 21868
rect 42308 21644 42532 21700
rect 42252 21606 42308 21644
rect 42700 21474 42756 21486
rect 42700 21422 42702 21474
rect 42754 21422 42756 21474
rect 42364 20692 42420 20702
rect 42364 20598 42420 20636
rect 42588 20690 42644 20702
rect 42588 20638 42590 20690
rect 42642 20638 42644 20690
rect 42476 20244 42532 20254
rect 42476 20150 42532 20188
rect 42028 20018 42308 20020
rect 42028 19966 42030 20018
rect 42082 19966 42308 20018
rect 42028 19964 42308 19966
rect 42028 19954 42084 19964
rect 41804 19058 41860 19068
rect 42252 19346 42308 19964
rect 42588 19796 42644 20638
rect 42588 19730 42644 19740
rect 42700 19572 42756 21422
rect 42924 20804 42980 20814
rect 42924 20710 42980 20748
rect 42252 19294 42254 19346
rect 42306 19294 42308 19346
rect 42252 19012 42308 19294
rect 42252 18946 42308 18956
rect 42476 19516 42756 19572
rect 42812 20578 42868 20590
rect 42812 20526 42814 20578
rect 42866 20526 42868 20578
rect 42476 18676 42532 19516
rect 42700 19348 42756 19358
rect 42700 19254 42756 19292
rect 42588 19236 42644 19246
rect 42588 19142 42644 19180
rect 42812 18900 42868 20526
rect 42924 20132 42980 20142
rect 43036 20132 43092 22428
rect 43148 22418 43204 22428
rect 43372 21586 43428 23548
rect 43596 23548 43764 23604
rect 43484 22932 43540 22942
rect 43484 22482 43540 22876
rect 43484 22430 43486 22482
rect 43538 22430 43540 22482
rect 43484 22418 43540 22430
rect 43596 22370 43652 23548
rect 43820 23492 43876 24892
rect 44156 24836 44212 25454
rect 44044 24724 44100 24734
rect 44156 24724 44212 24780
rect 44044 24722 44212 24724
rect 44044 24670 44046 24722
rect 44098 24670 44212 24722
rect 44044 24668 44212 24670
rect 44044 24658 44100 24668
rect 43932 23828 43988 23838
rect 43932 23734 43988 23772
rect 44044 23826 44100 23838
rect 44044 23774 44046 23826
rect 44098 23774 44100 23826
rect 44044 23716 44100 23774
rect 44044 23650 44100 23660
rect 44156 23604 44212 24668
rect 44156 23538 44212 23548
rect 44380 25172 44436 26238
rect 43596 22318 43598 22370
rect 43650 22318 43652 22370
rect 43596 22306 43652 22318
rect 43708 23436 43876 23492
rect 43372 21534 43374 21586
rect 43426 21534 43428 21586
rect 43372 21522 43428 21534
rect 43596 21924 43652 21934
rect 43596 20578 43652 21868
rect 43596 20526 43598 20578
rect 43650 20526 43652 20578
rect 43596 20356 43652 20526
rect 42924 20130 43092 20132
rect 42924 20078 42926 20130
rect 42978 20078 43092 20130
rect 42924 20076 43092 20078
rect 43372 20132 43428 20142
rect 42924 20066 42980 20076
rect 43372 20018 43428 20076
rect 43372 19966 43374 20018
rect 43426 19966 43428 20018
rect 43372 19954 43428 19966
rect 43596 19236 43652 20300
rect 43372 19180 43652 19236
rect 43708 19684 43764 23436
rect 44380 23154 44436 25116
rect 44380 23102 44382 23154
rect 44434 23102 44436 23154
rect 44380 23090 44436 23102
rect 43932 22932 43988 22942
rect 43932 22838 43988 22876
rect 44156 22258 44212 22270
rect 44156 22206 44158 22258
rect 44210 22206 44212 22258
rect 44044 22146 44100 22158
rect 44044 22094 44046 22146
rect 44098 22094 44100 22146
rect 44044 21698 44100 22094
rect 44044 21646 44046 21698
rect 44098 21646 44100 21698
rect 44044 21634 44100 21646
rect 44044 20916 44100 20926
rect 44044 20822 44100 20860
rect 44156 20356 44212 22206
rect 44044 20300 44212 20356
rect 43708 19234 43764 19628
rect 43708 19182 43710 19234
rect 43762 19182 43764 19234
rect 42924 19124 42980 19134
rect 42980 19068 43092 19124
rect 42924 19030 42980 19068
rect 42812 18834 42868 18844
rect 42588 18676 42644 18686
rect 42476 18620 42588 18676
rect 40796 17612 40964 17668
rect 40572 17500 40852 17556
rect 39676 17220 39732 17230
rect 39676 17106 39732 17164
rect 39676 17054 39678 17106
rect 39730 17054 39732 17106
rect 39676 17042 39732 17054
rect 39452 16930 39508 16940
rect 39340 16818 39396 16828
rect 39228 15988 39284 15998
rect 39228 15894 39284 15932
rect 39116 15486 39118 15538
rect 39170 15486 39172 15538
rect 39116 15474 39172 15486
rect 39004 15374 39006 15426
rect 39058 15374 39060 15426
rect 38668 14532 38724 14542
rect 38668 13524 38724 14476
rect 38780 14420 38836 14430
rect 38780 14326 38836 14364
rect 39004 14308 39060 15374
rect 39788 15428 39844 15438
rect 39788 15314 39844 15372
rect 39788 15262 39790 15314
rect 39842 15262 39844 15314
rect 39788 15148 39844 15262
rect 39116 15092 39172 15102
rect 39676 15092 39844 15148
rect 39116 15090 39284 15092
rect 39116 15038 39118 15090
rect 39170 15038 39284 15090
rect 39116 15036 39284 15038
rect 39116 15026 39172 15036
rect 39004 14242 39060 14252
rect 38780 13972 38836 13982
rect 38780 13878 38836 13916
rect 39228 13970 39284 15036
rect 39228 13918 39230 13970
rect 39282 13918 39284 13970
rect 39228 13906 39284 13918
rect 39564 14980 39620 14990
rect 39004 13748 39060 13758
rect 39564 13748 39620 14924
rect 39676 14756 39732 15092
rect 39900 14980 39956 17500
rect 40348 17442 40404 17454
rect 40348 17390 40350 17442
rect 40402 17390 40404 17442
rect 40124 17108 40180 17118
rect 40348 17108 40404 17390
rect 40180 17052 40404 17108
rect 40796 17444 40852 17500
rect 40124 17014 40180 17052
rect 40348 16884 40404 16894
rect 40236 16100 40292 16110
rect 40012 15316 40068 15326
rect 40012 15222 40068 15260
rect 40236 15148 40292 16044
rect 40348 15538 40404 16828
rect 40796 16882 40852 17388
rect 40796 16830 40798 16882
rect 40850 16830 40852 16882
rect 40796 16818 40852 16830
rect 40908 16660 40964 17612
rect 41244 17612 41412 17668
rect 41468 18450 41524 18462
rect 41468 18398 41470 18450
rect 41522 18398 41524 18450
rect 41468 17666 41524 18398
rect 42140 18452 42196 18462
rect 42140 18358 42196 18396
rect 41468 17614 41470 17666
rect 41522 17614 41524 17666
rect 41132 16882 41188 16894
rect 41132 16830 41134 16882
rect 41186 16830 41188 16882
rect 40908 16594 40964 16604
rect 41020 16658 41076 16670
rect 41020 16606 41022 16658
rect 41074 16606 41076 16658
rect 41020 16436 41076 16606
rect 40684 16380 41076 16436
rect 40684 15876 40740 16380
rect 41132 16324 41188 16830
rect 40684 15810 40740 15820
rect 40796 16268 41188 16324
rect 40348 15486 40350 15538
rect 40402 15486 40404 15538
rect 40348 15474 40404 15486
rect 40460 15316 40516 15326
rect 40236 15092 40404 15148
rect 39900 14914 39956 14924
rect 40236 14868 40292 14878
rect 39676 14700 40180 14756
rect 39676 14306 39732 14700
rect 39788 14532 39844 14542
rect 39788 14530 40068 14532
rect 39788 14478 39790 14530
rect 39842 14478 40068 14530
rect 39788 14476 40068 14478
rect 39788 14466 39844 14476
rect 39676 14254 39678 14306
rect 39730 14254 39732 14306
rect 39676 14242 39732 14254
rect 39900 14308 39956 14318
rect 39676 13748 39732 13758
rect 39564 13746 39732 13748
rect 39564 13694 39678 13746
rect 39730 13694 39732 13746
rect 39564 13692 39732 13694
rect 39004 13654 39060 13692
rect 39676 13682 39732 13692
rect 38892 13636 38948 13646
rect 38892 13542 38948 13580
rect 38668 12290 38724 13468
rect 39900 13076 39956 14252
rect 40012 13412 40068 14476
rect 40124 13970 40180 14700
rect 40236 14530 40292 14812
rect 40236 14478 40238 14530
rect 40290 14478 40292 14530
rect 40236 14466 40292 14478
rect 40348 14308 40404 15092
rect 40124 13918 40126 13970
rect 40178 13918 40180 13970
rect 40124 13906 40180 13918
rect 40236 14252 40404 14308
rect 40236 13970 40292 14252
rect 40236 13918 40238 13970
rect 40290 13918 40292 13970
rect 40236 13906 40292 13918
rect 40348 13972 40404 13982
rect 40460 13972 40516 15260
rect 40796 14420 40852 16268
rect 40908 15988 40964 15998
rect 40908 14642 40964 15932
rect 41020 15876 41076 15886
rect 41020 15314 41076 15820
rect 41020 15262 41022 15314
rect 41074 15262 41076 15314
rect 41020 15250 41076 15262
rect 41244 15148 41300 17612
rect 41468 17602 41524 17614
rect 41580 18004 41636 18014
rect 41356 17108 41412 17118
rect 41356 17014 41412 17052
rect 41580 17108 41636 17948
rect 41804 17780 41860 17790
rect 41804 17666 41860 17724
rect 41804 17614 41806 17666
rect 41858 17614 41860 17666
rect 41804 17602 41860 17614
rect 41580 17042 41636 17052
rect 41692 17442 41748 17454
rect 41692 17390 41694 17442
rect 41746 17390 41748 17442
rect 41692 16996 41748 17390
rect 41580 15428 41636 15438
rect 41580 15314 41636 15372
rect 41580 15262 41582 15314
rect 41634 15262 41636 15314
rect 41580 15250 41636 15262
rect 40908 14590 40910 14642
rect 40962 14590 40964 14642
rect 40908 14578 40964 14590
rect 41020 15092 41300 15148
rect 41692 15092 41748 16940
rect 42588 17442 42644 18620
rect 42924 18564 42980 18574
rect 42924 18450 42980 18508
rect 42924 18398 42926 18450
rect 42978 18398 42980 18450
rect 42924 18386 42980 18398
rect 43036 18228 43092 19068
rect 42924 18172 43092 18228
rect 43148 19122 43204 19134
rect 43372 19124 43428 19180
rect 43148 19070 43150 19122
rect 43202 19070 43204 19122
rect 43148 19012 43204 19070
rect 42588 17390 42590 17442
rect 42642 17390 42644 17442
rect 41804 16882 41860 16894
rect 41804 16830 41806 16882
rect 41858 16830 41860 16882
rect 41804 16100 41860 16830
rect 42028 16884 42084 16894
rect 42364 16884 42420 16894
rect 42028 16790 42084 16828
rect 42140 16882 42420 16884
rect 42140 16830 42366 16882
rect 42418 16830 42420 16882
rect 42140 16828 42420 16830
rect 41804 16034 41860 16044
rect 41916 16770 41972 16782
rect 41916 16718 41918 16770
rect 41970 16718 41972 16770
rect 41916 15988 41972 16718
rect 41916 15922 41972 15932
rect 42028 16660 42084 16670
rect 42028 15426 42084 16604
rect 42028 15374 42030 15426
rect 42082 15374 42084 15426
rect 42028 15362 42084 15374
rect 40796 14364 40964 14420
rect 40348 13970 40516 13972
rect 40348 13918 40350 13970
rect 40402 13918 40516 13970
rect 40348 13916 40516 13918
rect 40348 13906 40404 13916
rect 40796 13860 40852 13870
rect 40012 13356 40404 13412
rect 40348 13186 40404 13356
rect 40348 13134 40350 13186
rect 40402 13134 40404 13186
rect 40348 13122 40404 13134
rect 40012 13076 40068 13086
rect 38668 12238 38670 12290
rect 38722 12238 38724 12290
rect 38668 12226 38724 12238
rect 39564 13074 40068 13076
rect 39564 13022 40014 13074
rect 40066 13022 40068 13074
rect 39564 13020 40068 13022
rect 38892 12180 38948 12190
rect 38892 12086 38948 12124
rect 39564 12180 39620 13020
rect 40012 13010 40068 13020
rect 40796 12962 40852 13804
rect 40796 12910 40798 12962
rect 40850 12910 40852 12962
rect 40796 12898 40852 12910
rect 40460 12850 40516 12862
rect 40460 12798 40462 12850
rect 40514 12798 40516 12850
rect 40236 12404 40292 12414
rect 40236 12310 40292 12348
rect 39564 12086 39620 12124
rect 38556 11666 38612 11676
rect 39340 11732 39396 11742
rect 38668 11618 38724 11630
rect 38668 11566 38670 11618
rect 38722 11566 38724 11618
rect 38668 11508 38724 11566
rect 38332 11218 38388 11228
rect 38444 11452 38724 11508
rect 37884 3378 37940 3388
rect 37996 9772 38276 9828
rect 38332 10610 38388 10622
rect 38332 10558 38334 10610
rect 38386 10558 38388 10610
rect 37996 3442 38052 9772
rect 38108 9602 38164 9614
rect 38108 9550 38110 9602
rect 38162 9550 38164 9602
rect 38108 9492 38164 9550
rect 38332 9492 38388 10558
rect 38108 9426 38164 9436
rect 38220 9436 38388 9492
rect 38220 5012 38276 9436
rect 38332 9268 38388 9278
rect 38332 9042 38388 9212
rect 38444 9156 38500 11452
rect 39228 11396 39284 11406
rect 39116 11394 39284 11396
rect 39116 11342 39230 11394
rect 39282 11342 39284 11394
rect 39116 11340 39284 11342
rect 38780 11284 38836 11294
rect 38780 10722 38836 11228
rect 38780 10670 38782 10722
rect 38834 10670 38836 10722
rect 38556 10164 38612 10174
rect 38556 9938 38612 10108
rect 38780 10164 38836 10670
rect 38780 10098 38836 10108
rect 38556 9886 38558 9938
rect 38610 9886 38612 9938
rect 38556 9874 38612 9886
rect 38892 9826 38948 9838
rect 38892 9774 38894 9826
rect 38946 9774 38948 9826
rect 38892 9604 38948 9774
rect 38780 9548 38892 9604
rect 38780 9266 38836 9548
rect 38892 9538 38948 9548
rect 38780 9214 38782 9266
rect 38834 9214 38836 9266
rect 38780 9202 38836 9214
rect 38444 9090 38500 9100
rect 38332 8990 38334 9042
rect 38386 8990 38388 9042
rect 38332 8978 38388 8990
rect 38220 4946 38276 4956
rect 38444 4226 38500 4238
rect 38444 4174 38446 4226
rect 38498 4174 38500 4226
rect 37996 3390 37998 3442
rect 38050 3390 38052 3442
rect 37996 3378 38052 3390
rect 38220 3554 38276 3566
rect 38220 3502 38222 3554
rect 38274 3502 38276 3554
rect 38220 2548 38276 3502
rect 38444 3388 38500 4174
rect 38668 3444 38724 3454
rect 38556 3442 38724 3444
rect 38556 3390 38670 3442
rect 38722 3390 38724 3442
rect 38556 3388 38724 3390
rect 38444 3332 38612 3388
rect 38668 3378 38724 3388
rect 39004 3444 39060 3454
rect 39116 3444 39172 11340
rect 39228 11330 39284 11340
rect 39340 9826 39396 11676
rect 40348 11620 40404 11630
rect 39900 11508 39956 11518
rect 39900 11396 39956 11452
rect 39788 11394 39956 11396
rect 39788 11342 39902 11394
rect 39954 11342 39956 11394
rect 39788 11340 39956 11342
rect 39676 11284 39732 11294
rect 39676 11190 39732 11228
rect 39676 10836 39732 10846
rect 39788 10836 39844 11340
rect 39900 11330 39956 11340
rect 40236 11170 40292 11182
rect 40236 11118 40238 11170
rect 40290 11118 40292 11170
rect 39676 10834 39844 10836
rect 39676 10782 39678 10834
rect 39730 10782 39844 10834
rect 39676 10780 39844 10782
rect 40012 11060 40068 11070
rect 40236 11060 40292 11118
rect 40068 11004 40292 11060
rect 39676 10770 39732 10780
rect 39340 9774 39342 9826
rect 39394 9774 39396 9826
rect 39340 9762 39396 9774
rect 39228 9268 39284 9278
rect 39228 9174 39284 9212
rect 39676 9156 39732 9166
rect 39676 9062 39732 9100
rect 39564 8818 39620 8830
rect 39564 8766 39566 8818
rect 39618 8766 39620 8818
rect 39564 7586 39620 8766
rect 40012 8428 40068 11004
rect 40124 9714 40180 9726
rect 40124 9662 40126 9714
rect 40178 9662 40180 9714
rect 40124 9268 40180 9662
rect 40236 9268 40292 9278
rect 40124 9266 40292 9268
rect 40124 9214 40238 9266
rect 40290 9214 40292 9266
rect 40124 9212 40292 9214
rect 40236 9202 40292 9212
rect 40348 9154 40404 11564
rect 40460 11506 40516 12798
rect 40908 12740 40964 14364
rect 40796 12738 40964 12740
rect 40796 12686 40910 12738
rect 40962 12686 40964 12738
rect 40796 12684 40964 12686
rect 40460 11454 40462 11506
rect 40514 11454 40516 11506
rect 40460 11442 40516 11454
rect 40572 12180 40628 12190
rect 40460 11284 40516 11294
rect 40572 11284 40628 12124
rect 40460 11282 40628 11284
rect 40460 11230 40462 11282
rect 40514 11230 40628 11282
rect 40460 11228 40628 11230
rect 40460 11218 40516 11228
rect 40796 11172 40852 12684
rect 40908 12674 40964 12684
rect 40908 11284 40964 11294
rect 40908 11190 40964 11228
rect 40796 11106 40852 11116
rect 40348 9102 40350 9154
rect 40402 9102 40404 9154
rect 40348 9090 40404 9102
rect 40908 9604 40964 9614
rect 40908 9266 40964 9548
rect 40908 9214 40910 9266
rect 40962 9214 40964 9266
rect 39900 8372 40068 8428
rect 40236 9044 40292 9054
rect 39900 8370 39956 8372
rect 39900 8318 39902 8370
rect 39954 8318 39956 8370
rect 39900 8306 39956 8318
rect 39564 7534 39566 7586
rect 39618 7534 39620 7586
rect 39564 7522 39620 7534
rect 39004 3442 39172 3444
rect 39004 3390 39006 3442
rect 39058 3390 39172 3442
rect 39004 3388 39172 3390
rect 39676 4226 39732 4238
rect 39676 4174 39678 4226
rect 39730 4174 39732 4226
rect 39676 3444 39732 4174
rect 39900 3444 39956 3454
rect 39676 3442 39956 3444
rect 39676 3390 39902 3442
rect 39954 3390 39956 3442
rect 39676 3388 39956 3390
rect 39004 3378 39060 3388
rect 38556 2772 38612 3332
rect 36316 2492 36708 2548
rect 36988 2492 37380 2548
rect 37660 2492 38276 2548
rect 38332 2716 38612 2772
rect 36316 800 36372 2492
rect 36988 800 37044 2492
rect 37660 800 37716 2492
rect 38332 800 38388 2716
rect 39676 800 39732 3388
rect 39900 3378 39956 3388
rect 40236 3442 40292 8988
rect 40908 8428 40964 9214
rect 40348 8372 40404 8382
rect 40348 7474 40404 8316
rect 40684 8372 40964 8428
rect 40684 8370 40740 8372
rect 40684 8318 40686 8370
rect 40738 8318 40740 8370
rect 40684 8306 40740 8318
rect 40348 7422 40350 7474
rect 40402 7422 40404 7474
rect 40348 7410 40404 7422
rect 40236 3390 40238 3442
rect 40290 3390 40292 3442
rect 40236 3378 40292 3390
rect 40348 4226 40404 4238
rect 40348 4174 40350 4226
rect 40402 4174 40404 4226
rect 40348 3444 40404 4174
rect 40572 3444 40628 3454
rect 40348 3442 40628 3444
rect 40348 3390 40574 3442
rect 40626 3390 40628 3442
rect 40348 3388 40628 3390
rect 40348 800 40404 3388
rect 40572 3378 40628 3388
rect 40908 3444 40964 3454
rect 41020 3444 41076 15092
rect 41692 15026 41748 15036
rect 41916 15316 41972 15326
rect 41916 15202 41972 15260
rect 41916 15150 41918 15202
rect 41970 15150 41972 15202
rect 41580 14868 41636 14878
rect 41468 13972 41524 13982
rect 41132 13860 41188 13870
rect 41188 13804 41300 13860
rect 41132 13794 41188 13804
rect 41132 13634 41188 13646
rect 41132 13582 41134 13634
rect 41186 13582 41188 13634
rect 41132 12962 41188 13582
rect 41132 12910 41134 12962
rect 41186 12910 41188 12962
rect 41132 12898 41188 12910
rect 41244 12740 41300 13804
rect 41468 13746 41524 13916
rect 41468 13694 41470 13746
rect 41522 13694 41524 13746
rect 41468 13682 41524 13694
rect 41468 12964 41524 12974
rect 41580 12964 41636 14812
rect 41916 13858 41972 15150
rect 42140 13970 42196 16828
rect 42364 16818 42420 16828
rect 42140 13918 42142 13970
rect 42194 13918 42196 13970
rect 42140 13906 42196 13918
rect 42364 15092 42420 15102
rect 42364 13970 42420 15036
rect 42364 13918 42366 13970
rect 42418 13918 42420 13970
rect 42364 13906 42420 13918
rect 42476 13972 42532 13982
rect 41916 13806 41918 13858
rect 41970 13806 41972 13858
rect 41916 13794 41972 13806
rect 42476 13858 42532 13916
rect 42476 13806 42478 13858
rect 42530 13806 42532 13858
rect 42476 13794 42532 13806
rect 41468 12962 41636 12964
rect 41468 12910 41470 12962
rect 41522 12910 41636 12962
rect 41468 12908 41636 12910
rect 41468 12898 41524 12908
rect 41132 12684 41300 12740
rect 41132 12402 41188 12684
rect 41132 12350 41134 12402
rect 41186 12350 41188 12402
rect 41132 12338 41188 12350
rect 41244 12180 41300 12190
rect 41468 12180 41524 12190
rect 41300 12178 41524 12180
rect 41300 12126 41470 12178
rect 41522 12126 41524 12178
rect 41300 12124 41524 12126
rect 41132 10836 41188 10846
rect 41244 10836 41300 12124
rect 41468 12114 41524 12124
rect 41468 11620 41524 11630
rect 41468 11526 41524 11564
rect 41132 10834 41300 10836
rect 41132 10782 41134 10834
rect 41186 10782 41300 10834
rect 41132 10780 41300 10782
rect 41356 11394 41412 11406
rect 41356 11342 41358 11394
rect 41410 11342 41412 11394
rect 41132 10770 41188 10780
rect 41356 9044 41412 11342
rect 41580 10500 41636 12908
rect 42140 12852 42196 12862
rect 42140 12850 42308 12852
rect 42140 12798 42142 12850
rect 42194 12798 42308 12850
rect 42140 12796 42308 12798
rect 42140 12786 42196 12796
rect 42140 11394 42196 11406
rect 42140 11342 42142 11394
rect 42194 11342 42196 11394
rect 42140 11172 42196 11342
rect 42140 11106 42196 11116
rect 42252 10834 42308 12796
rect 42588 12404 42644 17390
rect 42812 17444 42868 17454
rect 42812 17106 42868 17388
rect 42812 17054 42814 17106
rect 42866 17054 42868 17106
rect 42812 16660 42868 17054
rect 42812 16594 42868 16604
rect 42812 16098 42868 16110
rect 42812 16046 42814 16098
rect 42866 16046 42868 16098
rect 42700 15540 42756 15550
rect 42812 15540 42868 16046
rect 42700 15538 42868 15540
rect 42700 15486 42702 15538
rect 42754 15486 42868 15538
rect 42700 15484 42868 15486
rect 42700 15204 42756 15484
rect 42700 15138 42756 15148
rect 42924 13748 42980 18172
rect 43036 17780 43092 17790
rect 43148 17780 43204 18956
rect 43092 17724 43204 17780
rect 43260 19068 43428 19124
rect 43036 17686 43092 17724
rect 43036 15314 43092 15326
rect 43036 15262 43038 15314
rect 43090 15262 43092 15314
rect 43036 14868 43092 15262
rect 43260 15148 43316 19068
rect 43484 19010 43540 19022
rect 43484 18958 43486 19010
rect 43538 18958 43540 19010
rect 43372 18900 43428 18910
rect 43484 18900 43540 18958
rect 43428 18844 43540 18900
rect 43596 19010 43652 19022
rect 43596 18958 43598 19010
rect 43650 18958 43652 19010
rect 43372 18834 43428 18844
rect 43596 18564 43652 18958
rect 43596 18498 43652 18508
rect 43372 18452 43428 18462
rect 43372 17556 43428 18396
rect 43708 18340 43764 19182
rect 43820 19906 43876 19918
rect 43820 19854 43822 19906
rect 43874 19854 43876 19906
rect 43820 18676 43876 19854
rect 44044 19794 44100 20300
rect 44492 20188 44548 27244
rect 44716 26908 44772 33964
rect 44828 33954 44884 33964
rect 46060 33346 46116 38612
rect 46844 37938 46900 37950
rect 46844 37886 46846 37938
rect 46898 37886 46900 37938
rect 46732 37828 46788 37838
rect 46396 37826 46788 37828
rect 46396 37774 46734 37826
rect 46786 37774 46788 37826
rect 46396 37772 46788 37774
rect 46172 36482 46228 36494
rect 46172 36430 46174 36482
rect 46226 36430 46228 36482
rect 46172 35588 46228 36430
rect 46284 35924 46340 35934
rect 46284 35830 46340 35868
rect 46396 35922 46452 37772
rect 46732 37762 46788 37772
rect 46396 35870 46398 35922
rect 46450 35870 46452 35922
rect 46396 35858 46452 35870
rect 46508 37156 46564 37166
rect 46508 35922 46564 37100
rect 46844 37156 46900 37886
rect 46844 37090 46900 37100
rect 46508 35870 46510 35922
rect 46562 35870 46564 35922
rect 46508 35858 46564 35870
rect 46844 35812 46900 35822
rect 46956 35812 47012 38612
rect 47180 38050 47236 40348
rect 47292 39506 47348 42252
rect 47516 42084 47572 42094
rect 47628 42084 47684 42364
rect 47516 42082 47684 42084
rect 47516 42030 47518 42082
rect 47570 42030 47684 42082
rect 47516 42028 47684 42030
rect 47516 42018 47572 42028
rect 47740 40516 47796 43374
rect 47852 42756 47908 42766
rect 47852 42662 47908 42700
rect 48076 42194 48132 43652
rect 48188 43538 48244 43550
rect 48188 43486 48190 43538
rect 48242 43486 48244 43538
rect 48188 42756 48244 43486
rect 48188 42662 48244 42700
rect 48412 42754 48468 43652
rect 48860 43538 48916 43550
rect 48860 43486 48862 43538
rect 48914 43486 48916 43538
rect 48412 42702 48414 42754
rect 48466 42702 48468 42754
rect 48412 42690 48468 42702
rect 48748 43204 48804 43214
rect 48748 42754 48804 43148
rect 48748 42702 48750 42754
rect 48802 42702 48804 42754
rect 48748 42690 48804 42702
rect 48076 42142 48078 42194
rect 48130 42142 48132 42194
rect 48076 42130 48132 42142
rect 48524 42530 48580 42542
rect 48524 42478 48526 42530
rect 48578 42478 48580 42530
rect 48524 40516 48580 42478
rect 48860 41412 48916 43486
rect 49084 42754 49140 43652
rect 49532 43426 49588 43438
rect 49532 43374 49534 43426
rect 49586 43374 49588 43426
rect 49532 42866 49588 43374
rect 49532 42814 49534 42866
rect 49586 42814 49588 42866
rect 49532 42802 49588 42814
rect 49084 42702 49086 42754
rect 49138 42702 49140 42754
rect 49084 42690 49140 42702
rect 49308 42532 49364 42542
rect 48636 41356 48916 41412
rect 48972 42530 49364 42532
rect 48972 42478 49310 42530
rect 49362 42478 49364 42530
rect 48972 42476 49364 42478
rect 48636 41298 48692 41356
rect 48636 41246 48638 41298
rect 48690 41246 48692 41298
rect 48636 41234 48692 41246
rect 47740 40460 47908 40516
rect 47740 40292 47796 40302
rect 47740 39730 47796 40236
rect 47740 39678 47742 39730
rect 47794 39678 47796 39730
rect 47740 39666 47796 39678
rect 47292 39454 47294 39506
rect 47346 39454 47348 39506
rect 47292 39442 47348 39454
rect 47628 39396 47684 39406
rect 47628 39302 47684 39340
rect 47516 38052 47572 38062
rect 47180 37998 47182 38050
rect 47234 37998 47236 38050
rect 47180 37986 47236 37998
rect 47292 38050 47572 38052
rect 47292 37998 47518 38050
rect 47570 37998 47572 38050
rect 47292 37996 47572 37998
rect 46844 35810 47012 35812
rect 46844 35758 46846 35810
rect 46898 35758 47012 35810
rect 46844 35756 47012 35758
rect 46844 35746 46900 35756
rect 46172 35522 46228 35532
rect 46620 35698 46676 35710
rect 46620 35646 46622 35698
rect 46674 35646 46676 35698
rect 46396 35476 46452 35486
rect 46396 34914 46452 35420
rect 46396 34862 46398 34914
rect 46450 34862 46452 34914
rect 46396 34850 46452 34862
rect 46508 34356 46564 34366
rect 46620 34356 46676 35646
rect 47068 35028 47124 35038
rect 47292 35028 47348 37996
rect 47516 37986 47572 37996
rect 47068 35026 47348 35028
rect 47068 34974 47070 35026
rect 47122 34974 47348 35026
rect 47068 34972 47348 34974
rect 47404 37826 47460 37838
rect 47404 37774 47406 37826
rect 47458 37774 47460 37826
rect 47068 34962 47124 34972
rect 46508 34354 46676 34356
rect 46508 34302 46510 34354
rect 46562 34302 46676 34354
rect 46508 34300 46676 34302
rect 46844 34692 46900 34702
rect 46508 34290 46564 34300
rect 46060 33294 46062 33346
rect 46114 33294 46116 33346
rect 46060 33282 46116 33294
rect 46284 34242 46340 34254
rect 46284 34190 46286 34242
rect 46338 34190 46340 34242
rect 46284 33460 46340 34190
rect 46284 33348 46340 33404
rect 46732 34244 46788 34254
rect 46396 33348 46452 33358
rect 46284 33346 46452 33348
rect 46284 33294 46398 33346
rect 46450 33294 46452 33346
rect 46284 33292 46452 33294
rect 46396 33282 46452 33292
rect 44940 33124 44996 33134
rect 44940 30212 44996 33068
rect 46284 33124 46340 33134
rect 46284 33030 46340 33068
rect 46284 32450 46340 32462
rect 46284 32398 46286 32450
rect 46338 32398 46340 32450
rect 46284 32004 46340 32398
rect 45500 31948 46340 32004
rect 45500 31890 45556 31948
rect 45500 31838 45502 31890
rect 45554 31838 45556 31890
rect 45500 31826 45556 31838
rect 45612 31780 45668 31790
rect 45612 31778 46228 31780
rect 45612 31726 45614 31778
rect 45666 31726 46228 31778
rect 45612 31724 46228 31726
rect 45612 31714 45668 31724
rect 45164 31668 45220 31678
rect 45164 31556 45220 31612
rect 45052 31554 45220 31556
rect 45052 31502 45166 31554
rect 45218 31502 45220 31554
rect 45052 31500 45220 31502
rect 45052 30324 45108 31500
rect 45164 31490 45220 31500
rect 45388 31554 45444 31566
rect 45388 31502 45390 31554
rect 45442 31502 45444 31554
rect 45388 31332 45444 31502
rect 45836 31556 45892 31566
rect 45836 31554 46004 31556
rect 45836 31502 45838 31554
rect 45890 31502 46004 31554
rect 45836 31500 46004 31502
rect 45836 31490 45892 31500
rect 45388 31276 45780 31332
rect 45724 31218 45780 31276
rect 45724 31166 45726 31218
rect 45778 31166 45780 31218
rect 45724 31154 45780 31166
rect 45164 30996 45220 31006
rect 45164 30902 45220 30940
rect 45612 30994 45668 31006
rect 45612 30942 45614 30994
rect 45666 30942 45668 30994
rect 45052 30258 45108 30268
rect 45164 30772 45220 30782
rect 44940 28642 44996 30156
rect 44940 28590 44942 28642
rect 44994 28590 44996 28642
rect 44940 28578 44996 28590
rect 45052 30098 45108 30110
rect 45052 30046 45054 30098
rect 45106 30046 45108 30098
rect 45052 28642 45108 30046
rect 45164 29764 45220 30716
rect 45612 30548 45668 30942
rect 45836 30994 45892 31006
rect 45836 30942 45838 30994
rect 45890 30942 45892 30994
rect 45836 30884 45892 30942
rect 45948 30996 46004 31500
rect 46172 31218 46228 31724
rect 46508 31778 46564 31790
rect 46508 31726 46510 31778
rect 46562 31726 46564 31778
rect 46508 31668 46564 31726
rect 46508 31602 46564 31612
rect 46172 31166 46174 31218
rect 46226 31166 46228 31218
rect 46172 31154 46228 31166
rect 46284 31554 46340 31566
rect 46284 31502 46286 31554
rect 46338 31502 46340 31554
rect 46284 31220 46340 31502
rect 46732 31332 46788 34188
rect 46844 34242 46900 34636
rect 47404 34354 47460 37774
rect 47628 37828 47684 37838
rect 47628 37734 47684 37772
rect 47740 37826 47796 37838
rect 47740 37774 47742 37826
rect 47794 37774 47796 37826
rect 47740 37492 47796 37774
rect 47740 37426 47796 37436
rect 47852 37156 47908 40460
rect 48524 40450 48580 40460
rect 48636 40404 48692 40414
rect 48748 40404 48804 41356
rect 48692 40402 48804 40404
rect 48692 40350 48750 40402
rect 48802 40350 48804 40402
rect 48692 40348 48804 40350
rect 48636 39618 48692 40348
rect 48748 40338 48804 40348
rect 48860 40516 48916 40526
rect 48636 39566 48638 39618
rect 48690 39566 48692 39618
rect 48636 39554 48692 39566
rect 48524 37938 48580 37950
rect 48524 37886 48526 37938
rect 48578 37886 48580 37938
rect 48412 37828 48468 37838
rect 48412 37734 48468 37772
rect 48076 37492 48132 37502
rect 47628 37100 47908 37156
rect 47964 37156 48020 37166
rect 47628 35698 47684 37100
rect 47964 37062 48020 37100
rect 47964 36260 48020 36270
rect 47964 35922 48020 36204
rect 47964 35870 47966 35922
rect 48018 35870 48020 35922
rect 47964 35858 48020 35870
rect 48076 35924 48132 37436
rect 48524 37268 48580 37886
rect 48524 37202 48580 37212
rect 48860 37266 48916 40460
rect 48972 38668 49028 42476
rect 49308 42466 49364 42476
rect 49532 42532 49588 42542
rect 49532 42438 49588 42476
rect 49308 42084 49364 42094
rect 49308 41990 49364 42028
rect 49532 42082 49588 42094
rect 49532 42030 49534 42082
rect 49586 42030 49588 42082
rect 49084 41972 49140 41982
rect 49084 41878 49140 41916
rect 49420 41858 49476 41870
rect 49420 41806 49422 41858
rect 49474 41806 49476 41858
rect 49196 41188 49252 41198
rect 49196 41094 49252 41132
rect 49196 40964 49252 40974
rect 49084 39060 49140 39070
rect 49084 38966 49140 39004
rect 49196 39058 49252 40908
rect 49420 40516 49476 41806
rect 49532 41412 49588 42030
rect 49532 41346 49588 41356
rect 49532 40516 49588 40526
rect 49420 40514 49588 40516
rect 49420 40462 49534 40514
rect 49586 40462 49588 40514
rect 49420 40460 49588 40462
rect 49532 40450 49588 40460
rect 49196 39006 49198 39058
rect 49250 39006 49252 39058
rect 49196 38994 49252 39006
rect 49308 39506 49364 39518
rect 49308 39454 49310 39506
rect 49362 39454 49364 39506
rect 49308 39058 49364 39454
rect 49308 39006 49310 39058
rect 49362 39006 49364 39058
rect 49308 38994 49364 39006
rect 49644 38946 49700 43652
rect 49868 42868 49924 53676
rect 50540 53666 50596 53676
rect 50204 53618 50260 53630
rect 50204 53566 50206 53618
rect 50258 53566 50260 53618
rect 50204 53284 50260 53566
rect 50316 53620 50372 53630
rect 50316 53526 50372 53564
rect 50876 53620 50932 53630
rect 50876 53526 50932 53564
rect 50556 53340 50820 53350
rect 50612 53284 50660 53340
rect 50716 53284 50764 53340
rect 50556 53274 50820 53284
rect 50092 52724 50148 52734
rect 50204 52724 50260 53228
rect 50148 52668 50260 52724
rect 50092 52658 50148 52668
rect 50556 51772 50820 51782
rect 50612 51716 50660 51772
rect 50716 51716 50764 51772
rect 50556 51706 50820 51716
rect 49980 50594 50036 50606
rect 49980 50542 49982 50594
rect 50034 50542 50036 50594
rect 49980 50372 50036 50542
rect 49980 50306 50036 50316
rect 51660 50372 51716 54462
rect 50556 50204 50820 50214
rect 50612 50148 50660 50204
rect 50716 50148 50764 50204
rect 50556 50138 50820 50148
rect 51660 49922 51716 50316
rect 51660 49870 51662 49922
rect 51714 49870 51716 49922
rect 51660 49858 51716 49870
rect 49980 49140 50036 49150
rect 49980 49138 50484 49140
rect 49980 49086 49982 49138
rect 50034 49086 50484 49138
rect 49980 49084 50484 49086
rect 49980 49074 50036 49084
rect 50428 49026 50484 49084
rect 50428 48974 50430 49026
rect 50482 48974 50484 49026
rect 50428 48962 50484 48974
rect 50316 48804 50372 48814
rect 50316 48710 50372 48748
rect 50556 48636 50820 48646
rect 50612 48580 50660 48636
rect 50716 48580 50764 48636
rect 50556 48570 50820 48580
rect 50556 47068 50820 47078
rect 50612 47012 50660 47068
rect 50716 47012 50764 47068
rect 50556 47002 50820 47012
rect 51100 45892 51156 45902
rect 50556 45500 50820 45510
rect 50612 45444 50660 45500
rect 50716 45444 50764 45500
rect 50556 45434 50820 45444
rect 50556 43932 50820 43942
rect 50612 43876 50660 43932
rect 50716 43876 50764 43932
rect 50556 43866 50820 43876
rect 50652 43764 50708 43774
rect 49868 42802 49924 42812
rect 50204 42868 50260 42878
rect 50204 42774 50260 42812
rect 50652 42866 50708 43708
rect 50652 42814 50654 42866
rect 50706 42814 50708 42866
rect 50652 42802 50708 42814
rect 49756 42754 49812 42766
rect 49756 42702 49758 42754
rect 49810 42702 49812 42754
rect 49756 41970 49812 42702
rect 50540 42532 50596 42570
rect 50540 42466 50596 42476
rect 50556 42364 50820 42374
rect 50612 42308 50660 42364
rect 50716 42308 50764 42364
rect 50556 42298 50820 42308
rect 50316 42084 50372 42094
rect 50372 42028 50484 42084
rect 50316 42018 50372 42028
rect 49756 41918 49758 41970
rect 49810 41918 49812 41970
rect 49756 39060 49812 41918
rect 49756 38994 49812 39004
rect 49644 38894 49646 38946
rect 49698 38894 49700 38946
rect 49644 38882 49700 38894
rect 49420 38836 49476 38846
rect 49420 38834 49588 38836
rect 49420 38782 49422 38834
rect 49474 38782 49588 38834
rect 49420 38780 49588 38782
rect 49420 38770 49476 38780
rect 49532 38668 49588 38780
rect 48972 38612 49476 38668
rect 49532 38612 49812 38668
rect 49308 37492 49364 37502
rect 49308 37398 49364 37436
rect 48860 37214 48862 37266
rect 48914 37214 48916 37266
rect 48860 37202 48916 37214
rect 48972 37266 49028 37278
rect 48972 37214 48974 37266
rect 49026 37214 49028 37266
rect 48748 36370 48804 36382
rect 48748 36318 48750 36370
rect 48802 36318 48804 36370
rect 48076 35830 48132 35868
rect 48188 36036 48244 36046
rect 47628 35646 47630 35698
rect 47682 35646 47684 35698
rect 47628 35634 47684 35646
rect 47740 35698 47796 35710
rect 47740 35646 47742 35698
rect 47794 35646 47796 35698
rect 47740 34916 47796 35646
rect 47740 34850 47796 34860
rect 47964 35586 48020 35598
rect 47964 35534 47966 35586
rect 48018 35534 48020 35586
rect 47404 34302 47406 34354
rect 47458 34302 47460 34354
rect 47404 34290 47460 34302
rect 47516 34692 47572 34702
rect 46844 34190 46846 34242
rect 46898 34190 46900 34242
rect 46844 34178 46900 34190
rect 47516 34132 47572 34636
rect 47628 34356 47684 34366
rect 47628 34262 47684 34300
rect 47964 34244 48020 35534
rect 48188 34692 48244 35980
rect 48748 35698 48804 36318
rect 48972 36036 49028 37214
rect 49196 37266 49252 37278
rect 49196 37214 49198 37266
rect 49250 37214 49252 37266
rect 48748 35646 48750 35698
rect 48802 35646 48804 35698
rect 48748 35476 48804 35646
rect 48748 35410 48804 35420
rect 48860 35980 49028 36036
rect 49084 37154 49140 37166
rect 49084 37102 49086 37154
rect 49138 37102 49140 37154
rect 48860 35140 48916 35980
rect 49084 35924 49140 37102
rect 49196 36708 49252 37214
rect 49196 36642 49252 36652
rect 49308 37268 49364 37278
rect 49084 35858 49140 35868
rect 49308 35812 49364 37212
rect 49420 36148 49476 38612
rect 49420 36092 49700 36148
rect 49420 35924 49476 35934
rect 49476 35868 49588 35924
rect 49420 35858 49476 35868
rect 48188 34626 48244 34636
rect 48636 35084 48916 35140
rect 49196 35756 49364 35812
rect 49532 35810 49588 35868
rect 49532 35758 49534 35810
rect 49586 35758 49588 35810
rect 47964 34178 48020 34188
rect 48188 34356 48244 34366
rect 47740 34132 47796 34142
rect 47516 34130 47796 34132
rect 47516 34078 47742 34130
rect 47794 34078 47796 34130
rect 47516 34076 47796 34078
rect 47068 33684 47124 33694
rect 47068 32562 47124 33628
rect 47740 33348 47796 34076
rect 48188 34020 48244 34300
rect 48188 33954 48244 33964
rect 48188 33796 48244 33806
rect 48076 33572 48132 33582
rect 48188 33572 48244 33740
rect 48636 33796 48692 35084
rect 49196 35026 49252 35756
rect 49532 35746 49588 35758
rect 49644 35588 49700 36092
rect 49196 34974 49198 35026
rect 49250 34974 49252 35026
rect 49196 34962 49252 34974
rect 49420 35532 49700 35588
rect 48860 34916 48916 34926
rect 48636 33730 48692 33740
rect 48748 34130 48804 34142
rect 48748 34078 48750 34130
rect 48802 34078 48804 34130
rect 48748 33684 48804 34078
rect 48748 33618 48804 33628
rect 48076 33570 48244 33572
rect 48076 33518 48078 33570
rect 48130 33518 48244 33570
rect 48076 33516 48244 33518
rect 48860 33570 48916 34860
rect 48860 33518 48862 33570
rect 48914 33518 48916 33570
rect 48076 33506 48132 33516
rect 48860 33506 48916 33518
rect 49420 33570 49476 35532
rect 49532 34244 49588 34254
rect 49532 34150 49588 34188
rect 49420 33518 49422 33570
rect 49474 33518 49476 33570
rect 49420 33506 49476 33518
rect 49532 33460 49588 33470
rect 47964 33348 48020 33358
rect 47740 33292 47964 33348
rect 47964 33254 48020 33292
rect 48748 33348 48804 33358
rect 48748 33254 48804 33292
rect 49532 33346 49588 33404
rect 49532 33294 49534 33346
rect 49586 33294 49588 33346
rect 49532 33282 49588 33294
rect 49756 33346 49812 38612
rect 50428 36932 50484 42028
rect 50988 41412 51044 41422
rect 50988 41318 51044 41356
rect 51100 41300 51156 45836
rect 51660 44324 51716 44334
rect 51660 43764 51716 44268
rect 51660 43426 51716 43708
rect 51660 43374 51662 43426
rect 51714 43374 51716 43426
rect 51660 43362 51716 43374
rect 52108 43316 52164 59724
rect 52332 58996 52388 59006
rect 52220 56980 52276 56990
rect 52220 44548 52276 56924
rect 52332 48356 52388 58940
rect 52332 48290 52388 48300
rect 57932 47570 57988 47582
rect 57932 47518 57934 47570
rect 57986 47518 57988 47570
rect 55580 47460 55636 47470
rect 55468 47458 55636 47460
rect 55468 47406 55582 47458
rect 55634 47406 55636 47458
rect 55468 47404 55636 47406
rect 53452 46674 53508 46686
rect 53452 46622 53454 46674
rect 53506 46622 53508 46674
rect 53228 46564 53284 46574
rect 53452 46564 53508 46622
rect 53228 46562 53508 46564
rect 53228 46510 53230 46562
rect 53282 46510 53508 46562
rect 53228 46508 53508 46510
rect 52220 44482 52276 44492
rect 52668 45890 52724 45902
rect 52668 45838 52670 45890
rect 52722 45838 52724 45890
rect 52108 43250 52164 43260
rect 51660 42084 51716 42094
rect 51100 41298 51380 41300
rect 51100 41246 51102 41298
rect 51154 41246 51380 41298
rect 51100 41244 51380 41246
rect 51100 41234 51156 41244
rect 50556 40796 50820 40806
rect 50612 40740 50660 40796
rect 50716 40740 50764 40796
rect 50556 40730 50820 40740
rect 51324 40740 51380 41244
rect 51548 41188 51604 41198
rect 51660 41188 51716 42028
rect 52668 42084 52724 45838
rect 53228 42980 53284 46508
rect 55356 46452 55412 46462
rect 55356 46358 55412 46396
rect 55020 46002 55076 46014
rect 55020 45950 55022 46002
rect 55074 45950 55076 46002
rect 55020 45780 55076 45950
rect 55020 45714 55076 45724
rect 53228 42914 53284 42924
rect 52668 42018 52724 42028
rect 53788 42756 53844 42766
rect 52108 41972 52164 41982
rect 51548 41186 51828 41188
rect 51548 41134 51550 41186
rect 51602 41134 51828 41186
rect 51548 41132 51828 41134
rect 51548 41122 51604 41132
rect 51436 40964 51492 40974
rect 51436 40870 51492 40908
rect 51324 40684 51716 40740
rect 51660 40290 51716 40684
rect 51660 40238 51662 40290
rect 51714 40238 51716 40290
rect 51660 40226 51716 40238
rect 51772 40068 51828 41132
rect 52108 40292 52164 41916
rect 53452 41970 53508 41982
rect 53452 41918 53454 41970
rect 53506 41918 53508 41970
rect 53228 41860 53284 41870
rect 53452 41860 53508 41918
rect 53228 41858 53508 41860
rect 53228 41806 53230 41858
rect 53282 41806 53508 41858
rect 53228 41804 53508 41806
rect 53228 41524 53284 41804
rect 53228 41458 53284 41468
rect 52108 40226 52164 40236
rect 52668 41186 52724 41198
rect 52668 41134 52670 41186
rect 52722 41134 52724 41186
rect 51436 40012 51828 40068
rect 51436 39730 51492 40012
rect 51436 39678 51438 39730
rect 51490 39678 51492 39730
rect 51436 39666 51492 39678
rect 50556 39228 50820 39238
rect 50612 39172 50660 39228
rect 50716 39172 50764 39228
rect 50556 39162 50820 39172
rect 52668 38948 52724 41134
rect 53452 40404 53508 40414
rect 53452 40310 53508 40348
rect 53788 40180 53844 42700
rect 55468 41972 55524 47404
rect 55580 47394 55636 47404
rect 57820 46002 57876 46014
rect 57820 45950 57822 46002
rect 57874 45950 57876 46002
rect 55580 45892 55636 45902
rect 55580 45798 55636 45836
rect 57820 44436 57876 45950
rect 57932 45108 57988 47518
rect 57932 45042 57988 45052
rect 57820 44370 57876 44380
rect 57932 44434 57988 44446
rect 57932 44382 57934 44434
rect 57986 44382 57988 44434
rect 55580 44324 55636 44334
rect 55580 44230 55636 44268
rect 57932 43764 57988 44382
rect 57932 43698 57988 43708
rect 57932 43092 57988 43102
rect 57932 42978 57988 43036
rect 57932 42926 57934 42978
rect 57986 42926 57988 42978
rect 57932 42914 57988 42926
rect 55580 42756 55636 42766
rect 55580 42662 55636 42700
rect 55468 41906 55524 41916
rect 57932 42420 57988 42430
rect 55356 41748 55412 41758
rect 55356 41654 55412 41692
rect 57932 41410 57988 42364
rect 57932 41358 57934 41410
rect 57986 41358 57988 41410
rect 57932 41346 57988 41358
rect 55020 41298 55076 41310
rect 55020 41246 55022 41298
rect 55074 41246 55076 41298
rect 55020 40404 55076 41246
rect 55580 41188 55636 41198
rect 55020 40338 55076 40348
rect 55468 41186 55636 41188
rect 55468 41134 55582 41186
rect 55634 41134 55636 41186
rect 55468 41132 55636 41134
rect 53788 40114 53844 40124
rect 55356 40178 55412 40190
rect 55356 40126 55358 40178
rect 55410 40126 55412 40178
rect 55356 39732 55412 40126
rect 55356 39666 55412 39676
rect 55468 39844 55524 41132
rect 55580 41122 55636 41132
rect 55356 39508 55412 39518
rect 55468 39508 55524 39788
rect 57932 41076 57988 41086
rect 57932 39842 57988 41020
rect 57932 39790 57934 39842
rect 57986 39790 57988 39842
rect 57932 39778 57988 39790
rect 55580 39620 55636 39630
rect 55580 39526 55636 39564
rect 55356 39506 55524 39508
rect 55356 39454 55358 39506
rect 55410 39454 55524 39506
rect 55356 39452 55524 39454
rect 55356 39442 55412 39452
rect 52668 38882 52724 38892
rect 57932 39060 57988 39070
rect 53452 38834 53508 38846
rect 53452 38782 53454 38834
rect 53506 38782 53508 38834
rect 53228 38724 53284 38734
rect 53452 38724 53508 38782
rect 53228 38722 53508 38724
rect 53228 38670 53230 38722
rect 53282 38670 53508 38722
rect 53228 38668 53508 38670
rect 53228 38164 53284 38668
rect 55356 38612 55412 38622
rect 55356 38518 55412 38556
rect 57932 38274 57988 39004
rect 57932 38222 57934 38274
rect 57986 38222 57988 38274
rect 57932 38210 57988 38222
rect 53228 38098 53284 38108
rect 55356 38052 55412 38062
rect 55580 38052 55636 38062
rect 55412 38050 55636 38052
rect 55412 37998 55582 38050
rect 55634 37998 55636 38050
rect 55412 37996 55636 37998
rect 55356 37958 55412 37996
rect 55580 37986 55636 37996
rect 57932 37716 57988 37726
rect 50556 37660 50820 37670
rect 50612 37604 50660 37660
rect 50716 37604 50764 37660
rect 50556 37594 50820 37604
rect 53452 37268 53508 37278
rect 53452 37174 53508 37212
rect 50316 36876 50484 36932
rect 52668 37156 52724 37166
rect 49868 35700 49924 35710
rect 49868 35364 49924 35644
rect 50316 35476 50372 36876
rect 50428 36708 50484 36718
rect 50428 36614 50484 36652
rect 52108 36484 52164 36494
rect 50540 36372 50596 36382
rect 50428 36370 50596 36372
rect 50428 36318 50542 36370
rect 50594 36318 50596 36370
rect 50428 36316 50596 36318
rect 50428 35588 50484 36316
rect 50540 36306 50596 36316
rect 50988 36370 51044 36382
rect 50988 36318 50990 36370
rect 51042 36318 51044 36370
rect 50876 36260 50932 36270
rect 50876 36166 50932 36204
rect 50556 36092 50820 36102
rect 50612 36036 50660 36092
rect 50716 36036 50764 36092
rect 50556 36026 50820 36036
rect 50540 35588 50596 35598
rect 50428 35532 50540 35588
rect 50540 35522 50596 35532
rect 50316 35420 50484 35476
rect 49868 35298 49924 35308
rect 50428 33572 50484 35420
rect 50556 34524 50820 34534
rect 50612 34468 50660 34524
rect 50716 34468 50764 34524
rect 50556 34458 50820 34468
rect 50988 34020 51044 36318
rect 52108 36258 52164 36428
rect 52108 36206 52110 36258
rect 52162 36206 52164 36258
rect 52108 35812 52164 36206
rect 52108 35746 52164 35756
rect 51660 35588 51716 35598
rect 51660 35494 51716 35532
rect 50988 33954 51044 33964
rect 51660 34020 51716 34030
rect 51660 33926 51716 33964
rect 50540 33572 50596 33582
rect 50428 33570 50596 33572
rect 50428 33518 50542 33570
rect 50594 33518 50596 33570
rect 50428 33516 50596 33518
rect 50540 33506 50596 33516
rect 49756 33294 49758 33346
rect 49810 33294 49812 33346
rect 49756 33282 49812 33294
rect 50092 33460 50148 33470
rect 50092 33346 50148 33404
rect 50092 33294 50094 33346
rect 50146 33294 50148 33346
rect 50092 33282 50148 33294
rect 50652 33460 50708 33470
rect 50652 33346 50708 33404
rect 50652 33294 50654 33346
rect 50706 33294 50708 33346
rect 50652 33282 50708 33294
rect 47740 33124 47796 33134
rect 48076 33124 48132 33134
rect 47740 33122 48132 33124
rect 47740 33070 47742 33122
rect 47794 33070 48078 33122
rect 48130 33070 48132 33122
rect 47740 33068 48132 33070
rect 47740 33058 47796 33068
rect 47068 32510 47070 32562
rect 47122 32510 47124 32562
rect 47068 31780 47124 32510
rect 47628 31780 47684 31790
rect 47068 31778 47684 31780
rect 47068 31726 47630 31778
rect 47682 31726 47684 31778
rect 47068 31724 47684 31726
rect 46956 31556 47012 31566
rect 46956 31554 47124 31556
rect 46956 31502 46958 31554
rect 47010 31502 47124 31554
rect 46956 31500 47124 31502
rect 46956 31490 47012 31500
rect 46732 31276 47012 31332
rect 46284 31154 46340 31164
rect 46396 31052 46900 31108
rect 46396 30996 46452 31052
rect 45948 30940 46452 30996
rect 45836 30660 45892 30828
rect 46508 30884 46564 30894
rect 46732 30884 46788 30894
rect 46508 30790 46564 30828
rect 46620 30882 46788 30884
rect 46620 30830 46734 30882
rect 46786 30830 46788 30882
rect 46620 30828 46788 30830
rect 45612 30482 45668 30492
rect 45724 30604 45892 30660
rect 45612 30212 45668 30222
rect 45724 30212 45780 30604
rect 45500 30210 45780 30212
rect 45500 30158 45614 30210
rect 45666 30158 45780 30210
rect 45500 30156 45780 30158
rect 45948 30548 46004 30558
rect 45948 30210 46004 30492
rect 46620 30548 46676 30828
rect 46732 30818 46788 30828
rect 45948 30158 45950 30210
rect 46002 30158 46004 30210
rect 45388 30098 45444 30110
rect 45388 30046 45390 30098
rect 45442 30046 45444 30098
rect 45276 29988 45332 29998
rect 45276 29894 45332 29932
rect 45164 29708 45332 29764
rect 45052 28590 45054 28642
rect 45106 28590 45108 28642
rect 45052 27636 45108 28590
rect 45164 28530 45220 28542
rect 45164 28478 45166 28530
rect 45218 28478 45220 28530
rect 45164 28084 45220 28478
rect 45164 28018 45220 28028
rect 45276 27858 45332 29708
rect 45388 29652 45444 30046
rect 45388 29586 45444 29596
rect 45500 28420 45556 30156
rect 45612 30146 45668 30156
rect 45948 30146 46004 30158
rect 46060 30324 46116 30334
rect 45836 29986 45892 29998
rect 45836 29934 45838 29986
rect 45890 29934 45892 29986
rect 45836 29204 45892 29934
rect 45836 29138 45892 29148
rect 45948 29988 46004 29998
rect 45948 28866 46004 29932
rect 46060 29204 46116 30268
rect 46172 30100 46228 30110
rect 46172 29428 46228 30044
rect 46172 29334 46228 29372
rect 46284 30098 46340 30110
rect 46284 30046 46286 30098
rect 46338 30046 46340 30098
rect 46060 29138 46116 29148
rect 45948 28814 45950 28866
rect 46002 28814 46004 28866
rect 45948 28802 46004 28814
rect 45612 28644 45668 28654
rect 46284 28644 46340 30046
rect 46508 29652 46564 29662
rect 46508 29558 46564 29596
rect 46620 29650 46676 30492
rect 46732 30436 46788 30446
rect 46844 30436 46900 31052
rect 46732 30434 46900 30436
rect 46732 30382 46734 30434
rect 46786 30382 46900 30434
rect 46732 30380 46900 30382
rect 46732 30370 46788 30380
rect 46844 30212 46900 30222
rect 46844 30118 46900 30156
rect 46732 30100 46788 30110
rect 46732 30006 46788 30044
rect 46844 29876 46900 29886
rect 46620 29598 46622 29650
rect 46674 29598 46676 29650
rect 46620 29586 46676 29598
rect 46732 29652 46788 29662
rect 46844 29652 46900 29820
rect 46732 29650 46900 29652
rect 46732 29598 46734 29650
rect 46786 29598 46900 29650
rect 46732 29596 46900 29598
rect 46732 29586 46788 29596
rect 46956 29428 47012 31276
rect 47068 30884 47124 31500
rect 47292 31554 47348 31566
rect 47292 31502 47294 31554
rect 47346 31502 47348 31554
rect 47180 30884 47236 30894
rect 47068 30882 47236 30884
rect 47068 30830 47182 30882
rect 47234 30830 47236 30882
rect 47068 30828 47236 30830
rect 47180 30436 47236 30828
rect 47180 30370 47236 30380
rect 47292 30100 47348 31502
rect 47628 31108 47684 31724
rect 48076 31220 48132 33068
rect 48860 33122 48916 33134
rect 48860 33070 48862 33122
rect 48914 33070 48916 33122
rect 48860 32452 48916 33070
rect 49420 33122 49476 33134
rect 49420 33070 49422 33122
rect 49474 33070 49476 33122
rect 48860 32386 48916 32396
rect 49196 32452 49252 32462
rect 49196 32358 49252 32396
rect 49420 31892 49476 33070
rect 49420 31826 49476 31836
rect 49980 33122 50036 33134
rect 50540 33124 50596 33134
rect 49980 33070 49982 33122
rect 50034 33070 50036 33122
rect 48412 31668 48468 31678
rect 48412 31666 48916 31668
rect 48412 31614 48414 31666
rect 48466 31614 48916 31666
rect 48412 31612 48916 31614
rect 48412 31602 48468 31612
rect 48076 31154 48132 31164
rect 48636 31220 48692 31230
rect 47404 30996 47460 31006
rect 47404 30902 47460 30940
rect 47628 30772 47684 31052
rect 47852 30996 47908 31006
rect 47628 30706 47684 30716
rect 47740 30994 47908 30996
rect 47740 30942 47854 30994
rect 47906 30942 47908 30994
rect 47740 30940 47908 30942
rect 47292 30034 47348 30044
rect 47628 30322 47684 30334
rect 47628 30270 47630 30322
rect 47682 30270 47684 30322
rect 47628 29652 47684 30270
rect 47740 29876 47796 30940
rect 47852 30930 47908 30940
rect 48076 30994 48132 31006
rect 48076 30942 48078 30994
rect 48130 30942 48132 30994
rect 47964 30882 48020 30894
rect 47964 30830 47966 30882
rect 48018 30830 48020 30882
rect 47740 29810 47796 29820
rect 47852 30210 47908 30222
rect 47852 30158 47854 30210
rect 47906 30158 47908 30210
rect 47852 30100 47908 30158
rect 47964 30212 48020 30830
rect 47964 30146 48020 30156
rect 47628 29596 47796 29652
rect 47404 29540 47460 29550
rect 47404 29446 47460 29484
rect 45612 28642 46340 28644
rect 45612 28590 45614 28642
rect 45666 28590 46286 28642
rect 46338 28590 46340 28642
rect 45612 28588 46340 28590
rect 45612 28578 45668 28588
rect 46284 28578 46340 28588
rect 46396 29372 47012 29428
rect 47180 29426 47236 29438
rect 47180 29374 47182 29426
rect 47234 29374 47236 29426
rect 46060 28420 46116 28430
rect 45500 28418 46116 28420
rect 45500 28366 46062 28418
rect 46114 28366 46116 28418
rect 45500 28364 46116 28366
rect 46060 28354 46116 28364
rect 45724 28084 45780 28094
rect 45780 28028 46004 28084
rect 45724 27990 45780 28028
rect 45276 27806 45278 27858
rect 45330 27806 45332 27858
rect 45276 27794 45332 27806
rect 45388 27972 45444 27982
rect 45052 27570 45108 27580
rect 45388 27076 45444 27916
rect 45724 27076 45780 27086
rect 45388 27074 45780 27076
rect 45388 27022 45390 27074
rect 45442 27022 45726 27074
rect 45778 27022 45780 27074
rect 45388 27020 45780 27022
rect 45388 27010 45444 27020
rect 45724 27010 45780 27020
rect 44604 26852 44772 26908
rect 44828 26962 44884 26974
rect 44828 26910 44830 26962
rect 44882 26910 44884 26962
rect 44604 23604 44660 26852
rect 44828 26066 44884 26910
rect 45836 26962 45892 26974
rect 45836 26910 45838 26962
rect 45890 26910 45892 26962
rect 44940 26852 44996 26862
rect 44940 26758 44996 26796
rect 45612 26852 45668 26862
rect 44828 26014 44830 26066
rect 44882 26014 44884 26066
rect 44828 26002 44884 26014
rect 44940 26290 44996 26302
rect 44940 26238 44942 26290
rect 44994 26238 44996 26290
rect 44828 25506 44884 25518
rect 44828 25454 44830 25506
rect 44882 25454 44884 25506
rect 44828 24836 44884 25454
rect 44828 24770 44884 24780
rect 44940 25284 44996 26238
rect 45276 26290 45332 26302
rect 45276 26238 45278 26290
rect 45330 26238 45332 26290
rect 45276 26068 45332 26238
rect 45276 26002 45332 26012
rect 45612 25618 45668 26796
rect 45612 25566 45614 25618
rect 45666 25566 45668 25618
rect 45612 25554 45668 25566
rect 45836 26852 45892 26910
rect 45948 26908 46004 28028
rect 46172 27188 46228 27198
rect 46060 27076 46116 27114
rect 46060 27010 46116 27020
rect 46172 27074 46228 27132
rect 46172 27022 46174 27074
rect 46226 27022 46228 27074
rect 45948 26852 46116 26908
rect 44716 24612 44772 24622
rect 44716 24518 44772 24556
rect 44604 23548 44772 23604
rect 44604 23380 44660 23390
rect 44604 23154 44660 23324
rect 44604 23102 44606 23154
rect 44658 23102 44660 23154
rect 44604 21924 44660 23102
rect 44604 21858 44660 21868
rect 44044 19742 44046 19794
rect 44098 19742 44100 19794
rect 44044 19730 44100 19742
rect 44380 20132 44548 20188
rect 44380 19908 44436 20132
rect 44492 20020 44548 20030
rect 44492 19926 44548 19964
rect 44380 19460 44436 19852
rect 44044 19404 44436 19460
rect 44044 19124 44100 19404
rect 44716 19236 44772 23548
rect 44940 23492 44996 25228
rect 45836 25172 45892 26796
rect 45836 25106 45892 25116
rect 44940 23426 44996 23436
rect 45836 23492 45892 23502
rect 45892 23436 46004 23492
rect 45836 23426 45892 23436
rect 45276 23268 45332 23278
rect 44940 23156 44996 23166
rect 44940 23062 44996 23100
rect 45164 23154 45220 23166
rect 45164 23102 45166 23154
rect 45218 23102 45220 23154
rect 44828 22372 44884 22382
rect 44828 22278 44884 22316
rect 45052 22146 45108 22158
rect 45052 22094 45054 22146
rect 45106 22094 45108 22146
rect 45052 22036 45108 22094
rect 45052 19348 45108 21980
rect 45164 22148 45220 23102
rect 45276 22482 45332 23212
rect 45276 22430 45278 22482
rect 45330 22430 45332 22482
rect 45276 22418 45332 22430
rect 45836 23156 45892 23166
rect 45500 22372 45556 22382
rect 45388 22370 45556 22372
rect 45388 22318 45502 22370
rect 45554 22318 45556 22370
rect 45388 22316 45556 22318
rect 45276 22148 45332 22158
rect 45164 22092 45276 22148
rect 45164 20018 45220 22092
rect 45276 22054 45332 22092
rect 45164 19966 45166 20018
rect 45218 19966 45220 20018
rect 45164 19954 45220 19966
rect 45276 20916 45332 20926
rect 45388 20916 45444 22316
rect 45500 22306 45556 22316
rect 45836 22146 45892 23100
rect 45948 23154 46004 23436
rect 45948 23102 45950 23154
rect 46002 23102 46004 23154
rect 45948 23090 46004 23102
rect 45836 22094 45838 22146
rect 45890 22094 45892 22146
rect 45836 22082 45892 22094
rect 45948 22258 46004 22270
rect 45948 22206 45950 22258
rect 46002 22206 46004 22258
rect 45948 22148 46004 22206
rect 45948 22082 46004 22092
rect 45276 20914 45444 20916
rect 45276 20862 45278 20914
rect 45330 20862 45444 20914
rect 45276 20860 45444 20862
rect 45948 21028 46004 21038
rect 44044 19058 44100 19068
rect 44604 19180 44772 19236
rect 44828 19292 45108 19348
rect 43932 19012 43988 19022
rect 43932 18918 43988 18956
rect 43820 18610 43876 18620
rect 43596 18284 43764 18340
rect 43596 17778 43652 18284
rect 44604 18004 44660 19180
rect 44716 19012 44772 19022
rect 44716 18918 44772 18956
rect 44604 17938 44660 17948
rect 43596 17726 43598 17778
rect 43650 17726 43652 17778
rect 43596 17714 43652 17726
rect 43932 17780 43988 17790
rect 43932 17686 43988 17724
rect 44716 17668 44772 17678
rect 43372 17220 43428 17500
rect 44268 17666 44772 17668
rect 44268 17614 44718 17666
rect 44770 17614 44772 17666
rect 44268 17612 44772 17614
rect 43372 17164 43876 17220
rect 43372 16994 43428 17164
rect 43372 16942 43374 16994
rect 43426 16942 43428 16994
rect 43372 16930 43428 16942
rect 43708 16996 43764 17006
rect 43484 16770 43540 16782
rect 43484 16718 43486 16770
rect 43538 16718 43540 16770
rect 43484 16100 43540 16718
rect 43484 16034 43540 16044
rect 43036 14802 43092 14812
rect 43148 15092 43316 15148
rect 43708 15148 43764 16940
rect 43820 15652 43876 17164
rect 43932 16996 43988 17006
rect 44268 16996 44324 17612
rect 44716 17602 44772 17612
rect 44828 17444 44884 19292
rect 44940 19124 44996 19134
rect 44940 19030 44996 19068
rect 45052 19122 45108 19134
rect 45052 19070 45054 19122
rect 45106 19070 45108 19122
rect 45052 18340 45108 19070
rect 45276 18452 45332 20860
rect 45388 20580 45444 20590
rect 45388 19908 45444 20524
rect 45836 20578 45892 20590
rect 45836 20526 45838 20578
rect 45890 20526 45892 20578
rect 45500 20356 45556 20366
rect 45836 20356 45892 20526
rect 45556 20300 45892 20356
rect 45500 20290 45556 20300
rect 45612 20130 45668 20300
rect 45612 20078 45614 20130
rect 45666 20078 45668 20130
rect 45612 20066 45668 20078
rect 45388 19852 45668 19908
rect 45500 19236 45556 19246
rect 45500 18564 45556 19180
rect 45500 18498 45556 18508
rect 45276 18386 45332 18396
rect 45052 18338 45220 18340
rect 45052 18286 45054 18338
rect 45106 18286 45220 18338
rect 45052 18284 45220 18286
rect 45052 18274 45108 18284
rect 45052 17444 45108 17454
rect 44828 17442 45108 17444
rect 44828 17390 45054 17442
rect 45106 17390 45108 17442
rect 44828 17388 45108 17390
rect 45052 17332 45108 17388
rect 45052 17266 45108 17276
rect 43932 16994 44324 16996
rect 43932 16942 43934 16994
rect 43986 16942 44270 16994
rect 44322 16942 44324 16994
rect 43932 16940 44324 16942
rect 43932 16930 43988 16940
rect 44268 16930 44324 16940
rect 44940 17108 44996 17118
rect 44828 16884 44884 16894
rect 44828 16098 44884 16828
rect 44940 16882 44996 17052
rect 44940 16830 44942 16882
rect 44994 16830 44996 16882
rect 44940 16818 44996 16830
rect 45164 16772 45220 18284
rect 45276 17442 45332 17454
rect 45276 17390 45278 17442
rect 45330 17390 45332 17442
rect 45276 16996 45332 17390
rect 45388 17444 45444 17454
rect 45388 17350 45444 17388
rect 45500 17442 45556 17454
rect 45500 17390 45502 17442
rect 45554 17390 45556 17442
rect 45276 16930 45332 16940
rect 45164 16678 45220 16716
rect 44828 16046 44830 16098
rect 44882 16046 44884 16098
rect 44828 16034 44884 16046
rect 45052 16100 45108 16110
rect 45052 16006 45108 16044
rect 45500 16098 45556 17390
rect 45612 17332 45668 19852
rect 45836 19794 45892 19806
rect 45836 19742 45838 19794
rect 45890 19742 45892 19794
rect 45724 18452 45780 18462
rect 45836 18452 45892 19742
rect 45948 18788 46004 20972
rect 46060 20804 46116 26852
rect 46172 26514 46228 27022
rect 46396 26908 46452 29372
rect 46508 29204 46564 29214
rect 47180 29204 47236 29374
rect 47628 29426 47684 29438
rect 47628 29374 47630 29426
rect 47682 29374 47684 29426
rect 47516 29204 47572 29214
rect 47180 29202 47572 29204
rect 47180 29150 47518 29202
rect 47570 29150 47572 29202
rect 47180 29148 47572 29150
rect 46508 28084 46564 29148
rect 47516 29138 47572 29148
rect 47628 28868 47684 29374
rect 47404 28812 47684 28868
rect 46956 28642 47012 28654
rect 46956 28590 46958 28642
rect 47010 28590 47012 28642
rect 46956 28532 47012 28590
rect 47180 28532 47236 28542
rect 46956 28530 47236 28532
rect 46956 28478 47182 28530
rect 47234 28478 47236 28530
rect 46956 28476 47236 28478
rect 46508 28082 46676 28084
rect 46508 28030 46510 28082
rect 46562 28030 46676 28082
rect 46508 28028 46676 28030
rect 46508 28018 46564 28028
rect 46172 26462 46174 26514
rect 46226 26462 46228 26514
rect 46172 26450 46228 26462
rect 46284 26852 46452 26908
rect 46508 27074 46564 27086
rect 46508 27022 46510 27074
rect 46562 27022 46564 27074
rect 46508 26852 46564 27022
rect 46172 23044 46228 23054
rect 46172 22372 46228 22988
rect 46172 22278 46228 22316
rect 46172 21588 46228 21598
rect 46172 21474 46228 21532
rect 46172 21422 46174 21474
rect 46226 21422 46228 21474
rect 46172 21410 46228 21422
rect 46284 21028 46340 26852
rect 46508 26786 46564 26796
rect 46620 26516 46676 28028
rect 46844 27748 46900 27758
rect 46844 27298 46900 27692
rect 46844 27246 46846 27298
rect 46898 27246 46900 27298
rect 46844 27234 46900 27246
rect 46732 27188 46788 27198
rect 46732 26962 46788 27132
rect 46732 26910 46734 26962
rect 46786 26910 46788 26962
rect 46732 26898 46788 26910
rect 46844 26516 46900 26526
rect 46620 26514 46900 26516
rect 46620 26462 46846 26514
rect 46898 26462 46900 26514
rect 46620 26460 46900 26462
rect 46844 26450 46900 26460
rect 46620 26178 46676 26190
rect 46620 26126 46622 26178
rect 46674 26126 46676 26178
rect 46620 25956 46676 26126
rect 46620 25890 46676 25900
rect 46844 25172 46900 25182
rect 46844 24610 46900 25116
rect 46956 25060 47012 28476
rect 47180 28466 47236 28476
rect 47292 28420 47348 28430
rect 47404 28420 47460 28812
rect 47516 28644 47572 28654
rect 47740 28644 47796 29596
rect 47852 29650 47908 30044
rect 47852 29598 47854 29650
rect 47906 29598 47908 29650
rect 47852 29586 47908 29598
rect 48076 29652 48132 30942
rect 48076 29586 48132 29596
rect 48412 30324 48468 30334
rect 48412 30098 48468 30268
rect 48412 30046 48414 30098
rect 48466 30046 48468 30098
rect 48412 29652 48468 30046
rect 48412 29586 48468 29596
rect 47964 29540 48020 29550
rect 47852 28756 47908 28766
rect 47964 28756 48020 29484
rect 47908 28700 48020 28756
rect 47852 28662 47908 28700
rect 47516 28642 47796 28644
rect 47516 28590 47518 28642
rect 47570 28590 47796 28642
rect 47516 28588 47796 28590
rect 47516 28578 47572 28588
rect 47292 28418 47460 28420
rect 47292 28366 47294 28418
rect 47346 28366 47460 28418
rect 47292 28364 47460 28366
rect 47292 26908 47348 28364
rect 48076 27860 48132 27870
rect 48076 27766 48132 27804
rect 47964 27748 48020 27758
rect 47964 27654 48020 27692
rect 47404 27186 47460 27198
rect 47404 27134 47406 27186
rect 47458 27134 47460 27186
rect 47404 27076 47460 27134
rect 47404 27010 47460 27020
rect 47740 27188 47796 27198
rect 47740 27074 47796 27132
rect 48524 27188 48580 27198
rect 48524 27094 48580 27132
rect 47740 27022 47742 27074
rect 47794 27022 47796 27074
rect 47740 27010 47796 27022
rect 47068 26852 47348 26908
rect 48188 26964 48244 27002
rect 47068 26292 47124 26852
rect 47180 26516 47236 26526
rect 47740 26516 47796 26526
rect 48076 26516 48132 26526
rect 47180 26514 47908 26516
rect 47180 26462 47182 26514
rect 47234 26462 47742 26514
rect 47794 26462 47908 26514
rect 47180 26460 47908 26462
rect 47180 26450 47236 26460
rect 47740 26450 47796 26460
rect 47068 26226 47124 26236
rect 47740 26292 47796 26302
rect 47740 25618 47796 26236
rect 47852 26180 47908 26460
rect 48076 26422 48132 26460
rect 48188 26514 48244 26908
rect 48188 26462 48190 26514
rect 48242 26462 48244 26514
rect 48188 26450 48244 26462
rect 47964 26402 48020 26414
rect 47964 26350 47966 26402
rect 48018 26350 48020 26402
rect 47964 26292 48020 26350
rect 48412 26404 48468 26414
rect 48076 26292 48132 26302
rect 47964 26236 48076 26292
rect 48076 26226 48132 26236
rect 47852 26124 48020 26180
rect 47740 25566 47742 25618
rect 47794 25566 47796 25618
rect 47740 25554 47796 25566
rect 46956 24994 47012 25004
rect 47852 24722 47908 24734
rect 47852 24670 47854 24722
rect 47906 24670 47908 24722
rect 46844 24558 46846 24610
rect 46898 24558 46900 24610
rect 46844 24546 46900 24558
rect 47292 24610 47348 24622
rect 47292 24558 47294 24610
rect 47346 24558 47348 24610
rect 47292 23940 47348 24558
rect 47292 23874 47348 23884
rect 46844 23828 46900 23838
rect 46396 23380 46452 23390
rect 46396 23154 46452 23324
rect 46396 23102 46398 23154
rect 46450 23102 46452 23154
rect 46396 23090 46452 23102
rect 46844 23154 46900 23772
rect 46956 23828 47012 23838
rect 47852 23828 47908 24670
rect 47964 24612 48020 26124
rect 48076 25956 48132 25966
rect 48076 24946 48132 25900
rect 48076 24894 48078 24946
rect 48130 24894 48132 24946
rect 48076 24882 48132 24894
rect 48188 24836 48244 24846
rect 48188 24742 48244 24780
rect 47964 24556 48244 24612
rect 46956 23826 47124 23828
rect 46956 23774 46958 23826
rect 47010 23774 47124 23826
rect 46956 23772 47124 23774
rect 46956 23762 47012 23772
rect 46844 23102 46846 23154
rect 46898 23102 46900 23154
rect 46844 23090 46900 23102
rect 47068 23604 47124 23772
rect 47852 23762 47908 23772
rect 47068 22370 47124 23548
rect 47852 23268 47908 23278
rect 47852 23174 47908 23212
rect 47964 23268 48020 23278
rect 47964 23266 48132 23268
rect 47964 23214 47966 23266
rect 48018 23214 48132 23266
rect 47964 23212 48132 23214
rect 47964 23202 48020 23212
rect 47292 23156 47348 23166
rect 47292 23062 47348 23100
rect 47516 23154 47572 23166
rect 47516 23102 47518 23154
rect 47570 23102 47572 23154
rect 47404 23042 47460 23054
rect 47404 22990 47406 23042
rect 47458 22990 47460 23042
rect 47404 22596 47460 22990
rect 47516 22932 47572 23102
rect 47964 22932 48020 22942
rect 47516 22930 48020 22932
rect 47516 22878 47966 22930
rect 48018 22878 48020 22930
rect 47516 22876 48020 22878
rect 47964 22866 48020 22876
rect 47404 22540 47908 22596
rect 47852 22482 47908 22540
rect 47852 22430 47854 22482
rect 47906 22430 47908 22482
rect 47852 22418 47908 22430
rect 47068 22318 47070 22370
rect 47122 22318 47124 22370
rect 46508 22148 46564 22158
rect 46508 21810 46564 22092
rect 46620 22146 46676 22158
rect 46620 22094 46622 22146
rect 46674 22094 46676 22146
rect 46620 22036 46676 22094
rect 46620 21970 46676 21980
rect 46508 21758 46510 21810
rect 46562 21758 46564 21810
rect 46508 21746 46564 21758
rect 46844 21588 46900 21598
rect 46844 21494 46900 21532
rect 46284 20962 46340 20972
rect 46060 20748 46564 20804
rect 46284 20580 46340 20590
rect 46284 20578 46452 20580
rect 46284 20526 46286 20578
rect 46338 20526 46452 20578
rect 46284 20524 46452 20526
rect 46284 20514 46340 20524
rect 46284 20020 46340 20030
rect 46060 19908 46116 19918
rect 46060 19814 46116 19852
rect 46172 19122 46228 19134
rect 46172 19070 46174 19122
rect 46226 19070 46228 19122
rect 45948 18732 46116 18788
rect 45724 18450 45892 18452
rect 45724 18398 45726 18450
rect 45778 18398 45892 18450
rect 45724 18396 45892 18398
rect 45948 18562 46004 18574
rect 45948 18510 45950 18562
rect 46002 18510 46004 18562
rect 45724 18228 45780 18396
rect 45724 18162 45780 18172
rect 45948 17780 46004 18510
rect 45724 17724 46004 17780
rect 45724 17556 45780 17724
rect 45724 17462 45780 17500
rect 45836 17556 45892 17566
rect 46060 17556 46116 18732
rect 46172 18452 46228 19070
rect 46284 19122 46340 19964
rect 46396 19794 46452 20524
rect 46396 19742 46398 19794
rect 46450 19742 46452 19794
rect 46396 19730 46452 19742
rect 46508 20244 46564 20748
rect 46844 20580 46900 20590
rect 46844 20486 46900 20524
rect 46284 19070 46286 19122
rect 46338 19070 46340 19122
rect 46284 18676 46340 19070
rect 46396 19236 46452 19246
rect 46508 19236 46564 20188
rect 46844 20130 46900 20142
rect 46844 20078 46846 20130
rect 46898 20078 46900 20130
rect 46396 19234 46564 19236
rect 46396 19182 46398 19234
rect 46450 19182 46564 19234
rect 46396 19180 46564 19182
rect 46620 19794 46676 19806
rect 46620 19742 46622 19794
rect 46674 19742 46676 19794
rect 46396 19012 46452 19180
rect 46396 18946 46452 18956
rect 46620 18676 46676 19742
rect 46844 19012 46900 20078
rect 46956 19794 47012 19806
rect 46956 19742 46958 19794
rect 47010 19742 47012 19794
rect 46956 19124 47012 19742
rect 47068 19236 47124 22318
rect 47516 22372 47572 22382
rect 47516 21810 47572 22316
rect 47516 21758 47518 21810
rect 47570 21758 47572 21810
rect 47516 21746 47572 21758
rect 47852 21812 47908 21822
rect 48076 21812 48132 23212
rect 47852 21810 48132 21812
rect 47852 21758 47854 21810
rect 47906 21758 48132 21810
rect 47852 21756 48132 21758
rect 47852 21746 47908 21756
rect 47292 21698 47348 21710
rect 47292 21646 47294 21698
rect 47346 21646 47348 21698
rect 47180 21586 47236 21598
rect 47180 21534 47182 21586
rect 47234 21534 47236 21586
rect 47180 20580 47236 21534
rect 47292 21588 47348 21646
rect 47292 21522 47348 21532
rect 47852 20804 47908 20814
rect 47404 20748 47796 20804
rect 47180 20514 47236 20524
rect 47292 20580 47348 20590
rect 47404 20580 47460 20748
rect 47740 20690 47796 20748
rect 47852 20710 47908 20748
rect 47740 20638 47742 20690
rect 47794 20638 47796 20690
rect 47740 20626 47796 20638
rect 47292 20578 47460 20580
rect 47292 20526 47294 20578
rect 47346 20526 47460 20578
rect 47292 20524 47460 20526
rect 47516 20578 47572 20590
rect 47516 20526 47518 20578
rect 47570 20526 47572 20578
rect 47292 19908 47348 20524
rect 47404 20244 47460 20254
rect 47516 20244 47572 20526
rect 47404 20242 47572 20244
rect 47404 20190 47406 20242
rect 47458 20190 47572 20242
rect 47404 20188 47572 20190
rect 47404 20178 47460 20188
rect 47740 20132 48020 20188
rect 47740 20130 47796 20132
rect 47740 20078 47742 20130
rect 47794 20078 47796 20130
rect 47740 20066 47796 20078
rect 47292 19842 47348 19852
rect 47628 20018 47684 20030
rect 47628 19966 47630 20018
rect 47682 19966 47684 20018
rect 47628 19684 47684 19966
rect 47628 19618 47684 19628
rect 47852 20018 47908 20030
rect 47852 19966 47854 20018
rect 47906 19966 47908 20018
rect 47740 19348 47796 19358
rect 47628 19292 47740 19348
rect 47180 19236 47236 19246
rect 47068 19234 47236 19236
rect 47068 19182 47182 19234
rect 47234 19182 47236 19234
rect 47068 19180 47236 19182
rect 47180 19170 47236 19180
rect 46956 19068 47124 19124
rect 46844 19010 47012 19012
rect 46844 18958 46846 19010
rect 46898 18958 47012 19010
rect 46844 18956 47012 18958
rect 46844 18946 46900 18956
rect 46284 18620 46452 18676
rect 46620 18620 46788 18676
rect 46396 18564 46452 18620
rect 46396 18508 46676 18564
rect 46284 18452 46340 18462
rect 46172 18450 46340 18452
rect 46172 18398 46286 18450
rect 46338 18398 46340 18450
rect 46172 18396 46340 18398
rect 46284 18340 46340 18396
rect 46284 18274 46340 18284
rect 46620 18450 46676 18508
rect 46620 18398 46622 18450
rect 46674 18398 46676 18450
rect 46620 18116 46676 18398
rect 46732 18338 46788 18620
rect 46732 18286 46734 18338
rect 46786 18286 46788 18338
rect 46732 18274 46788 18286
rect 46844 18564 46900 18574
rect 46844 18228 46900 18508
rect 46956 18452 47012 18956
rect 47068 18676 47124 19068
rect 47068 18610 47124 18620
rect 47404 18452 47460 18462
rect 46956 18450 47460 18452
rect 46956 18398 47406 18450
rect 47458 18398 47460 18450
rect 46956 18396 47460 18398
rect 47404 18386 47460 18396
rect 47516 18340 47572 18350
rect 47516 18228 47572 18284
rect 46844 18172 47236 18228
rect 46620 18060 46788 18116
rect 46620 17892 46676 17902
rect 46732 17892 46788 18060
rect 46956 18004 47012 18014
rect 46732 17836 46900 17892
rect 46396 17780 46452 17790
rect 46396 17686 46452 17724
rect 45836 17554 46116 17556
rect 45836 17502 45838 17554
rect 45890 17502 46116 17554
rect 45836 17500 46116 17502
rect 45836 17490 45892 17500
rect 45612 17276 45780 17332
rect 45500 16046 45502 16098
rect 45554 16046 45556 16098
rect 45500 16034 45556 16046
rect 45612 16772 45668 16782
rect 45612 16658 45668 16716
rect 45612 16606 45614 16658
rect 45666 16606 45668 16658
rect 45612 16100 45668 16606
rect 45612 16034 45668 16044
rect 44940 15874 44996 15886
rect 44940 15822 44942 15874
rect 44994 15822 44996 15874
rect 43820 15596 44100 15652
rect 43932 15428 43988 15438
rect 43820 15372 43932 15428
rect 43820 15314 43876 15372
rect 43932 15362 43988 15372
rect 43820 15262 43822 15314
rect 43874 15262 43876 15314
rect 43820 15250 43876 15262
rect 43708 15092 43988 15148
rect 43036 14644 43092 14654
rect 43036 13972 43092 14588
rect 43036 13878 43092 13916
rect 42924 13692 43092 13748
rect 42588 12310 42644 12348
rect 42812 12178 42868 12190
rect 42812 12126 42814 12178
rect 42866 12126 42868 12178
rect 42812 12068 42868 12126
rect 42812 11620 42868 12012
rect 42476 11564 42868 11620
rect 42476 11172 42532 11564
rect 42588 11396 42644 11406
rect 42644 11340 42756 11396
rect 42588 11302 42644 11340
rect 42476 11116 42644 11172
rect 42252 10782 42254 10834
rect 42306 10782 42308 10834
rect 42252 10770 42308 10782
rect 41580 10434 41636 10444
rect 41916 10612 41972 10622
rect 41916 10498 41972 10556
rect 41916 10446 41918 10498
rect 41970 10446 41972 10498
rect 41916 9268 41972 10446
rect 42364 10500 42420 10510
rect 42364 10498 42532 10500
rect 42364 10446 42366 10498
rect 42418 10446 42532 10498
rect 42364 10444 42532 10446
rect 42364 10434 42420 10444
rect 42364 10276 42420 10286
rect 42252 10220 42364 10276
rect 42252 9938 42308 10220
rect 42364 10210 42420 10220
rect 42252 9886 42254 9938
rect 42306 9886 42308 9938
rect 42252 9874 42308 9886
rect 41916 9202 41972 9212
rect 41356 8978 41412 8988
rect 42364 9044 42420 9054
rect 42364 8950 42420 8988
rect 41468 8930 41524 8942
rect 41468 8878 41470 8930
rect 41522 8878 41524 8930
rect 41468 8260 41524 8878
rect 42476 8482 42532 10444
rect 42588 9826 42644 11116
rect 42588 9774 42590 9826
rect 42642 9774 42644 9826
rect 42588 9762 42644 9774
rect 42476 8430 42478 8482
rect 42530 8430 42532 8482
rect 42476 8418 42532 8430
rect 42700 8370 42756 11340
rect 42924 11394 42980 11406
rect 42924 11342 42926 11394
rect 42978 11342 42980 11394
rect 42812 10276 42868 10286
rect 42812 9828 42868 10220
rect 42924 9940 42980 11342
rect 43036 11394 43092 13692
rect 43148 12068 43204 15092
rect 43484 14308 43540 14318
rect 43484 14214 43540 14252
rect 43484 13972 43540 13982
rect 43484 13878 43540 13916
rect 43932 13636 43988 15092
rect 44044 14642 44100 15596
rect 44940 15428 44996 15822
rect 44940 15362 44996 15372
rect 45164 15204 45220 15214
rect 45724 15148 45780 17276
rect 46060 17108 46116 17500
rect 45836 16994 45892 17006
rect 45836 16942 45838 16994
rect 45890 16942 45892 16994
rect 45836 16100 45892 16942
rect 46060 16772 46116 17052
rect 46284 17444 46340 17454
rect 46284 16994 46340 17388
rect 46396 17220 46452 17230
rect 46396 17108 46452 17164
rect 46620 17108 46676 17836
rect 46732 17442 46788 17454
rect 46732 17390 46734 17442
rect 46786 17390 46788 17442
rect 46732 17332 46788 17390
rect 46732 17266 46788 17276
rect 46396 17106 46676 17108
rect 46396 17054 46398 17106
rect 46450 17054 46676 17106
rect 46396 17052 46676 17054
rect 46396 17042 46452 17052
rect 46284 16942 46286 16994
rect 46338 16942 46340 16994
rect 46284 16930 46340 16942
rect 46620 16884 46676 16894
rect 46620 16790 46676 16828
rect 46060 16716 46340 16772
rect 45948 16660 46004 16670
rect 45948 16658 46228 16660
rect 45948 16606 45950 16658
rect 46002 16606 46228 16658
rect 45948 16604 46228 16606
rect 45948 16594 46004 16604
rect 45836 16098 46004 16100
rect 45836 16046 45838 16098
rect 45890 16046 46004 16098
rect 45836 16044 46004 16046
rect 45836 16034 45892 16044
rect 44044 14590 44046 14642
rect 44098 14590 44100 14642
rect 44044 14578 44100 14590
rect 44828 14644 44884 14654
rect 44828 14530 44884 14588
rect 44828 14478 44830 14530
rect 44882 14478 44884 14530
rect 44828 14466 44884 14478
rect 45164 14530 45220 15148
rect 45500 15092 45780 15148
rect 45948 15202 46004 16044
rect 45948 15150 45950 15202
rect 46002 15150 46004 15202
rect 45948 15138 46004 15150
rect 46060 15876 46116 15886
rect 45500 14644 45556 15092
rect 45500 14550 45556 14588
rect 45164 14478 45166 14530
rect 45218 14478 45220 14530
rect 45164 14466 45220 14478
rect 45948 14418 46004 14430
rect 45948 14366 45950 14418
rect 46002 14366 46004 14418
rect 44940 14306 44996 14318
rect 44940 14254 44942 14306
rect 44994 14254 44996 14306
rect 44940 14084 44996 14254
rect 44492 14028 44996 14084
rect 44492 13972 44548 14028
rect 43820 13634 43988 13636
rect 43820 13582 43934 13634
rect 43986 13582 43988 13634
rect 43820 13580 43988 13582
rect 43260 12068 43316 12078
rect 43148 12012 43260 12068
rect 43260 11974 43316 12012
rect 43036 11342 43038 11394
rect 43090 11342 43092 11394
rect 43036 10276 43092 11342
rect 43036 10210 43092 10220
rect 43596 10164 43652 10174
rect 43036 9940 43092 9950
rect 42924 9938 43428 9940
rect 42924 9886 43038 9938
rect 43090 9886 43428 9938
rect 42924 9884 43428 9886
rect 43036 9874 43092 9884
rect 42812 9772 42980 9828
rect 42924 9156 42980 9772
rect 42924 9100 43204 9156
rect 43036 8932 43092 8942
rect 42700 8318 42702 8370
rect 42754 8318 42756 8370
rect 42700 8306 42756 8318
rect 42812 8930 43092 8932
rect 42812 8878 43038 8930
rect 43090 8878 43092 8930
rect 42812 8876 43092 8878
rect 41804 8260 41860 8270
rect 41468 8194 41524 8204
rect 41692 8258 41860 8260
rect 41692 8206 41806 8258
rect 41858 8206 41860 8258
rect 41692 8204 41860 8206
rect 40908 3442 41076 3444
rect 40908 3390 40910 3442
rect 40962 3390 41076 3442
rect 40908 3388 41076 3390
rect 41132 4226 41188 4238
rect 41132 4174 41134 4226
rect 41186 4174 41188 4226
rect 41132 3444 41188 4174
rect 41244 3444 41300 3454
rect 41132 3442 41300 3444
rect 41132 3390 41246 3442
rect 41298 3390 41300 3442
rect 41132 3388 41300 3390
rect 40908 3378 40964 3388
rect 41244 2548 41300 3388
rect 41580 3444 41636 3454
rect 41692 3444 41748 8204
rect 41804 8194 41860 8204
rect 42364 8260 42420 8270
rect 42364 8166 42420 8204
rect 42812 7812 42868 8876
rect 43036 8866 43092 8876
rect 43148 8484 43204 9100
rect 42924 8428 43204 8484
rect 42924 8258 42980 8428
rect 42924 8206 42926 8258
rect 42978 8206 42980 8258
rect 42924 8194 42980 8206
rect 43372 8148 43428 9884
rect 43372 8082 43428 8092
rect 43596 8260 43652 10108
rect 42252 7756 42868 7812
rect 42252 7698 42308 7756
rect 42252 7646 42254 7698
rect 42306 7646 42308 7698
rect 42252 7634 42308 7646
rect 42924 7474 42980 7486
rect 42924 7422 42926 7474
rect 42978 7422 42980 7474
rect 42140 7362 42196 7374
rect 42140 7310 42142 7362
rect 42194 7310 42196 7362
rect 42140 7252 42196 7310
rect 42140 7186 42196 7196
rect 42588 6132 42644 6142
rect 42588 6038 42644 6076
rect 41580 3442 41748 3444
rect 41580 3390 41582 3442
rect 41634 3390 41748 3442
rect 41580 3388 41748 3390
rect 42364 3444 42420 3454
rect 42588 3444 42644 3454
rect 42364 3442 42644 3444
rect 42364 3390 42366 3442
rect 42418 3390 42590 3442
rect 42642 3390 42644 3442
rect 42364 3388 42644 3390
rect 41580 3378 41636 3388
rect 41020 2492 41300 2548
rect 41020 800 41076 2492
rect 42364 800 42420 3388
rect 42588 3378 42644 3388
rect 42924 3442 42980 7422
rect 43372 7476 43428 7486
rect 43596 7476 43652 8204
rect 43820 8258 43876 13580
rect 43932 13570 43988 13580
rect 44268 13970 44548 13972
rect 44268 13918 44494 13970
rect 44546 13918 44548 13970
rect 44268 13916 44548 13918
rect 44268 13074 44324 13916
rect 44492 13906 44548 13916
rect 45612 13748 45668 13758
rect 45948 13748 46004 14366
rect 45668 13692 46004 13748
rect 46060 14418 46116 15820
rect 46172 15652 46228 16604
rect 46284 16324 46340 16716
rect 46284 16268 46788 16324
rect 46284 16210 46340 16268
rect 46284 16158 46286 16210
rect 46338 16158 46340 16210
rect 46284 16146 46340 16158
rect 46732 16212 46788 16268
rect 46620 16100 46676 16110
rect 46620 16006 46676 16044
rect 46732 15986 46788 16156
rect 46732 15934 46734 15986
rect 46786 15934 46788 15986
rect 46732 15922 46788 15934
rect 46172 15596 46676 15652
rect 46620 15314 46676 15596
rect 46620 15262 46622 15314
rect 46674 15262 46676 15314
rect 46620 15250 46676 15262
rect 46508 15204 46564 15242
rect 46508 15138 46564 15148
rect 46732 15090 46788 15102
rect 46732 15038 46734 15090
rect 46786 15038 46788 15090
rect 46284 14532 46340 14542
rect 46620 14532 46676 14542
rect 46284 14530 46676 14532
rect 46284 14478 46286 14530
rect 46338 14478 46622 14530
rect 46674 14478 46676 14530
rect 46284 14476 46676 14478
rect 46284 14466 46340 14476
rect 46620 14466 46676 14476
rect 46060 14366 46062 14418
rect 46114 14366 46116 14418
rect 45612 13654 45668 13692
rect 44268 13022 44270 13074
rect 44322 13022 44324 13074
rect 44268 13010 44324 13022
rect 44604 13076 44660 13086
rect 43932 12852 43988 12862
rect 43932 12404 43988 12796
rect 43932 12402 44324 12404
rect 43932 12350 43934 12402
rect 43986 12350 44324 12402
rect 43932 12348 44324 12350
rect 43932 12338 43988 12348
rect 44268 12290 44324 12348
rect 44604 12402 44660 13020
rect 45500 13076 45556 13086
rect 45500 12982 45556 13020
rect 45836 12962 45892 12974
rect 45836 12910 45838 12962
rect 45890 12910 45892 12962
rect 45724 12404 45780 12414
rect 44604 12350 44606 12402
rect 44658 12350 44660 12402
rect 44604 12338 44660 12350
rect 44828 12348 45220 12404
rect 44268 12238 44270 12290
rect 44322 12238 44324 12290
rect 44268 12226 44324 12238
rect 44380 12292 44436 12302
rect 44380 12290 44548 12292
rect 44380 12238 44382 12290
rect 44434 12238 44548 12290
rect 44380 12236 44548 12238
rect 44380 12226 44436 12236
rect 44492 12180 44548 12236
rect 44828 12180 44884 12348
rect 45052 12180 45108 12190
rect 44492 12124 44884 12180
rect 44940 12178 45108 12180
rect 44940 12126 45054 12178
rect 45106 12126 45108 12178
rect 44940 12124 45108 12126
rect 44380 12068 44436 12078
rect 44268 12012 44380 12068
rect 44156 11620 44212 11630
rect 44156 10164 44212 11564
rect 44268 11172 44324 12012
rect 44380 12002 44436 12012
rect 44380 11396 44436 11406
rect 44828 11396 44884 11406
rect 44436 11340 44548 11396
rect 44380 11330 44436 11340
rect 44380 11172 44436 11182
rect 44268 11170 44436 11172
rect 44268 11118 44382 11170
rect 44434 11118 44436 11170
rect 44268 11116 44436 11118
rect 44380 11106 44436 11116
rect 44156 10098 44212 10108
rect 44380 9940 44436 9950
rect 44492 9940 44548 11340
rect 44828 11302 44884 11340
rect 44940 10724 44996 12124
rect 45052 12114 45108 12124
rect 44380 9938 44548 9940
rect 44380 9886 44382 9938
rect 44434 9886 44548 9938
rect 44380 9884 44548 9886
rect 44716 10668 44996 10724
rect 45164 11394 45220 12348
rect 45500 12180 45556 12190
rect 45276 12178 45556 12180
rect 45276 12126 45502 12178
rect 45554 12126 45556 12178
rect 45276 12124 45556 12126
rect 45276 11620 45332 12124
rect 45500 12114 45556 12124
rect 45724 12066 45780 12348
rect 45724 12014 45726 12066
rect 45778 12014 45780 12066
rect 45276 11554 45332 11564
rect 45388 11954 45444 11966
rect 45388 11902 45390 11954
rect 45442 11902 45444 11954
rect 45388 11396 45444 11902
rect 45164 11342 45166 11394
rect 45218 11342 45220 11394
rect 44380 9874 44436 9884
rect 44716 8428 44772 10668
rect 43820 8206 43822 8258
rect 43874 8206 43876 8258
rect 43372 7474 43652 7476
rect 43372 7422 43374 7474
rect 43426 7422 43652 7474
rect 43372 7420 43652 7422
rect 43372 7410 43428 7420
rect 43148 7252 43204 7262
rect 43148 7158 43204 7196
rect 43372 5908 43428 5918
rect 43372 5906 43540 5908
rect 43372 5854 43374 5906
rect 43426 5854 43540 5906
rect 43372 5852 43540 5854
rect 43372 5842 43428 5852
rect 43372 4226 43428 4238
rect 43372 4174 43374 4226
rect 43426 4174 43428 4226
rect 42924 3390 42926 3442
rect 42978 3390 42980 3442
rect 42924 3378 42980 3390
rect 43036 3444 43092 3454
rect 43036 800 43092 3388
rect 43372 3444 43428 4174
rect 43484 3444 43540 5852
rect 43596 5906 43652 7420
rect 43708 7700 43764 7710
rect 43708 7362 43764 7644
rect 43820 7474 43876 8206
rect 44380 8372 44772 8428
rect 44828 10500 44884 10510
rect 44828 9826 44884 10444
rect 44828 9774 44830 9826
rect 44882 9774 44884 9826
rect 44828 9044 44884 9774
rect 44828 8428 44884 8988
rect 45164 8932 45220 11342
rect 45276 11340 45444 11396
rect 45276 10948 45332 11340
rect 45500 11284 45556 11294
rect 45500 11190 45556 11228
rect 45388 11172 45444 11182
rect 45388 11078 45444 11116
rect 45276 10892 45556 10948
rect 45500 9154 45556 10892
rect 45612 9714 45668 9726
rect 45612 9662 45614 9714
rect 45666 9662 45668 9714
rect 45612 9266 45668 9662
rect 45612 9214 45614 9266
rect 45666 9214 45668 9266
rect 45612 9202 45668 9214
rect 45500 9102 45502 9154
rect 45554 9102 45556 9154
rect 45500 9090 45556 9102
rect 45724 9044 45780 12014
rect 45836 12404 45892 12910
rect 45948 12404 46004 12414
rect 45836 12348 45948 12404
rect 45836 11172 45892 12348
rect 45948 12338 46004 12348
rect 46060 12180 46116 14366
rect 46732 13860 46788 15038
rect 46844 13972 46900 17836
rect 46956 17106 47012 17948
rect 47180 17332 47236 18172
rect 47292 18172 47572 18228
rect 47292 17666 47348 18172
rect 47628 17892 47684 19292
rect 47740 19282 47796 19292
rect 47852 18674 47908 19966
rect 47964 19346 48020 20132
rect 47964 19294 47966 19346
rect 48018 19294 48020 19346
rect 47964 19282 48020 19294
rect 48076 19348 48132 21756
rect 48076 19282 48132 19292
rect 48188 19124 48244 24556
rect 48412 21252 48468 26348
rect 48412 21186 48468 21196
rect 48524 26180 48580 26190
rect 48524 21028 48580 26124
rect 47852 18622 47854 18674
rect 47906 18622 47908 18674
rect 47852 18610 47908 18622
rect 47964 19068 48244 19124
rect 48300 20972 48580 21028
rect 48300 20914 48356 20972
rect 48300 20862 48302 20914
rect 48354 20862 48356 20914
rect 47292 17614 47294 17666
rect 47346 17614 47348 17666
rect 47292 17602 47348 17614
rect 47516 17836 47628 17892
rect 47404 17556 47460 17566
rect 47404 17462 47460 17500
rect 47180 17276 47460 17332
rect 46956 17054 46958 17106
rect 47010 17054 47012 17106
rect 46956 17042 47012 17054
rect 47404 17106 47460 17276
rect 47404 17054 47406 17106
rect 47458 17054 47460 17106
rect 47404 17042 47460 17054
rect 47516 16884 47572 17836
rect 47628 17826 47684 17836
rect 47740 18450 47796 18462
rect 47740 18398 47742 18450
rect 47794 18398 47796 18450
rect 47740 17668 47796 18398
rect 47740 17602 47796 17612
rect 47628 17444 47684 17454
rect 47628 17350 47684 17388
rect 47964 17442 48020 19068
rect 48076 18676 48132 18686
rect 48076 18452 48132 18620
rect 48076 18450 48244 18452
rect 48076 18398 48078 18450
rect 48130 18398 48244 18450
rect 48076 18396 48244 18398
rect 48076 18386 48132 18396
rect 48188 18004 48244 18396
rect 48300 18340 48356 20862
rect 48300 18274 48356 18284
rect 48188 17948 48468 18004
rect 48412 17892 48468 17948
rect 48188 17668 48244 17678
rect 48188 17574 48244 17612
rect 48412 17666 48468 17836
rect 48412 17614 48414 17666
rect 48466 17614 48468 17666
rect 48412 17602 48468 17614
rect 47964 17390 47966 17442
rect 48018 17390 48020 17442
rect 47404 16828 47572 16884
rect 47292 16212 47348 16222
rect 47292 16118 47348 16156
rect 46956 15876 47012 15886
rect 46956 15874 47236 15876
rect 46956 15822 46958 15874
rect 47010 15822 47236 15874
rect 46956 15820 47236 15822
rect 46956 15810 47012 15820
rect 47180 15316 47236 15820
rect 47404 15428 47460 16828
rect 47852 16772 47908 16782
rect 47740 16770 47908 16772
rect 47740 16718 47854 16770
rect 47906 16718 47908 16770
rect 47740 16716 47908 16718
rect 47740 16212 47796 16716
rect 47852 16706 47908 16716
rect 47740 16146 47796 16156
rect 47628 16098 47684 16110
rect 47628 16046 47630 16098
rect 47682 16046 47684 16098
rect 47628 15764 47684 16046
rect 47628 15698 47684 15708
rect 47852 16098 47908 16110
rect 47852 16046 47854 16098
rect 47906 16046 47908 16098
rect 47852 15540 47908 16046
rect 47404 15362 47460 15372
rect 47516 15484 47852 15540
rect 47292 15316 47348 15326
rect 47180 15314 47348 15316
rect 47180 15262 47294 15314
rect 47346 15262 47348 15314
rect 47180 15260 47348 15262
rect 47292 15250 47348 15260
rect 47516 14642 47572 15484
rect 47852 15474 47908 15484
rect 47964 15316 48020 17390
rect 48076 17556 48132 17566
rect 48076 15988 48132 17500
rect 48300 17442 48356 17454
rect 48300 17390 48302 17442
rect 48354 17390 48356 17442
rect 48300 17108 48356 17390
rect 48300 17042 48356 17052
rect 48412 16660 48468 16670
rect 48412 16100 48468 16604
rect 48412 16006 48468 16044
rect 48076 15652 48132 15932
rect 48188 15876 48244 15886
rect 48188 15874 48356 15876
rect 48188 15822 48190 15874
rect 48242 15822 48356 15874
rect 48188 15820 48356 15822
rect 48188 15810 48244 15820
rect 48076 15596 48244 15652
rect 48076 15428 48132 15438
rect 48076 15334 48132 15372
rect 47516 14590 47518 14642
rect 47570 14590 47572 14642
rect 47516 14578 47572 14590
rect 47852 15260 48020 15316
rect 47068 14532 47124 14542
rect 47068 14438 47124 14476
rect 47852 13972 47908 15260
rect 47964 15092 48020 15102
rect 47964 14530 48020 15036
rect 47964 14478 47966 14530
rect 48018 14478 48020 14530
rect 47964 14466 48020 14478
rect 48188 14308 48244 15596
rect 46844 13916 47348 13972
rect 46620 13804 46732 13860
rect 45836 11106 45892 11116
rect 45948 12178 46116 12180
rect 45948 12126 46062 12178
rect 46114 12126 46116 12178
rect 45948 12124 46116 12126
rect 45948 11060 46004 12124
rect 46060 12114 46116 12124
rect 46172 13746 46228 13758
rect 46172 13694 46174 13746
rect 46226 13694 46228 13746
rect 46172 11506 46228 13694
rect 46284 13524 46340 13534
rect 46284 12962 46340 13468
rect 46284 12910 46286 12962
rect 46338 12910 46340 12962
rect 46284 12898 46340 12910
rect 46620 12962 46676 13804
rect 46732 13766 46788 13804
rect 47068 13746 47124 13758
rect 47068 13694 47070 13746
rect 47122 13694 47124 13746
rect 46732 13636 46788 13646
rect 47068 13636 47124 13694
rect 46732 13542 46788 13580
rect 46844 13580 47068 13636
rect 46844 13524 46900 13580
rect 47068 13570 47124 13580
rect 46844 13186 46900 13468
rect 46844 13134 46846 13186
rect 46898 13134 46900 13186
rect 46844 13122 46900 13134
rect 46620 12910 46622 12962
rect 46674 12910 46676 12962
rect 46620 12898 46676 12910
rect 47180 12852 47236 12862
rect 47180 12758 47236 12796
rect 46172 11454 46174 11506
rect 46226 11454 46228 11506
rect 46172 11442 46228 11454
rect 46508 12404 46564 12414
rect 46508 11508 46564 12348
rect 47292 12178 47348 13916
rect 47852 13878 47908 13916
rect 47964 14252 48244 14308
rect 47628 13860 47684 13870
rect 47628 13766 47684 13804
rect 47404 13746 47460 13758
rect 47404 13694 47406 13746
rect 47458 13694 47460 13746
rect 47404 13636 47460 13694
rect 47404 13570 47460 13580
rect 47516 13634 47572 13646
rect 47516 13582 47518 13634
rect 47570 13582 47572 13634
rect 47516 12962 47572 13582
rect 47516 12910 47518 12962
rect 47570 12910 47572 12962
rect 47516 12898 47572 12910
rect 47740 12852 47796 12862
rect 47740 12758 47796 12796
rect 47292 12126 47294 12178
rect 47346 12126 47348 12178
rect 46508 11506 46676 11508
rect 46508 11454 46510 11506
rect 46562 11454 46676 11506
rect 46508 11452 46676 11454
rect 46508 11442 46564 11452
rect 46060 11284 46116 11294
rect 46060 11190 46116 11228
rect 45948 11004 46228 11060
rect 45052 8930 45220 8932
rect 45052 8878 45166 8930
rect 45218 8878 45220 8930
rect 45052 8876 45220 8878
rect 44828 8372 44996 8428
rect 43820 7422 43822 7474
rect 43874 7422 43876 7474
rect 43820 7410 43876 7422
rect 44268 8148 44324 8158
rect 43708 7310 43710 7362
rect 43762 7310 43764 7362
rect 43708 6132 43764 7310
rect 44268 7364 44324 8092
rect 44268 7298 44324 7308
rect 43764 6076 43876 6132
rect 43708 6066 43764 6076
rect 43596 5854 43598 5906
rect 43650 5854 43652 5906
rect 43596 5842 43652 5854
rect 43820 5794 43876 6076
rect 43820 5742 43822 5794
rect 43874 5742 43876 5794
rect 43820 5730 43876 5742
rect 44044 4226 44100 4238
rect 44044 4174 44046 4226
rect 44098 4174 44100 4226
rect 43596 3444 43652 3454
rect 43484 3442 43652 3444
rect 43484 3390 43598 3442
rect 43650 3390 43652 3442
rect 43484 3388 43652 3390
rect 43372 3378 43428 3388
rect 43596 3378 43652 3388
rect 43932 3444 43988 3454
rect 44044 3444 44100 4174
rect 44268 3444 44324 3454
rect 44044 3442 44324 3444
rect 44044 3390 44270 3442
rect 44322 3390 44324 3442
rect 44044 3388 44324 3390
rect 44380 3444 44436 8372
rect 44940 8258 44996 8372
rect 44940 8206 44942 8258
rect 44994 8206 44996 8258
rect 44940 8194 44996 8206
rect 44716 7476 44772 7486
rect 45052 7476 45108 8876
rect 45164 8866 45220 8876
rect 45612 8988 45780 9044
rect 45612 7700 45668 8988
rect 46060 8930 46116 8942
rect 46060 8878 46062 8930
rect 46114 8878 46116 8930
rect 45948 8818 46004 8830
rect 45948 8766 45950 8818
rect 46002 8766 46004 8818
rect 45948 8428 46004 8766
rect 45724 8372 46004 8428
rect 45724 8370 45780 8372
rect 45724 8318 45726 8370
rect 45778 8318 45780 8370
rect 45724 8306 45780 8318
rect 45724 7700 45780 7710
rect 45668 7698 45780 7700
rect 45668 7646 45726 7698
rect 45778 7646 45780 7698
rect 45668 7644 45780 7646
rect 45612 7606 45668 7644
rect 45724 7634 45780 7644
rect 44716 7474 45108 7476
rect 44716 7422 44718 7474
rect 44770 7422 45108 7474
rect 44716 7420 45108 7422
rect 45276 7588 45332 7598
rect 44492 5908 44548 5918
rect 44716 5908 44772 7420
rect 45164 7364 45220 7374
rect 45164 7270 45220 7308
rect 45164 7028 45220 7038
rect 44492 5906 44772 5908
rect 44492 5854 44494 5906
rect 44546 5854 44772 5906
rect 44492 5852 44772 5854
rect 45052 6972 45164 7028
rect 44492 5842 44548 5852
rect 45052 5682 45108 6972
rect 45164 6962 45220 6972
rect 45276 5906 45332 7532
rect 45612 7364 45668 7374
rect 45612 6018 45668 7308
rect 46060 7028 46116 8878
rect 46172 8372 46228 11004
rect 46508 10612 46564 10622
rect 46508 10518 46564 10556
rect 46620 9266 46676 11452
rect 47292 9940 47348 12126
rect 47628 12738 47684 12750
rect 47628 12686 47630 12738
rect 47682 12686 47684 12738
rect 47404 12068 47460 12078
rect 47628 12068 47684 12686
rect 47852 12404 47908 12414
rect 47852 12290 47908 12348
rect 47964 12402 48020 14252
rect 47964 12350 47966 12402
rect 48018 12350 48020 12402
rect 47964 12338 48020 12350
rect 48188 12962 48244 12974
rect 48188 12910 48190 12962
rect 48242 12910 48244 12962
rect 48188 12402 48244 12910
rect 48300 12740 48356 15820
rect 48636 15148 48692 31164
rect 48860 30322 48916 31612
rect 48860 30270 48862 30322
rect 48914 30270 48916 30322
rect 48860 30258 48916 30270
rect 49084 30994 49140 31006
rect 49084 30942 49086 30994
rect 49138 30942 49140 30994
rect 48748 30212 48804 30222
rect 48748 30118 48804 30156
rect 48972 29988 49028 29998
rect 48972 29894 49028 29932
rect 48860 29428 48916 29438
rect 48860 29316 48916 29372
rect 49084 29316 49140 30942
rect 49868 30324 49924 30334
rect 49868 30230 49924 30268
rect 49420 30212 49476 30222
rect 49420 30118 49476 30156
rect 49644 30210 49700 30222
rect 49644 30158 49646 30210
rect 49698 30158 49700 30210
rect 48860 29314 49140 29316
rect 48860 29262 48862 29314
rect 48914 29262 49140 29314
rect 48860 29260 49140 29262
rect 49644 29876 49700 30158
rect 48748 27860 48804 27870
rect 48748 27766 48804 27804
rect 48748 26292 48804 26302
rect 48748 26178 48804 26236
rect 48748 26126 48750 26178
rect 48802 26126 48804 26178
rect 48748 24834 48804 26126
rect 48748 24782 48750 24834
rect 48802 24782 48804 24834
rect 48748 24770 48804 24782
rect 48860 23940 48916 29260
rect 49532 27970 49588 27982
rect 49532 27918 49534 27970
rect 49586 27918 49588 27970
rect 49308 27858 49364 27870
rect 49308 27806 49310 27858
rect 49362 27806 49364 27858
rect 48972 26964 49028 26974
rect 49308 26908 49364 27806
rect 48972 26852 49364 26908
rect 48972 26290 49028 26852
rect 48972 26238 48974 26290
rect 49026 26238 49028 26290
rect 48972 26226 49028 26238
rect 49532 26292 49588 27918
rect 49644 27746 49700 29820
rect 49980 29428 50036 33070
rect 50428 33122 50596 33124
rect 50428 33070 50542 33122
rect 50594 33070 50596 33122
rect 50428 33068 50596 33070
rect 50428 30436 50484 33068
rect 50540 33058 50596 33068
rect 50556 32956 50820 32966
rect 50612 32900 50660 32956
rect 50716 32900 50764 32956
rect 50556 32890 50820 32900
rect 50540 31892 50596 31902
rect 50540 31556 50596 31836
rect 52668 31778 52724 37100
rect 55356 37044 55412 37054
rect 55356 36950 55412 36988
rect 55580 36932 55636 36942
rect 55020 36594 55076 36606
rect 55020 36542 55022 36594
rect 55074 36542 55076 36594
rect 52780 36484 52836 36494
rect 52780 36390 52836 36428
rect 53452 35698 53508 35710
rect 53452 35646 53454 35698
rect 53506 35646 53508 35698
rect 53228 35588 53284 35598
rect 53452 35588 53508 35646
rect 55020 35700 55076 36542
rect 55580 36482 55636 36876
rect 57932 36706 57988 37660
rect 57932 36654 57934 36706
rect 57986 36654 57988 36706
rect 57932 36642 57988 36654
rect 55580 36430 55582 36482
rect 55634 36430 55636 36482
rect 55580 36418 55636 36430
rect 55020 35634 55076 35644
rect 55244 36372 55300 36382
rect 53228 35586 53508 35588
rect 53228 35534 53230 35586
rect 53282 35534 53508 35586
rect 53228 35532 53508 35534
rect 53228 35476 53284 35532
rect 53228 35410 53284 35420
rect 55244 35140 55300 36316
rect 55468 35588 55524 35598
rect 55244 35074 55300 35084
rect 55356 35474 55412 35486
rect 55356 35422 55358 35474
rect 55410 35422 55412 35474
rect 55356 35028 55412 35422
rect 55356 34962 55412 34972
rect 55244 34692 55300 34702
rect 53452 34130 53508 34142
rect 53452 34078 53454 34130
rect 53506 34078 53508 34130
rect 53452 34020 53508 34078
rect 53452 33954 53508 33964
rect 53452 33684 53508 33694
rect 52668 31726 52670 31778
rect 52722 31726 52724 31778
rect 52668 31714 52724 31726
rect 53228 32788 53284 32798
rect 50540 31500 50932 31556
rect 50556 31388 50820 31398
rect 50612 31332 50660 31388
rect 50716 31332 50764 31388
rect 50556 31322 50820 31332
rect 50764 31108 50820 31118
rect 50764 31014 50820 31052
rect 50428 30380 50596 30436
rect 50428 30212 50484 30222
rect 50428 30118 50484 30156
rect 50204 29988 50260 29998
rect 50540 29988 50596 30380
rect 50764 30100 50820 30110
rect 50876 30100 50932 31500
rect 50820 30044 50932 30100
rect 51324 31108 51380 31118
rect 50204 29894 50260 29932
rect 50428 29932 50596 29988
rect 50652 29988 50708 30026
rect 50764 30006 50820 30044
rect 50316 29876 50372 29886
rect 49980 29372 50260 29428
rect 49644 27694 49646 27746
rect 49698 27694 49700 27746
rect 49644 27682 49700 27694
rect 50092 27858 50148 27870
rect 50092 27806 50094 27858
rect 50146 27806 50148 27858
rect 49756 26964 49812 26974
rect 49644 26516 49700 26526
rect 49644 26422 49700 26460
rect 49756 26514 49812 26908
rect 49756 26462 49758 26514
rect 49810 26462 49812 26514
rect 49756 26450 49812 26462
rect 50092 26514 50148 27806
rect 50092 26462 50094 26514
rect 50146 26462 50148 26514
rect 50092 26450 50148 26462
rect 49868 26292 49924 26302
rect 49532 26226 49588 26236
rect 49756 26290 49924 26292
rect 49756 26238 49870 26290
rect 49922 26238 49924 26290
rect 49756 26236 49924 26238
rect 49308 26068 49364 26078
rect 49756 26068 49812 26236
rect 49868 26226 49924 26236
rect 49308 26066 49812 26068
rect 49308 26014 49310 26066
rect 49362 26014 49812 26066
rect 49308 26012 49812 26014
rect 49308 26002 49364 26012
rect 50204 24948 50260 29372
rect 50316 27970 50372 29820
rect 50316 27918 50318 27970
rect 50370 27918 50372 27970
rect 50316 25956 50372 27918
rect 50428 27970 50484 29932
rect 50652 29922 50708 29932
rect 50556 29820 50820 29830
rect 50612 29764 50660 29820
rect 50716 29764 50764 29820
rect 50556 29754 50820 29764
rect 50556 28252 50820 28262
rect 50612 28196 50660 28252
rect 50716 28196 50764 28252
rect 50556 28186 50820 28196
rect 50428 27918 50430 27970
rect 50482 27918 50484 27970
rect 50428 27188 50484 27918
rect 50428 27122 50484 27132
rect 51324 27074 51380 31052
rect 53228 30212 53284 32732
rect 53452 32562 53508 33628
rect 53452 32510 53454 32562
rect 53506 32510 53508 32562
rect 53452 32498 53508 32510
rect 55020 31890 55076 31902
rect 55020 31838 55022 31890
rect 55074 31838 55076 31890
rect 55020 30996 55076 31838
rect 55020 30930 55076 30940
rect 53452 30212 53508 30222
rect 53228 30210 53508 30212
rect 53228 30158 53230 30210
rect 53282 30158 53454 30210
rect 53506 30158 53508 30210
rect 53228 30156 53508 30158
rect 53228 30146 53284 30156
rect 53452 30146 53508 30156
rect 55244 28756 55300 34636
rect 55356 33908 55412 33918
rect 55356 33814 55412 33852
rect 55356 33236 55412 33246
rect 55356 33142 55412 33180
rect 55356 32340 55412 32350
rect 55356 32246 55412 32284
rect 55468 31948 55524 35532
rect 56588 35140 56644 35150
rect 56588 35046 56644 35084
rect 55580 34916 55636 34926
rect 55580 34822 55636 34860
rect 57932 34356 57988 34366
rect 57932 33570 57988 34300
rect 57932 33518 57934 33570
rect 57986 33518 57988 33570
rect 57932 33506 57988 33518
rect 55580 33348 55636 33358
rect 55580 33254 55636 33292
rect 57932 33012 57988 33022
rect 55468 31892 55636 31948
rect 55580 31778 55636 31892
rect 57932 31890 57988 32956
rect 57932 31838 57934 31890
rect 57986 31838 57988 31890
rect 57932 31826 57988 31838
rect 55580 31726 55582 31778
rect 55634 31726 55636 31778
rect 55580 31714 55636 31726
rect 57932 31668 57988 31678
rect 55356 30324 55412 30334
rect 55356 30230 55412 30268
rect 57932 28866 57988 31612
rect 57932 28814 57934 28866
rect 57986 28814 57988 28866
rect 57932 28802 57988 28814
rect 55356 28756 55412 28766
rect 55244 28754 55636 28756
rect 55244 28702 55358 28754
rect 55410 28702 55636 28754
rect 55244 28700 55636 28702
rect 55356 28662 55412 28700
rect 55580 28642 55636 28700
rect 55580 28590 55582 28642
rect 55634 28590 55636 28642
rect 55580 28578 55636 28590
rect 51324 27022 51326 27074
rect 51378 27022 51380 27074
rect 51324 27010 51380 27022
rect 50652 26964 50708 26974
rect 50652 26870 50708 26908
rect 50556 26684 50820 26694
rect 50612 26628 50660 26684
rect 50716 26628 50764 26684
rect 50556 26618 50820 26628
rect 50316 25890 50372 25900
rect 57036 26068 57092 26078
rect 50556 25116 50820 25126
rect 50612 25060 50660 25116
rect 50716 25060 50764 25116
rect 50556 25050 50820 25060
rect 49868 24892 50260 24948
rect 57036 24948 57092 26012
rect 57596 25396 57652 25406
rect 57596 25302 57652 25340
rect 58156 25396 58212 25406
rect 57820 25284 57876 25294
rect 57820 25190 57876 25228
rect 49868 24836 49924 24892
rect 57036 24882 57092 24892
rect 57820 24948 57876 24958
rect 57820 24854 57876 24892
rect 58156 24948 58212 25340
rect 58156 24882 58212 24892
rect 49420 24724 49476 24734
rect 49420 24630 49476 24668
rect 48860 23874 48916 23884
rect 48972 24610 49028 24622
rect 48972 24558 48974 24610
rect 49026 24558 49028 24610
rect 48748 23044 48804 23054
rect 48748 22950 48804 22988
rect 48972 22372 49028 24558
rect 49420 23828 49476 23838
rect 49420 23154 49476 23772
rect 49868 23828 49924 24780
rect 50652 24834 50708 24846
rect 50652 24782 50654 24834
rect 50706 24782 50708 24834
rect 49420 23102 49422 23154
rect 49474 23102 49476 23154
rect 49420 23090 49476 23102
rect 49644 23604 49700 23614
rect 49644 23154 49700 23548
rect 49868 23492 49924 23772
rect 49868 23426 49924 23436
rect 49980 24722 50036 24734
rect 49980 24670 49982 24722
rect 50034 24670 50036 24722
rect 49980 23378 50036 24670
rect 50540 24724 50596 24734
rect 50540 24630 50596 24668
rect 50428 24500 50484 24510
rect 50316 24498 50484 24500
rect 50316 24446 50430 24498
rect 50482 24446 50484 24498
rect 50316 24444 50484 24446
rect 50092 23940 50148 23950
rect 50092 23846 50148 23884
rect 50204 23716 50260 23726
rect 49980 23326 49982 23378
rect 50034 23326 50036 23378
rect 49980 23314 50036 23326
rect 50092 23660 50204 23716
rect 49644 23102 49646 23154
rect 49698 23102 49700 23154
rect 49644 23090 49700 23102
rect 49980 22484 50036 22494
rect 50092 22484 50148 23660
rect 50204 23650 50260 23660
rect 50316 23604 50372 24444
rect 50428 24434 50484 24444
rect 50652 23938 50708 24782
rect 58156 24722 58212 24734
rect 58156 24670 58158 24722
rect 58210 24670 58212 24722
rect 57596 24612 57652 24622
rect 58156 24612 58212 24670
rect 57596 24610 58212 24612
rect 57596 24558 57598 24610
rect 57650 24558 58212 24610
rect 57596 24556 58212 24558
rect 57596 24546 57652 24556
rect 58156 24276 58212 24556
rect 58156 24210 58212 24220
rect 50652 23886 50654 23938
rect 50706 23886 50708 23938
rect 50428 23828 50484 23838
rect 50428 23734 50484 23772
rect 50652 23716 50708 23886
rect 50652 23650 50708 23660
rect 50988 23940 51044 23950
rect 50204 23492 50260 23502
rect 50204 23378 50260 23436
rect 50204 23326 50206 23378
rect 50258 23326 50260 23378
rect 50204 23314 50260 23326
rect 49980 22482 50148 22484
rect 49980 22430 49982 22482
rect 50034 22430 50148 22482
rect 49980 22428 50148 22430
rect 50316 23266 50372 23548
rect 50556 23548 50820 23558
rect 50612 23492 50660 23548
rect 50716 23492 50764 23548
rect 50556 23482 50820 23492
rect 50316 23214 50318 23266
rect 50370 23214 50372 23266
rect 49980 22418 50036 22428
rect 48972 22306 49028 22316
rect 50316 22148 50372 23214
rect 50092 22092 50372 22148
rect 49644 21252 49700 21262
rect 48860 19906 48916 19918
rect 48860 19854 48862 19906
rect 48914 19854 48916 19906
rect 48860 19684 48916 19854
rect 48860 19618 48916 19628
rect 48748 18340 48804 18350
rect 48748 18246 48804 18284
rect 48972 17892 49028 17902
rect 48972 17798 49028 17836
rect 48748 17668 48804 17678
rect 48748 16884 48804 17612
rect 48860 17444 48916 17454
rect 49308 17444 49364 17454
rect 48860 17106 48916 17388
rect 48860 17054 48862 17106
rect 48914 17054 48916 17106
rect 48860 17042 48916 17054
rect 49084 17442 49364 17444
rect 49084 17390 49310 17442
rect 49362 17390 49364 17442
rect 49084 17388 49364 17390
rect 49084 17106 49140 17388
rect 49308 17378 49364 17388
rect 49084 17054 49086 17106
rect 49138 17054 49140 17106
rect 49084 17042 49140 17054
rect 49308 17108 49364 17118
rect 49308 17014 49364 17052
rect 49644 17108 49700 21196
rect 50092 20804 50148 22092
rect 50556 21980 50820 21990
rect 50612 21924 50660 21980
rect 50716 21924 50764 21980
rect 50556 21914 50820 21924
rect 50092 19346 50148 20748
rect 50556 20412 50820 20422
rect 50612 20356 50660 20412
rect 50716 20356 50764 20412
rect 50556 20346 50820 20356
rect 50092 19294 50094 19346
rect 50146 19294 50148 19346
rect 50092 19282 50148 19294
rect 50556 18844 50820 18854
rect 50612 18788 50660 18844
rect 50716 18788 50764 18844
rect 50556 18778 50820 18788
rect 49756 18340 49812 18350
rect 49756 17780 49812 18284
rect 50876 18338 50932 18350
rect 50876 18286 50878 18338
rect 50930 18286 50932 18338
rect 50204 17780 50260 17790
rect 49756 17778 50260 17780
rect 49756 17726 49758 17778
rect 49810 17726 50206 17778
rect 50258 17726 50260 17778
rect 49756 17724 50260 17726
rect 49756 17714 49812 17724
rect 50204 17714 50260 17724
rect 50556 17276 50820 17286
rect 50612 17220 50660 17276
rect 50716 17220 50764 17276
rect 50556 17210 50820 17220
rect 49756 17108 49812 17118
rect 49644 17106 49812 17108
rect 49644 17054 49758 17106
rect 49810 17054 49812 17106
rect 49644 17052 49812 17054
rect 49196 16996 49252 17006
rect 49196 16902 49252 16940
rect 48748 16828 48916 16884
rect 48748 15876 48804 15886
rect 48748 15782 48804 15820
rect 48524 15092 48692 15148
rect 48748 15540 48804 15550
rect 48412 13636 48468 13646
rect 48412 12962 48468 13580
rect 48524 13300 48580 15092
rect 48524 13234 48580 13244
rect 48636 14418 48692 14430
rect 48636 14366 48638 14418
rect 48690 14366 48692 14418
rect 48524 13076 48580 13086
rect 48636 13076 48692 14366
rect 48748 13970 48804 15484
rect 48860 15538 48916 16828
rect 49084 16324 49140 16334
rect 49084 16322 49364 16324
rect 49084 16270 49086 16322
rect 49138 16270 49364 16322
rect 49084 16268 49364 16270
rect 49084 16258 49140 16268
rect 48972 15876 49028 15886
rect 48972 15782 49028 15820
rect 49196 15874 49252 15886
rect 49196 15822 49198 15874
rect 49250 15822 49252 15874
rect 48860 15486 48862 15538
rect 48914 15486 48916 15538
rect 48860 15474 48916 15486
rect 48748 13918 48750 13970
rect 48802 13918 48804 13970
rect 48748 13906 48804 13918
rect 48972 15314 49028 15326
rect 48972 15262 48974 15314
rect 49026 15262 49028 15314
rect 48972 15204 49028 15262
rect 48972 13748 49028 15148
rect 49196 15148 49252 15822
rect 49308 15314 49364 16268
rect 49532 16100 49588 16110
rect 49644 16100 49700 17052
rect 49756 17042 49812 17052
rect 50876 16996 50932 18286
rect 50876 16930 50932 16940
rect 49980 16212 50036 16222
rect 49980 16118 50036 16156
rect 49532 16098 49700 16100
rect 49532 16046 49534 16098
rect 49586 16046 49700 16098
rect 49532 16044 49700 16046
rect 49756 16100 49812 16110
rect 50428 16100 50484 16110
rect 49420 15988 49476 15998
rect 49420 15894 49476 15932
rect 49532 15876 49588 16044
rect 49532 15810 49588 15820
rect 49756 15538 49812 16044
rect 49756 15486 49758 15538
rect 49810 15486 49812 15538
rect 49756 15474 49812 15486
rect 50316 16044 50428 16100
rect 49308 15262 49310 15314
rect 49362 15262 49364 15314
rect 49308 15250 49364 15262
rect 50316 15316 50372 16044
rect 50428 16006 50484 16044
rect 50556 15708 50820 15718
rect 50612 15652 50660 15708
rect 50716 15652 50764 15708
rect 50556 15642 50820 15652
rect 50428 15540 50484 15550
rect 50988 15540 51044 23884
rect 58156 23826 58212 23838
rect 58156 23774 58158 23826
rect 58210 23774 58212 23826
rect 57596 23714 57652 23726
rect 57596 23662 57598 23714
rect 57650 23662 57652 23714
rect 57596 23604 57652 23662
rect 57820 23716 57876 23726
rect 57820 23622 57876 23660
rect 57596 23538 57652 23548
rect 58156 23604 58212 23774
rect 58156 23538 58212 23548
rect 57596 22260 57652 22270
rect 57596 22166 57652 22204
rect 58156 22260 58212 22270
rect 57820 22148 57876 22158
rect 57820 22054 57876 22092
rect 53788 21924 53844 21934
rect 53788 20132 53844 21868
rect 58156 21588 58212 22204
rect 58156 21522 58212 21532
rect 53788 20066 53844 20076
rect 50428 15538 51044 15540
rect 50428 15486 50430 15538
rect 50482 15486 51044 15538
rect 50428 15484 51044 15486
rect 50428 15474 50484 15484
rect 50316 15260 50820 15316
rect 50316 15148 50372 15260
rect 49196 15092 49364 15148
rect 49308 14308 49364 15092
rect 48972 13654 49028 13692
rect 49084 14252 49364 14308
rect 49420 15092 49476 15102
rect 48860 13636 48916 13646
rect 48860 13542 48916 13580
rect 48524 13074 48692 13076
rect 48524 13022 48526 13074
rect 48578 13022 48692 13074
rect 48524 13020 48692 13022
rect 48860 13300 48916 13310
rect 48524 13010 48580 13020
rect 48412 12910 48414 12962
rect 48466 12910 48468 12962
rect 48412 12898 48468 12910
rect 48636 12740 48692 12750
rect 48300 12738 48692 12740
rect 48300 12686 48638 12738
rect 48690 12686 48692 12738
rect 48300 12684 48692 12686
rect 48636 12674 48692 12684
rect 48188 12350 48190 12402
rect 48242 12350 48244 12402
rect 48188 12338 48244 12350
rect 48860 12404 48916 13244
rect 49084 12962 49140 14252
rect 49196 13972 49252 13982
rect 49196 13878 49252 13916
rect 49420 13524 49476 15036
rect 49868 15092 50372 15148
rect 49868 14532 49924 15092
rect 50764 14642 50820 15260
rect 50988 15314 51044 15484
rect 50988 15262 50990 15314
rect 51042 15262 51044 15314
rect 50988 15250 51044 15262
rect 51660 18450 51716 18462
rect 51660 18398 51662 18450
rect 51714 18398 51716 18450
rect 51660 15092 51716 18398
rect 51660 15026 51716 15036
rect 52780 15202 52836 15214
rect 52780 15150 52782 15202
rect 52834 15150 52836 15202
rect 52780 15092 52836 15150
rect 52780 15026 52836 15036
rect 50764 14590 50766 14642
rect 50818 14590 50820 14642
rect 50764 14578 50820 14590
rect 49868 13970 49924 14476
rect 50556 14140 50820 14150
rect 50612 14084 50660 14140
rect 50716 14084 50764 14140
rect 50556 14074 50820 14084
rect 49868 13918 49870 13970
rect 49922 13918 49924 13970
rect 49868 13906 49924 13918
rect 49084 12910 49086 12962
rect 49138 12910 49140 12962
rect 49084 12898 49140 12910
rect 49308 13468 49476 13524
rect 48860 12310 48916 12348
rect 47852 12238 47854 12290
rect 47906 12238 47908 12290
rect 47852 12226 47908 12238
rect 47628 12012 48692 12068
rect 47404 11974 47460 12012
rect 48636 11506 48692 12012
rect 48636 11454 48638 11506
rect 48690 11454 48692 11506
rect 48636 11442 48692 11454
rect 49308 11394 49364 13468
rect 49420 13300 49476 13310
rect 49420 13074 49476 13244
rect 49420 13022 49422 13074
rect 49474 13022 49476 13074
rect 49420 13010 49476 13022
rect 50556 12572 50820 12582
rect 50612 12516 50660 12572
rect 50716 12516 50764 12572
rect 50556 12506 50820 12516
rect 49308 11342 49310 11394
rect 49362 11342 49364 11394
rect 49308 11330 49364 11342
rect 50556 11004 50820 11014
rect 50612 10948 50660 11004
rect 50716 10948 50764 11004
rect 50556 10938 50820 10948
rect 47740 9940 47796 9950
rect 47292 9938 47796 9940
rect 47292 9886 47742 9938
rect 47794 9886 47796 9938
rect 47292 9884 47796 9886
rect 47740 9874 47796 9884
rect 50556 9436 50820 9446
rect 50612 9380 50660 9436
rect 50716 9380 50764 9436
rect 50556 9370 50820 9380
rect 46620 9214 46622 9266
rect 46674 9214 46676 9266
rect 46620 9202 46676 9214
rect 46172 7588 46228 8316
rect 47852 8372 47908 8382
rect 47852 8278 47908 8316
rect 50556 7868 50820 7878
rect 50612 7812 50660 7868
rect 50716 7812 50764 7868
rect 50556 7802 50820 7812
rect 46172 7522 46228 7532
rect 46060 6962 46116 6972
rect 50556 6300 50820 6310
rect 50612 6244 50660 6300
rect 50716 6244 50764 6300
rect 50556 6234 50820 6244
rect 45612 5966 45614 6018
rect 45666 5966 45668 6018
rect 45612 5954 45668 5966
rect 45276 5854 45278 5906
rect 45330 5854 45332 5906
rect 45276 5842 45332 5854
rect 45052 5630 45054 5682
rect 45106 5630 45108 5682
rect 45052 5618 45108 5630
rect 50556 4732 50820 4742
rect 50612 4676 50660 4732
rect 50716 4676 50764 4732
rect 50556 4666 50820 4676
rect 44604 3444 44660 3454
rect 44380 3442 44660 3444
rect 44380 3390 44606 3442
rect 44658 3390 44660 3442
rect 44380 3388 44660 3390
rect 43932 3350 43988 3388
rect 44268 2548 44324 3388
rect 44604 3378 44660 3388
rect 50556 3164 50820 3174
rect 50612 3108 50660 3164
rect 50716 3108 50764 3164
rect 50556 3098 50820 3108
rect 43708 2492 44324 2548
rect 43708 800 43764 2492
rect 0 0 112 800
rect 672 0 784 800
rect 1344 0 1456 800
rect 2016 0 2128 800
rect 2688 0 2800 800
rect 3360 0 3472 800
rect 4032 0 4144 800
rect 4704 0 4816 800
rect 5376 0 5488 800
rect 6048 0 6160 800
rect 6720 0 6832 800
rect 7392 0 7504 800
rect 8064 0 8176 800
rect 8736 0 8848 800
rect 9408 0 9520 800
rect 12768 0 12880 800
rect 16128 0 16240 800
rect 16800 0 16912 800
rect 18144 0 18256 800
rect 18816 0 18928 800
rect 19488 0 19600 800
rect 20160 0 20272 800
rect 20832 0 20944 800
rect 22848 0 22960 800
rect 23520 0 23632 800
rect 24192 0 24304 800
rect 25536 0 25648 800
rect 26208 0 26320 800
rect 26880 0 26992 800
rect 27552 0 27664 800
rect 28896 0 29008 800
rect 29568 0 29680 800
rect 30240 0 30352 800
rect 30912 0 31024 800
rect 32928 0 33040 800
rect 33600 0 33712 800
rect 34272 0 34384 800
rect 35616 0 35728 800
rect 36288 0 36400 800
rect 36960 0 37072 800
rect 37632 0 37744 800
rect 38304 0 38416 800
rect 39648 0 39760 800
rect 40320 0 40432 800
rect 40992 0 41104 800
rect 42336 0 42448 800
rect 43008 0 43120 800
rect 43680 0 43792 800
<< via2 >>
rect 19836 76858 19892 76860
rect 19836 76806 19838 76858
rect 19838 76806 19890 76858
rect 19890 76806 19892 76858
rect 19836 76804 19892 76806
rect 19940 76858 19996 76860
rect 19940 76806 19942 76858
rect 19942 76806 19994 76858
rect 19994 76806 19996 76858
rect 19940 76804 19996 76806
rect 20044 76858 20100 76860
rect 20044 76806 20046 76858
rect 20046 76806 20098 76858
rect 20098 76806 20100 76858
rect 20044 76804 20100 76806
rect 50556 76858 50612 76860
rect 50556 76806 50558 76858
rect 50558 76806 50610 76858
rect 50610 76806 50612 76858
rect 50556 76804 50612 76806
rect 50660 76858 50716 76860
rect 50660 76806 50662 76858
rect 50662 76806 50714 76858
rect 50714 76806 50716 76858
rect 50660 76804 50716 76806
rect 50764 76858 50820 76860
rect 50764 76806 50766 76858
rect 50766 76806 50818 76858
rect 50818 76806 50820 76858
rect 50764 76804 50820 76806
rect 4476 76074 4532 76076
rect 4476 76022 4478 76074
rect 4478 76022 4530 76074
rect 4530 76022 4532 76074
rect 4476 76020 4532 76022
rect 4580 76074 4636 76076
rect 4580 76022 4582 76074
rect 4582 76022 4634 76074
rect 4634 76022 4636 76074
rect 4580 76020 4636 76022
rect 4684 76074 4740 76076
rect 4684 76022 4686 76074
rect 4686 76022 4738 76074
rect 4738 76022 4740 76074
rect 4684 76020 4740 76022
rect 35196 76074 35252 76076
rect 35196 76022 35198 76074
rect 35198 76022 35250 76074
rect 35250 76022 35252 76074
rect 35196 76020 35252 76022
rect 35300 76074 35356 76076
rect 35300 76022 35302 76074
rect 35302 76022 35354 76074
rect 35354 76022 35356 76074
rect 35300 76020 35356 76022
rect 35404 76074 35460 76076
rect 35404 76022 35406 76074
rect 35406 76022 35458 76074
rect 35458 76022 35460 76074
rect 35404 76020 35460 76022
rect 19836 75290 19892 75292
rect 19836 75238 19838 75290
rect 19838 75238 19890 75290
rect 19890 75238 19892 75290
rect 19836 75236 19892 75238
rect 19940 75290 19996 75292
rect 19940 75238 19942 75290
rect 19942 75238 19994 75290
rect 19994 75238 19996 75290
rect 19940 75236 19996 75238
rect 20044 75290 20100 75292
rect 20044 75238 20046 75290
rect 20046 75238 20098 75290
rect 20098 75238 20100 75290
rect 20044 75236 20100 75238
rect 50556 75290 50612 75292
rect 50556 75238 50558 75290
rect 50558 75238 50610 75290
rect 50610 75238 50612 75290
rect 50556 75236 50612 75238
rect 50660 75290 50716 75292
rect 50660 75238 50662 75290
rect 50662 75238 50714 75290
rect 50714 75238 50716 75290
rect 50660 75236 50716 75238
rect 50764 75290 50820 75292
rect 50764 75238 50766 75290
rect 50766 75238 50818 75290
rect 50818 75238 50820 75290
rect 50764 75236 50820 75238
rect 4476 74506 4532 74508
rect 4476 74454 4478 74506
rect 4478 74454 4530 74506
rect 4530 74454 4532 74506
rect 4476 74452 4532 74454
rect 4580 74506 4636 74508
rect 4580 74454 4582 74506
rect 4582 74454 4634 74506
rect 4634 74454 4636 74506
rect 4580 74452 4636 74454
rect 4684 74506 4740 74508
rect 4684 74454 4686 74506
rect 4686 74454 4738 74506
rect 4738 74454 4740 74506
rect 4684 74452 4740 74454
rect 35196 74506 35252 74508
rect 35196 74454 35198 74506
rect 35198 74454 35250 74506
rect 35250 74454 35252 74506
rect 35196 74452 35252 74454
rect 35300 74506 35356 74508
rect 35300 74454 35302 74506
rect 35302 74454 35354 74506
rect 35354 74454 35356 74506
rect 35300 74452 35356 74454
rect 35404 74506 35460 74508
rect 35404 74454 35406 74506
rect 35406 74454 35458 74506
rect 35458 74454 35460 74506
rect 35404 74452 35460 74454
rect 19836 73722 19892 73724
rect 19836 73670 19838 73722
rect 19838 73670 19890 73722
rect 19890 73670 19892 73722
rect 19836 73668 19892 73670
rect 19940 73722 19996 73724
rect 19940 73670 19942 73722
rect 19942 73670 19994 73722
rect 19994 73670 19996 73722
rect 19940 73668 19996 73670
rect 20044 73722 20100 73724
rect 20044 73670 20046 73722
rect 20046 73670 20098 73722
rect 20098 73670 20100 73722
rect 20044 73668 20100 73670
rect 50556 73722 50612 73724
rect 50556 73670 50558 73722
rect 50558 73670 50610 73722
rect 50610 73670 50612 73722
rect 50556 73668 50612 73670
rect 50660 73722 50716 73724
rect 50660 73670 50662 73722
rect 50662 73670 50714 73722
rect 50714 73670 50716 73722
rect 50660 73668 50716 73670
rect 50764 73722 50820 73724
rect 50764 73670 50766 73722
rect 50766 73670 50818 73722
rect 50818 73670 50820 73722
rect 50764 73668 50820 73670
rect 4476 72938 4532 72940
rect 4476 72886 4478 72938
rect 4478 72886 4530 72938
rect 4530 72886 4532 72938
rect 4476 72884 4532 72886
rect 4580 72938 4636 72940
rect 4580 72886 4582 72938
rect 4582 72886 4634 72938
rect 4634 72886 4636 72938
rect 4580 72884 4636 72886
rect 4684 72938 4740 72940
rect 4684 72886 4686 72938
rect 4686 72886 4738 72938
rect 4738 72886 4740 72938
rect 4684 72884 4740 72886
rect 35196 72938 35252 72940
rect 35196 72886 35198 72938
rect 35198 72886 35250 72938
rect 35250 72886 35252 72938
rect 35196 72884 35252 72886
rect 35300 72938 35356 72940
rect 35300 72886 35302 72938
rect 35302 72886 35354 72938
rect 35354 72886 35356 72938
rect 35300 72884 35356 72886
rect 35404 72938 35460 72940
rect 35404 72886 35406 72938
rect 35406 72886 35458 72938
rect 35458 72886 35460 72938
rect 35404 72884 35460 72886
rect 19836 72154 19892 72156
rect 19836 72102 19838 72154
rect 19838 72102 19890 72154
rect 19890 72102 19892 72154
rect 19836 72100 19892 72102
rect 19940 72154 19996 72156
rect 19940 72102 19942 72154
rect 19942 72102 19994 72154
rect 19994 72102 19996 72154
rect 19940 72100 19996 72102
rect 20044 72154 20100 72156
rect 20044 72102 20046 72154
rect 20046 72102 20098 72154
rect 20098 72102 20100 72154
rect 20044 72100 20100 72102
rect 50556 72154 50612 72156
rect 50556 72102 50558 72154
rect 50558 72102 50610 72154
rect 50610 72102 50612 72154
rect 50556 72100 50612 72102
rect 50660 72154 50716 72156
rect 50660 72102 50662 72154
rect 50662 72102 50714 72154
rect 50714 72102 50716 72154
rect 50660 72100 50716 72102
rect 50764 72154 50820 72156
rect 50764 72102 50766 72154
rect 50766 72102 50818 72154
rect 50818 72102 50820 72154
rect 50764 72100 50820 72102
rect 4476 71370 4532 71372
rect 4476 71318 4478 71370
rect 4478 71318 4530 71370
rect 4530 71318 4532 71370
rect 4476 71316 4532 71318
rect 4580 71370 4636 71372
rect 4580 71318 4582 71370
rect 4582 71318 4634 71370
rect 4634 71318 4636 71370
rect 4580 71316 4636 71318
rect 4684 71370 4740 71372
rect 4684 71318 4686 71370
rect 4686 71318 4738 71370
rect 4738 71318 4740 71370
rect 4684 71316 4740 71318
rect 35196 71370 35252 71372
rect 35196 71318 35198 71370
rect 35198 71318 35250 71370
rect 35250 71318 35252 71370
rect 35196 71316 35252 71318
rect 35300 71370 35356 71372
rect 35300 71318 35302 71370
rect 35302 71318 35354 71370
rect 35354 71318 35356 71370
rect 35300 71316 35356 71318
rect 35404 71370 35460 71372
rect 35404 71318 35406 71370
rect 35406 71318 35458 71370
rect 35458 71318 35460 71370
rect 35404 71316 35460 71318
rect 4172 70588 4228 70644
rect 1708 54348 1764 54404
rect 2492 54402 2548 54404
rect 2492 54350 2494 54402
rect 2494 54350 2546 54402
rect 2546 54350 2548 54402
rect 2492 54348 2548 54350
rect 1708 53788 1764 53844
rect 1708 53116 1764 53172
rect 1596 53004 1652 53060
rect 1484 50540 1540 50596
rect 1484 43596 1540 43652
rect 2044 53058 2100 53060
rect 2044 53006 2046 53058
rect 2046 53006 2098 53058
rect 2098 53006 2100 53058
rect 2044 53004 2100 53006
rect 1708 52444 1764 52500
rect 1708 51772 1764 51828
rect 1708 51100 1764 51156
rect 1820 50316 1876 50372
rect 1820 49756 1876 49812
rect 1708 49644 1764 49700
rect 2044 50652 2100 50708
rect 1708 49084 1764 49140
rect 1708 46396 1764 46452
rect 2044 49196 2100 49252
rect 1932 48412 1988 48468
rect 1932 48018 1988 48020
rect 1932 47966 1934 48018
rect 1934 47966 1986 48018
rect 1986 47966 1988 48018
rect 1932 47964 1988 47966
rect 1932 47068 1988 47124
rect 2044 46786 2100 46788
rect 2044 46734 2046 46786
rect 2046 46734 2098 46786
rect 2098 46734 2100 46786
rect 2044 46732 2100 46734
rect 1820 45052 1876 45108
rect 1708 44940 1764 44996
rect 2044 45666 2100 45668
rect 2044 45614 2046 45666
rect 2046 45614 2098 45666
rect 2098 45614 2100 45666
rect 2044 45612 2100 45614
rect 2044 45218 2100 45220
rect 2044 45166 2046 45218
rect 2046 45166 2098 45218
rect 2098 45166 2100 45218
rect 2044 45164 2100 45166
rect 1932 44828 1988 44884
rect 1708 44380 1764 44436
rect 2044 44098 2100 44100
rect 2044 44046 2046 44098
rect 2046 44046 2098 44098
rect 2098 44046 2100 44098
rect 2044 44044 2100 44046
rect 1708 43708 1764 43764
rect 2492 53116 2548 53172
rect 2492 52444 2548 52500
rect 2492 51772 2548 51828
rect 2380 50482 2436 50484
rect 2380 50430 2382 50482
rect 2382 50430 2434 50482
rect 2434 50430 2436 50482
rect 2380 50428 2436 50430
rect 2940 51100 2996 51156
rect 2716 50540 2772 50596
rect 3164 50482 3220 50484
rect 3164 50430 3166 50482
rect 3166 50430 3218 50482
rect 3218 50430 3220 50482
rect 3164 50428 3220 50430
rect 2492 50316 2548 50372
rect 2492 49698 2548 49700
rect 2492 49646 2494 49698
rect 2494 49646 2546 49698
rect 2546 49646 2548 49698
rect 2492 49644 2548 49646
rect 2380 45778 2436 45780
rect 2380 45726 2382 45778
rect 2382 45726 2434 45778
rect 2434 45726 2436 45778
rect 2380 45724 2436 45726
rect 2268 45052 2324 45108
rect 2492 44994 2548 44996
rect 2492 44942 2494 44994
rect 2494 44942 2546 44994
rect 2546 44942 2548 44994
rect 2492 44940 2548 44942
rect 2716 44380 2772 44436
rect 2492 43708 2548 43764
rect 2156 43372 2212 43428
rect 1932 43314 1988 43316
rect 1932 43262 1934 43314
rect 1934 43262 1986 43314
rect 1986 43262 1988 43314
rect 1932 43260 1988 43262
rect 2940 46396 2996 46452
rect 3164 45778 3220 45780
rect 3164 45726 3166 45778
rect 3166 45726 3218 45778
rect 3218 45726 3220 45778
rect 3164 45724 3220 45726
rect 3388 44492 3444 44548
rect 2828 42812 2884 42868
rect 1708 42364 1764 42420
rect 2492 42364 2548 42420
rect 2044 42252 2100 42308
rect 2044 41916 2100 41972
rect 1708 41692 1764 41748
rect 2492 41692 2548 41748
rect 1596 41356 1652 41412
rect 1708 41074 1764 41076
rect 1708 41022 1710 41074
rect 1710 41022 1762 41074
rect 1762 41022 1764 41074
rect 1708 41020 1764 41022
rect 2044 40962 2100 40964
rect 2044 40910 2046 40962
rect 2046 40910 2098 40962
rect 2098 40910 2100 40962
rect 2044 40908 2100 40910
rect 2492 41020 2548 41076
rect 2716 41074 2772 41076
rect 2716 41022 2718 41074
rect 2718 41022 2770 41074
rect 2770 41022 2772 41074
rect 2716 41020 2772 41022
rect 2380 40348 2436 40404
rect 2044 40236 2100 40292
rect 1708 39676 1764 39732
rect 19836 70586 19892 70588
rect 19836 70534 19838 70586
rect 19838 70534 19890 70586
rect 19890 70534 19892 70586
rect 19836 70532 19892 70534
rect 19940 70586 19996 70588
rect 19940 70534 19942 70586
rect 19942 70534 19994 70586
rect 19994 70534 19996 70586
rect 19940 70532 19996 70534
rect 20044 70586 20100 70588
rect 20044 70534 20046 70586
rect 20046 70534 20098 70586
rect 20098 70534 20100 70586
rect 20044 70532 20100 70534
rect 31612 70476 31668 70532
rect 33180 70476 33236 70532
rect 22876 69916 22932 69972
rect 4476 69802 4532 69804
rect 4476 69750 4478 69802
rect 4478 69750 4530 69802
rect 4530 69750 4532 69802
rect 4476 69748 4532 69750
rect 4580 69802 4636 69804
rect 4580 69750 4582 69802
rect 4582 69750 4634 69802
rect 4634 69750 4636 69802
rect 4580 69748 4636 69750
rect 4684 69802 4740 69804
rect 4684 69750 4686 69802
rect 4686 69750 4738 69802
rect 4738 69750 4740 69802
rect 4684 69748 4740 69750
rect 23884 69970 23940 69972
rect 23884 69918 23886 69970
rect 23886 69918 23938 69970
rect 23938 69918 23940 69970
rect 23884 69916 23940 69918
rect 19836 69018 19892 69020
rect 19836 68966 19838 69018
rect 19838 68966 19890 69018
rect 19890 68966 19892 69018
rect 19836 68964 19892 68966
rect 19940 69018 19996 69020
rect 19940 68966 19942 69018
rect 19942 68966 19994 69018
rect 19994 68966 19996 69018
rect 19940 68964 19996 68966
rect 20044 69018 20100 69020
rect 20044 68966 20046 69018
rect 20046 68966 20098 69018
rect 20098 68966 20100 69018
rect 20044 68964 20100 68966
rect 22204 68908 22260 68964
rect 22988 68908 23044 68964
rect 25340 69410 25396 69412
rect 25340 69358 25342 69410
rect 25342 69358 25394 69410
rect 25394 69358 25396 69410
rect 25340 69356 25396 69358
rect 25340 68908 25396 68964
rect 4476 68234 4532 68236
rect 4476 68182 4478 68234
rect 4478 68182 4530 68234
rect 4530 68182 4532 68234
rect 4476 68180 4532 68182
rect 4580 68234 4636 68236
rect 4580 68182 4582 68234
rect 4582 68182 4634 68234
rect 4634 68182 4636 68234
rect 4580 68180 4636 68182
rect 4684 68234 4740 68236
rect 4684 68182 4686 68234
rect 4686 68182 4738 68234
rect 4738 68182 4740 68234
rect 4684 68180 4740 68182
rect 20748 68124 20804 68180
rect 21308 68124 21364 68180
rect 19852 67788 19908 67844
rect 19836 67450 19892 67452
rect 19836 67398 19838 67450
rect 19838 67398 19890 67450
rect 19890 67398 19892 67450
rect 19836 67396 19892 67398
rect 19940 67450 19996 67452
rect 19940 67398 19942 67450
rect 19942 67398 19994 67450
rect 19994 67398 19996 67450
rect 19940 67396 19996 67398
rect 20044 67450 20100 67452
rect 20044 67398 20046 67450
rect 20046 67398 20098 67450
rect 20098 67398 20100 67450
rect 20044 67396 20100 67398
rect 20524 67282 20580 67284
rect 20524 67230 20526 67282
rect 20526 67230 20578 67282
rect 20578 67230 20580 67282
rect 20524 67228 20580 67230
rect 14252 66780 14308 66836
rect 4476 66666 4532 66668
rect 4476 66614 4478 66666
rect 4478 66614 4530 66666
rect 4530 66614 4532 66666
rect 4476 66612 4532 66614
rect 4580 66666 4636 66668
rect 4580 66614 4582 66666
rect 4582 66614 4634 66666
rect 4634 66614 4636 66666
rect 4580 66612 4636 66614
rect 4684 66666 4740 66668
rect 4684 66614 4686 66666
rect 4686 66614 4738 66666
rect 4738 66614 4740 66666
rect 4684 66612 4740 66614
rect 4476 65098 4532 65100
rect 4476 65046 4478 65098
rect 4478 65046 4530 65098
rect 4530 65046 4532 65098
rect 4476 65044 4532 65046
rect 4580 65098 4636 65100
rect 4580 65046 4582 65098
rect 4582 65046 4634 65098
rect 4634 65046 4636 65098
rect 4580 65044 4636 65046
rect 4684 65098 4740 65100
rect 4684 65046 4686 65098
rect 4686 65046 4738 65098
rect 4738 65046 4740 65098
rect 4684 65044 4740 65046
rect 10108 64764 10164 64820
rect 12684 65378 12740 65380
rect 12684 65326 12686 65378
rect 12686 65326 12738 65378
rect 12738 65326 12740 65378
rect 12684 65324 12740 65326
rect 10556 63756 10612 63812
rect 4476 63530 4532 63532
rect 4476 63478 4478 63530
rect 4478 63478 4530 63530
rect 4530 63478 4532 63530
rect 4476 63476 4532 63478
rect 4580 63530 4636 63532
rect 4580 63478 4582 63530
rect 4582 63478 4634 63530
rect 4634 63478 4636 63530
rect 4580 63476 4636 63478
rect 4684 63530 4740 63532
rect 4684 63478 4686 63530
rect 4686 63478 4738 63530
rect 4738 63478 4740 63530
rect 4684 63476 4740 63478
rect 11564 63922 11620 63924
rect 11564 63870 11566 63922
rect 11566 63870 11618 63922
rect 11618 63870 11620 63922
rect 11564 63868 11620 63870
rect 11452 63308 11508 63364
rect 12460 64034 12516 64036
rect 12460 63982 12462 64034
rect 12462 63982 12514 64034
rect 12514 63982 12516 64034
rect 12460 63980 12516 63982
rect 11900 63868 11956 63924
rect 4476 61962 4532 61964
rect 4476 61910 4478 61962
rect 4478 61910 4530 61962
rect 4530 61910 4532 61962
rect 4476 61908 4532 61910
rect 4580 61962 4636 61964
rect 4580 61910 4582 61962
rect 4582 61910 4634 61962
rect 4634 61910 4636 61962
rect 4580 61908 4636 61910
rect 4684 61962 4740 61964
rect 4684 61910 4686 61962
rect 4686 61910 4738 61962
rect 4738 61910 4740 61962
rect 4684 61908 4740 61910
rect 4476 60394 4532 60396
rect 4476 60342 4478 60394
rect 4478 60342 4530 60394
rect 4530 60342 4532 60394
rect 4476 60340 4532 60342
rect 4580 60394 4636 60396
rect 4580 60342 4582 60394
rect 4582 60342 4634 60394
rect 4634 60342 4636 60394
rect 4580 60340 4636 60342
rect 4684 60394 4740 60396
rect 4684 60342 4686 60394
rect 4686 60342 4738 60394
rect 4738 60342 4740 60394
rect 4684 60340 4740 60342
rect 4476 58826 4532 58828
rect 4476 58774 4478 58826
rect 4478 58774 4530 58826
rect 4530 58774 4532 58826
rect 4476 58772 4532 58774
rect 4580 58826 4636 58828
rect 4580 58774 4582 58826
rect 4582 58774 4634 58826
rect 4634 58774 4636 58826
rect 4580 58772 4636 58774
rect 4684 58826 4740 58828
rect 4684 58774 4686 58826
rect 4686 58774 4738 58826
rect 4738 58774 4740 58826
rect 4684 58772 4740 58774
rect 6188 58492 6244 58548
rect 4476 57258 4532 57260
rect 4476 57206 4478 57258
rect 4478 57206 4530 57258
rect 4530 57206 4532 57258
rect 4476 57204 4532 57206
rect 4580 57258 4636 57260
rect 4580 57206 4582 57258
rect 4582 57206 4634 57258
rect 4634 57206 4636 57258
rect 4580 57204 4636 57206
rect 4684 57258 4740 57260
rect 4684 57206 4686 57258
rect 4686 57206 4738 57258
rect 4738 57206 4740 57258
rect 4684 57204 4740 57206
rect 6860 56924 6916 56980
rect 4476 55690 4532 55692
rect 4476 55638 4478 55690
rect 4478 55638 4530 55690
rect 4530 55638 4532 55690
rect 4476 55636 4532 55638
rect 4580 55690 4636 55692
rect 4580 55638 4582 55690
rect 4582 55638 4634 55690
rect 4634 55638 4636 55690
rect 4580 55636 4636 55638
rect 4684 55690 4740 55692
rect 4684 55638 4686 55690
rect 4686 55638 4738 55690
rect 4738 55638 4740 55690
rect 4684 55636 4740 55638
rect 6412 56252 6468 56308
rect 7084 56252 7140 56308
rect 9996 62188 10052 62244
rect 10668 61570 10724 61572
rect 10668 61518 10670 61570
rect 10670 61518 10722 61570
rect 10722 61518 10724 61570
rect 10668 61516 10724 61518
rect 11452 62524 11508 62580
rect 11676 62524 11732 62580
rect 10332 61292 10388 61348
rect 10892 60956 10948 61012
rect 12572 63922 12628 63924
rect 12572 63870 12574 63922
rect 12574 63870 12626 63922
rect 12626 63870 12628 63922
rect 12572 63868 12628 63870
rect 12460 63810 12516 63812
rect 12460 63758 12462 63810
rect 12462 63758 12514 63810
rect 12514 63758 12516 63810
rect 12460 63756 12516 63758
rect 13132 64764 13188 64820
rect 14028 65660 14084 65716
rect 13916 65324 13972 65380
rect 14028 64482 14084 64484
rect 14028 64430 14030 64482
rect 14030 64430 14082 64482
rect 14082 64430 14084 64482
rect 14028 64428 14084 64430
rect 13804 64204 13860 64260
rect 13020 63922 13076 63924
rect 13020 63870 13022 63922
rect 13022 63870 13074 63922
rect 13074 63870 13076 63922
rect 13020 63868 13076 63870
rect 13692 63922 13748 63924
rect 13692 63870 13694 63922
rect 13694 63870 13746 63922
rect 13746 63870 13748 63922
rect 13692 63868 13748 63870
rect 13468 63756 13524 63812
rect 12572 63362 12628 63364
rect 12572 63310 12574 63362
rect 12574 63310 12626 63362
rect 12626 63310 12628 63362
rect 12572 63308 12628 63310
rect 12908 62578 12964 62580
rect 12908 62526 12910 62578
rect 12910 62526 12962 62578
rect 12962 62526 12964 62578
rect 12908 62524 12964 62526
rect 12460 62242 12516 62244
rect 12460 62190 12462 62242
rect 12462 62190 12514 62242
rect 12514 62190 12516 62242
rect 12460 62188 12516 62190
rect 13020 62188 13076 62244
rect 11900 62076 11956 62132
rect 11900 61570 11956 61572
rect 11900 61518 11902 61570
rect 11902 61518 11954 61570
rect 11954 61518 11956 61570
rect 11900 61516 11956 61518
rect 11788 61346 11844 61348
rect 11788 61294 11790 61346
rect 11790 61294 11842 61346
rect 11842 61294 11844 61346
rect 11788 61292 11844 61294
rect 11676 60956 11732 61012
rect 12572 61516 12628 61572
rect 13916 64034 13972 64036
rect 13916 63982 13918 64034
rect 13918 63982 13970 64034
rect 13970 63982 13972 64034
rect 13916 63980 13972 63982
rect 15260 66834 15316 66836
rect 15260 66782 15262 66834
rect 15262 66782 15314 66834
rect 15314 66782 15316 66834
rect 15260 66780 15316 66782
rect 14924 65660 14980 65716
rect 14364 64764 14420 64820
rect 14476 64540 14532 64596
rect 15260 65436 15316 65492
rect 16380 65714 16436 65716
rect 16380 65662 16382 65714
rect 16382 65662 16434 65714
rect 16434 65662 16436 65714
rect 16380 65660 16436 65662
rect 16492 65602 16548 65604
rect 16492 65550 16494 65602
rect 16494 65550 16546 65602
rect 16546 65550 16548 65602
rect 16492 65548 16548 65550
rect 21084 67058 21140 67060
rect 21084 67006 21086 67058
rect 21086 67006 21138 67058
rect 21138 67006 21140 67058
rect 21084 67004 21140 67006
rect 20188 66050 20244 66052
rect 20188 65998 20190 66050
rect 20190 65998 20242 66050
rect 20242 65998 20244 66050
rect 20188 65996 20244 65998
rect 19836 65882 19892 65884
rect 19836 65830 19838 65882
rect 19838 65830 19890 65882
rect 19890 65830 19892 65882
rect 19836 65828 19892 65830
rect 19940 65882 19996 65884
rect 19940 65830 19942 65882
rect 19942 65830 19994 65882
rect 19994 65830 19996 65882
rect 19940 65828 19996 65830
rect 20044 65882 20100 65884
rect 20044 65830 20046 65882
rect 20046 65830 20098 65882
rect 20098 65830 20100 65882
rect 20044 65828 20100 65830
rect 17500 65548 17556 65604
rect 18508 65602 18564 65604
rect 18508 65550 18510 65602
rect 18510 65550 18562 65602
rect 18562 65550 18564 65602
rect 18508 65548 18564 65550
rect 15036 64540 15092 64596
rect 14924 64034 14980 64036
rect 14924 63982 14926 64034
rect 14926 63982 14978 64034
rect 14978 63982 14980 64034
rect 14924 63980 14980 63982
rect 14700 63756 14756 63812
rect 15148 64428 15204 64484
rect 15372 64092 15428 64148
rect 15596 64204 15652 64260
rect 15932 63980 15988 64036
rect 16380 64876 16436 64932
rect 17388 64540 17444 64596
rect 16380 64428 16436 64484
rect 16156 64316 16212 64372
rect 15260 63756 15316 63812
rect 12908 61346 12964 61348
rect 12908 61294 12910 61346
rect 12910 61294 12962 61346
rect 12962 61294 12964 61346
rect 12908 61292 12964 61294
rect 12796 61010 12852 61012
rect 12796 60958 12798 61010
rect 12798 60958 12850 61010
rect 12850 60958 12852 61010
rect 12796 60956 12852 60958
rect 13132 60786 13188 60788
rect 13132 60734 13134 60786
rect 13134 60734 13186 60786
rect 13186 60734 13188 60786
rect 13132 60732 13188 60734
rect 13580 60732 13636 60788
rect 13916 60732 13972 60788
rect 9660 58546 9716 58548
rect 9660 58494 9662 58546
rect 9662 58494 9714 58546
rect 9714 58494 9716 58546
rect 9660 58492 9716 58494
rect 9548 57820 9604 57876
rect 8988 56978 9044 56980
rect 8988 56926 8990 56978
rect 8990 56926 9042 56978
rect 9042 56926 9044 56978
rect 8988 56924 9044 56926
rect 9100 56754 9156 56756
rect 9100 56702 9102 56754
rect 9102 56702 9154 56754
rect 9154 56702 9156 56754
rect 9100 56700 9156 56702
rect 8876 56588 8932 56644
rect 9324 56364 9380 56420
rect 6972 56082 7028 56084
rect 6972 56030 6974 56082
rect 6974 56030 7026 56082
rect 7026 56030 7028 56082
rect 6972 56028 7028 56030
rect 6636 55804 6692 55860
rect 4476 54122 4532 54124
rect 4476 54070 4478 54122
rect 4478 54070 4530 54122
rect 4530 54070 4532 54122
rect 4476 54068 4532 54070
rect 4580 54122 4636 54124
rect 4580 54070 4582 54122
rect 4582 54070 4634 54122
rect 4634 54070 4636 54122
rect 4580 54068 4636 54070
rect 4684 54122 4740 54124
rect 4684 54070 4686 54122
rect 4686 54070 4738 54122
rect 4738 54070 4740 54122
rect 4684 54068 4740 54070
rect 5292 53788 5348 53844
rect 6636 53842 6692 53844
rect 6636 53790 6638 53842
rect 6638 53790 6690 53842
rect 6690 53790 6692 53842
rect 6636 53788 6692 53790
rect 6636 53506 6692 53508
rect 6636 53454 6638 53506
rect 6638 53454 6690 53506
rect 6690 53454 6692 53506
rect 6636 53452 6692 53454
rect 6748 53004 6804 53060
rect 4476 52554 4532 52556
rect 4476 52502 4478 52554
rect 4478 52502 4530 52554
rect 4530 52502 4532 52554
rect 4476 52500 4532 52502
rect 4580 52554 4636 52556
rect 4580 52502 4582 52554
rect 4582 52502 4634 52554
rect 4634 52502 4636 52554
rect 4580 52500 4636 52502
rect 4684 52554 4740 52556
rect 4684 52502 4686 52554
rect 4686 52502 4738 52554
rect 4738 52502 4740 52554
rect 4684 52500 4740 52502
rect 6524 52332 6580 52388
rect 5292 52220 5348 52276
rect 6636 52274 6692 52276
rect 6636 52222 6638 52274
rect 6638 52222 6690 52274
rect 6690 52222 6692 52274
rect 6636 52220 6692 52222
rect 8092 56028 8148 56084
rect 7868 55858 7924 55860
rect 7868 55806 7870 55858
rect 7870 55806 7922 55858
rect 7922 55806 7924 55858
rect 7868 55804 7924 55806
rect 7644 54738 7700 54740
rect 7644 54686 7646 54738
rect 7646 54686 7698 54738
rect 7698 54686 7700 54738
rect 7644 54684 7700 54686
rect 9660 56588 9716 56644
rect 10444 57650 10500 57652
rect 10444 57598 10446 57650
rect 10446 57598 10498 57650
rect 10498 57598 10500 57650
rect 10444 57596 10500 57598
rect 10220 56642 10276 56644
rect 10220 56590 10222 56642
rect 10222 56590 10274 56642
rect 10274 56590 10276 56642
rect 10220 56588 10276 56590
rect 10332 56364 10388 56420
rect 10444 56700 10500 56756
rect 9548 56028 9604 56084
rect 10108 56082 10164 56084
rect 10108 56030 10110 56082
rect 10110 56030 10162 56082
rect 10162 56030 10164 56082
rect 10108 56028 10164 56030
rect 8652 54738 8708 54740
rect 8652 54686 8654 54738
rect 8654 54686 8706 54738
rect 8706 54686 8708 54738
rect 8652 54684 8708 54686
rect 6972 53116 7028 53172
rect 4476 50986 4532 50988
rect 4476 50934 4478 50986
rect 4478 50934 4530 50986
rect 4530 50934 4532 50986
rect 4476 50932 4532 50934
rect 4580 50986 4636 50988
rect 4580 50934 4582 50986
rect 4582 50934 4634 50986
rect 4634 50934 4636 50986
rect 4580 50932 4636 50934
rect 4684 50986 4740 50988
rect 4684 50934 4686 50986
rect 4686 50934 4738 50986
rect 4738 50934 4740 50986
rect 4684 50932 4740 50934
rect 4476 49418 4532 49420
rect 4476 49366 4478 49418
rect 4478 49366 4530 49418
rect 4530 49366 4532 49418
rect 4476 49364 4532 49366
rect 4580 49418 4636 49420
rect 4580 49366 4582 49418
rect 4582 49366 4634 49418
rect 4634 49366 4636 49418
rect 4580 49364 4636 49366
rect 4684 49418 4740 49420
rect 4684 49366 4686 49418
rect 4686 49366 4738 49418
rect 4738 49366 4740 49418
rect 4684 49364 4740 49366
rect 8092 53506 8148 53508
rect 8092 53454 8094 53506
rect 8094 53454 8146 53506
rect 8146 53454 8148 53506
rect 8092 53452 8148 53454
rect 8428 53170 8484 53172
rect 8428 53118 8430 53170
rect 8430 53118 8482 53170
rect 8482 53118 8484 53170
rect 8428 53116 8484 53118
rect 9436 53676 9492 53732
rect 8652 53116 8708 53172
rect 7756 53058 7812 53060
rect 7756 53006 7758 53058
rect 7758 53006 7810 53058
rect 7810 53006 7812 53058
rect 7756 53004 7812 53006
rect 8316 52892 8372 52948
rect 8092 52386 8148 52388
rect 8092 52334 8094 52386
rect 8094 52334 8146 52386
rect 8146 52334 8148 52386
rect 8092 52332 8148 52334
rect 4844 49084 4900 49140
rect 5404 50652 5460 50708
rect 4284 48860 4340 48916
rect 4732 48914 4788 48916
rect 4732 48862 4734 48914
rect 4734 48862 4786 48914
rect 4786 48862 4788 48914
rect 4732 48860 4788 48862
rect 4476 47850 4532 47852
rect 4476 47798 4478 47850
rect 4478 47798 4530 47850
rect 4530 47798 4532 47850
rect 4476 47796 4532 47798
rect 4580 47850 4636 47852
rect 4580 47798 4582 47850
rect 4582 47798 4634 47850
rect 4634 47798 4636 47850
rect 4580 47796 4636 47798
rect 4684 47850 4740 47852
rect 4684 47798 4686 47850
rect 4686 47798 4738 47850
rect 4738 47798 4740 47850
rect 4684 47796 4740 47798
rect 4844 47404 4900 47460
rect 4620 46956 4676 47012
rect 4476 46282 4532 46284
rect 4476 46230 4478 46282
rect 4478 46230 4530 46282
rect 4530 46230 4532 46282
rect 4476 46228 4532 46230
rect 4580 46282 4636 46284
rect 4580 46230 4582 46282
rect 4582 46230 4634 46282
rect 4634 46230 4636 46282
rect 4580 46228 4636 46230
rect 4684 46282 4740 46284
rect 4684 46230 4686 46282
rect 4686 46230 4738 46282
rect 4738 46230 4740 46282
rect 4684 46228 4740 46230
rect 4476 44714 4532 44716
rect 4476 44662 4478 44714
rect 4478 44662 4530 44714
rect 4530 44662 4532 44714
rect 4476 44660 4532 44662
rect 4580 44714 4636 44716
rect 4580 44662 4582 44714
rect 4582 44662 4634 44714
rect 4634 44662 4636 44714
rect 4580 44660 4636 44662
rect 4684 44714 4740 44716
rect 4684 44662 4686 44714
rect 4686 44662 4738 44714
rect 4738 44662 4740 44714
rect 4684 44660 4740 44662
rect 5292 46956 5348 47012
rect 5292 46562 5348 46564
rect 5292 46510 5294 46562
rect 5294 46510 5346 46562
rect 5346 46510 5348 46562
rect 5292 46508 5348 46510
rect 7084 50482 7140 50484
rect 7084 50430 7086 50482
rect 7086 50430 7138 50482
rect 7138 50430 7140 50482
rect 7084 50428 7140 50430
rect 5628 49084 5684 49140
rect 6412 48412 6468 48468
rect 6300 47964 6356 48020
rect 5852 46956 5908 47012
rect 7308 50428 7364 50484
rect 7868 50428 7924 50484
rect 7196 49980 7252 50036
rect 7756 50316 7812 50372
rect 7420 48748 7476 48804
rect 6860 47964 6916 48020
rect 6412 46844 6468 46900
rect 5404 46284 5460 46340
rect 7084 48466 7140 48468
rect 7084 48414 7086 48466
rect 7086 48414 7138 48466
rect 7138 48414 7140 48466
rect 7084 48412 7140 48414
rect 7196 48354 7252 48356
rect 7196 48302 7198 48354
rect 7198 48302 7250 48354
rect 7250 48302 7252 48354
rect 7196 48300 7252 48302
rect 8316 50316 8372 50372
rect 8764 50428 8820 50484
rect 9436 50482 9492 50484
rect 9436 50430 9438 50482
rect 9438 50430 9490 50482
rect 9490 50430 9492 50482
rect 9436 50428 9492 50430
rect 10780 56364 10836 56420
rect 11340 57596 11396 57652
rect 13020 58492 13076 58548
rect 10892 56028 10948 56084
rect 12236 57820 12292 57876
rect 10668 55132 10724 55188
rect 12796 57650 12852 57652
rect 12796 57598 12798 57650
rect 12798 57598 12850 57650
rect 12850 57598 12852 57650
rect 12796 57596 12852 57598
rect 13804 58380 13860 58436
rect 13468 57820 13524 57876
rect 14476 61292 14532 61348
rect 14364 58210 14420 58212
rect 14364 58158 14366 58210
rect 14366 58158 14418 58210
rect 14418 58158 14420 58210
rect 14364 58156 14420 58158
rect 13692 56754 13748 56756
rect 13692 56702 13694 56754
rect 13694 56702 13746 56754
rect 13746 56702 13748 56754
rect 13692 56700 13748 56702
rect 11452 55186 11508 55188
rect 11452 55134 11454 55186
rect 11454 55134 11506 55186
rect 11506 55134 11508 55186
rect 11452 55132 11508 55134
rect 11228 54236 11284 54292
rect 10556 53730 10612 53732
rect 10556 53678 10558 53730
rect 10558 53678 10610 53730
rect 10610 53678 10612 53730
rect 10556 53676 10612 53678
rect 13468 55410 13524 55412
rect 13468 55358 13470 55410
rect 13470 55358 13522 55410
rect 13522 55358 13524 55410
rect 13468 55356 13524 55358
rect 12460 54236 12516 54292
rect 11676 53170 11732 53172
rect 11676 53118 11678 53170
rect 11678 53118 11730 53170
rect 11730 53118 11732 53170
rect 11676 53116 11732 53118
rect 12684 53004 12740 53060
rect 9660 52892 9716 52948
rect 11116 52892 11172 52948
rect 12012 52946 12068 52948
rect 12012 52894 12014 52946
rect 12014 52894 12066 52946
rect 12066 52894 12068 52946
rect 12012 52892 12068 52894
rect 11452 52162 11508 52164
rect 11452 52110 11454 52162
rect 11454 52110 11506 52162
rect 11506 52110 11508 52162
rect 11452 52108 11508 52110
rect 9772 50540 9828 50596
rect 12572 52162 12628 52164
rect 12572 52110 12574 52162
rect 12574 52110 12626 52162
rect 12626 52110 12628 52162
rect 12572 52108 12628 52110
rect 11788 51436 11844 51492
rect 10108 50764 10164 50820
rect 9884 50428 9940 50484
rect 8316 49980 8372 50036
rect 7756 48354 7812 48356
rect 7756 48302 7758 48354
rect 7758 48302 7810 48354
rect 7810 48302 7812 48354
rect 7756 48300 7812 48302
rect 7420 47964 7476 48020
rect 7756 46844 7812 46900
rect 9996 50316 10052 50372
rect 8540 49138 8596 49140
rect 8540 49086 8542 49138
rect 8542 49086 8594 49138
rect 8594 49086 8596 49138
rect 8540 49084 8596 49086
rect 8428 48860 8484 48916
rect 8652 48354 8708 48356
rect 8652 48302 8654 48354
rect 8654 48302 8706 48354
rect 8706 48302 8708 48354
rect 8652 48300 8708 48302
rect 9660 49810 9716 49812
rect 9660 49758 9662 49810
rect 9662 49758 9714 49810
rect 9714 49758 9716 49810
rect 9660 49756 9716 49758
rect 8988 49138 9044 49140
rect 8988 49086 8990 49138
rect 8990 49086 9042 49138
rect 9042 49086 9044 49138
rect 8988 49084 9044 49086
rect 11228 50540 11284 50596
rect 10892 50482 10948 50484
rect 10892 50430 10894 50482
rect 10894 50430 10946 50482
rect 10946 50430 10948 50482
rect 10892 50428 10948 50430
rect 10332 49698 10388 49700
rect 10332 49646 10334 49698
rect 10334 49646 10386 49698
rect 10386 49646 10388 49698
rect 10332 49644 10388 49646
rect 10556 48860 10612 48916
rect 8876 48802 8932 48804
rect 8876 48750 8878 48802
rect 8878 48750 8930 48802
rect 8930 48750 8932 48802
rect 8876 48748 8932 48750
rect 8988 48300 9044 48356
rect 8428 46844 8484 46900
rect 8092 46562 8148 46564
rect 8092 46510 8094 46562
rect 8094 46510 8146 46562
rect 8146 46510 8148 46562
rect 8092 46508 8148 46510
rect 7980 46172 8036 46228
rect 6524 45778 6580 45780
rect 6524 45726 6526 45778
rect 6526 45726 6578 45778
rect 6578 45726 6580 45778
rect 6524 45724 6580 45726
rect 5180 44604 5236 44660
rect 6636 45612 6692 45668
rect 7532 45778 7588 45780
rect 7532 45726 7534 45778
rect 7534 45726 7586 45778
rect 7586 45726 7588 45778
rect 7532 45724 7588 45726
rect 6860 45500 6916 45556
rect 7644 45666 7700 45668
rect 7644 45614 7646 45666
rect 7646 45614 7698 45666
rect 7698 45614 7700 45666
rect 7644 45612 7700 45614
rect 7756 45500 7812 45556
rect 8428 45778 8484 45780
rect 8428 45726 8430 45778
rect 8430 45726 8482 45778
rect 8482 45726 8484 45778
rect 8428 45724 8484 45726
rect 7980 45276 8036 45332
rect 8092 45500 8148 45556
rect 7420 44156 7476 44212
rect 6412 43708 6468 43764
rect 6636 44044 6692 44100
rect 4476 43146 4532 43148
rect 4476 43094 4478 43146
rect 4478 43094 4530 43146
rect 4530 43094 4532 43146
rect 4476 43092 4532 43094
rect 4580 43146 4636 43148
rect 4580 43094 4582 43146
rect 4582 43094 4634 43146
rect 4634 43094 4636 43146
rect 4580 43092 4636 43094
rect 4684 43146 4740 43148
rect 4684 43094 4686 43146
rect 4686 43094 4738 43146
rect 4738 43094 4740 43146
rect 4684 43092 4740 43094
rect 4844 42924 4900 42980
rect 7644 43708 7700 43764
rect 8764 45724 8820 45780
rect 8652 45330 8708 45332
rect 8652 45278 8654 45330
rect 8654 45278 8706 45330
rect 8706 45278 8708 45330
rect 8652 45276 8708 45278
rect 10108 48354 10164 48356
rect 10108 48302 10110 48354
rect 10110 48302 10162 48354
rect 10162 48302 10164 48354
rect 10108 48300 10164 48302
rect 9548 46396 9604 46452
rect 10108 48076 10164 48132
rect 10556 47180 10612 47236
rect 10220 46396 10276 46452
rect 10332 46956 10388 47012
rect 8988 45778 9044 45780
rect 8988 45726 8990 45778
rect 8990 45726 9042 45778
rect 9042 45726 9044 45778
rect 8988 45724 9044 45726
rect 9548 45724 9604 45780
rect 8876 45500 8932 45556
rect 9772 45164 9828 45220
rect 9660 44828 9716 44884
rect 8988 44210 9044 44212
rect 8988 44158 8990 44210
rect 8990 44158 9042 44210
rect 9042 44158 9044 44210
rect 8988 44156 9044 44158
rect 9548 43820 9604 43876
rect 9324 42866 9380 42868
rect 9324 42814 9326 42866
rect 9326 42814 9378 42866
rect 9378 42814 9380 42866
rect 9324 42812 9380 42814
rect 6636 41804 6692 41860
rect 4476 41578 4532 41580
rect 4476 41526 4478 41578
rect 4478 41526 4530 41578
rect 4530 41526 4532 41578
rect 4476 41524 4532 41526
rect 4580 41578 4636 41580
rect 4580 41526 4582 41578
rect 4582 41526 4634 41578
rect 4634 41526 4636 41578
rect 4580 41524 4636 41526
rect 4684 41578 4740 41580
rect 4684 41526 4686 41578
rect 4686 41526 4738 41578
rect 4738 41526 4740 41578
rect 4684 41524 4740 41526
rect 4172 40572 4228 40628
rect 9436 40572 9492 40628
rect 3164 40348 3220 40404
rect 9436 40348 9492 40404
rect 4476 40010 4532 40012
rect 4476 39958 4478 40010
rect 4478 39958 4530 40010
rect 4530 39958 4532 40010
rect 4476 39956 4532 39958
rect 4580 40010 4636 40012
rect 4580 39958 4582 40010
rect 4582 39958 4634 40010
rect 4634 39958 4636 40010
rect 4580 39956 4636 39958
rect 4684 40010 4740 40012
rect 4684 39958 4686 40010
rect 4686 39958 4738 40010
rect 4738 39958 4740 40010
rect 4684 39956 4740 39958
rect 5852 39900 5908 39956
rect 2940 39676 2996 39732
rect 4284 39788 4340 39844
rect 2044 39506 2100 39508
rect 2044 39454 2046 39506
rect 2046 39454 2098 39506
rect 2098 39454 2100 39506
rect 2044 39452 2100 39454
rect 1708 39004 1764 39060
rect 2492 39004 2548 39060
rect 1932 38610 1988 38612
rect 1932 38558 1934 38610
rect 1934 38558 1986 38610
rect 1986 38558 1988 38610
rect 1932 38556 1988 38558
rect 4476 38442 4532 38444
rect 4476 38390 4478 38442
rect 4478 38390 4530 38442
rect 4530 38390 4532 38442
rect 4476 38388 4532 38390
rect 4580 38442 4636 38444
rect 4580 38390 4582 38442
rect 4582 38390 4634 38442
rect 4634 38390 4636 38442
rect 4580 38388 4636 38390
rect 4684 38442 4740 38444
rect 4684 38390 4686 38442
rect 4686 38390 4738 38442
rect 4738 38390 4740 38442
rect 4684 38388 4740 38390
rect 2044 37826 2100 37828
rect 2044 37774 2046 37826
rect 2046 37774 2098 37826
rect 2098 37774 2100 37826
rect 2044 37772 2100 37774
rect 1708 37660 1764 37716
rect 2492 37660 2548 37716
rect 2716 37660 2772 37716
rect 1708 36988 1764 37044
rect 1932 36594 1988 36596
rect 1932 36542 1934 36594
rect 1934 36542 1986 36594
rect 1986 36542 1988 36594
rect 1932 36540 1988 36542
rect 2044 35810 2100 35812
rect 2044 35758 2046 35810
rect 2046 35758 2098 35810
rect 2098 35758 2100 35810
rect 2044 35756 2100 35758
rect 1708 35698 1764 35700
rect 1708 35646 1710 35698
rect 1710 35646 1762 35698
rect 1762 35646 1764 35698
rect 1708 35644 1764 35646
rect 2492 36988 2548 37044
rect 4476 36874 4532 36876
rect 4476 36822 4478 36874
rect 4478 36822 4530 36874
rect 4530 36822 4532 36874
rect 4476 36820 4532 36822
rect 4580 36874 4636 36876
rect 4580 36822 4582 36874
rect 4582 36822 4634 36874
rect 4634 36822 4636 36874
rect 4580 36820 4636 36822
rect 4684 36874 4740 36876
rect 4684 36822 4686 36874
rect 4686 36822 4738 36874
rect 4738 36822 4740 36874
rect 4684 36820 4740 36822
rect 4844 36876 4900 36932
rect 4172 36482 4228 36484
rect 4172 36430 4174 36482
rect 4174 36430 4226 36482
rect 4226 36430 4228 36482
rect 4172 36428 4228 36430
rect 4844 36428 4900 36484
rect 2156 35532 2212 35588
rect 2380 34972 2436 35028
rect 2492 35644 2548 35700
rect 4476 35306 4532 35308
rect 4476 35254 4478 35306
rect 4478 35254 4530 35306
rect 4530 35254 4532 35306
rect 4476 35252 4532 35254
rect 4580 35306 4636 35308
rect 4580 35254 4582 35306
rect 4582 35254 4634 35306
rect 4634 35254 4636 35306
rect 4580 35252 4636 35254
rect 4684 35306 4740 35308
rect 4684 35254 4686 35306
rect 4686 35254 4738 35306
rect 4738 35254 4740 35306
rect 4684 35252 4740 35254
rect 3164 34972 3220 35028
rect 2044 34690 2100 34692
rect 2044 34638 2046 34690
rect 2046 34638 2098 34690
rect 2098 34638 2100 34690
rect 2044 34636 2100 34638
rect 1708 34300 1764 34356
rect 2940 34300 2996 34356
rect 4284 33964 4340 34020
rect 4732 34018 4788 34020
rect 4732 33966 4734 34018
rect 4734 33966 4786 34018
rect 4786 33966 4788 34018
rect 4732 33964 4788 33966
rect 1932 33906 1988 33908
rect 1932 33854 1934 33906
rect 1934 33854 1986 33906
rect 1986 33854 1988 33906
rect 1932 33852 1988 33854
rect 4476 33738 4532 33740
rect 4476 33686 4478 33738
rect 4478 33686 4530 33738
rect 4530 33686 4532 33738
rect 4476 33684 4532 33686
rect 4580 33738 4636 33740
rect 4580 33686 4582 33738
rect 4582 33686 4634 33738
rect 4634 33686 4636 33738
rect 4580 33684 4636 33686
rect 4684 33738 4740 33740
rect 4684 33686 4686 33738
rect 4686 33686 4738 33738
rect 4738 33686 4740 33738
rect 4684 33684 4740 33686
rect 2044 33122 2100 33124
rect 2044 33070 2046 33122
rect 2046 33070 2098 33122
rect 2098 33070 2100 33122
rect 2044 33068 2100 33070
rect 1708 32956 1764 33012
rect 2492 32956 2548 33012
rect 5068 32956 5124 33012
rect 1708 32284 1764 32340
rect 1932 31890 1988 31892
rect 1932 31838 1934 31890
rect 1934 31838 1986 31890
rect 1986 31838 1988 31890
rect 1932 31836 1988 31838
rect 2492 32284 2548 32340
rect 4476 32170 4532 32172
rect 4476 32118 4478 32170
rect 4478 32118 4530 32170
rect 4530 32118 4532 32170
rect 4476 32116 4532 32118
rect 4580 32170 4636 32172
rect 4580 32118 4582 32170
rect 4582 32118 4634 32170
rect 4634 32118 4636 32170
rect 4580 32116 4636 32118
rect 4684 32170 4740 32172
rect 4684 32118 4686 32170
rect 4686 32118 4738 32170
rect 4738 32118 4740 32170
rect 4684 32116 4740 32118
rect 4172 31778 4228 31780
rect 4172 31726 4174 31778
rect 4174 31726 4226 31778
rect 4226 31726 4228 31778
rect 4172 31724 4228 31726
rect 4844 31724 4900 31780
rect 2044 31500 2100 31556
rect 2044 31218 2100 31220
rect 2044 31166 2046 31218
rect 2046 31166 2098 31218
rect 2098 31166 2100 31218
rect 2044 31164 2100 31166
rect 6748 39564 6804 39620
rect 6748 37660 6804 37716
rect 8428 37996 8484 38052
rect 9100 38050 9156 38052
rect 9100 37998 9102 38050
rect 9102 37998 9154 38050
rect 9154 37998 9156 38050
rect 9100 37996 9156 37998
rect 9212 36988 9268 37044
rect 9100 35420 9156 35476
rect 5852 31164 5908 31220
rect 1708 30994 1764 30996
rect 1708 30942 1710 30994
rect 1710 30942 1762 30994
rect 1762 30942 1764 30994
rect 1708 30940 1764 30942
rect 2380 30828 2436 30884
rect 2044 30492 2100 30548
rect 2380 30268 2436 30324
rect 2492 30940 2548 30996
rect 3164 30882 3220 30884
rect 3164 30830 3166 30882
rect 3166 30830 3218 30882
rect 3218 30830 3220 30882
rect 3164 30828 3220 30830
rect 4476 30602 4532 30604
rect 4476 30550 4478 30602
rect 4478 30550 4530 30602
rect 4530 30550 4532 30602
rect 4476 30548 4532 30550
rect 4580 30602 4636 30604
rect 4580 30550 4582 30602
rect 4582 30550 4634 30602
rect 4634 30550 4636 30602
rect 4580 30548 4636 30550
rect 4684 30602 4740 30604
rect 4684 30550 4686 30602
rect 4686 30550 4738 30602
rect 4738 30550 4740 30602
rect 4684 30548 4740 30550
rect 2716 30380 2772 30436
rect 10444 46284 10500 46340
rect 10892 49196 10948 49252
rect 10668 46002 10724 46004
rect 10668 45950 10670 46002
rect 10670 45950 10722 46002
rect 10722 45950 10724 46002
rect 10668 45948 10724 45950
rect 10780 45890 10836 45892
rect 10780 45838 10782 45890
rect 10782 45838 10834 45890
rect 10834 45838 10836 45890
rect 10780 45836 10836 45838
rect 10220 44268 10276 44324
rect 9772 43148 9828 43204
rect 9884 43596 9940 43652
rect 10444 43426 10500 43428
rect 10444 43374 10446 43426
rect 10446 43374 10498 43426
rect 10498 43374 10500 43426
rect 10444 43372 10500 43374
rect 10220 42866 10276 42868
rect 10220 42814 10222 42866
rect 10222 42814 10274 42866
rect 10274 42814 10276 42866
rect 10220 42812 10276 42814
rect 10220 42530 10276 42532
rect 10220 42478 10222 42530
rect 10222 42478 10274 42530
rect 10274 42478 10276 42530
rect 10220 42476 10276 42478
rect 9996 42140 10052 42196
rect 9884 41916 9940 41972
rect 9884 41746 9940 41748
rect 9884 41694 9886 41746
rect 9886 41694 9938 41746
rect 9938 41694 9940 41746
rect 9884 41692 9940 41694
rect 9772 41020 9828 41076
rect 9772 38668 9828 38724
rect 10444 42028 10500 42084
rect 10108 41356 10164 41412
rect 10556 41858 10612 41860
rect 10556 41806 10558 41858
rect 10558 41806 10610 41858
rect 10610 41806 10612 41858
rect 10556 41804 10612 41806
rect 10444 41356 10500 41412
rect 10444 39618 10500 39620
rect 10444 39566 10446 39618
rect 10446 39566 10498 39618
rect 10498 39566 10500 39618
rect 10444 39564 10500 39566
rect 13580 53058 13636 53060
rect 13580 53006 13582 53058
rect 13582 53006 13634 53058
rect 13634 53006 13636 53058
rect 13580 53004 13636 53006
rect 13916 52780 13972 52836
rect 13804 52668 13860 52724
rect 13020 52162 13076 52164
rect 13020 52110 13022 52162
rect 13022 52110 13074 52162
rect 13074 52110 13076 52162
rect 13020 52108 13076 52110
rect 12236 50764 12292 50820
rect 12348 50540 12404 50596
rect 12908 50594 12964 50596
rect 12908 50542 12910 50594
rect 12910 50542 12962 50594
rect 12962 50542 12964 50594
rect 12908 50540 12964 50542
rect 13132 50540 13188 50596
rect 12796 50482 12852 50484
rect 12796 50430 12798 50482
rect 12798 50430 12850 50482
rect 12850 50430 12852 50482
rect 12796 50428 12852 50430
rect 11788 49756 11844 49812
rect 12012 50316 12068 50372
rect 11452 49196 11508 49252
rect 11228 48972 11284 49028
rect 11116 48130 11172 48132
rect 11116 48078 11118 48130
rect 11118 48078 11170 48130
rect 11170 48078 11172 48130
rect 11116 48076 11172 48078
rect 11676 48748 11732 48804
rect 13468 50482 13524 50484
rect 13468 50430 13470 50482
rect 13470 50430 13522 50482
rect 13522 50430 13524 50482
rect 13468 50428 13524 50430
rect 13132 50316 13188 50372
rect 13692 52108 13748 52164
rect 14476 56642 14532 56644
rect 14476 56590 14478 56642
rect 14478 56590 14530 56642
rect 14530 56590 14532 56642
rect 14476 56588 14532 56590
rect 16268 64146 16324 64148
rect 16268 64094 16270 64146
rect 16270 64094 16322 64146
rect 16322 64094 16324 64146
rect 16268 64092 16324 64094
rect 16604 64204 16660 64260
rect 16604 63922 16660 63924
rect 16604 63870 16606 63922
rect 16606 63870 16658 63922
rect 16658 63870 16660 63922
rect 16604 63868 16660 63870
rect 17388 63922 17444 63924
rect 17388 63870 17390 63922
rect 17390 63870 17442 63922
rect 17442 63870 17444 63922
rect 17388 63868 17444 63870
rect 17724 65490 17780 65492
rect 17724 65438 17726 65490
rect 17726 65438 17778 65490
rect 17778 65438 17780 65490
rect 17724 65436 17780 65438
rect 17836 64876 17892 64932
rect 17948 64764 18004 64820
rect 19964 64764 20020 64820
rect 17612 64316 17668 64372
rect 15036 62188 15092 62244
rect 15932 62242 15988 62244
rect 15932 62190 15934 62242
rect 15934 62190 15986 62242
rect 15986 62190 15988 62242
rect 15932 62188 15988 62190
rect 16156 60898 16212 60900
rect 16156 60846 16158 60898
rect 16158 60846 16210 60898
rect 16210 60846 16212 60898
rect 16156 60844 16212 60846
rect 16044 60732 16100 60788
rect 17500 63084 17556 63140
rect 17388 60844 17444 60900
rect 17948 64204 18004 64260
rect 19836 64314 19892 64316
rect 19836 64262 19838 64314
rect 19838 64262 19890 64314
rect 19890 64262 19892 64314
rect 19836 64260 19892 64262
rect 19940 64314 19996 64316
rect 19940 64262 19942 64314
rect 19942 64262 19994 64314
rect 19994 64262 19996 64314
rect 19940 64260 19996 64262
rect 20044 64314 20100 64316
rect 20044 64262 20046 64314
rect 20046 64262 20098 64314
rect 20098 64262 20100 64314
rect 20044 64260 20100 64262
rect 20524 66892 20580 66948
rect 22876 68124 22932 68180
rect 21868 67842 21924 67844
rect 21868 67790 21870 67842
rect 21870 67790 21922 67842
rect 21922 67790 21924 67842
rect 21868 67788 21924 67790
rect 22428 67788 22484 67844
rect 21308 67730 21364 67732
rect 21308 67678 21310 67730
rect 21310 67678 21362 67730
rect 21362 67678 21364 67730
rect 21308 67676 21364 67678
rect 21980 67730 22036 67732
rect 21980 67678 21982 67730
rect 21982 67678 22034 67730
rect 22034 67678 22036 67730
rect 21980 67676 22036 67678
rect 22092 67618 22148 67620
rect 22092 67566 22094 67618
rect 22094 67566 22146 67618
rect 22146 67566 22148 67618
rect 22092 67564 22148 67566
rect 22204 67340 22260 67396
rect 21308 66892 21364 66948
rect 21420 66386 21476 66388
rect 21420 66334 21422 66386
rect 21422 66334 21474 66386
rect 21474 66334 21476 66386
rect 21420 66332 21476 66334
rect 20524 65996 20580 66052
rect 18732 63138 18788 63140
rect 18732 63086 18734 63138
rect 18734 63086 18786 63138
rect 18786 63086 18788 63138
rect 18732 63084 18788 63086
rect 19740 63138 19796 63140
rect 19740 63086 19742 63138
rect 19742 63086 19794 63138
rect 19794 63086 19796 63138
rect 19740 63084 19796 63086
rect 21420 65996 21476 66052
rect 17948 62578 18004 62580
rect 17948 62526 17950 62578
rect 17950 62526 18002 62578
rect 18002 62526 18004 62578
rect 17948 62524 18004 62526
rect 18508 62524 18564 62580
rect 17724 61516 17780 61572
rect 16604 60786 16660 60788
rect 16604 60734 16606 60786
rect 16606 60734 16658 60786
rect 16658 60734 16660 60786
rect 16604 60732 16660 60734
rect 15708 60508 15764 60564
rect 14700 59724 14756 59780
rect 15708 59778 15764 59780
rect 15708 59726 15710 59778
rect 15710 59726 15762 59778
rect 15762 59726 15764 59778
rect 15708 59724 15764 59726
rect 16492 59890 16548 59892
rect 16492 59838 16494 59890
rect 16494 59838 16546 59890
rect 16546 59838 16548 59890
rect 16492 59836 16548 59838
rect 14924 58546 14980 58548
rect 14924 58494 14926 58546
rect 14926 58494 14978 58546
rect 14978 58494 14980 58546
rect 14924 58492 14980 58494
rect 14812 58434 14868 58436
rect 14812 58382 14814 58434
rect 14814 58382 14866 58434
rect 14866 58382 14868 58434
rect 14812 58380 14868 58382
rect 15484 58434 15540 58436
rect 15484 58382 15486 58434
rect 15486 58382 15538 58434
rect 15538 58382 15540 58434
rect 15484 58380 15540 58382
rect 15260 58044 15316 58100
rect 14924 57820 14980 57876
rect 15148 56700 15204 56756
rect 14140 52556 14196 52612
rect 13916 50428 13972 50484
rect 14028 51436 14084 51492
rect 12796 49810 12852 49812
rect 12796 49758 12798 49810
rect 12798 49758 12850 49810
rect 12850 49758 12852 49810
rect 12796 49756 12852 49758
rect 12012 48748 12068 48804
rect 13580 49644 13636 49700
rect 12572 49196 12628 49252
rect 12796 48802 12852 48804
rect 12796 48750 12798 48802
rect 12798 48750 12850 48802
rect 12850 48750 12852 48802
rect 12796 48748 12852 48750
rect 12460 48130 12516 48132
rect 12460 48078 12462 48130
rect 12462 48078 12514 48130
rect 12514 48078 12516 48130
rect 12460 48076 12516 48078
rect 12908 48188 12964 48244
rect 13692 48914 13748 48916
rect 13692 48862 13694 48914
rect 13694 48862 13746 48914
rect 13746 48862 13748 48914
rect 13692 48860 13748 48862
rect 11228 46956 11284 47012
rect 11676 47234 11732 47236
rect 11676 47182 11678 47234
rect 11678 47182 11730 47234
rect 11730 47182 11732 47234
rect 11676 47180 11732 47182
rect 12236 47180 12292 47236
rect 12124 46732 12180 46788
rect 11564 46396 11620 46452
rect 11340 45948 11396 46004
rect 11116 45890 11172 45892
rect 11116 45838 11118 45890
rect 11118 45838 11170 45890
rect 11170 45838 11172 45890
rect 11116 45836 11172 45838
rect 11228 45778 11284 45780
rect 11228 45726 11230 45778
rect 11230 45726 11282 45778
rect 11282 45726 11284 45778
rect 11228 45724 11284 45726
rect 11116 44492 11172 44548
rect 11340 43708 11396 43764
rect 11004 42476 11060 42532
rect 11900 44434 11956 44436
rect 11900 44382 11902 44434
rect 11902 44382 11954 44434
rect 11954 44382 11956 44434
rect 11900 44380 11956 44382
rect 11900 44156 11956 44212
rect 11452 43596 11508 43652
rect 11676 43538 11732 43540
rect 11676 43486 11678 43538
rect 11678 43486 11730 43538
rect 11730 43486 11732 43538
rect 11676 43484 11732 43486
rect 11900 43372 11956 43428
rect 12124 44044 12180 44100
rect 13916 49026 13972 49028
rect 13916 48974 13918 49026
rect 13918 48974 13970 49026
rect 13970 48974 13972 49026
rect 13916 48972 13972 48974
rect 14700 52780 14756 52836
rect 14588 52668 14644 52724
rect 14588 52162 14644 52164
rect 14588 52110 14590 52162
rect 14590 52110 14642 52162
rect 14642 52110 14644 52162
rect 14588 52108 14644 52110
rect 14588 50706 14644 50708
rect 14588 50654 14590 50706
rect 14590 50654 14642 50706
rect 14642 50654 14644 50706
rect 14588 50652 14644 50654
rect 15596 56588 15652 56644
rect 15932 56252 15988 56308
rect 16492 58322 16548 58324
rect 16492 58270 16494 58322
rect 16494 58270 16546 58322
rect 16546 58270 16548 58322
rect 16492 58268 16548 58270
rect 16828 60620 16884 60676
rect 17388 60562 17444 60564
rect 17388 60510 17390 60562
rect 17390 60510 17442 60562
rect 17442 60510 17444 60562
rect 17388 60508 17444 60510
rect 16828 59836 16884 59892
rect 16828 59106 16884 59108
rect 16828 59054 16830 59106
rect 16830 59054 16882 59106
rect 16882 59054 16884 59106
rect 16828 59052 16884 59054
rect 16044 58044 16100 58100
rect 15148 56140 15204 56196
rect 15260 55356 15316 55412
rect 15148 54626 15204 54628
rect 15148 54574 15150 54626
rect 15150 54574 15202 54626
rect 15202 54574 15204 54626
rect 15148 54572 15204 54574
rect 18284 61292 18340 61348
rect 17948 60786 18004 60788
rect 17948 60734 17950 60786
rect 17950 60734 18002 60786
rect 18002 60734 18004 60786
rect 17948 60732 18004 60734
rect 17836 60620 17892 60676
rect 17164 59052 17220 59108
rect 17276 58210 17332 58212
rect 17276 58158 17278 58210
rect 17278 58158 17330 58210
rect 17330 58158 17332 58210
rect 17276 58156 17332 58158
rect 17612 58434 17668 58436
rect 17612 58382 17614 58434
rect 17614 58382 17666 58434
rect 17666 58382 17668 58434
rect 17612 58380 17668 58382
rect 17500 58322 17556 58324
rect 17500 58270 17502 58322
rect 17502 58270 17554 58322
rect 17554 58270 17556 58322
rect 17500 58268 17556 58270
rect 20188 62914 20244 62916
rect 20188 62862 20190 62914
rect 20190 62862 20242 62914
rect 20242 62862 20244 62914
rect 20188 62860 20244 62862
rect 19836 62746 19892 62748
rect 19836 62694 19838 62746
rect 19838 62694 19890 62746
rect 19890 62694 19892 62746
rect 19836 62692 19892 62694
rect 19940 62746 19996 62748
rect 19940 62694 19942 62746
rect 19942 62694 19994 62746
rect 19994 62694 19996 62746
rect 19940 62692 19996 62694
rect 20044 62746 20100 62748
rect 20044 62694 20046 62746
rect 20046 62694 20098 62746
rect 20098 62694 20100 62746
rect 20044 62692 20100 62694
rect 18844 61292 18900 61348
rect 18956 61180 19012 61236
rect 19836 61178 19892 61180
rect 19836 61126 19838 61178
rect 19838 61126 19890 61178
rect 19890 61126 19892 61178
rect 19836 61124 19892 61126
rect 19940 61178 19996 61180
rect 19940 61126 19942 61178
rect 19942 61126 19994 61178
rect 19994 61126 19996 61178
rect 19940 61124 19996 61126
rect 20044 61178 20100 61180
rect 20044 61126 20046 61178
rect 20046 61126 20098 61178
rect 20098 61126 20100 61178
rect 20044 61124 20100 61126
rect 19740 60956 19796 61012
rect 19516 60786 19572 60788
rect 19516 60734 19518 60786
rect 19518 60734 19570 60786
rect 19570 60734 19572 60786
rect 19516 60732 19572 60734
rect 19404 60620 19460 60676
rect 19180 59836 19236 59892
rect 18732 58828 18788 58884
rect 17836 58210 17892 58212
rect 17836 58158 17838 58210
rect 17838 58158 17890 58210
rect 17890 58158 17892 58210
rect 17836 58156 17892 58158
rect 16940 57596 16996 57652
rect 16268 54124 16324 54180
rect 16380 53788 16436 53844
rect 16716 56194 16772 56196
rect 16716 56142 16718 56194
rect 16718 56142 16770 56194
rect 16770 56142 16772 56194
rect 16716 56140 16772 56142
rect 16492 54626 16548 54628
rect 16492 54574 16494 54626
rect 16494 54574 16546 54626
rect 16546 54574 16548 54626
rect 16492 54572 16548 54574
rect 16156 53452 16212 53508
rect 15372 52556 15428 52612
rect 15484 52668 15540 52724
rect 14700 50316 14756 50372
rect 14252 49980 14308 50036
rect 14700 49026 14756 49028
rect 14700 48974 14702 49026
rect 14702 48974 14754 49026
rect 14754 48974 14756 49026
rect 14700 48972 14756 48974
rect 14476 47682 14532 47684
rect 14476 47630 14478 47682
rect 14478 47630 14530 47682
rect 14530 47630 14532 47682
rect 14476 47628 14532 47630
rect 15596 52780 15652 52836
rect 15596 49980 15652 50036
rect 16604 54124 16660 54180
rect 16604 53506 16660 53508
rect 16604 53454 16606 53506
rect 16606 53454 16658 53506
rect 16658 53454 16660 53506
rect 16604 53452 16660 53454
rect 18620 57932 18676 57988
rect 18508 57090 18564 57092
rect 18508 57038 18510 57090
rect 18510 57038 18562 57090
rect 18562 57038 18564 57090
rect 18508 57036 18564 57038
rect 17388 56306 17444 56308
rect 17388 56254 17390 56306
rect 17390 56254 17442 56306
rect 17442 56254 17444 56306
rect 17388 56252 17444 56254
rect 18396 56754 18452 56756
rect 18396 56702 18398 56754
rect 18398 56702 18450 56754
rect 18450 56702 18452 56754
rect 18396 56700 18452 56702
rect 16716 52946 16772 52948
rect 16716 52894 16718 52946
rect 16718 52894 16770 52946
rect 16770 52894 16772 52946
rect 16716 52892 16772 52894
rect 16604 52556 16660 52612
rect 16604 52108 16660 52164
rect 16492 51436 16548 51492
rect 15708 50652 15764 50708
rect 15484 49756 15540 49812
rect 15820 50428 15876 50484
rect 16828 51490 16884 51492
rect 16828 51438 16830 51490
rect 16830 51438 16882 51490
rect 16882 51438 16884 51490
rect 16828 51436 16884 51438
rect 18396 55468 18452 55524
rect 16940 50428 16996 50484
rect 17052 51996 17108 52052
rect 16604 50316 16660 50372
rect 16268 50034 16324 50036
rect 16268 49982 16270 50034
rect 16270 49982 16322 50034
rect 16322 49982 16324 50034
rect 16268 49980 16324 49982
rect 17164 50540 17220 50596
rect 17388 55074 17444 55076
rect 17388 55022 17390 55074
rect 17390 55022 17442 55074
rect 17442 55022 17444 55074
rect 17388 55020 17444 55022
rect 18956 56364 19012 56420
rect 19180 58828 19236 58884
rect 19180 58156 19236 58212
rect 19068 56924 19124 56980
rect 19628 60002 19684 60004
rect 19628 59950 19630 60002
rect 19630 59950 19682 60002
rect 19682 59950 19684 60002
rect 19628 59948 19684 59950
rect 19964 60732 20020 60788
rect 20300 60786 20356 60788
rect 20300 60734 20302 60786
rect 20302 60734 20354 60786
rect 20354 60734 20356 60786
rect 20300 60732 20356 60734
rect 20860 61010 20916 61012
rect 20860 60958 20862 61010
rect 20862 60958 20914 61010
rect 20914 60958 20916 61010
rect 20860 60956 20916 60958
rect 21308 63084 21364 63140
rect 21308 62860 21364 62916
rect 21308 61570 21364 61572
rect 21308 61518 21310 61570
rect 21310 61518 21362 61570
rect 21362 61518 21364 61570
rect 21308 61516 21364 61518
rect 21868 66332 21924 66388
rect 22876 67340 22932 67396
rect 22428 66780 22484 66836
rect 21756 65324 21812 65380
rect 22876 66780 22932 66836
rect 21644 63026 21700 63028
rect 21644 62974 21646 63026
rect 21646 62974 21698 63026
rect 21698 62974 21700 63026
rect 21644 62972 21700 62974
rect 23100 67340 23156 67396
rect 23324 67116 23380 67172
rect 23436 68012 23492 68068
rect 23772 67618 23828 67620
rect 23772 67566 23774 67618
rect 23774 67566 23826 67618
rect 23826 67566 23828 67618
rect 23772 67564 23828 67566
rect 24668 67788 24724 67844
rect 24892 67730 24948 67732
rect 24892 67678 24894 67730
rect 24894 67678 24946 67730
rect 24946 67678 24948 67730
rect 24892 67676 24948 67678
rect 24332 67564 24388 67620
rect 23996 67452 24052 67508
rect 24444 67452 24500 67508
rect 23548 67340 23604 67396
rect 24668 67340 24724 67396
rect 23100 67058 23156 67060
rect 23100 67006 23102 67058
rect 23102 67006 23154 67058
rect 23154 67006 23156 67058
rect 23100 67004 23156 67006
rect 23100 65436 23156 65492
rect 22876 65212 22932 65268
rect 22204 63308 22260 63364
rect 22428 63420 22484 63476
rect 22092 62748 22148 62804
rect 20636 60396 20692 60452
rect 19852 59724 19908 59780
rect 19836 59610 19892 59612
rect 19836 59558 19838 59610
rect 19838 59558 19890 59610
rect 19890 59558 19892 59610
rect 19836 59556 19892 59558
rect 19940 59610 19996 59612
rect 19940 59558 19942 59610
rect 19942 59558 19994 59610
rect 19994 59558 19996 59610
rect 19940 59556 19996 59558
rect 20044 59610 20100 59612
rect 20044 59558 20046 59610
rect 20046 59558 20098 59610
rect 20098 59558 20100 59610
rect 20044 59556 20100 59558
rect 20524 60002 20580 60004
rect 20524 59950 20526 60002
rect 20526 59950 20578 60002
rect 20578 59950 20580 60002
rect 20524 59948 20580 59950
rect 20748 59890 20804 59892
rect 20748 59838 20750 59890
rect 20750 59838 20802 59890
rect 20802 59838 20804 59890
rect 20748 59836 20804 59838
rect 19740 59330 19796 59332
rect 19740 59278 19742 59330
rect 19742 59278 19794 59330
rect 19794 59278 19796 59330
rect 19740 59276 19796 59278
rect 20076 59164 20132 59220
rect 20748 59218 20804 59220
rect 20748 59166 20750 59218
rect 20750 59166 20802 59218
rect 20802 59166 20804 59218
rect 20748 59164 20804 59166
rect 19852 58434 19908 58436
rect 19852 58382 19854 58434
rect 19854 58382 19906 58434
rect 19906 58382 19908 58434
rect 19852 58380 19908 58382
rect 19404 57932 19460 57988
rect 20300 58210 20356 58212
rect 20300 58158 20302 58210
rect 20302 58158 20354 58210
rect 20354 58158 20356 58210
rect 20300 58156 20356 58158
rect 19836 58042 19892 58044
rect 19836 57990 19838 58042
rect 19838 57990 19890 58042
rect 19890 57990 19892 58042
rect 19836 57988 19892 57990
rect 19940 58042 19996 58044
rect 19940 57990 19942 58042
rect 19942 57990 19994 58042
rect 19994 57990 19996 58042
rect 19940 57988 19996 57990
rect 20044 58042 20100 58044
rect 20044 57990 20046 58042
rect 20046 57990 20098 58042
rect 20098 57990 20100 58042
rect 20188 58044 20244 58100
rect 20044 57988 20100 57990
rect 20636 58380 20692 58436
rect 20748 58322 20804 58324
rect 20748 58270 20750 58322
rect 20750 58270 20802 58322
rect 20802 58270 20804 58322
rect 20748 58268 20804 58270
rect 19628 57036 19684 57092
rect 20300 57090 20356 57092
rect 20300 57038 20302 57090
rect 20302 57038 20354 57090
rect 20354 57038 20356 57090
rect 20300 57036 20356 57038
rect 21084 57762 21140 57764
rect 21084 57710 21086 57762
rect 21086 57710 21138 57762
rect 21138 57710 21140 57762
rect 21084 57708 21140 57710
rect 21532 60396 21588 60452
rect 21532 60060 21588 60116
rect 21420 59836 21476 59892
rect 22316 62914 22372 62916
rect 22316 62862 22318 62914
rect 22318 62862 22370 62914
rect 22370 62862 22372 62914
rect 22316 62860 22372 62862
rect 22428 61516 22484 61572
rect 22204 61404 22260 61460
rect 21756 61010 21812 61012
rect 21756 60958 21758 61010
rect 21758 60958 21810 61010
rect 21810 60958 21812 61010
rect 21756 60956 21812 60958
rect 21644 59948 21700 60004
rect 22652 63756 22708 63812
rect 22764 63420 22820 63476
rect 23212 65324 23268 65380
rect 22988 64146 23044 64148
rect 22988 64094 22990 64146
rect 22990 64094 23042 64146
rect 23042 64094 23044 64146
rect 22988 64092 23044 64094
rect 22876 63308 22932 63364
rect 22764 62748 22820 62804
rect 22092 60786 22148 60788
rect 22092 60734 22094 60786
rect 22094 60734 22146 60786
rect 22146 60734 22148 60786
rect 22092 60732 22148 60734
rect 22652 60898 22708 60900
rect 22652 60846 22654 60898
rect 22654 60846 22706 60898
rect 22706 60846 22708 60898
rect 22652 60844 22708 60846
rect 22204 60060 22260 60116
rect 23100 63026 23156 63028
rect 23100 62974 23102 63026
rect 23102 62974 23154 63026
rect 23154 62974 23156 63026
rect 23100 62972 23156 62974
rect 23100 62300 23156 62356
rect 23436 65212 23492 65268
rect 23324 63698 23380 63700
rect 23324 63646 23326 63698
rect 23326 63646 23378 63698
rect 23378 63646 23380 63698
rect 23324 63644 23380 63646
rect 23548 64428 23604 64484
rect 23548 63138 23604 63140
rect 23548 63086 23550 63138
rect 23550 63086 23602 63138
rect 23602 63086 23604 63138
rect 23548 63084 23604 63086
rect 23996 67170 24052 67172
rect 23996 67118 23998 67170
rect 23998 67118 24050 67170
rect 24050 67118 24052 67170
rect 23996 67116 24052 67118
rect 24220 66892 24276 66948
rect 24332 66780 24388 66836
rect 27804 69356 27860 69412
rect 26124 67842 26180 67844
rect 26124 67790 26126 67842
rect 26126 67790 26178 67842
rect 26178 67790 26180 67842
rect 26124 67788 26180 67790
rect 28028 67842 28084 67844
rect 28028 67790 28030 67842
rect 28030 67790 28082 67842
rect 28082 67790 28084 67842
rect 28028 67788 28084 67790
rect 26348 67676 26404 67732
rect 25564 67618 25620 67620
rect 25564 67566 25566 67618
rect 25566 67566 25618 67618
rect 25618 67566 25620 67618
rect 25564 67564 25620 67566
rect 25788 67618 25844 67620
rect 25788 67566 25790 67618
rect 25790 67566 25842 67618
rect 25842 67566 25844 67618
rect 25788 67564 25844 67566
rect 29708 70028 29764 70084
rect 29036 69298 29092 69300
rect 29036 69246 29038 69298
rect 29038 69246 29090 69298
rect 29090 69246 29092 69298
rect 29036 69244 29092 69246
rect 29260 69186 29316 69188
rect 29260 69134 29262 69186
rect 29262 69134 29314 69186
rect 29314 69134 29316 69186
rect 29260 69132 29316 69134
rect 29708 68908 29764 68964
rect 29372 68796 29428 68852
rect 29932 69020 29988 69076
rect 30044 68796 30100 68852
rect 28364 67564 28420 67620
rect 26236 67228 26292 67284
rect 28364 67116 28420 67172
rect 24444 65660 24500 65716
rect 24780 66050 24836 66052
rect 24780 65998 24782 66050
rect 24782 65998 24834 66050
rect 24834 65998 24836 66050
rect 24780 65996 24836 65998
rect 25452 66162 25508 66164
rect 25452 66110 25454 66162
rect 25454 66110 25506 66162
rect 25506 66110 25508 66162
rect 25452 66108 25508 66110
rect 24556 64204 24612 64260
rect 25228 65772 25284 65828
rect 25564 65996 25620 66052
rect 25676 65772 25732 65828
rect 25004 65660 25060 65716
rect 24444 64092 24500 64148
rect 23660 62524 23716 62580
rect 22764 60732 22820 60788
rect 21532 59500 21588 59556
rect 22652 59778 22708 59780
rect 22652 59726 22654 59778
rect 22654 59726 22706 59778
rect 22706 59726 22708 59778
rect 22652 59724 22708 59726
rect 20636 57036 20692 57092
rect 21532 58546 21588 58548
rect 21532 58494 21534 58546
rect 21534 58494 21586 58546
rect 21586 58494 21588 58546
rect 21532 58492 21588 58494
rect 21420 58044 21476 58100
rect 19516 56812 19572 56868
rect 19404 56754 19460 56756
rect 19404 56702 19406 56754
rect 19406 56702 19458 56754
rect 19458 56702 19460 56754
rect 19404 56700 19460 56702
rect 18956 55804 19012 55860
rect 18396 55074 18452 55076
rect 18396 55022 18398 55074
rect 18398 55022 18450 55074
rect 18450 55022 18452 55074
rect 18396 55020 18452 55022
rect 18620 55244 18676 55300
rect 17500 54124 17556 54180
rect 17948 53730 18004 53732
rect 17948 53678 17950 53730
rect 17950 53678 18002 53730
rect 18002 53678 18004 53730
rect 17948 53676 18004 53678
rect 18060 53116 18116 53172
rect 17500 52108 17556 52164
rect 17948 51772 18004 51828
rect 18172 52834 18228 52836
rect 18172 52782 18174 52834
rect 18174 52782 18226 52834
rect 18226 52782 18228 52834
rect 18172 52780 18228 52782
rect 18732 52108 18788 52164
rect 18172 51996 18228 52052
rect 17388 51436 17444 51492
rect 17276 50092 17332 50148
rect 17500 50764 17556 50820
rect 18620 51938 18676 51940
rect 18620 51886 18622 51938
rect 18622 51886 18674 51938
rect 18674 51886 18676 51938
rect 18620 51884 18676 51886
rect 18844 51772 18900 51828
rect 18844 51436 18900 51492
rect 18396 50764 18452 50820
rect 18060 50540 18116 50596
rect 19180 52892 19236 52948
rect 19068 51548 19124 51604
rect 19836 56474 19892 56476
rect 19836 56422 19838 56474
rect 19838 56422 19890 56474
rect 19890 56422 19892 56474
rect 19836 56420 19892 56422
rect 19940 56474 19996 56476
rect 19940 56422 19942 56474
rect 19942 56422 19994 56474
rect 19994 56422 19996 56474
rect 19940 56420 19996 56422
rect 20044 56474 20100 56476
rect 20044 56422 20046 56474
rect 20046 56422 20098 56474
rect 20098 56422 20100 56474
rect 20044 56420 20100 56422
rect 20300 55244 20356 55300
rect 19852 55132 19908 55188
rect 19404 55020 19460 55076
rect 19404 51884 19460 51940
rect 16492 49810 16548 49812
rect 16492 49758 16494 49810
rect 16494 49758 16546 49810
rect 16546 49758 16548 49810
rect 16492 49756 16548 49758
rect 15260 48972 15316 49028
rect 14924 46172 14980 46228
rect 15036 48748 15092 48804
rect 12796 45724 12852 45780
rect 12684 45052 12740 45108
rect 12572 44940 12628 44996
rect 12460 44828 12516 44884
rect 12684 44828 12740 44884
rect 12460 44044 12516 44100
rect 12348 43932 12404 43988
rect 12236 43708 12292 43764
rect 13020 44940 13076 44996
rect 12796 44156 12852 44212
rect 12796 43932 12852 43988
rect 12796 43708 12852 43764
rect 12348 43650 12404 43652
rect 12348 43598 12350 43650
rect 12350 43598 12402 43650
rect 12402 43598 12404 43650
rect 12348 43596 12404 43598
rect 12236 43538 12292 43540
rect 12236 43486 12238 43538
rect 12238 43486 12290 43538
rect 12290 43486 12292 43538
rect 12236 43484 12292 43486
rect 12124 43260 12180 43316
rect 12012 42588 12068 42644
rect 13244 44882 13300 44884
rect 13244 44830 13246 44882
rect 13246 44830 13298 44882
rect 13298 44830 13300 44882
rect 13244 44828 13300 44830
rect 13244 44156 13300 44212
rect 12908 43372 12964 43428
rect 13020 43314 13076 43316
rect 13020 43262 13022 43314
rect 13022 43262 13074 43314
rect 13074 43262 13076 43314
rect 13020 43260 13076 43262
rect 13580 44994 13636 44996
rect 13580 44942 13582 44994
rect 13582 44942 13634 44994
rect 13634 44942 13636 44994
rect 13580 44940 13636 44942
rect 13692 43708 13748 43764
rect 14476 45778 14532 45780
rect 14476 45726 14478 45778
rect 14478 45726 14530 45778
rect 14530 45726 14532 45778
rect 14476 45724 14532 45726
rect 14364 45052 14420 45108
rect 14476 44940 14532 44996
rect 14028 43260 14084 43316
rect 13916 42642 13972 42644
rect 13916 42590 13918 42642
rect 13918 42590 13970 42642
rect 13970 42590 13972 42642
rect 13916 42588 13972 42590
rect 10892 41692 10948 41748
rect 10780 41410 10836 41412
rect 10780 41358 10782 41410
rect 10782 41358 10834 41410
rect 10834 41358 10836 41410
rect 10780 41356 10836 41358
rect 11564 41074 11620 41076
rect 11564 41022 11566 41074
rect 11566 41022 11618 41074
rect 11618 41022 11620 41074
rect 11564 41020 11620 41022
rect 12236 41074 12292 41076
rect 12236 41022 12238 41074
rect 12238 41022 12290 41074
rect 12290 41022 12292 41074
rect 12236 41020 12292 41022
rect 12684 41020 12740 41076
rect 11228 39900 11284 39956
rect 11004 39618 11060 39620
rect 11004 39566 11006 39618
rect 11006 39566 11058 39618
rect 11058 39566 11060 39618
rect 11004 39564 11060 39566
rect 10556 39452 10612 39508
rect 10668 38722 10724 38724
rect 10668 38670 10670 38722
rect 10670 38670 10722 38722
rect 10722 38670 10724 38722
rect 10668 38668 10724 38670
rect 10780 38220 10836 38276
rect 11228 37996 11284 38052
rect 11900 39340 11956 39396
rect 11676 38108 11732 38164
rect 10220 37042 10276 37044
rect 10220 36990 10222 37042
rect 10222 36990 10274 37042
rect 10274 36990 10276 37042
rect 10220 36988 10276 36990
rect 10108 35474 10164 35476
rect 10108 35422 10110 35474
rect 10110 35422 10162 35474
rect 10162 35422 10164 35474
rect 10108 35420 10164 35422
rect 11788 37996 11844 38052
rect 11788 37378 11844 37380
rect 11788 37326 11790 37378
rect 11790 37326 11842 37378
rect 11842 37326 11844 37378
rect 11788 37324 11844 37326
rect 11900 37212 11956 37268
rect 11004 35756 11060 35812
rect 10332 35420 10388 35476
rect 10220 33852 10276 33908
rect 10780 35698 10836 35700
rect 10780 35646 10782 35698
rect 10782 35646 10834 35698
rect 10834 35646 10836 35698
rect 10780 35644 10836 35646
rect 9996 32284 10052 32340
rect 9548 31164 9604 31220
rect 8988 30716 9044 30772
rect 10108 31500 10164 31556
rect 11116 35474 11172 35476
rect 11116 35422 11118 35474
rect 11118 35422 11170 35474
rect 11170 35422 11172 35474
rect 11116 35420 11172 35422
rect 11340 35420 11396 35476
rect 11228 35026 11284 35028
rect 11228 34974 11230 35026
rect 11230 34974 11282 35026
rect 11282 34974 11284 35026
rect 11228 34972 11284 34974
rect 12684 40572 12740 40628
rect 13916 39788 13972 39844
rect 12908 39676 12964 39732
rect 13580 39730 13636 39732
rect 13580 39678 13582 39730
rect 13582 39678 13634 39730
rect 13634 39678 13636 39730
rect 13580 39676 13636 39678
rect 12684 38668 12740 38724
rect 13468 39394 13524 39396
rect 13468 39342 13470 39394
rect 13470 39342 13522 39394
rect 13522 39342 13524 39394
rect 13468 39340 13524 39342
rect 14028 39394 14084 39396
rect 14028 39342 14030 39394
rect 14030 39342 14082 39394
rect 14082 39342 14084 39394
rect 14028 39340 14084 39342
rect 13468 38274 13524 38276
rect 13468 38222 13470 38274
rect 13470 38222 13522 38274
rect 13522 38222 13524 38274
rect 13468 38220 13524 38222
rect 14028 38722 14084 38724
rect 14028 38670 14030 38722
rect 14030 38670 14082 38722
rect 14082 38670 14084 38722
rect 14028 38668 14084 38670
rect 14364 38668 14420 38724
rect 14252 38556 14308 38612
rect 12236 37212 12292 37268
rect 12012 34860 12068 34916
rect 13468 37324 13524 37380
rect 13692 37212 13748 37268
rect 16492 48972 16548 49028
rect 16940 49420 16996 49476
rect 16828 48354 16884 48356
rect 16828 48302 16830 48354
rect 16830 48302 16882 48354
rect 16882 48302 16884 48354
rect 16828 48300 16884 48302
rect 15708 48130 15764 48132
rect 15708 48078 15710 48130
rect 15710 48078 15762 48130
rect 15762 48078 15764 48130
rect 15708 48076 15764 48078
rect 15820 47628 15876 47684
rect 16044 47346 16100 47348
rect 16044 47294 16046 47346
rect 16046 47294 16098 47346
rect 16098 47294 16100 47346
rect 16044 47292 16100 47294
rect 16268 47570 16324 47572
rect 16268 47518 16270 47570
rect 16270 47518 16322 47570
rect 16322 47518 16324 47570
rect 16268 47516 16324 47518
rect 16268 47180 16324 47236
rect 17836 49586 17892 49588
rect 17836 49534 17838 49586
rect 17838 49534 17890 49586
rect 17890 49534 17892 49586
rect 17836 49532 17892 49534
rect 18284 49026 18340 49028
rect 18284 48974 18286 49026
rect 18286 48974 18338 49026
rect 18338 48974 18340 49026
rect 18284 48972 18340 48974
rect 17724 48860 17780 48916
rect 17388 48354 17444 48356
rect 17388 48302 17390 48354
rect 17390 48302 17442 48354
rect 17442 48302 17444 48354
rect 17388 48300 17444 48302
rect 17388 47180 17444 47236
rect 16604 45276 16660 45332
rect 15932 43708 15988 43764
rect 15708 41020 15764 41076
rect 15036 39900 15092 39956
rect 15260 39564 15316 39620
rect 16940 43932 16996 43988
rect 16828 43484 16884 43540
rect 16604 43260 16660 43316
rect 16828 40684 16884 40740
rect 17164 46002 17220 46004
rect 17164 45950 17166 46002
rect 17166 45950 17218 46002
rect 17218 45950 17220 46002
rect 17164 45948 17220 45950
rect 17052 40236 17108 40292
rect 16268 40012 16324 40068
rect 15036 39116 15092 39172
rect 14588 39058 14644 39060
rect 14588 39006 14590 39058
rect 14590 39006 14642 39058
rect 14642 39006 14644 39058
rect 14588 39004 14644 39006
rect 15260 39058 15316 39060
rect 15260 39006 15262 39058
rect 15262 39006 15314 39058
rect 15314 39006 15316 39058
rect 15260 39004 15316 39006
rect 14476 38332 14532 38388
rect 14588 38108 14644 38164
rect 14364 37436 14420 37492
rect 15596 38610 15652 38612
rect 15596 38558 15598 38610
rect 15598 38558 15650 38610
rect 15650 38558 15652 38610
rect 15596 38556 15652 38558
rect 15708 38220 15764 38276
rect 15708 38050 15764 38052
rect 15708 37998 15710 38050
rect 15710 37998 15762 38050
rect 15762 37998 15764 38050
rect 15708 37996 15764 37998
rect 15484 37884 15540 37940
rect 15372 37436 15428 37492
rect 16828 39730 16884 39732
rect 16828 39678 16830 39730
rect 16830 39678 16882 39730
rect 16882 39678 16884 39730
rect 16828 39676 16884 39678
rect 15820 37436 15876 37492
rect 17052 39340 17108 39396
rect 15932 39116 15988 39172
rect 15372 36092 15428 36148
rect 12348 35420 12404 35476
rect 12124 34690 12180 34692
rect 12124 34638 12126 34690
rect 12126 34638 12178 34690
rect 12178 34638 12180 34690
rect 12124 34636 12180 34638
rect 11788 34130 11844 34132
rect 11788 34078 11790 34130
rect 11790 34078 11842 34130
rect 11842 34078 11844 34130
rect 11788 34076 11844 34078
rect 11116 33906 11172 33908
rect 11116 33854 11118 33906
rect 11118 33854 11170 33906
rect 11170 33854 11172 33906
rect 11116 33852 11172 33854
rect 11116 32508 11172 32564
rect 11788 33068 11844 33124
rect 12012 32338 12068 32340
rect 12012 32286 12014 32338
rect 12014 32286 12066 32338
rect 12066 32286 12068 32338
rect 12012 32284 12068 32286
rect 10556 30994 10612 30996
rect 10556 30942 10558 30994
rect 10558 30942 10610 30994
rect 10610 30942 10612 30994
rect 10556 30940 10612 30942
rect 10332 30770 10388 30772
rect 10332 30718 10334 30770
rect 10334 30718 10386 30770
rect 10386 30718 10388 30770
rect 10332 30716 10388 30718
rect 11340 32172 11396 32228
rect 10780 30716 10836 30772
rect 9996 30604 10052 30660
rect 1708 29596 1764 29652
rect 2940 29596 2996 29652
rect 2044 29538 2100 29540
rect 2044 29486 2046 29538
rect 2046 29486 2098 29538
rect 2098 29486 2100 29538
rect 2044 29484 2100 29486
rect 1708 28924 1764 28980
rect 2492 28924 2548 28980
rect 4476 29034 4532 29036
rect 4476 28982 4478 29034
rect 4478 28982 4530 29034
rect 4530 28982 4532 29034
rect 4476 28980 4532 28982
rect 4580 29034 4636 29036
rect 4580 28982 4582 29034
rect 4582 28982 4634 29034
rect 4634 28982 4636 29034
rect 4580 28980 4636 28982
rect 4684 29034 4740 29036
rect 4684 28982 4686 29034
rect 4686 28982 4738 29034
rect 4738 28982 4740 29034
rect 4684 28980 4740 28982
rect 2044 28588 2100 28644
rect 1708 28252 1764 28308
rect 2492 28252 2548 28308
rect 8316 28588 8372 28644
rect 2044 27970 2100 27972
rect 2044 27918 2046 27970
rect 2046 27918 2098 27970
rect 2098 27918 2100 27970
rect 2044 27916 2100 27918
rect 1708 27580 1764 27636
rect 2492 27580 2548 27636
rect 2716 27580 2772 27636
rect 1708 26962 1764 26964
rect 1708 26910 1710 26962
rect 1710 26910 1762 26962
rect 1762 26910 1764 26962
rect 1708 26908 1764 26910
rect 2044 26850 2100 26852
rect 2044 26798 2046 26850
rect 2046 26798 2098 26850
rect 2098 26798 2100 26850
rect 2044 26796 2100 26798
rect 2380 26796 2436 26852
rect 2156 26684 2212 26740
rect 2492 26908 2548 26964
rect 4476 27466 4532 27468
rect 4476 27414 4478 27466
rect 4478 27414 4530 27466
rect 4530 27414 4532 27466
rect 4476 27412 4532 27414
rect 4580 27466 4636 27468
rect 4580 27414 4582 27466
rect 4582 27414 4634 27466
rect 4634 27414 4636 27466
rect 4580 27412 4636 27414
rect 4684 27466 4740 27468
rect 4684 27414 4686 27466
rect 4686 27414 4738 27466
rect 4738 27414 4740 27466
rect 4684 27412 4740 27414
rect 8316 27356 8372 27412
rect 10108 30044 10164 30100
rect 10556 29426 10612 29428
rect 10556 29374 10558 29426
rect 10558 29374 10610 29426
rect 10610 29374 10612 29426
rect 10556 29372 10612 29374
rect 10780 29260 10836 29316
rect 8988 29148 9044 29204
rect 10332 29202 10388 29204
rect 10332 29150 10334 29202
rect 10334 29150 10386 29202
rect 10386 29150 10388 29202
rect 10332 29148 10388 29150
rect 9996 28812 10052 28868
rect 3164 26796 3220 26852
rect 6524 26908 6580 26964
rect 2380 26236 2436 26292
rect 1708 26124 1764 26180
rect 2940 26178 2996 26180
rect 2940 26126 2942 26178
rect 2942 26126 2994 26178
rect 2994 26126 2996 26178
rect 2940 26124 2996 26126
rect 4476 25898 4532 25900
rect 4476 25846 4478 25898
rect 4478 25846 4530 25898
rect 4530 25846 4532 25898
rect 4476 25844 4532 25846
rect 4580 25898 4636 25900
rect 4580 25846 4582 25898
rect 4582 25846 4634 25898
rect 4634 25846 4636 25898
rect 4580 25844 4636 25846
rect 4684 25898 4740 25900
rect 4684 25846 4686 25898
rect 4686 25846 4738 25898
rect 4738 25846 4740 25898
rect 4684 25844 4740 25846
rect 1708 25564 1764 25620
rect 8428 26908 8484 26964
rect 8988 27916 9044 27972
rect 2044 25452 2100 25508
rect 1708 24892 1764 24948
rect 2492 24892 2548 24948
rect 1708 24220 1764 24276
rect 2044 23826 2100 23828
rect 2044 23774 2046 23826
rect 2046 23774 2098 23826
rect 2098 23774 2100 23826
rect 2044 23772 2100 23774
rect 1708 23548 1764 23604
rect 1708 22876 1764 22932
rect 8316 24780 8372 24836
rect 11676 31948 11732 32004
rect 13020 34972 13076 35028
rect 12908 34690 12964 34692
rect 12908 34638 12910 34690
rect 12910 34638 12962 34690
rect 12962 34638 12964 34690
rect 12908 34636 12964 34638
rect 15260 35308 15316 35364
rect 12460 32396 12516 32452
rect 12124 30940 12180 30996
rect 12348 31500 12404 31556
rect 11676 30716 11732 30772
rect 11228 29596 11284 29652
rect 11340 29372 11396 29428
rect 12236 29260 12292 29316
rect 11788 28588 11844 28644
rect 13580 34130 13636 34132
rect 13580 34078 13582 34130
rect 13582 34078 13634 34130
rect 13634 34078 13636 34130
rect 13580 34076 13636 34078
rect 13580 32562 13636 32564
rect 13580 32510 13582 32562
rect 13582 32510 13634 32562
rect 13634 32510 13636 32562
rect 13580 32508 13636 32510
rect 13468 32396 13524 32452
rect 14924 33852 14980 33908
rect 14700 33516 14756 33572
rect 15036 33404 15092 33460
rect 17052 39116 17108 39172
rect 16044 39058 16100 39060
rect 16044 39006 16046 39058
rect 16046 39006 16098 39058
rect 16098 39006 16100 39058
rect 16044 39004 16100 39006
rect 18060 48914 18116 48916
rect 18060 48862 18062 48914
rect 18062 48862 18114 48914
rect 18114 48862 18116 48914
rect 18060 48860 18116 48862
rect 18172 48636 18228 48692
rect 18844 48748 18900 48804
rect 18508 47852 18564 47908
rect 18620 48636 18676 48692
rect 17948 47516 18004 47572
rect 18060 47740 18116 47796
rect 17724 45388 17780 45444
rect 17612 44322 17668 44324
rect 17612 44270 17614 44322
rect 17614 44270 17666 44322
rect 17666 44270 17668 44322
rect 17612 44268 17668 44270
rect 19068 47852 19124 47908
rect 19292 51266 19348 51268
rect 19292 51214 19294 51266
rect 19294 51214 19346 51266
rect 19346 51214 19348 51266
rect 19292 51212 19348 51214
rect 19836 54906 19892 54908
rect 19836 54854 19838 54906
rect 19838 54854 19890 54906
rect 19890 54854 19892 54906
rect 19836 54852 19892 54854
rect 19940 54906 19996 54908
rect 19940 54854 19942 54906
rect 19942 54854 19994 54906
rect 19994 54854 19996 54906
rect 19940 54852 19996 54854
rect 20044 54906 20100 54908
rect 20044 54854 20046 54906
rect 20046 54854 20098 54906
rect 20098 54854 20100 54906
rect 20044 54852 20100 54854
rect 20300 55074 20356 55076
rect 20300 55022 20302 55074
rect 20302 55022 20354 55074
rect 20354 55022 20356 55074
rect 20300 55020 20356 55022
rect 20524 55356 20580 55412
rect 20748 56028 20804 56084
rect 20636 55244 20692 55300
rect 20524 55186 20580 55188
rect 20524 55134 20526 55186
rect 20526 55134 20578 55186
rect 20578 55134 20580 55186
rect 20524 55132 20580 55134
rect 20076 53452 20132 53508
rect 19836 53338 19892 53340
rect 19836 53286 19838 53338
rect 19838 53286 19890 53338
rect 19890 53286 19892 53338
rect 19836 53284 19892 53286
rect 19940 53338 19996 53340
rect 19940 53286 19942 53338
rect 19942 53286 19994 53338
rect 19994 53286 19996 53338
rect 19940 53284 19996 53286
rect 20044 53338 20100 53340
rect 20044 53286 20046 53338
rect 20046 53286 20098 53338
rect 20098 53286 20100 53338
rect 20044 53284 20100 53286
rect 20748 53004 20804 53060
rect 19964 52108 20020 52164
rect 20300 52332 20356 52388
rect 19836 51770 19892 51772
rect 19836 51718 19838 51770
rect 19838 51718 19890 51770
rect 19890 51718 19892 51770
rect 19836 51716 19892 51718
rect 19940 51770 19996 51772
rect 19940 51718 19942 51770
rect 19942 51718 19994 51770
rect 19994 51718 19996 51770
rect 19940 51716 19996 51718
rect 20044 51770 20100 51772
rect 20044 51718 20046 51770
rect 20046 51718 20098 51770
rect 20098 51718 20100 51770
rect 20044 51716 20100 51718
rect 19740 51602 19796 51604
rect 19740 51550 19742 51602
rect 19742 51550 19794 51602
rect 19794 51550 19796 51602
rect 19740 51548 19796 51550
rect 19964 51490 20020 51492
rect 19964 51438 19966 51490
rect 19966 51438 20018 51490
rect 20018 51438 20020 51490
rect 19964 51436 20020 51438
rect 20524 52780 20580 52836
rect 21532 58268 21588 58324
rect 21644 57036 21700 57092
rect 21756 59164 21812 59220
rect 21308 56866 21364 56868
rect 21308 56814 21310 56866
rect 21310 56814 21362 56866
rect 21362 56814 21364 56866
rect 21308 56812 21364 56814
rect 21644 56812 21700 56868
rect 21420 56754 21476 56756
rect 21420 56702 21422 56754
rect 21422 56702 21474 56754
rect 21474 56702 21476 56754
rect 21420 56700 21476 56702
rect 21980 58492 22036 58548
rect 21868 57148 21924 57204
rect 22428 59500 22484 59556
rect 21756 56700 21812 56756
rect 22988 61068 23044 61124
rect 23100 61010 23156 61012
rect 23100 60958 23102 61010
rect 23102 60958 23154 61010
rect 23154 60958 23156 61010
rect 23100 60956 23156 60958
rect 23212 60898 23268 60900
rect 23212 60846 23214 60898
rect 23214 60846 23266 60898
rect 23266 60846 23268 60898
rect 23212 60844 23268 60846
rect 23100 60732 23156 60788
rect 22988 59500 23044 59556
rect 22764 59218 22820 59220
rect 22764 59166 22766 59218
rect 22766 59166 22818 59218
rect 22818 59166 22820 59218
rect 22764 59164 22820 59166
rect 22988 59052 23044 59108
rect 22876 58828 22932 58884
rect 22428 57708 22484 57764
rect 22988 57372 23044 57428
rect 22428 57036 22484 57092
rect 22092 56866 22148 56868
rect 22092 56814 22094 56866
rect 22094 56814 22146 56866
rect 22146 56814 22148 56866
rect 22092 56812 22148 56814
rect 21980 55468 22036 55524
rect 21308 55356 21364 55412
rect 21308 53730 21364 53732
rect 21308 53678 21310 53730
rect 21310 53678 21362 53730
rect 21362 53678 21364 53730
rect 21308 53676 21364 53678
rect 20972 53058 21028 53060
rect 20972 53006 20974 53058
rect 20974 53006 21026 53058
rect 21026 53006 21028 53058
rect 20972 53004 21028 53006
rect 21196 52946 21252 52948
rect 21196 52894 21198 52946
rect 21198 52894 21250 52946
rect 21250 52894 21252 52946
rect 21196 52892 21252 52894
rect 20972 52668 21028 52724
rect 20748 52556 20804 52612
rect 21420 52274 21476 52276
rect 21420 52222 21422 52274
rect 21422 52222 21474 52274
rect 21474 52222 21476 52274
rect 21420 52220 21476 52222
rect 20524 51602 20580 51604
rect 20524 51550 20526 51602
rect 20526 51550 20578 51602
rect 20578 51550 20580 51602
rect 20524 51548 20580 51550
rect 21196 51490 21252 51492
rect 21196 51438 21198 51490
rect 21198 51438 21250 51490
rect 21250 51438 21252 51490
rect 21196 51436 21252 51438
rect 20300 51212 20356 51268
rect 20636 51100 20692 51156
rect 19516 50764 19572 50820
rect 18508 47404 18564 47460
rect 18284 45330 18340 45332
rect 18284 45278 18286 45330
rect 18286 45278 18338 45330
rect 18338 45278 18340 45330
rect 18284 45276 18340 45278
rect 18172 45218 18228 45220
rect 18172 45166 18174 45218
rect 18174 45166 18226 45218
rect 18226 45166 18228 45218
rect 18172 45164 18228 45166
rect 17836 44044 17892 44100
rect 17500 43932 17556 43988
rect 17724 43596 17780 43652
rect 18396 43596 18452 43652
rect 18172 43538 18228 43540
rect 18172 43486 18174 43538
rect 18174 43486 18226 43538
rect 18226 43486 18228 43538
rect 18172 43484 18228 43486
rect 19180 45612 19236 45668
rect 18956 45330 19012 45332
rect 18956 45278 18958 45330
rect 18958 45278 19010 45330
rect 19010 45278 19012 45330
rect 18956 45276 19012 45278
rect 19292 45276 19348 45332
rect 20636 50876 20692 50932
rect 20188 50652 20244 50708
rect 20076 50428 20132 50484
rect 19836 50202 19892 50204
rect 19836 50150 19838 50202
rect 19838 50150 19890 50202
rect 19890 50150 19892 50202
rect 19836 50148 19892 50150
rect 19940 50202 19996 50204
rect 19940 50150 19942 50202
rect 19942 50150 19994 50202
rect 19994 50150 19996 50202
rect 19940 50148 19996 50150
rect 20044 50202 20100 50204
rect 20044 50150 20046 50202
rect 20046 50150 20098 50202
rect 20098 50150 20100 50202
rect 20044 50148 20100 50150
rect 20076 49698 20132 49700
rect 20076 49646 20078 49698
rect 20078 49646 20130 49698
rect 20130 49646 20132 49698
rect 20076 49644 20132 49646
rect 20748 50594 20804 50596
rect 20748 50542 20750 50594
rect 20750 50542 20802 50594
rect 20802 50542 20804 50594
rect 20748 50540 20804 50542
rect 20412 49644 20468 49700
rect 20748 49308 20804 49364
rect 19836 48634 19892 48636
rect 19836 48582 19838 48634
rect 19838 48582 19890 48634
rect 19890 48582 19892 48634
rect 19836 48580 19892 48582
rect 19940 48634 19996 48636
rect 19940 48582 19942 48634
rect 19942 48582 19994 48634
rect 19994 48582 19996 48634
rect 19940 48580 19996 48582
rect 20044 48634 20100 48636
rect 20044 48582 20046 48634
rect 20046 48582 20098 48634
rect 20098 48582 20100 48634
rect 20044 48580 20100 48582
rect 21420 50988 21476 51044
rect 21420 50764 21476 50820
rect 22092 53842 22148 53844
rect 22092 53790 22094 53842
rect 22094 53790 22146 53842
rect 22146 53790 22148 53842
rect 22092 53788 22148 53790
rect 21868 53452 21924 53508
rect 22316 55244 22372 55300
rect 21868 52668 21924 52724
rect 21644 52108 21700 52164
rect 21868 51378 21924 51380
rect 21868 51326 21870 51378
rect 21870 51326 21922 51378
rect 21922 51326 21924 51378
rect 21868 51324 21924 51326
rect 22204 52892 22260 52948
rect 22876 56812 22932 56868
rect 22652 56754 22708 56756
rect 22652 56702 22654 56754
rect 22654 56702 22706 56754
rect 22706 56702 22708 56754
rect 22652 56700 22708 56702
rect 23324 58940 23380 58996
rect 23212 57932 23268 57988
rect 24332 63810 24388 63812
rect 24332 63758 24334 63810
rect 24334 63758 24386 63810
rect 24386 63758 24388 63810
rect 24332 63756 24388 63758
rect 23884 61068 23940 61124
rect 23772 60956 23828 61012
rect 24220 62860 24276 62916
rect 24332 63138 24388 63140
rect 24332 63086 24334 63138
rect 24334 63086 24386 63138
rect 24386 63086 24388 63138
rect 24332 63084 24388 63086
rect 23996 60844 24052 60900
rect 23884 60002 23940 60004
rect 23884 59950 23886 60002
rect 23886 59950 23938 60002
rect 23938 59950 23940 60002
rect 23884 59948 23940 59950
rect 23996 59724 24052 59780
rect 23996 59388 24052 59444
rect 23772 58716 23828 58772
rect 23772 57820 23828 57876
rect 23436 57596 23492 57652
rect 23100 56700 23156 56756
rect 22540 56082 22596 56084
rect 22540 56030 22542 56082
rect 22542 56030 22594 56082
rect 22594 56030 22596 56082
rect 22540 56028 22596 56030
rect 22092 51548 22148 51604
rect 22988 55244 23044 55300
rect 23660 57372 23716 57428
rect 23548 57260 23604 57316
rect 23884 57036 23940 57092
rect 24220 61740 24276 61796
rect 25788 65714 25844 65716
rect 25788 65662 25790 65714
rect 25790 65662 25842 65714
rect 25842 65662 25844 65714
rect 25788 65660 25844 65662
rect 25340 65548 25396 65604
rect 25228 65324 25284 65380
rect 25116 63644 25172 63700
rect 25564 63756 25620 63812
rect 25228 63308 25284 63364
rect 24780 62860 24836 62916
rect 25340 61740 25396 61796
rect 25340 60844 25396 60900
rect 25228 60508 25284 60564
rect 24332 59724 24388 59780
rect 24892 59948 24948 60004
rect 24556 59442 24612 59444
rect 24556 59390 24558 59442
rect 24558 59390 24610 59442
rect 24610 59390 24612 59442
rect 24556 59388 24612 59390
rect 24444 59164 24500 59220
rect 24108 57596 24164 57652
rect 24220 58716 24276 58772
rect 24556 58994 24612 58996
rect 24556 58942 24558 58994
rect 24558 58942 24610 58994
rect 24610 58942 24612 58994
rect 24556 58940 24612 58942
rect 24668 58716 24724 58772
rect 24668 58380 24724 58436
rect 24556 57874 24612 57876
rect 24556 57822 24558 57874
rect 24558 57822 24610 57874
rect 24610 57822 24612 57874
rect 24556 57820 24612 57822
rect 24668 57036 24724 57092
rect 23996 56476 24052 56532
rect 23548 56028 23604 56084
rect 24220 56866 24276 56868
rect 24220 56814 24222 56866
rect 24222 56814 24274 56866
rect 24274 56814 24276 56866
rect 24220 56812 24276 56814
rect 22988 53170 23044 53172
rect 22988 53118 22990 53170
rect 22990 53118 23042 53170
rect 23042 53118 23044 53170
rect 22988 53116 23044 53118
rect 23324 53676 23380 53732
rect 22764 52946 22820 52948
rect 22764 52894 22766 52946
rect 22766 52894 22818 52946
rect 22818 52894 22820 52946
rect 22764 52892 22820 52894
rect 22764 52220 22820 52276
rect 23212 52892 23268 52948
rect 22652 51548 22708 51604
rect 23100 52050 23156 52052
rect 23100 51998 23102 52050
rect 23102 51998 23154 52050
rect 23154 51998 23156 52050
rect 23100 51996 23156 51998
rect 24332 56754 24388 56756
rect 24332 56702 24334 56754
rect 24334 56702 24386 56754
rect 24386 56702 24388 56754
rect 24332 56700 24388 56702
rect 24444 56588 24500 56644
rect 24444 56306 24500 56308
rect 24444 56254 24446 56306
rect 24446 56254 24498 56306
rect 24498 56254 24500 56306
rect 24444 56252 24500 56254
rect 24220 54684 24276 54740
rect 25564 63308 25620 63364
rect 25900 65548 25956 65604
rect 26236 66274 26292 66276
rect 26236 66222 26238 66274
rect 26238 66222 26290 66274
rect 26290 66222 26292 66274
rect 26236 66220 26292 66222
rect 26124 66162 26180 66164
rect 26124 66110 26126 66162
rect 26126 66110 26178 66162
rect 26178 66110 26180 66162
rect 26124 66108 26180 66110
rect 26012 65324 26068 65380
rect 26124 65660 26180 65716
rect 26572 65490 26628 65492
rect 26572 65438 26574 65490
rect 26574 65438 26626 65490
rect 26626 65438 26628 65490
rect 26572 65436 26628 65438
rect 26012 63922 26068 63924
rect 26012 63870 26014 63922
rect 26014 63870 26066 63922
rect 26066 63870 26068 63922
rect 26012 63868 26068 63870
rect 25900 63756 25956 63812
rect 26460 64482 26516 64484
rect 26460 64430 26462 64482
rect 26462 64430 26514 64482
rect 26514 64430 26516 64482
rect 26460 64428 26516 64430
rect 26348 64316 26404 64372
rect 25676 61068 25732 61124
rect 25452 59500 25508 59556
rect 25788 59276 25844 59332
rect 24892 57484 24948 57540
rect 24892 57260 24948 57316
rect 25228 58828 25284 58884
rect 25340 57932 25396 57988
rect 25228 57650 25284 57652
rect 25228 57598 25230 57650
rect 25230 57598 25282 57650
rect 25282 57598 25284 57650
rect 25228 57596 25284 57598
rect 26460 64204 26516 64260
rect 27020 66444 27076 66500
rect 29708 67452 29764 67508
rect 29260 67282 29316 67284
rect 29260 67230 29262 67282
rect 29262 67230 29314 67282
rect 29314 67230 29316 67282
rect 29260 67228 29316 67230
rect 29148 67170 29204 67172
rect 29148 67118 29150 67170
rect 29150 67118 29202 67170
rect 29202 67118 29204 67170
rect 29148 67116 29204 67118
rect 28588 67004 28644 67060
rect 27804 66274 27860 66276
rect 27804 66222 27806 66274
rect 27806 66222 27858 66274
rect 27858 66222 27860 66274
rect 27804 66220 27860 66222
rect 26908 65996 26964 66052
rect 27244 66050 27300 66052
rect 27244 65998 27246 66050
rect 27246 65998 27298 66050
rect 27298 65998 27300 66050
rect 27244 65996 27300 65998
rect 27468 65436 27524 65492
rect 27468 64706 27524 64708
rect 27468 64654 27470 64706
rect 27470 64654 27522 64706
rect 27522 64654 27524 64706
rect 27468 64652 27524 64654
rect 27244 64316 27300 64372
rect 27356 64540 27412 64596
rect 27356 64204 27412 64260
rect 27020 64092 27076 64148
rect 27468 63868 27524 63924
rect 28252 66220 28308 66276
rect 27804 64540 27860 64596
rect 28140 63756 28196 63812
rect 26012 62914 26068 62916
rect 26012 62862 26014 62914
rect 26014 62862 26066 62914
rect 26066 62862 26068 62914
rect 26012 62860 26068 62862
rect 27132 62972 27188 63028
rect 26012 61964 26068 62020
rect 26572 62076 26628 62132
rect 28700 66220 28756 66276
rect 29484 67228 29540 67284
rect 29260 66220 29316 66276
rect 28364 65324 28420 65380
rect 29260 65996 29316 66052
rect 28588 64316 28644 64372
rect 28924 64204 28980 64260
rect 28588 64146 28644 64148
rect 28588 64094 28590 64146
rect 28590 64094 28642 64146
rect 28642 64094 28644 64146
rect 28588 64092 28644 64094
rect 26236 60508 26292 60564
rect 26348 61068 26404 61124
rect 26012 60284 26068 60340
rect 26236 60226 26292 60228
rect 26236 60174 26238 60226
rect 26238 60174 26290 60226
rect 26290 60174 26292 60226
rect 26236 60172 26292 60174
rect 26012 59836 26068 59892
rect 26236 59330 26292 59332
rect 26236 59278 26238 59330
rect 26238 59278 26290 59330
rect 26290 59278 26292 59330
rect 26236 59276 26292 59278
rect 26012 59164 26068 59220
rect 25676 57932 25732 57988
rect 25788 57820 25844 57876
rect 25452 57260 25508 57316
rect 25676 57148 25732 57204
rect 25340 56642 25396 56644
rect 25340 56590 25342 56642
rect 25342 56590 25394 56642
rect 25394 56590 25396 56642
rect 25340 56588 25396 56590
rect 25228 56306 25284 56308
rect 25228 56254 25230 56306
rect 25230 56254 25282 56306
rect 25282 56254 25284 56306
rect 25228 56252 25284 56254
rect 24220 53116 24276 53172
rect 23996 52946 24052 52948
rect 23996 52894 23998 52946
rect 23998 52894 24050 52946
rect 24050 52894 24052 52946
rect 23996 52892 24052 52894
rect 23548 52274 23604 52276
rect 23548 52222 23550 52274
rect 23550 52222 23602 52274
rect 23602 52222 23604 52274
rect 23548 52220 23604 52222
rect 22876 51490 22932 51492
rect 22876 51438 22878 51490
rect 22878 51438 22930 51490
rect 22930 51438 22932 51490
rect 22876 51436 22932 51438
rect 23436 51996 23492 52052
rect 22204 51100 22260 51156
rect 21196 49308 21252 49364
rect 22092 50540 22148 50596
rect 22316 50764 22372 50820
rect 23212 51490 23268 51492
rect 23212 51438 23214 51490
rect 23214 51438 23266 51490
rect 23266 51438 23268 51490
rect 23212 51436 23268 51438
rect 23324 51378 23380 51380
rect 23324 51326 23326 51378
rect 23326 51326 23378 51378
rect 23378 51326 23380 51378
rect 23324 51324 23380 51326
rect 23436 50988 23492 51044
rect 23324 50764 23380 50820
rect 23996 52444 24052 52500
rect 23772 51548 23828 51604
rect 23772 51378 23828 51380
rect 23772 51326 23774 51378
rect 23774 51326 23826 51378
rect 23826 51326 23828 51378
rect 23772 51324 23828 51326
rect 23660 50482 23716 50484
rect 23660 50430 23662 50482
rect 23662 50430 23714 50482
rect 23714 50430 23716 50482
rect 23660 50428 23716 50430
rect 24220 52668 24276 52724
rect 24892 54572 24948 54628
rect 24556 54460 24612 54516
rect 24444 53730 24500 53732
rect 24444 53678 24446 53730
rect 24446 53678 24498 53730
rect 24498 53678 24500 53730
rect 24444 53676 24500 53678
rect 24668 54236 24724 54292
rect 24780 53900 24836 53956
rect 24444 52892 24500 52948
rect 24220 52162 24276 52164
rect 24220 52110 24222 52162
rect 24222 52110 24274 52162
rect 24274 52110 24276 52162
rect 24220 52108 24276 52110
rect 24220 51378 24276 51380
rect 24220 51326 24222 51378
rect 24222 51326 24274 51378
rect 24274 51326 24276 51378
rect 24220 51324 24276 51326
rect 19628 47180 19684 47236
rect 20076 47292 20132 47348
rect 19836 47066 19892 47068
rect 19836 47014 19838 47066
rect 19838 47014 19890 47066
rect 19890 47014 19892 47066
rect 19836 47012 19892 47014
rect 19940 47066 19996 47068
rect 19940 47014 19942 47066
rect 19942 47014 19994 47066
rect 19994 47014 19996 47066
rect 19940 47012 19996 47014
rect 20044 47066 20100 47068
rect 20044 47014 20046 47066
rect 20046 47014 20098 47066
rect 20098 47014 20100 47066
rect 20044 47012 20100 47014
rect 20076 45612 20132 45668
rect 21532 48242 21588 48244
rect 21532 48190 21534 48242
rect 21534 48190 21586 48242
rect 21586 48190 21588 48242
rect 21532 48188 21588 48190
rect 20972 48076 21028 48132
rect 20972 47292 21028 47348
rect 21084 47628 21140 47684
rect 20636 46562 20692 46564
rect 20636 46510 20638 46562
rect 20638 46510 20690 46562
rect 20690 46510 20692 46562
rect 20636 46508 20692 46510
rect 20748 45948 20804 46004
rect 19836 45498 19892 45500
rect 19836 45446 19838 45498
rect 19838 45446 19890 45498
rect 19890 45446 19892 45498
rect 19836 45444 19892 45446
rect 19940 45498 19996 45500
rect 19940 45446 19942 45498
rect 19942 45446 19994 45498
rect 19994 45446 19996 45498
rect 19940 45444 19996 45446
rect 20044 45498 20100 45500
rect 20044 45446 20046 45498
rect 20046 45446 20098 45498
rect 20098 45446 20100 45498
rect 20044 45444 20100 45446
rect 18844 45164 18900 45220
rect 18620 43932 18676 43988
rect 18732 44044 18788 44100
rect 18172 43260 18228 43316
rect 17836 42028 17892 42084
rect 17836 40684 17892 40740
rect 17388 39676 17444 39732
rect 17500 39564 17556 39620
rect 17948 39900 18004 39956
rect 16380 36652 16436 36708
rect 16828 37436 16884 37492
rect 16492 36540 16548 36596
rect 16716 36540 16772 36596
rect 16492 35644 16548 35700
rect 16940 35644 16996 35700
rect 16716 35308 16772 35364
rect 15708 34300 15764 34356
rect 15260 33516 15316 33572
rect 15484 33516 15540 33572
rect 14028 32172 14084 32228
rect 12684 31948 12740 32004
rect 15596 32450 15652 32452
rect 15596 32398 15598 32450
rect 15598 32398 15650 32450
rect 15650 32398 15652 32450
rect 15596 32396 15652 32398
rect 14700 32284 14756 32340
rect 14476 31778 14532 31780
rect 14476 31726 14478 31778
rect 14478 31726 14530 31778
rect 14530 31726 14532 31778
rect 14476 31724 14532 31726
rect 14140 31666 14196 31668
rect 14140 31614 14142 31666
rect 14142 31614 14194 31666
rect 14194 31614 14196 31666
rect 14140 31612 14196 31614
rect 12684 31554 12740 31556
rect 12684 31502 12686 31554
rect 12686 31502 12738 31554
rect 12738 31502 12740 31554
rect 12684 31500 12740 31502
rect 13692 31554 13748 31556
rect 13692 31502 13694 31554
rect 13694 31502 13746 31554
rect 13746 31502 13748 31554
rect 13692 31500 13748 31502
rect 14028 31388 14084 31444
rect 12796 30882 12852 30884
rect 12796 30830 12798 30882
rect 12798 30830 12850 30882
rect 12850 30830 12852 30882
rect 12796 30828 12852 30830
rect 15372 31778 15428 31780
rect 15372 31726 15374 31778
rect 15374 31726 15426 31778
rect 15426 31726 15428 31778
rect 15372 31724 15428 31726
rect 15036 31554 15092 31556
rect 15036 31502 15038 31554
rect 15038 31502 15090 31554
rect 15090 31502 15092 31554
rect 15036 31500 15092 31502
rect 16828 35138 16884 35140
rect 16828 35086 16830 35138
rect 16830 35086 16882 35138
rect 16882 35086 16884 35138
rect 16828 35084 16884 35086
rect 16380 34860 16436 34916
rect 16156 34354 16212 34356
rect 16156 34302 16158 34354
rect 16158 34302 16210 34354
rect 16210 34302 16212 34354
rect 16156 34300 16212 34302
rect 16156 33906 16212 33908
rect 16156 33854 16158 33906
rect 16158 33854 16210 33906
rect 16210 33854 16212 33906
rect 16156 33852 16212 33854
rect 16268 33516 16324 33572
rect 16940 33234 16996 33236
rect 16940 33182 16942 33234
rect 16942 33182 16994 33234
rect 16994 33182 16996 33234
rect 16940 33180 16996 33182
rect 17500 38050 17556 38052
rect 17500 37998 17502 38050
rect 17502 37998 17554 38050
rect 17554 37998 17556 38050
rect 17500 37996 17556 37998
rect 17388 37938 17444 37940
rect 17388 37886 17390 37938
rect 17390 37886 17442 37938
rect 17442 37886 17444 37938
rect 17388 37884 17444 37886
rect 17836 37996 17892 38052
rect 18060 37884 18116 37940
rect 17500 36876 17556 36932
rect 17388 35698 17444 35700
rect 17388 35646 17390 35698
rect 17390 35646 17442 35698
rect 17442 35646 17444 35698
rect 17388 35644 17444 35646
rect 17612 35420 17668 35476
rect 17724 36540 17780 36596
rect 17948 37436 18004 37492
rect 18060 37100 18116 37156
rect 17164 34914 17220 34916
rect 17164 34862 17166 34914
rect 17166 34862 17218 34914
rect 17218 34862 17220 34914
rect 17164 34860 17220 34862
rect 17612 33404 17668 33460
rect 15820 31778 15876 31780
rect 15820 31726 15822 31778
rect 15822 31726 15874 31778
rect 15874 31726 15876 31778
rect 15820 31724 15876 31726
rect 16044 31612 16100 31668
rect 15596 31388 15652 31444
rect 14028 30828 14084 30884
rect 13020 30156 13076 30212
rect 12796 29426 12852 29428
rect 12796 29374 12798 29426
rect 12798 29374 12850 29426
rect 12850 29374 12852 29426
rect 12796 29372 12852 29374
rect 12796 28028 12852 28084
rect 12348 27804 12404 27860
rect 12572 27692 12628 27748
rect 12124 27244 12180 27300
rect 11228 27186 11284 27188
rect 11228 27134 11230 27186
rect 11230 27134 11282 27186
rect 11282 27134 11284 27186
rect 11228 27132 11284 27134
rect 11116 26460 11172 26516
rect 12012 26460 12068 26516
rect 11676 26348 11732 26404
rect 11340 26012 11396 26068
rect 8988 24668 9044 24724
rect 6300 24610 6356 24612
rect 6300 24558 6302 24610
rect 6302 24558 6354 24610
rect 6354 24558 6356 24610
rect 6300 24556 6356 24558
rect 2492 24220 2548 24276
rect 4476 24330 4532 24332
rect 4476 24278 4478 24330
rect 4478 24278 4530 24330
rect 4530 24278 4532 24330
rect 4476 24276 4532 24278
rect 4580 24330 4636 24332
rect 4580 24278 4582 24330
rect 4582 24278 4634 24330
rect 4634 24278 4636 24330
rect 4580 24276 4636 24278
rect 4684 24330 4740 24332
rect 4684 24278 4686 24330
rect 4686 24278 4738 24330
rect 4738 24278 4740 24330
rect 4684 24276 4740 24278
rect 6972 23826 7028 23828
rect 6972 23774 6974 23826
rect 6974 23774 7026 23826
rect 7026 23774 7028 23826
rect 6972 23772 7028 23774
rect 2492 23548 2548 23604
rect 7644 23938 7700 23940
rect 7644 23886 7646 23938
rect 7646 23886 7698 23938
rect 7698 23886 7700 23938
rect 7644 23884 7700 23886
rect 8764 24610 8820 24612
rect 8764 24558 8766 24610
rect 8766 24558 8818 24610
rect 8818 24558 8820 24610
rect 8764 24556 8820 24558
rect 10444 25506 10500 25508
rect 10444 25454 10446 25506
rect 10446 25454 10498 25506
rect 10498 25454 10500 25506
rect 10444 25452 10500 25454
rect 10220 24946 10276 24948
rect 10220 24894 10222 24946
rect 10222 24894 10274 24946
rect 10274 24894 10276 24946
rect 10220 24892 10276 24894
rect 10108 24780 10164 24836
rect 9324 23884 9380 23940
rect 8092 23772 8148 23828
rect 7756 23548 7812 23604
rect 7196 23436 7252 23492
rect 2156 23100 2212 23156
rect 2492 22876 2548 22932
rect 4476 22762 4532 22764
rect 4476 22710 4478 22762
rect 4478 22710 4530 22762
rect 4530 22710 4532 22762
rect 4476 22708 4532 22710
rect 4580 22762 4636 22764
rect 4580 22710 4582 22762
rect 4582 22710 4634 22762
rect 4634 22710 4636 22762
rect 4580 22708 4636 22710
rect 4684 22762 4740 22764
rect 4684 22710 4686 22762
rect 4686 22710 4738 22762
rect 4738 22710 4740 22762
rect 4684 22708 4740 22710
rect 2044 22316 2100 22372
rect 1708 22258 1764 22260
rect 1708 22206 1710 22258
rect 1710 22206 1762 22258
rect 1762 22206 1764 22258
rect 1708 22204 1764 22206
rect 2044 21698 2100 21700
rect 2044 21646 2046 21698
rect 2046 21646 2098 21698
rect 2098 21646 2100 21698
rect 2044 21644 2100 21646
rect 2380 21756 2436 21812
rect 2492 22204 2548 22260
rect 2156 21532 2212 21588
rect 1708 21420 1764 21476
rect 1708 20860 1764 20916
rect 1708 20188 1764 20244
rect 2044 20130 2100 20132
rect 2044 20078 2046 20130
rect 2046 20078 2098 20130
rect 2098 20078 2100 20130
rect 2044 20076 2100 20078
rect 1708 19516 1764 19572
rect 2044 18284 2100 18340
rect 1708 18172 1764 18228
rect 1708 17554 1764 17556
rect 1708 17502 1710 17554
rect 1710 17502 1762 17554
rect 1762 17502 1764 17554
rect 1708 17500 1764 17502
rect 2044 17442 2100 17444
rect 2044 17390 2046 17442
rect 2046 17390 2098 17442
rect 2098 17390 2100 17442
rect 2044 17388 2100 17390
rect 2492 20188 2548 20244
rect 3164 21756 3220 21812
rect 2940 21474 2996 21476
rect 2940 21422 2942 21474
rect 2942 21422 2994 21474
rect 2994 21422 2996 21474
rect 2940 21420 2996 21422
rect 4476 21194 4532 21196
rect 4476 21142 4478 21194
rect 4478 21142 4530 21194
rect 4530 21142 4532 21194
rect 4476 21140 4532 21142
rect 4580 21194 4636 21196
rect 4580 21142 4582 21194
rect 4582 21142 4634 21194
rect 4634 21142 4636 21194
rect 4580 21140 4636 21142
rect 4684 21194 4740 21196
rect 4684 21142 4686 21194
rect 4686 21142 4738 21194
rect 4738 21142 4740 21194
rect 4684 21140 4740 21142
rect 6076 23042 6132 23044
rect 6076 22990 6078 23042
rect 6078 22990 6130 23042
rect 6130 22990 6132 23042
rect 6076 22988 6132 22990
rect 6972 22988 7028 23044
rect 7084 22482 7140 22484
rect 7084 22430 7086 22482
rect 7086 22430 7138 22482
rect 7138 22430 7140 22482
rect 7084 22428 7140 22430
rect 7756 22428 7812 22484
rect 8764 23772 8820 23828
rect 8428 22428 8484 22484
rect 2716 19740 2772 19796
rect 6524 21586 6580 21588
rect 6524 21534 6526 21586
rect 6526 21534 6578 21586
rect 6578 21534 6580 21586
rect 6524 21532 6580 21534
rect 7868 21586 7924 21588
rect 7868 21534 7870 21586
rect 7870 21534 7922 21586
rect 7922 21534 7924 21586
rect 7868 21532 7924 21534
rect 9212 23548 9268 23604
rect 8988 22428 9044 22484
rect 9996 23660 10052 23716
rect 9660 23548 9716 23604
rect 9772 23154 9828 23156
rect 9772 23102 9774 23154
rect 9774 23102 9826 23154
rect 9826 23102 9828 23154
rect 9772 23100 9828 23102
rect 11228 24892 11284 24948
rect 10332 23436 10388 23492
rect 11116 24556 11172 24612
rect 11788 24722 11844 24724
rect 11788 24670 11790 24722
rect 11790 24670 11842 24722
rect 11842 24670 11844 24722
rect 11788 24668 11844 24670
rect 11676 24556 11732 24612
rect 11228 23996 11284 24052
rect 11788 23884 11844 23940
rect 11228 23660 11284 23716
rect 14028 29596 14084 29652
rect 14252 29372 14308 29428
rect 13692 29314 13748 29316
rect 13692 29262 13694 29314
rect 13694 29262 13746 29314
rect 13746 29262 13748 29314
rect 13692 29260 13748 29262
rect 13580 29148 13636 29204
rect 14252 29148 14308 29204
rect 13468 28812 13524 28868
rect 13468 28642 13524 28644
rect 13468 28590 13470 28642
rect 13470 28590 13522 28642
rect 13522 28590 13524 28642
rect 13468 28588 13524 28590
rect 14252 28642 14308 28644
rect 14252 28590 14254 28642
rect 14254 28590 14306 28642
rect 14306 28590 14308 28642
rect 14252 28588 14308 28590
rect 12796 27244 12852 27300
rect 15036 28530 15092 28532
rect 15036 28478 15038 28530
rect 15038 28478 15090 28530
rect 15090 28478 15092 28530
rect 15036 28476 15092 28478
rect 14364 28082 14420 28084
rect 14364 28030 14366 28082
rect 14366 28030 14418 28082
rect 14418 28030 14420 28082
rect 14364 28028 14420 28030
rect 14924 28028 14980 28084
rect 12572 27132 12628 27188
rect 12124 24050 12180 24052
rect 12124 23998 12126 24050
rect 12126 23998 12178 24050
rect 12178 23998 12180 24050
rect 12124 23996 12180 23998
rect 12124 23772 12180 23828
rect 13692 27580 13748 27636
rect 13020 26348 13076 26404
rect 12796 25676 12852 25732
rect 12908 25004 12964 25060
rect 12348 23660 12404 23716
rect 12236 23100 12292 23156
rect 6860 21308 6916 21364
rect 6300 20636 6356 20692
rect 6748 20972 6804 21028
rect 2492 19516 2548 19572
rect 4476 19626 4532 19628
rect 4476 19574 4478 19626
rect 4478 19574 4530 19626
rect 4530 19574 4532 19626
rect 4476 19572 4532 19574
rect 4580 19626 4636 19628
rect 4580 19574 4582 19626
rect 4582 19574 4634 19626
rect 4634 19574 4636 19626
rect 4580 19572 4636 19574
rect 4684 19626 4740 19628
rect 4684 19574 4686 19626
rect 4686 19574 4738 19626
rect 4738 19574 4740 19626
rect 4684 19572 4740 19574
rect 10108 22370 10164 22372
rect 10108 22318 10110 22370
rect 10110 22318 10162 22370
rect 10162 22318 10164 22370
rect 10108 22316 10164 22318
rect 11788 22482 11844 22484
rect 11788 22430 11790 22482
rect 11790 22430 11842 22482
rect 11842 22430 11844 22482
rect 11788 22428 11844 22430
rect 11004 22092 11060 22148
rect 9212 21532 9268 21588
rect 8988 21420 9044 21476
rect 8988 20914 9044 20916
rect 8988 20862 8990 20914
rect 8990 20862 9042 20914
rect 9042 20862 9044 20914
rect 8988 20860 9044 20862
rect 9996 21980 10052 22036
rect 9660 21474 9716 21476
rect 9660 21422 9662 21474
rect 9662 21422 9714 21474
rect 9714 21422 9716 21474
rect 9660 21420 9716 21422
rect 9548 21362 9604 21364
rect 9548 21310 9550 21362
rect 9550 21310 9602 21362
rect 9602 21310 9604 21362
rect 9548 21308 9604 21310
rect 9212 20748 9268 20804
rect 9324 20690 9380 20692
rect 9324 20638 9326 20690
rect 9326 20638 9378 20690
rect 9378 20638 9380 20690
rect 9324 20636 9380 20638
rect 7980 19852 8036 19908
rect 7196 19628 7252 19684
rect 6076 18396 6132 18452
rect 6524 18284 6580 18340
rect 2492 18172 2548 18228
rect 4476 18058 4532 18060
rect 4476 18006 4478 18058
rect 4478 18006 4530 18058
rect 4530 18006 4532 18058
rect 4476 18004 4532 18006
rect 4580 18058 4636 18060
rect 4580 18006 4582 18058
rect 4582 18006 4634 18058
rect 4634 18006 4636 18058
rect 4580 18004 4636 18006
rect 4684 18058 4740 18060
rect 4684 18006 4686 18058
rect 4686 18006 4738 18058
rect 4738 18006 4740 18058
rect 6972 18060 7028 18116
rect 7084 18396 7140 18452
rect 4684 18004 4740 18006
rect 2156 17276 2212 17332
rect 2492 17500 2548 17556
rect 2716 17554 2772 17556
rect 2716 17502 2718 17554
rect 2718 17502 2770 17554
rect 2770 17502 2772 17554
rect 2716 17500 2772 17502
rect 7868 19068 7924 19124
rect 8988 19906 9044 19908
rect 8988 19854 8990 19906
rect 8990 19854 9042 19906
rect 9042 19854 9044 19906
rect 8988 19852 9044 19854
rect 8764 19068 8820 19124
rect 8876 18620 8932 18676
rect 8316 18396 8372 18452
rect 8204 18284 8260 18340
rect 7868 18172 7924 18228
rect 7420 17500 7476 17556
rect 2380 16828 2436 16884
rect 3164 16828 3220 16884
rect 5180 17388 5236 17444
rect 2044 16716 2100 16772
rect 4476 16490 4532 16492
rect 4476 16438 4478 16490
rect 4478 16438 4530 16490
rect 4530 16438 4532 16490
rect 4476 16436 4532 16438
rect 4580 16490 4636 16492
rect 4580 16438 4582 16490
rect 4582 16438 4634 16490
rect 4634 16438 4636 16490
rect 4580 16436 4636 16438
rect 4684 16490 4740 16492
rect 4684 16438 4686 16490
rect 4686 16438 4738 16490
rect 4738 16438 4740 16490
rect 4684 16436 4740 16438
rect 1820 16210 1876 16212
rect 1820 16158 1822 16210
rect 1822 16158 1874 16210
rect 1874 16158 1876 16210
rect 1820 16156 1876 16158
rect 4476 14922 4532 14924
rect 4476 14870 4478 14922
rect 4478 14870 4530 14922
rect 4530 14870 4532 14922
rect 4476 14868 4532 14870
rect 4580 14922 4636 14924
rect 4580 14870 4582 14922
rect 4582 14870 4634 14922
rect 4634 14870 4636 14922
rect 4580 14868 4636 14870
rect 4684 14922 4740 14924
rect 4684 14870 4686 14922
rect 4686 14870 4738 14922
rect 4738 14870 4740 14922
rect 4684 14868 4740 14870
rect 9548 20076 9604 20132
rect 9660 19234 9716 19236
rect 9660 19182 9662 19234
rect 9662 19182 9714 19234
rect 9714 19182 9716 19234
rect 9660 19180 9716 19182
rect 8988 16828 9044 16884
rect 9548 18060 9604 18116
rect 8876 16770 8932 16772
rect 8876 16718 8878 16770
rect 8878 16718 8930 16770
rect 8930 16718 8932 16770
rect 8876 16716 8932 16718
rect 8764 16604 8820 16660
rect 5180 14476 5236 14532
rect 9884 18620 9940 18676
rect 11228 21980 11284 22036
rect 13580 26908 13636 26964
rect 13468 25730 13524 25732
rect 13468 25678 13470 25730
rect 13470 25678 13522 25730
rect 13522 25678 13524 25730
rect 13468 25676 13524 25678
rect 14028 27020 14084 27076
rect 14140 27244 14196 27300
rect 14476 27020 14532 27076
rect 12908 23772 12964 23828
rect 13692 23826 13748 23828
rect 13692 23774 13694 23826
rect 13694 23774 13746 23826
rect 13746 23774 13748 23826
rect 13692 23772 13748 23774
rect 13020 23154 13076 23156
rect 13020 23102 13022 23154
rect 13022 23102 13074 23154
rect 13074 23102 13076 23154
rect 13020 23100 13076 23102
rect 13468 23100 13524 23156
rect 13804 23324 13860 23380
rect 10108 21026 10164 21028
rect 10108 20974 10110 21026
rect 10110 20974 10162 21026
rect 10162 20974 10164 21026
rect 10108 20972 10164 20974
rect 10332 20914 10388 20916
rect 10332 20862 10334 20914
rect 10334 20862 10386 20914
rect 10386 20862 10388 20914
rect 10332 20860 10388 20862
rect 10556 20802 10612 20804
rect 10556 20750 10558 20802
rect 10558 20750 10610 20802
rect 10610 20750 10612 20802
rect 10556 20748 10612 20750
rect 9772 17724 9828 17780
rect 9884 18396 9940 18452
rect 11452 19852 11508 19908
rect 11004 19628 11060 19684
rect 10108 16716 10164 16772
rect 10220 16604 10276 16660
rect 11452 19068 11508 19124
rect 11340 18396 11396 18452
rect 10556 18338 10612 18340
rect 10556 18286 10558 18338
rect 10558 18286 10610 18338
rect 10610 18286 10612 18338
rect 10556 18284 10612 18286
rect 10444 18226 10500 18228
rect 10444 18174 10446 18226
rect 10446 18174 10498 18226
rect 10498 18174 10500 18226
rect 10444 18172 10500 18174
rect 11116 17778 11172 17780
rect 11116 17726 11118 17778
rect 11118 17726 11170 17778
rect 11170 17726 11172 17778
rect 11116 17724 11172 17726
rect 11116 17500 11172 17556
rect 10332 16492 10388 16548
rect 9772 14530 9828 14532
rect 9772 14478 9774 14530
rect 9774 14478 9826 14530
rect 9826 14478 9828 14530
rect 9772 14476 9828 14478
rect 13468 22146 13524 22148
rect 13468 22094 13470 22146
rect 13470 22094 13522 22146
rect 13522 22094 13524 22146
rect 13468 22092 13524 22094
rect 14252 25506 14308 25508
rect 14252 25454 14254 25506
rect 14254 25454 14306 25506
rect 14306 25454 14308 25506
rect 14252 25452 14308 25454
rect 15148 27692 15204 27748
rect 15372 28588 15428 28644
rect 15932 29314 15988 29316
rect 15932 29262 15934 29314
rect 15934 29262 15986 29314
rect 15986 29262 15988 29314
rect 15932 29260 15988 29262
rect 16044 29148 16100 29204
rect 16716 31890 16772 31892
rect 16716 31838 16718 31890
rect 16718 31838 16770 31890
rect 16770 31838 16772 31890
rect 16716 31836 16772 31838
rect 16604 31724 16660 31780
rect 16380 31500 16436 31556
rect 16604 31106 16660 31108
rect 16604 31054 16606 31106
rect 16606 31054 16658 31106
rect 16658 31054 16660 31106
rect 16604 31052 16660 31054
rect 16268 30716 16324 30772
rect 16716 29538 16772 29540
rect 16716 29486 16718 29538
rect 16718 29486 16770 29538
rect 16770 29486 16772 29538
rect 16716 29484 16772 29486
rect 16604 29202 16660 29204
rect 16604 29150 16606 29202
rect 16606 29150 16658 29202
rect 16658 29150 16660 29202
rect 16604 29148 16660 29150
rect 16156 28700 16212 28756
rect 16604 28700 16660 28756
rect 15820 28476 15876 28532
rect 15484 27074 15540 27076
rect 15484 27022 15486 27074
rect 15486 27022 15538 27074
rect 15538 27022 15540 27074
rect 15484 27020 15540 27022
rect 15596 27804 15652 27860
rect 14700 26348 14756 26404
rect 14924 26012 14980 26068
rect 14924 25676 14980 25732
rect 14700 25618 14756 25620
rect 14700 25566 14702 25618
rect 14702 25566 14754 25618
rect 14754 25566 14756 25618
rect 14700 25564 14756 25566
rect 14252 25004 14308 25060
rect 14588 24946 14644 24948
rect 14588 24894 14590 24946
rect 14590 24894 14642 24946
rect 14642 24894 14644 24946
rect 14588 24892 14644 24894
rect 14364 23378 14420 23380
rect 14364 23326 14366 23378
rect 14366 23326 14418 23378
rect 14418 23326 14420 23378
rect 14364 23324 14420 23326
rect 13916 21980 13972 22036
rect 11900 19234 11956 19236
rect 11900 19182 11902 19234
rect 11902 19182 11954 19234
rect 11954 19182 11956 19234
rect 11900 19180 11956 19182
rect 11452 17500 11508 17556
rect 11564 18508 11620 18564
rect 11340 17164 11396 17220
rect 11228 16828 11284 16884
rect 12236 20076 12292 20132
rect 11676 18396 11732 18452
rect 12348 19516 12404 19572
rect 12348 18508 12404 18564
rect 12684 19180 12740 19236
rect 12124 18060 12180 18116
rect 12348 17500 12404 17556
rect 12124 17164 12180 17220
rect 13468 20076 13524 20132
rect 13692 20076 13748 20132
rect 13132 19292 13188 19348
rect 13580 19404 13636 19460
rect 12908 19122 12964 19124
rect 12908 19070 12910 19122
rect 12910 19070 12962 19122
rect 12962 19070 12964 19122
rect 12908 19068 12964 19070
rect 12908 18060 12964 18116
rect 14252 21420 14308 21476
rect 13916 19740 13972 19796
rect 13692 18060 13748 18116
rect 14252 19628 14308 19684
rect 14364 18172 14420 18228
rect 14588 19740 14644 19796
rect 15372 26460 15428 26516
rect 15148 25676 15204 25732
rect 15372 25452 15428 25508
rect 17164 28754 17220 28756
rect 17164 28702 17166 28754
rect 17166 28702 17218 28754
rect 17218 28702 17220 28754
rect 17164 28700 17220 28702
rect 16716 28082 16772 28084
rect 16716 28030 16718 28082
rect 16718 28030 16770 28082
rect 16770 28030 16772 28082
rect 16716 28028 16772 28030
rect 15036 23884 15092 23940
rect 16268 26908 16324 26964
rect 15820 26012 15876 26068
rect 16156 26178 16212 26180
rect 16156 26126 16158 26178
rect 16158 26126 16210 26178
rect 16210 26126 16212 26178
rect 16156 26124 16212 26126
rect 15596 23660 15652 23716
rect 16940 26962 16996 26964
rect 16940 26910 16942 26962
rect 16942 26910 16994 26962
rect 16994 26910 16996 26962
rect 16940 26908 16996 26910
rect 16604 26460 16660 26516
rect 16492 26124 16548 26180
rect 17724 32508 17780 32564
rect 17500 31836 17556 31892
rect 18620 42530 18676 42532
rect 18620 42478 18622 42530
rect 18622 42478 18674 42530
rect 18674 42478 18676 42530
rect 18620 42476 18676 42478
rect 19292 44492 19348 44548
rect 19180 43538 19236 43540
rect 19180 43486 19182 43538
rect 19182 43486 19234 43538
rect 19234 43486 19236 43538
rect 19180 43484 19236 43486
rect 19404 43932 19460 43988
rect 19180 43148 19236 43204
rect 20188 44210 20244 44212
rect 20188 44158 20190 44210
rect 20190 44158 20242 44210
rect 20242 44158 20244 44210
rect 20188 44156 20244 44158
rect 20076 44098 20132 44100
rect 20076 44046 20078 44098
rect 20078 44046 20130 44098
rect 20130 44046 20132 44098
rect 20076 44044 20132 44046
rect 19836 43930 19892 43932
rect 19836 43878 19838 43930
rect 19838 43878 19890 43930
rect 19890 43878 19892 43930
rect 19836 43876 19892 43878
rect 19940 43930 19996 43932
rect 19940 43878 19942 43930
rect 19942 43878 19994 43930
rect 19994 43878 19996 43930
rect 19940 43876 19996 43878
rect 20044 43930 20100 43932
rect 20044 43878 20046 43930
rect 20046 43878 20098 43930
rect 20098 43878 20100 43930
rect 20044 43876 20100 43878
rect 20188 43708 20244 43764
rect 20636 45052 20692 45108
rect 20748 44210 20804 44212
rect 20748 44158 20750 44210
rect 20750 44158 20802 44210
rect 20802 44158 20804 44210
rect 20748 44156 20804 44158
rect 20524 43596 20580 43652
rect 20972 45388 21028 45444
rect 19740 43148 19796 43204
rect 20188 42924 20244 42980
rect 18844 42700 18900 42756
rect 19964 42754 20020 42756
rect 19964 42702 19966 42754
rect 19966 42702 20018 42754
rect 20018 42702 20020 42754
rect 19964 42700 20020 42702
rect 19836 42362 19892 42364
rect 19836 42310 19838 42362
rect 19838 42310 19890 42362
rect 19890 42310 19892 42362
rect 19836 42308 19892 42310
rect 19940 42362 19996 42364
rect 19940 42310 19942 42362
rect 19942 42310 19994 42362
rect 19994 42310 19996 42362
rect 19940 42308 19996 42310
rect 20044 42362 20100 42364
rect 20044 42310 20046 42362
rect 20046 42310 20098 42362
rect 20098 42310 20100 42362
rect 20044 42308 20100 42310
rect 18508 40572 18564 40628
rect 18284 40236 18340 40292
rect 18732 39676 18788 39732
rect 18284 38220 18340 38276
rect 18396 37100 18452 37156
rect 18284 36652 18340 36708
rect 18620 37100 18676 37156
rect 19964 41186 20020 41188
rect 19964 41134 19966 41186
rect 19966 41134 20018 41186
rect 20018 41134 20020 41186
rect 19964 41132 20020 41134
rect 19068 40572 19124 40628
rect 19852 40962 19908 40964
rect 19852 40910 19854 40962
rect 19854 40910 19906 40962
rect 19906 40910 19908 40962
rect 19852 40908 19908 40910
rect 19836 40794 19892 40796
rect 19836 40742 19838 40794
rect 19838 40742 19890 40794
rect 19890 40742 19892 40794
rect 19836 40740 19892 40742
rect 19940 40794 19996 40796
rect 19940 40742 19942 40794
rect 19942 40742 19994 40794
rect 19994 40742 19996 40794
rect 19940 40740 19996 40742
rect 20044 40794 20100 40796
rect 20044 40742 20046 40794
rect 20046 40742 20098 40794
rect 20098 40742 20100 40794
rect 20044 40740 20100 40742
rect 19628 40012 19684 40068
rect 20412 40572 20468 40628
rect 20188 39788 20244 39844
rect 19964 39730 20020 39732
rect 19964 39678 19966 39730
rect 19966 39678 20018 39730
rect 20018 39678 20020 39730
rect 19964 39676 20020 39678
rect 19516 39618 19572 39620
rect 19516 39566 19518 39618
rect 19518 39566 19570 39618
rect 19570 39566 19572 39618
rect 19516 39564 19572 39566
rect 19292 39116 19348 39172
rect 19836 39226 19892 39228
rect 19836 39174 19838 39226
rect 19838 39174 19890 39226
rect 19890 39174 19892 39226
rect 19836 39172 19892 39174
rect 19940 39226 19996 39228
rect 19940 39174 19942 39226
rect 19942 39174 19994 39226
rect 19994 39174 19996 39226
rect 19940 39172 19996 39174
rect 20044 39226 20100 39228
rect 20044 39174 20046 39226
rect 20046 39174 20098 39226
rect 20098 39174 20100 39226
rect 20044 39172 20100 39174
rect 19852 38556 19908 38612
rect 18844 37996 18900 38052
rect 19516 38332 19572 38388
rect 20524 38444 20580 38500
rect 19292 37660 19348 37716
rect 18956 37490 19012 37492
rect 18956 37438 18958 37490
rect 18958 37438 19010 37490
rect 19010 37438 19012 37490
rect 18956 37436 19012 37438
rect 19836 37658 19892 37660
rect 19836 37606 19838 37658
rect 19838 37606 19890 37658
rect 19890 37606 19892 37658
rect 19836 37604 19892 37606
rect 19940 37658 19996 37660
rect 19940 37606 19942 37658
rect 19942 37606 19994 37658
rect 19994 37606 19996 37658
rect 19940 37604 19996 37606
rect 20044 37658 20100 37660
rect 20044 37606 20046 37658
rect 20046 37606 20098 37658
rect 20098 37606 20100 37658
rect 20044 37604 20100 37606
rect 20076 37436 20132 37492
rect 20076 37266 20132 37268
rect 20076 37214 20078 37266
rect 20078 37214 20130 37266
rect 20130 37214 20132 37266
rect 20076 37212 20132 37214
rect 18844 36876 18900 36932
rect 20412 38050 20468 38052
rect 20412 37998 20414 38050
rect 20414 37998 20466 38050
rect 20466 37998 20468 38050
rect 20412 37996 20468 37998
rect 20188 36988 20244 37044
rect 20524 37436 20580 37492
rect 20524 36876 20580 36932
rect 18732 35532 18788 35588
rect 18060 33458 18116 33460
rect 18060 33406 18062 33458
rect 18062 33406 18114 33458
rect 18114 33406 18116 33458
rect 18060 33404 18116 33406
rect 18508 33516 18564 33572
rect 18956 35084 19012 35140
rect 19404 35810 19460 35812
rect 19404 35758 19406 35810
rect 19406 35758 19458 35810
rect 19458 35758 19460 35810
rect 19404 35756 19460 35758
rect 19404 35420 19460 35476
rect 18844 33346 18900 33348
rect 18844 33294 18846 33346
rect 18846 33294 18898 33346
rect 18898 33294 18900 33346
rect 18844 33292 18900 33294
rect 18508 32562 18564 32564
rect 18508 32510 18510 32562
rect 18510 32510 18562 32562
rect 18562 32510 18564 32562
rect 18508 32508 18564 32510
rect 18844 32396 18900 32452
rect 17836 31836 17892 31892
rect 19292 33404 19348 33460
rect 19180 31724 19236 31780
rect 17612 31500 17668 31556
rect 17500 31106 17556 31108
rect 17500 31054 17502 31106
rect 17502 31054 17554 31106
rect 17554 31054 17556 31106
rect 17500 31052 17556 31054
rect 17500 30770 17556 30772
rect 17500 30718 17502 30770
rect 17502 30718 17554 30770
rect 17554 30718 17556 30770
rect 17500 30716 17556 30718
rect 17500 28642 17556 28644
rect 17500 28590 17502 28642
rect 17502 28590 17554 28642
rect 17554 28590 17556 28642
rect 17500 28588 17556 28590
rect 17500 28082 17556 28084
rect 17500 28030 17502 28082
rect 17502 28030 17554 28082
rect 17554 28030 17556 28082
rect 17500 28028 17556 28030
rect 17612 27356 17668 27412
rect 18284 26908 18340 26964
rect 18508 26796 18564 26852
rect 17388 26236 17444 26292
rect 19836 36090 19892 36092
rect 19836 36038 19838 36090
rect 19838 36038 19890 36090
rect 19890 36038 19892 36090
rect 19836 36036 19892 36038
rect 19940 36090 19996 36092
rect 19940 36038 19942 36090
rect 19942 36038 19994 36090
rect 19994 36038 19996 36090
rect 19940 36036 19996 36038
rect 20044 36090 20100 36092
rect 20044 36038 20046 36090
rect 20046 36038 20098 36090
rect 20098 36038 20100 36090
rect 20044 36036 20100 36038
rect 19740 35532 19796 35588
rect 19836 34522 19892 34524
rect 19836 34470 19838 34522
rect 19838 34470 19890 34522
rect 19890 34470 19892 34522
rect 19836 34468 19892 34470
rect 19940 34522 19996 34524
rect 19940 34470 19942 34522
rect 19942 34470 19994 34522
rect 19994 34470 19996 34522
rect 19940 34468 19996 34470
rect 20044 34522 20100 34524
rect 20044 34470 20046 34522
rect 20046 34470 20098 34522
rect 20098 34470 20100 34522
rect 20044 34468 20100 34470
rect 19628 33346 19684 33348
rect 19628 33294 19630 33346
rect 19630 33294 19682 33346
rect 19682 33294 19684 33346
rect 19628 33292 19684 33294
rect 19852 33628 19908 33684
rect 20412 33628 20468 33684
rect 20412 33180 20468 33236
rect 19836 32954 19892 32956
rect 19836 32902 19838 32954
rect 19838 32902 19890 32954
rect 19890 32902 19892 32954
rect 19836 32900 19892 32902
rect 19940 32954 19996 32956
rect 19940 32902 19942 32954
rect 19942 32902 19994 32954
rect 19994 32902 19996 32954
rect 19940 32900 19996 32902
rect 20044 32954 20100 32956
rect 20044 32902 20046 32954
rect 20046 32902 20098 32954
rect 20098 32902 20100 32954
rect 20044 32900 20100 32902
rect 21756 48076 21812 48132
rect 21420 47516 21476 47572
rect 21756 47628 21812 47684
rect 21980 47516 22036 47572
rect 22428 48242 22484 48244
rect 22428 48190 22430 48242
rect 22430 48190 22482 48242
rect 22482 48190 22484 48242
rect 22428 48188 22484 48190
rect 22428 47516 22484 47572
rect 22092 46844 22148 46900
rect 21308 45612 21364 45668
rect 21420 45276 21476 45332
rect 21308 45052 21364 45108
rect 21532 44492 21588 44548
rect 21532 44098 21588 44100
rect 21532 44046 21534 44098
rect 21534 44046 21586 44098
rect 21586 44046 21588 44098
rect 21532 44044 21588 44046
rect 21756 46620 21812 46676
rect 22652 47458 22708 47460
rect 22652 47406 22654 47458
rect 22654 47406 22706 47458
rect 22706 47406 22708 47458
rect 22652 47404 22708 47406
rect 23772 48466 23828 48468
rect 23772 48414 23774 48466
rect 23774 48414 23826 48466
rect 23826 48414 23828 48466
rect 23772 48412 23828 48414
rect 23660 48076 23716 48132
rect 23100 47346 23156 47348
rect 23100 47294 23102 47346
rect 23102 47294 23154 47346
rect 23154 47294 23156 47346
rect 23100 47292 23156 47294
rect 22428 46844 22484 46900
rect 22428 46508 22484 46564
rect 22540 45890 22596 45892
rect 22540 45838 22542 45890
rect 22542 45838 22594 45890
rect 22594 45838 22596 45890
rect 22540 45836 22596 45838
rect 21756 45612 21812 45668
rect 22092 45666 22148 45668
rect 22092 45614 22094 45666
rect 22094 45614 22146 45666
rect 22146 45614 22148 45666
rect 22092 45612 22148 45614
rect 20748 42924 20804 42980
rect 21308 43260 21364 43316
rect 20748 40908 20804 40964
rect 20748 39788 20804 39844
rect 20748 39116 20804 39172
rect 20860 38892 20916 38948
rect 21084 42700 21140 42756
rect 21084 40626 21140 40628
rect 21084 40574 21086 40626
rect 21086 40574 21138 40626
rect 21138 40574 21140 40626
rect 21084 40572 21140 40574
rect 21644 43260 21700 43316
rect 21868 45388 21924 45444
rect 22092 44492 22148 44548
rect 22652 44322 22708 44324
rect 22652 44270 22654 44322
rect 22654 44270 22706 44322
rect 22706 44270 22708 44322
rect 22652 44268 22708 44270
rect 23660 47346 23716 47348
rect 23660 47294 23662 47346
rect 23662 47294 23714 47346
rect 23714 47294 23716 47346
rect 23660 47292 23716 47294
rect 23884 47180 23940 47236
rect 23548 46396 23604 46452
rect 23772 45890 23828 45892
rect 23772 45838 23774 45890
rect 23774 45838 23826 45890
rect 23826 45838 23828 45890
rect 23772 45836 23828 45838
rect 23324 45666 23380 45668
rect 23324 45614 23326 45666
rect 23326 45614 23378 45666
rect 23378 45614 23380 45666
rect 23324 45612 23380 45614
rect 23212 45106 23268 45108
rect 23212 45054 23214 45106
rect 23214 45054 23266 45106
rect 23266 45054 23268 45106
rect 23212 45052 23268 45054
rect 24332 49532 24388 49588
rect 24220 48412 24276 48468
rect 24220 47292 24276 47348
rect 23212 44268 23268 44324
rect 24108 44380 24164 44436
rect 22204 43260 22260 43316
rect 23100 42924 23156 42980
rect 21980 42866 22036 42868
rect 21980 42814 21982 42866
rect 21982 42814 22034 42866
rect 22034 42814 22036 42866
rect 21980 42812 22036 42814
rect 21644 42364 21700 42420
rect 21308 42028 21364 42084
rect 20972 38220 21028 38276
rect 21084 38892 21140 38948
rect 20860 37772 20916 37828
rect 20860 37154 20916 37156
rect 20860 37102 20862 37154
rect 20862 37102 20914 37154
rect 20914 37102 20916 37154
rect 20860 37100 20916 37102
rect 20972 36988 21028 37044
rect 22540 42364 22596 42420
rect 21980 41916 22036 41972
rect 22652 41804 22708 41860
rect 21532 41356 21588 41412
rect 21420 40908 21476 40964
rect 21980 41298 22036 41300
rect 21980 41246 21982 41298
rect 21982 41246 22034 41298
rect 22034 41246 22036 41298
rect 21980 41244 22036 41246
rect 24220 44210 24276 44212
rect 24220 44158 24222 44210
rect 24222 44158 24274 44210
rect 24274 44158 24276 44210
rect 24220 44156 24276 44158
rect 23324 43538 23380 43540
rect 23324 43486 23326 43538
rect 23326 43486 23378 43538
rect 23378 43486 23380 43538
rect 23324 43484 23380 43486
rect 23324 42924 23380 42980
rect 22988 41804 23044 41860
rect 22652 41074 22708 41076
rect 22652 41022 22654 41074
rect 22654 41022 22706 41074
rect 22706 41022 22708 41074
rect 22652 41020 22708 41022
rect 22988 41074 23044 41076
rect 22988 41022 22990 41074
rect 22990 41022 23042 41074
rect 23042 41022 23044 41074
rect 22988 41020 23044 41022
rect 23100 41132 23156 41188
rect 21868 40908 21924 40964
rect 23100 40626 23156 40628
rect 23100 40574 23102 40626
rect 23102 40574 23154 40626
rect 23154 40574 23156 40626
rect 23100 40572 23156 40574
rect 21532 39788 21588 39844
rect 21196 37212 21252 37268
rect 21308 37436 21364 37492
rect 20636 36652 20692 36708
rect 20636 36204 20692 36260
rect 20748 34802 20804 34804
rect 20748 34750 20750 34802
rect 20750 34750 20802 34802
rect 20802 34750 20804 34802
rect 20748 34748 20804 34750
rect 20636 33516 20692 33572
rect 19628 31778 19684 31780
rect 19628 31726 19630 31778
rect 19630 31726 19682 31778
rect 19682 31726 19684 31778
rect 19628 31724 19684 31726
rect 19836 31386 19892 31388
rect 19836 31334 19838 31386
rect 19838 31334 19890 31386
rect 19890 31334 19892 31386
rect 19836 31332 19892 31334
rect 19940 31386 19996 31388
rect 19940 31334 19942 31386
rect 19942 31334 19994 31386
rect 19994 31334 19996 31386
rect 19940 31332 19996 31334
rect 20044 31386 20100 31388
rect 20044 31334 20046 31386
rect 20046 31334 20098 31386
rect 20098 31334 20100 31386
rect 20044 31332 20100 31334
rect 19404 30322 19460 30324
rect 19404 30270 19406 30322
rect 19406 30270 19458 30322
rect 19458 30270 19460 30322
rect 19404 30268 19460 30270
rect 18956 30044 19012 30100
rect 18956 28700 19012 28756
rect 19068 29932 19124 29988
rect 20076 29932 20132 29988
rect 19836 29818 19892 29820
rect 19836 29766 19838 29818
rect 19838 29766 19890 29818
rect 19890 29766 19892 29818
rect 19836 29764 19892 29766
rect 19940 29818 19996 29820
rect 19940 29766 19942 29818
rect 19942 29766 19994 29818
rect 19994 29766 19996 29818
rect 19940 29764 19996 29766
rect 20044 29818 20100 29820
rect 20044 29766 20046 29818
rect 20046 29766 20098 29818
rect 20098 29766 20100 29818
rect 20044 29764 20100 29766
rect 19068 28588 19124 28644
rect 19628 28588 19684 28644
rect 19836 28250 19892 28252
rect 19836 28198 19838 28250
rect 19838 28198 19890 28250
rect 19890 28198 19892 28250
rect 19836 28196 19892 28198
rect 19940 28250 19996 28252
rect 19940 28198 19942 28250
rect 19942 28198 19994 28250
rect 19994 28198 19996 28250
rect 19940 28196 19996 28198
rect 20044 28250 20100 28252
rect 20044 28198 20046 28250
rect 20046 28198 20098 28250
rect 20098 28198 20100 28250
rect 20044 28196 20100 28198
rect 19852 27746 19908 27748
rect 19852 27694 19854 27746
rect 19854 27694 19906 27746
rect 19906 27694 19908 27746
rect 19852 27692 19908 27694
rect 17612 26572 17668 26628
rect 18732 26908 18788 26964
rect 18060 26290 18116 26292
rect 18060 26238 18062 26290
rect 18062 26238 18114 26290
rect 18114 26238 18116 26290
rect 18060 26236 18116 26238
rect 18508 26124 18564 26180
rect 17052 26012 17108 26068
rect 17948 26066 18004 26068
rect 17948 26014 17950 26066
rect 17950 26014 18002 26066
rect 18002 26014 18004 26066
rect 17948 26012 18004 26014
rect 18172 26012 18228 26068
rect 16828 25452 16884 25508
rect 18396 25618 18452 25620
rect 18396 25566 18398 25618
rect 18398 25566 18450 25618
rect 18450 25566 18452 25618
rect 18396 25564 18452 25566
rect 17724 24610 17780 24612
rect 17724 24558 17726 24610
rect 17726 24558 17778 24610
rect 17778 24558 17780 24610
rect 17724 24556 17780 24558
rect 17276 23938 17332 23940
rect 17276 23886 17278 23938
rect 17278 23886 17330 23938
rect 17330 23886 17332 23938
rect 17276 23884 17332 23886
rect 17724 23884 17780 23940
rect 16156 23324 16212 23380
rect 19068 26796 19124 26852
rect 18844 26572 18900 26628
rect 19068 26348 19124 26404
rect 19180 26684 19236 26740
rect 20076 26962 20132 26964
rect 20076 26910 20078 26962
rect 20078 26910 20130 26962
rect 20130 26910 20132 26962
rect 20076 26908 20132 26910
rect 20524 32620 20580 32676
rect 20412 28754 20468 28756
rect 20412 28702 20414 28754
rect 20414 28702 20466 28754
rect 20466 28702 20468 28754
rect 20412 28700 20468 28702
rect 19628 26572 19684 26628
rect 19836 26682 19892 26684
rect 19836 26630 19838 26682
rect 19838 26630 19890 26682
rect 19890 26630 19892 26682
rect 19836 26628 19892 26630
rect 19940 26682 19996 26684
rect 19940 26630 19942 26682
rect 19942 26630 19994 26682
rect 19994 26630 19996 26682
rect 19940 26628 19996 26630
rect 20044 26682 20100 26684
rect 20044 26630 20046 26682
rect 20046 26630 20098 26682
rect 20098 26630 20100 26682
rect 20044 26628 20100 26630
rect 19180 26124 19236 26180
rect 18732 25452 18788 25508
rect 20412 26290 20468 26292
rect 20412 26238 20414 26290
rect 20414 26238 20466 26290
rect 20466 26238 20468 26290
rect 20412 26236 20468 26238
rect 19740 25788 19796 25844
rect 19516 25564 19572 25620
rect 19404 25506 19460 25508
rect 19404 25454 19406 25506
rect 19406 25454 19458 25506
rect 19458 25454 19460 25506
rect 19404 25452 19460 25454
rect 20188 25228 20244 25284
rect 19836 25114 19892 25116
rect 19836 25062 19838 25114
rect 19838 25062 19890 25114
rect 19890 25062 19892 25114
rect 19836 25060 19892 25062
rect 19940 25114 19996 25116
rect 19940 25062 19942 25114
rect 19942 25062 19994 25114
rect 19994 25062 19996 25114
rect 19940 25060 19996 25062
rect 20044 25114 20100 25116
rect 20044 25062 20046 25114
rect 20046 25062 20098 25114
rect 20098 25062 20100 25114
rect 20044 25060 20100 25062
rect 19068 23884 19124 23940
rect 18508 23212 18564 23268
rect 14924 22876 14980 22932
rect 14812 20748 14868 20804
rect 14924 22428 14980 22484
rect 15148 21980 15204 22036
rect 18396 22370 18452 22372
rect 18396 22318 18398 22370
rect 18398 22318 18450 22370
rect 18450 22318 18452 22370
rect 18396 22316 18452 22318
rect 17724 21644 17780 21700
rect 18172 21810 18228 21812
rect 18172 21758 18174 21810
rect 18174 21758 18226 21810
rect 18226 21758 18228 21810
rect 18172 21756 18228 21758
rect 15036 20076 15092 20132
rect 15372 19964 15428 20020
rect 15708 19906 15764 19908
rect 15708 19854 15710 19906
rect 15710 19854 15762 19906
rect 15762 19854 15764 19906
rect 15708 19852 15764 19854
rect 15708 19628 15764 19684
rect 14588 19346 14644 19348
rect 14588 19294 14590 19346
rect 14590 19294 14642 19346
rect 14642 19294 14644 19346
rect 14588 19292 14644 19294
rect 15484 19292 15540 19348
rect 13692 17276 13748 17332
rect 15036 19180 15092 19236
rect 12796 15874 12852 15876
rect 12796 15822 12798 15874
rect 12798 15822 12850 15874
rect 12850 15822 12852 15874
rect 12796 15820 12852 15822
rect 13692 15820 13748 15876
rect 15148 15986 15204 15988
rect 15148 15934 15150 15986
rect 15150 15934 15202 15986
rect 15202 15934 15204 15986
rect 15148 15932 15204 15934
rect 14476 15314 14532 15316
rect 14476 15262 14478 15314
rect 14478 15262 14530 15314
rect 14530 15262 14532 15314
rect 14476 15260 14532 15262
rect 11228 14476 11284 14532
rect 11900 14530 11956 14532
rect 11900 14478 11902 14530
rect 11902 14478 11954 14530
rect 11954 14478 11956 14530
rect 11900 14476 11956 14478
rect 4476 13354 4532 13356
rect 4476 13302 4478 13354
rect 4478 13302 4530 13354
rect 4530 13302 4532 13354
rect 4476 13300 4532 13302
rect 4580 13354 4636 13356
rect 4580 13302 4582 13354
rect 4582 13302 4634 13354
rect 4634 13302 4636 13354
rect 4580 13300 4636 13302
rect 4684 13354 4740 13356
rect 4684 13302 4686 13354
rect 4686 13302 4738 13354
rect 4738 13302 4740 13354
rect 4684 13300 4740 13302
rect 4476 11786 4532 11788
rect 4476 11734 4478 11786
rect 4478 11734 4530 11786
rect 4530 11734 4532 11786
rect 4476 11732 4532 11734
rect 4580 11786 4636 11788
rect 4580 11734 4582 11786
rect 4582 11734 4634 11786
rect 4634 11734 4636 11786
rect 4580 11732 4636 11734
rect 4684 11786 4740 11788
rect 4684 11734 4686 11786
rect 4686 11734 4738 11786
rect 4738 11734 4740 11786
rect 4684 11732 4740 11734
rect 4476 10218 4532 10220
rect 4476 10166 4478 10218
rect 4478 10166 4530 10218
rect 4530 10166 4532 10218
rect 4476 10164 4532 10166
rect 4580 10218 4636 10220
rect 4580 10166 4582 10218
rect 4582 10166 4634 10218
rect 4634 10166 4636 10218
rect 4580 10164 4636 10166
rect 4684 10218 4740 10220
rect 4684 10166 4686 10218
rect 4686 10166 4738 10218
rect 4738 10166 4740 10218
rect 4684 10164 4740 10166
rect 4476 8650 4532 8652
rect 4476 8598 4478 8650
rect 4478 8598 4530 8650
rect 4530 8598 4532 8650
rect 4476 8596 4532 8598
rect 4580 8650 4636 8652
rect 4580 8598 4582 8650
rect 4582 8598 4634 8650
rect 4634 8598 4636 8650
rect 4580 8596 4636 8598
rect 4684 8650 4740 8652
rect 4684 8598 4686 8650
rect 4686 8598 4738 8650
rect 4738 8598 4740 8650
rect 4684 8596 4740 8598
rect 16044 20636 16100 20692
rect 15596 18226 15652 18228
rect 15596 18174 15598 18226
rect 15598 18174 15650 18226
rect 15650 18174 15652 18226
rect 15596 18172 15652 18174
rect 16156 20802 16212 20804
rect 16156 20750 16158 20802
rect 16158 20750 16210 20802
rect 16210 20750 16212 20802
rect 16156 20748 16212 20750
rect 16044 20130 16100 20132
rect 16044 20078 16046 20130
rect 16046 20078 16098 20130
rect 16098 20078 16100 20130
rect 16044 20076 16100 20078
rect 16828 20860 16884 20916
rect 16716 20188 16772 20244
rect 16604 19964 16660 20020
rect 16604 19628 16660 19684
rect 16828 19458 16884 19460
rect 16828 19406 16830 19458
rect 16830 19406 16882 19458
rect 16882 19406 16884 19458
rect 16828 19404 16884 19406
rect 16940 19234 16996 19236
rect 16940 19182 16942 19234
rect 16942 19182 16994 19234
rect 16994 19182 16996 19234
rect 16940 19180 16996 19182
rect 16156 19068 16212 19124
rect 15932 18060 15988 18116
rect 16828 18956 16884 19012
rect 16268 18284 16324 18340
rect 16492 18450 16548 18452
rect 16492 18398 16494 18450
rect 16494 18398 16546 18450
rect 16546 18398 16548 18450
rect 16492 18396 16548 18398
rect 16380 18060 16436 18116
rect 16492 18172 16548 18228
rect 16492 17388 16548 17444
rect 16604 15932 16660 15988
rect 16380 15538 16436 15540
rect 16380 15486 16382 15538
rect 16382 15486 16434 15538
rect 16434 15486 16436 15538
rect 16380 15484 16436 15486
rect 4476 7082 4532 7084
rect 4476 7030 4478 7082
rect 4478 7030 4530 7082
rect 4530 7030 4532 7082
rect 4476 7028 4532 7030
rect 4580 7082 4636 7084
rect 4580 7030 4582 7082
rect 4582 7030 4634 7082
rect 4634 7030 4636 7082
rect 4580 7028 4636 7030
rect 4684 7082 4740 7084
rect 4684 7030 4686 7082
rect 4686 7030 4738 7082
rect 4738 7030 4740 7082
rect 4684 7028 4740 7030
rect 4476 5514 4532 5516
rect 4476 5462 4478 5514
rect 4478 5462 4530 5514
rect 4530 5462 4532 5514
rect 4476 5460 4532 5462
rect 4580 5514 4636 5516
rect 4580 5462 4582 5514
rect 4582 5462 4634 5514
rect 4634 5462 4636 5514
rect 4580 5460 4636 5462
rect 4684 5514 4740 5516
rect 4684 5462 4686 5514
rect 4686 5462 4738 5514
rect 4738 5462 4740 5514
rect 4684 5460 4740 5462
rect 4476 3946 4532 3948
rect 4476 3894 4478 3946
rect 4478 3894 4530 3946
rect 4530 3894 4532 3946
rect 4476 3892 4532 3894
rect 4580 3946 4636 3948
rect 4580 3894 4582 3946
rect 4582 3894 4634 3946
rect 4634 3894 4636 3946
rect 4580 3892 4636 3894
rect 4684 3946 4740 3948
rect 4684 3894 4686 3946
rect 4686 3894 4738 3946
rect 4738 3894 4740 3946
rect 4684 3892 4740 3894
rect 13468 3442 13524 3444
rect 13468 3390 13470 3442
rect 13470 3390 13522 3442
rect 13522 3390 13524 3442
rect 13468 3388 13524 3390
rect 17724 20860 17780 20916
rect 17612 20636 17668 20692
rect 17612 20076 17668 20132
rect 17388 19794 17444 19796
rect 17388 19742 17390 19794
rect 17390 19742 17442 19794
rect 17442 19742 17444 19794
rect 17388 19740 17444 19742
rect 17500 18956 17556 19012
rect 17388 18396 17444 18452
rect 17836 19628 17892 19684
rect 17724 19516 17780 19572
rect 20300 24444 20356 24500
rect 21308 36482 21364 36484
rect 21308 36430 21310 36482
rect 21310 36430 21362 36482
rect 21362 36430 21364 36482
rect 21308 36428 21364 36430
rect 21196 33516 21252 33572
rect 21420 35698 21476 35700
rect 21420 35646 21422 35698
rect 21422 35646 21474 35698
rect 21474 35646 21476 35698
rect 21420 35644 21476 35646
rect 21868 39116 21924 39172
rect 22764 40514 22820 40516
rect 22764 40462 22766 40514
rect 22766 40462 22818 40514
rect 22818 40462 22820 40514
rect 22764 40460 22820 40462
rect 23212 39730 23268 39732
rect 23212 39678 23214 39730
rect 23214 39678 23266 39730
rect 23266 39678 23268 39730
rect 23212 39676 23268 39678
rect 21756 38332 21812 38388
rect 22988 38332 23044 38388
rect 22092 38274 22148 38276
rect 22092 38222 22094 38274
rect 22094 38222 22146 38274
rect 22146 38222 22148 38274
rect 22092 38220 22148 38222
rect 21868 38108 21924 38164
rect 21644 37996 21700 38052
rect 23100 37996 23156 38052
rect 22092 37548 22148 37604
rect 21644 37154 21700 37156
rect 21644 37102 21646 37154
rect 21646 37102 21698 37154
rect 21698 37102 21700 37154
rect 21644 37100 21700 37102
rect 22204 37266 22260 37268
rect 22204 37214 22206 37266
rect 22206 37214 22258 37266
rect 22258 37214 22260 37266
rect 22204 37212 22260 37214
rect 23884 43538 23940 43540
rect 23884 43486 23886 43538
rect 23886 43486 23938 43538
rect 23938 43486 23940 43538
rect 23884 43484 23940 43486
rect 23772 42588 23828 42644
rect 24444 47234 24500 47236
rect 24444 47182 24446 47234
rect 24446 47182 24498 47234
rect 24498 47182 24500 47234
rect 24444 47180 24500 47182
rect 24444 45052 24500 45108
rect 24780 48412 24836 48468
rect 24892 52108 24948 52164
rect 24668 47852 24724 47908
rect 24780 48076 24836 48132
rect 25340 54908 25396 54964
rect 25564 55356 25620 55412
rect 25900 55132 25956 55188
rect 25452 54290 25508 54292
rect 25452 54238 25454 54290
rect 25454 54238 25506 54290
rect 25506 54238 25508 54290
rect 25452 54236 25508 54238
rect 25788 53452 25844 53508
rect 26236 59052 26292 59108
rect 26572 60956 26628 61012
rect 26572 60732 26628 60788
rect 26908 61346 26964 61348
rect 26908 61294 26910 61346
rect 26910 61294 26962 61346
rect 26962 61294 26964 61346
rect 26908 61292 26964 61294
rect 26796 60172 26852 60228
rect 26460 59388 26516 59444
rect 26908 60508 26964 60564
rect 27020 60284 27076 60340
rect 27468 61964 27524 62020
rect 27580 61852 27636 61908
rect 27916 61964 27972 62020
rect 28252 61740 28308 61796
rect 28476 62354 28532 62356
rect 28476 62302 28478 62354
rect 28478 62302 28530 62354
rect 28530 62302 28532 62354
rect 28476 62300 28532 62302
rect 28700 62076 28756 62132
rect 28812 63196 28868 63252
rect 28252 61292 28308 61348
rect 28476 61292 28532 61348
rect 27356 60674 27412 60676
rect 27356 60622 27358 60674
rect 27358 60622 27410 60674
rect 27410 60622 27412 60674
rect 27356 60620 27412 60622
rect 28252 60508 28308 60564
rect 28028 60226 28084 60228
rect 28028 60174 28030 60226
rect 28030 60174 28082 60226
rect 28082 60174 28084 60226
rect 28028 60172 28084 60174
rect 28700 60786 28756 60788
rect 28700 60734 28702 60786
rect 28702 60734 28754 60786
rect 28754 60734 28756 60786
rect 28700 60732 28756 60734
rect 28588 60674 28644 60676
rect 28588 60622 28590 60674
rect 28590 60622 28642 60674
rect 28642 60622 28644 60674
rect 28588 60620 28644 60622
rect 29372 65324 29428 65380
rect 29372 64706 29428 64708
rect 29372 64654 29374 64706
rect 29374 64654 29426 64706
rect 29426 64654 29428 64706
rect 29372 64652 29428 64654
rect 30044 67340 30100 67396
rect 30716 70082 30772 70084
rect 30716 70030 30718 70082
rect 30718 70030 30770 70082
rect 30770 70030 30772 70082
rect 30716 70028 30772 70030
rect 30380 69580 30436 69636
rect 31276 69634 31332 69636
rect 31276 69582 31278 69634
rect 31278 69582 31330 69634
rect 31330 69582 31332 69634
rect 31276 69580 31332 69582
rect 30380 67340 30436 67396
rect 30828 69186 30884 69188
rect 30828 69134 30830 69186
rect 30830 69134 30882 69186
rect 30882 69134 30884 69186
rect 30828 69132 30884 69134
rect 30604 67228 30660 67284
rect 30828 68908 30884 68964
rect 30156 67004 30212 67060
rect 30604 67058 30660 67060
rect 30604 67006 30606 67058
rect 30606 67006 30658 67058
rect 30658 67006 30660 67058
rect 30604 67004 30660 67006
rect 30044 66892 30100 66948
rect 30716 66892 30772 66948
rect 36428 70476 36484 70532
rect 31836 69298 31892 69300
rect 31836 69246 31838 69298
rect 31838 69246 31890 69298
rect 31890 69246 31892 69298
rect 31836 69244 31892 69246
rect 33292 69244 33348 69300
rect 31052 68572 31108 68628
rect 31164 67452 31220 67508
rect 31276 69132 31332 69188
rect 31612 69186 31668 69188
rect 31612 69134 31614 69186
rect 31614 69134 31666 69186
rect 31666 69134 31668 69186
rect 31612 69132 31668 69134
rect 33068 69020 33124 69076
rect 32844 68908 32900 68964
rect 32956 68626 33012 68628
rect 32956 68574 32958 68626
rect 32958 68574 33010 68626
rect 33010 68574 33012 68626
rect 32956 68572 33012 68574
rect 34412 69410 34468 69412
rect 34412 69358 34414 69410
rect 34414 69358 34466 69410
rect 34466 69358 34468 69410
rect 34412 69356 34468 69358
rect 34972 69298 35028 69300
rect 34972 69246 34974 69298
rect 34974 69246 35026 69298
rect 35026 69246 35028 69298
rect 34972 69244 35028 69246
rect 33964 69186 34020 69188
rect 33964 69134 33966 69186
rect 33966 69134 34018 69186
rect 34018 69134 34020 69186
rect 33964 69132 34020 69134
rect 34636 69186 34692 69188
rect 34636 69134 34638 69186
rect 34638 69134 34690 69186
rect 34690 69134 34692 69186
rect 34636 69132 34692 69134
rect 34188 69020 34244 69076
rect 33516 68850 33572 68852
rect 33516 68798 33518 68850
rect 33518 68798 33570 68850
rect 33570 68798 33572 68850
rect 33516 68796 33572 68798
rect 34972 68796 35028 68852
rect 35196 69802 35252 69804
rect 35196 69750 35198 69802
rect 35198 69750 35250 69802
rect 35250 69750 35252 69802
rect 35196 69748 35252 69750
rect 35300 69802 35356 69804
rect 35300 69750 35302 69802
rect 35302 69750 35354 69802
rect 35354 69750 35356 69802
rect 35300 69748 35356 69750
rect 35404 69802 35460 69804
rect 35404 69750 35406 69802
rect 35406 69750 35458 69802
rect 35458 69750 35460 69802
rect 35404 69748 35460 69750
rect 36428 69634 36484 69636
rect 36428 69582 36430 69634
rect 36430 69582 36482 69634
rect 36482 69582 36484 69634
rect 36428 69580 36484 69582
rect 36092 69356 36148 69412
rect 35084 68908 35140 68964
rect 34412 68738 34468 68740
rect 34412 68686 34414 68738
rect 34414 68686 34466 68738
rect 34466 68686 34468 68738
rect 34412 68684 34468 68686
rect 31500 68124 31556 68180
rect 32508 67116 32564 67172
rect 33068 67340 33124 67396
rect 32060 67004 32116 67060
rect 31052 66220 31108 66276
rect 30044 66050 30100 66052
rect 30044 65998 30046 66050
rect 30046 65998 30098 66050
rect 30098 65998 30100 66050
rect 30044 65996 30100 65998
rect 30156 65490 30212 65492
rect 30156 65438 30158 65490
rect 30158 65438 30210 65490
rect 30210 65438 30212 65490
rect 30156 65436 30212 65438
rect 30268 64652 30324 64708
rect 29484 64204 29540 64260
rect 29820 64316 29876 64372
rect 30156 64204 30212 64260
rect 30716 64316 30772 64372
rect 29372 64034 29428 64036
rect 29372 63982 29374 64034
rect 29374 63982 29426 64034
rect 29426 63982 29428 64034
rect 29372 63980 29428 63982
rect 29484 63810 29540 63812
rect 29484 63758 29486 63810
rect 29486 63758 29538 63810
rect 29538 63758 29540 63810
rect 29484 63756 29540 63758
rect 29484 62354 29540 62356
rect 29484 62302 29486 62354
rect 29486 62302 29538 62354
rect 29538 62302 29540 62354
rect 29484 62300 29540 62302
rect 29036 61740 29092 61796
rect 28924 61010 28980 61012
rect 28924 60958 28926 61010
rect 28926 60958 28978 61010
rect 28978 60958 28980 61010
rect 28924 60956 28980 60958
rect 29036 60508 29092 60564
rect 27132 59442 27188 59444
rect 27132 59390 27134 59442
rect 27134 59390 27186 59442
rect 27186 59390 27188 59442
rect 27132 59388 27188 59390
rect 26908 59276 26964 59332
rect 26684 58716 26740 58772
rect 26908 58434 26964 58436
rect 26908 58382 26910 58434
rect 26910 58382 26962 58434
rect 26962 58382 26964 58434
rect 26908 58380 26964 58382
rect 26124 57372 26180 57428
rect 26460 58156 26516 58212
rect 26572 57148 26628 57204
rect 26236 55356 26292 55412
rect 26124 54460 26180 54516
rect 26124 53900 26180 53956
rect 26012 53058 26068 53060
rect 26012 53006 26014 53058
rect 26014 53006 26066 53058
rect 26066 53006 26068 53058
rect 26012 53004 26068 53006
rect 25228 52780 25284 52836
rect 25340 52668 25396 52724
rect 25676 52556 25732 52612
rect 25116 51996 25172 52052
rect 25340 50316 25396 50372
rect 25228 49586 25284 49588
rect 25228 49534 25230 49586
rect 25230 49534 25282 49586
rect 25282 49534 25284 49586
rect 25228 49532 25284 49534
rect 27132 59218 27188 59220
rect 27132 59166 27134 59218
rect 27134 59166 27186 59218
rect 27186 59166 27188 59218
rect 27132 59164 27188 59166
rect 27692 59388 27748 59444
rect 27244 58716 27300 58772
rect 27804 59276 27860 59332
rect 27244 57538 27300 57540
rect 27244 57486 27246 57538
rect 27246 57486 27298 57538
rect 27298 57486 27300 57538
rect 27244 57484 27300 57486
rect 27356 55970 27412 55972
rect 27356 55918 27358 55970
rect 27358 55918 27410 55970
rect 27410 55918 27412 55970
rect 27356 55916 27412 55918
rect 26348 55298 26404 55300
rect 26348 55246 26350 55298
rect 26350 55246 26402 55298
rect 26402 55246 26404 55298
rect 26348 55244 26404 55246
rect 29260 61964 29316 62020
rect 29260 61458 29316 61460
rect 29260 61406 29262 61458
rect 29262 61406 29314 61458
rect 29314 61406 29316 61458
rect 29260 61404 29316 61406
rect 29596 61404 29652 61460
rect 30380 63980 30436 64036
rect 30044 62972 30100 63028
rect 30044 62188 30100 62244
rect 29932 61964 29988 62020
rect 29372 60732 29428 60788
rect 29148 59948 29204 60004
rect 27916 58716 27972 58772
rect 28028 58434 28084 58436
rect 28028 58382 28030 58434
rect 28030 58382 28082 58434
rect 28082 58382 28084 58434
rect 28028 58380 28084 58382
rect 29820 60732 29876 60788
rect 29596 60620 29652 60676
rect 30268 61964 30324 62020
rect 30716 62076 30772 62132
rect 31612 65996 31668 66052
rect 31164 63250 31220 63252
rect 31164 63198 31166 63250
rect 31166 63198 31218 63250
rect 31218 63198 31220 63250
rect 31164 63196 31220 63198
rect 31388 63980 31444 64036
rect 31164 62300 31220 62356
rect 31052 62188 31108 62244
rect 30828 61964 30884 62020
rect 30940 62076 30996 62132
rect 30604 61516 30660 61572
rect 30604 60956 30660 61012
rect 30156 60786 30212 60788
rect 30156 60734 30158 60786
rect 30158 60734 30210 60786
rect 30210 60734 30212 60786
rect 30156 60732 30212 60734
rect 28812 58380 28868 58436
rect 27916 57932 27972 57988
rect 28140 58322 28196 58324
rect 28140 58270 28142 58322
rect 28142 58270 28194 58322
rect 28194 58270 28196 58322
rect 28140 58268 28196 58270
rect 27804 55468 27860 55524
rect 28028 55916 28084 55972
rect 26460 54908 26516 54964
rect 26460 54738 26516 54740
rect 26460 54686 26462 54738
rect 26462 54686 26514 54738
rect 26514 54686 26516 54738
rect 26460 54684 26516 54686
rect 27244 55356 27300 55412
rect 26908 54460 26964 54516
rect 28252 58210 28308 58212
rect 28252 58158 28254 58210
rect 28254 58158 28306 58210
rect 28306 58158 28308 58210
rect 28252 58156 28308 58158
rect 28364 57820 28420 57876
rect 28588 57596 28644 57652
rect 31052 60732 31108 60788
rect 31052 60060 31108 60116
rect 30268 59052 30324 59108
rect 29820 58434 29876 58436
rect 29820 58382 29822 58434
rect 29822 58382 29874 58434
rect 29874 58382 29876 58434
rect 29820 58380 29876 58382
rect 30156 58434 30212 58436
rect 30156 58382 30158 58434
rect 30158 58382 30210 58434
rect 30210 58382 30212 58434
rect 30156 58380 30212 58382
rect 29932 58268 29988 58324
rect 31948 65490 32004 65492
rect 31948 65438 31950 65490
rect 31950 65438 32002 65490
rect 32002 65438 32004 65490
rect 31948 65436 32004 65438
rect 32620 65548 32676 65604
rect 32284 65436 32340 65492
rect 32508 65490 32564 65492
rect 32508 65438 32510 65490
rect 32510 65438 32562 65490
rect 32562 65438 32564 65490
rect 32508 65436 32564 65438
rect 32172 64428 32228 64484
rect 32396 64428 32452 64484
rect 31724 64204 31780 64260
rect 31948 64034 32004 64036
rect 31948 63982 31950 64034
rect 31950 63982 32002 64034
rect 32002 63982 32004 64034
rect 31948 63980 32004 63982
rect 31836 63868 31892 63924
rect 31612 62242 31668 62244
rect 31612 62190 31614 62242
rect 31614 62190 31666 62242
rect 31666 62190 31668 62242
rect 31612 62188 31668 62190
rect 32844 65324 32900 65380
rect 32396 62972 32452 63028
rect 32284 62242 32340 62244
rect 32284 62190 32286 62242
rect 32286 62190 32338 62242
rect 32338 62190 32340 62242
rect 32284 62188 32340 62190
rect 33404 67116 33460 67172
rect 33292 66050 33348 66052
rect 33292 65998 33294 66050
rect 33294 65998 33346 66050
rect 33346 65998 33348 66050
rect 33292 65996 33348 65998
rect 34748 66892 34804 66948
rect 34524 66444 34580 66500
rect 33404 65884 33460 65940
rect 33516 66050 33572 66052
rect 33516 65998 33518 66050
rect 33518 65998 33570 66050
rect 33570 65998 33572 66050
rect 33516 65996 33572 65998
rect 33404 65660 33460 65716
rect 33516 65548 33572 65604
rect 33740 65884 33796 65940
rect 33068 63868 33124 63924
rect 33628 65324 33684 65380
rect 33516 64146 33572 64148
rect 33516 64094 33518 64146
rect 33518 64094 33570 64146
rect 33570 64094 33572 64146
rect 33516 64092 33572 64094
rect 33628 64034 33684 64036
rect 33628 63982 33630 64034
rect 33630 63982 33682 64034
rect 33682 63982 33684 64034
rect 33628 63980 33684 63982
rect 33292 63922 33348 63924
rect 33292 63870 33294 63922
rect 33294 63870 33346 63922
rect 33346 63870 33348 63922
rect 33292 63868 33348 63870
rect 33068 62636 33124 62692
rect 32844 62188 32900 62244
rect 33180 62300 33236 62356
rect 32508 62076 32564 62132
rect 32732 61740 32788 61796
rect 31388 61570 31444 61572
rect 31388 61518 31390 61570
rect 31390 61518 31442 61570
rect 31442 61518 31444 61570
rect 31388 61516 31444 61518
rect 32172 61570 32228 61572
rect 32172 61518 32174 61570
rect 32174 61518 32226 61570
rect 32226 61518 32228 61570
rect 32172 61516 32228 61518
rect 31500 61458 31556 61460
rect 31500 61406 31502 61458
rect 31502 61406 31554 61458
rect 31554 61406 31556 61458
rect 31500 61404 31556 61406
rect 32508 61404 32564 61460
rect 31724 61180 31780 61236
rect 31500 61010 31556 61012
rect 31500 60958 31502 61010
rect 31502 60958 31554 61010
rect 31554 60958 31556 61010
rect 31500 60956 31556 60958
rect 30940 58546 30996 58548
rect 30940 58494 30942 58546
rect 30942 58494 30994 58546
rect 30994 58494 30996 58546
rect 30940 58492 30996 58494
rect 31500 58210 31556 58212
rect 31500 58158 31502 58210
rect 31502 58158 31554 58210
rect 31554 58158 31556 58210
rect 31500 58156 31556 58158
rect 29820 57484 29876 57540
rect 28588 55356 28644 55412
rect 28364 55132 28420 55188
rect 27916 55074 27972 55076
rect 27916 55022 27918 55074
rect 27918 55022 27970 55074
rect 27970 55022 27972 55074
rect 27916 55020 27972 55022
rect 27020 54796 27076 54852
rect 27916 54460 27972 54516
rect 27020 54348 27076 54404
rect 26684 53842 26740 53844
rect 26684 53790 26686 53842
rect 26686 53790 26738 53842
rect 26738 53790 26740 53842
rect 26684 53788 26740 53790
rect 27244 54124 27300 54180
rect 27132 53788 27188 53844
rect 26572 53506 26628 53508
rect 26572 53454 26574 53506
rect 26574 53454 26626 53506
rect 26626 53454 26628 53506
rect 26572 53452 26628 53454
rect 26684 53228 26740 53284
rect 26236 52668 26292 52724
rect 26348 52108 26404 52164
rect 26908 52892 26964 52948
rect 26460 52050 26516 52052
rect 26460 51998 26462 52050
rect 26462 51998 26514 52050
rect 26514 51998 26516 52050
rect 26460 51996 26516 51998
rect 26908 50652 26964 50708
rect 26236 50316 26292 50372
rect 26572 50370 26628 50372
rect 26572 50318 26574 50370
rect 26574 50318 26626 50370
rect 26626 50318 26628 50370
rect 26572 50316 26628 50318
rect 26348 49810 26404 49812
rect 26348 49758 26350 49810
rect 26350 49758 26402 49810
rect 26402 49758 26404 49810
rect 26348 49756 26404 49758
rect 25116 48076 25172 48132
rect 25228 47180 25284 47236
rect 25340 46674 25396 46676
rect 25340 46622 25342 46674
rect 25342 46622 25394 46674
rect 25394 46622 25396 46674
rect 25340 46620 25396 46622
rect 25788 46674 25844 46676
rect 25788 46622 25790 46674
rect 25790 46622 25842 46674
rect 25842 46622 25844 46674
rect 25788 46620 25844 46622
rect 25564 46508 25620 46564
rect 25228 46450 25284 46452
rect 25228 46398 25230 46450
rect 25230 46398 25282 46450
rect 25282 46398 25284 46450
rect 25228 46396 25284 46398
rect 24668 45276 24724 45332
rect 24892 45836 24948 45892
rect 24332 43708 24388 43764
rect 23884 42530 23940 42532
rect 23884 42478 23886 42530
rect 23886 42478 23938 42530
rect 23938 42478 23940 42530
rect 23884 42476 23940 42478
rect 23660 41916 23716 41972
rect 24332 42754 24388 42756
rect 24332 42702 24334 42754
rect 24334 42702 24386 42754
rect 24386 42702 24388 42754
rect 24332 42700 24388 42702
rect 23660 40908 23716 40964
rect 23436 40514 23492 40516
rect 23436 40462 23438 40514
rect 23438 40462 23490 40514
rect 23490 40462 23492 40514
rect 23436 40460 23492 40462
rect 23324 37996 23380 38052
rect 23324 37826 23380 37828
rect 23324 37774 23326 37826
rect 23326 37774 23378 37826
rect 23378 37774 23380 37826
rect 23324 37772 23380 37774
rect 22652 37266 22708 37268
rect 22652 37214 22654 37266
rect 22654 37214 22706 37266
rect 22706 37214 22708 37266
rect 22652 37212 22708 37214
rect 22540 37100 22596 37156
rect 22652 36540 22708 36596
rect 22428 36258 22484 36260
rect 22428 36206 22430 36258
rect 22430 36206 22482 36258
rect 22482 36206 22484 36258
rect 22428 36204 22484 36206
rect 21980 35644 22036 35700
rect 21868 35532 21924 35588
rect 22764 35644 22820 35700
rect 21756 34802 21812 34804
rect 21756 34750 21758 34802
rect 21758 34750 21810 34802
rect 21810 34750 21812 34802
rect 21756 34748 21812 34750
rect 21532 32620 21588 32676
rect 22652 33964 22708 34020
rect 21980 33458 22036 33460
rect 21980 33406 21982 33458
rect 21982 33406 22034 33458
rect 22034 33406 22036 33458
rect 21980 33404 22036 33406
rect 22428 33292 22484 33348
rect 23100 37100 23156 37156
rect 22988 35868 23044 35924
rect 23660 38892 23716 38948
rect 23660 38668 23716 38724
rect 23548 36540 23604 36596
rect 23548 35922 23604 35924
rect 23548 35870 23550 35922
rect 23550 35870 23602 35922
rect 23602 35870 23604 35922
rect 23548 35868 23604 35870
rect 23212 34972 23268 35028
rect 25788 46172 25844 46228
rect 25564 45276 25620 45332
rect 25340 45106 25396 45108
rect 25340 45054 25342 45106
rect 25342 45054 25394 45106
rect 25394 45054 25396 45106
rect 25340 45052 25396 45054
rect 25116 44492 25172 44548
rect 25116 43596 25172 43652
rect 25004 43148 25060 43204
rect 24556 42588 24612 42644
rect 24668 42476 24724 42532
rect 24556 42082 24612 42084
rect 24556 42030 24558 42082
rect 24558 42030 24610 42082
rect 24610 42030 24612 42082
rect 24556 42028 24612 42030
rect 24444 41804 24500 41860
rect 24780 42140 24836 42196
rect 24780 41468 24836 41524
rect 24444 41244 24500 41300
rect 23884 40626 23940 40628
rect 23884 40574 23886 40626
rect 23886 40574 23938 40626
rect 23938 40574 23940 40626
rect 23884 40572 23940 40574
rect 24332 40572 24388 40628
rect 24668 41020 24724 41076
rect 23884 40236 23940 40292
rect 24332 39676 24388 39732
rect 24668 39004 24724 39060
rect 24332 38780 24388 38836
rect 23884 38332 23940 38388
rect 24220 37996 24276 38052
rect 24108 37548 24164 37604
rect 24556 38722 24612 38724
rect 24556 38670 24558 38722
rect 24558 38670 24610 38722
rect 24610 38670 24612 38722
rect 24556 38668 24612 38670
rect 25004 41692 25060 41748
rect 26460 49138 26516 49140
rect 26460 49086 26462 49138
rect 26462 49086 26514 49138
rect 26514 49086 26516 49138
rect 26460 49084 26516 49086
rect 28364 54402 28420 54404
rect 28364 54350 28366 54402
rect 28366 54350 28418 54402
rect 28418 54350 28420 54402
rect 28364 54348 28420 54350
rect 27916 53842 27972 53844
rect 27916 53790 27918 53842
rect 27918 53790 27970 53842
rect 27970 53790 27972 53842
rect 27916 53788 27972 53790
rect 28028 53730 28084 53732
rect 28028 53678 28030 53730
rect 28030 53678 28082 53730
rect 28082 53678 28084 53730
rect 28028 53676 28084 53678
rect 27468 52946 27524 52948
rect 27468 52894 27470 52946
rect 27470 52894 27522 52946
rect 27522 52894 27524 52946
rect 27468 52892 27524 52894
rect 27916 52946 27972 52948
rect 27916 52894 27918 52946
rect 27918 52894 27970 52946
rect 27970 52894 27972 52946
rect 27916 52892 27972 52894
rect 27356 52834 27412 52836
rect 27356 52782 27358 52834
rect 27358 52782 27410 52834
rect 27410 52782 27412 52834
rect 27356 52780 27412 52782
rect 27244 52444 27300 52500
rect 27916 52444 27972 52500
rect 27244 52220 27300 52276
rect 26908 49756 26964 49812
rect 30156 57036 30212 57092
rect 29148 56924 29204 56980
rect 29148 55074 29204 55076
rect 29148 55022 29150 55074
rect 29150 55022 29202 55074
rect 29202 55022 29204 55074
rect 29148 55020 29204 55022
rect 29932 55356 29988 55412
rect 30044 55468 30100 55524
rect 29820 54908 29876 54964
rect 29148 54626 29204 54628
rect 29148 54574 29150 54626
rect 29150 54574 29202 54626
rect 29202 54574 29204 54626
rect 29148 54572 29204 54574
rect 28588 53900 28644 53956
rect 28252 53506 28308 53508
rect 28252 53454 28254 53506
rect 28254 53454 28306 53506
rect 28306 53454 28308 53506
rect 28252 53452 28308 53454
rect 28364 53170 28420 53172
rect 28364 53118 28366 53170
rect 28366 53118 28418 53170
rect 28418 53118 28420 53170
rect 28364 53116 28420 53118
rect 29036 53058 29092 53060
rect 29036 53006 29038 53058
rect 29038 53006 29090 53058
rect 29090 53006 29092 53058
rect 29036 53004 29092 53006
rect 28364 52722 28420 52724
rect 28364 52670 28366 52722
rect 28366 52670 28418 52722
rect 28418 52670 28420 52722
rect 28364 52668 28420 52670
rect 28252 52556 28308 52612
rect 28588 52274 28644 52276
rect 28588 52222 28590 52274
rect 28590 52222 28642 52274
rect 28642 52222 28644 52274
rect 28588 52220 28644 52222
rect 28812 52220 28868 52276
rect 29036 52668 29092 52724
rect 29932 54796 29988 54852
rect 29484 53676 29540 53732
rect 29148 52444 29204 52500
rect 29260 52892 29316 52948
rect 29148 52220 29204 52276
rect 28476 51996 28532 52052
rect 27468 50034 27524 50036
rect 27468 49982 27470 50034
rect 27470 49982 27522 50034
rect 27522 49982 27524 50034
rect 27468 49980 27524 49982
rect 28140 50034 28196 50036
rect 28140 49982 28142 50034
rect 28142 49982 28194 50034
rect 28194 49982 28196 50034
rect 28140 49980 28196 49982
rect 28252 50540 28308 50596
rect 27244 49810 27300 49812
rect 27244 49758 27246 49810
rect 27246 49758 27298 49810
rect 27298 49758 27300 49810
rect 27244 49756 27300 49758
rect 26684 49084 26740 49140
rect 26572 46956 26628 47012
rect 28700 49756 28756 49812
rect 26796 47404 26852 47460
rect 26908 48748 26964 48804
rect 26460 44098 26516 44100
rect 26460 44046 26462 44098
rect 26462 44046 26514 44098
rect 26514 44046 26516 44098
rect 26460 44044 26516 44046
rect 26348 43426 26404 43428
rect 26348 43374 26350 43426
rect 26350 43374 26402 43426
rect 26402 43374 26404 43426
rect 26348 43372 26404 43374
rect 26012 43148 26068 43204
rect 26348 43148 26404 43204
rect 25228 42642 25284 42644
rect 25228 42590 25230 42642
rect 25230 42590 25282 42642
rect 25282 42590 25284 42642
rect 25228 42588 25284 42590
rect 26012 42642 26068 42644
rect 26012 42590 26014 42642
rect 26014 42590 26066 42642
rect 26066 42590 26068 42642
rect 26012 42588 26068 42590
rect 26348 42530 26404 42532
rect 26348 42478 26350 42530
rect 26350 42478 26402 42530
rect 26402 42478 26404 42530
rect 26348 42476 26404 42478
rect 25228 42028 25284 42084
rect 25788 42252 25844 42308
rect 25116 41244 25172 41300
rect 25340 41804 25396 41860
rect 25116 40684 25172 40740
rect 25452 41692 25508 41748
rect 25452 41244 25508 41300
rect 25564 41020 25620 41076
rect 26796 43372 26852 43428
rect 26684 42588 26740 42644
rect 27244 48130 27300 48132
rect 27244 48078 27246 48130
rect 27246 48078 27298 48130
rect 27298 48078 27300 48130
rect 27244 48076 27300 48078
rect 27244 47740 27300 47796
rect 27132 46898 27188 46900
rect 27132 46846 27134 46898
rect 27134 46846 27186 46898
rect 27186 46846 27188 46898
rect 27132 46844 27188 46846
rect 27020 45724 27076 45780
rect 27132 44156 27188 44212
rect 27580 47292 27636 47348
rect 28028 47458 28084 47460
rect 28028 47406 28030 47458
rect 28030 47406 28082 47458
rect 28082 47406 28084 47458
rect 28028 47404 28084 47406
rect 28140 47292 28196 47348
rect 28252 47234 28308 47236
rect 28252 47182 28254 47234
rect 28254 47182 28306 47234
rect 28306 47182 28308 47234
rect 28252 47180 28308 47182
rect 27692 46898 27748 46900
rect 27692 46846 27694 46898
rect 27694 46846 27746 46898
rect 27746 46846 27748 46898
rect 27692 46844 27748 46846
rect 27580 46562 27636 46564
rect 27580 46510 27582 46562
rect 27582 46510 27634 46562
rect 27634 46510 27636 46562
rect 27580 46508 27636 46510
rect 28476 46956 28532 47012
rect 27916 46284 27972 46340
rect 27356 45724 27412 45780
rect 27468 44492 27524 44548
rect 28700 46844 28756 46900
rect 28700 46284 28756 46340
rect 28476 45778 28532 45780
rect 28476 45726 28478 45778
rect 28478 45726 28530 45778
rect 28530 45726 28532 45778
rect 28476 45724 28532 45726
rect 28700 45276 28756 45332
rect 28588 45218 28644 45220
rect 28588 45166 28590 45218
rect 28590 45166 28642 45218
rect 28642 45166 28644 45218
rect 28588 45164 28644 45166
rect 28364 44940 28420 44996
rect 26908 42476 26964 42532
rect 25452 40908 25508 40964
rect 25116 40236 25172 40292
rect 25452 40460 25508 40516
rect 25788 40514 25844 40516
rect 25788 40462 25790 40514
rect 25790 40462 25842 40514
rect 25842 40462 25844 40514
rect 25788 40460 25844 40462
rect 25452 39058 25508 39060
rect 25452 39006 25454 39058
rect 25454 39006 25506 39058
rect 25506 39006 25508 39058
rect 25452 39004 25508 39006
rect 25564 39340 25620 39396
rect 25004 37938 25060 37940
rect 25004 37886 25006 37938
rect 25006 37886 25058 37938
rect 25058 37886 25060 37938
rect 25004 37884 25060 37886
rect 24444 37436 24500 37492
rect 23996 35922 24052 35924
rect 23996 35870 23998 35922
rect 23998 35870 24050 35922
rect 24050 35870 24052 35922
rect 23996 35868 24052 35870
rect 24668 37266 24724 37268
rect 24668 37214 24670 37266
rect 24670 37214 24722 37266
rect 24722 37214 24724 37266
rect 24668 37212 24724 37214
rect 24892 36258 24948 36260
rect 24892 36206 24894 36258
rect 24894 36206 24946 36258
rect 24946 36206 24948 36258
rect 24892 36204 24948 36206
rect 24892 35308 24948 35364
rect 24556 35084 24612 35140
rect 25452 37266 25508 37268
rect 25452 37214 25454 37266
rect 25454 37214 25506 37266
rect 25506 37214 25508 37266
rect 25452 37212 25508 37214
rect 25340 37100 25396 37156
rect 25676 37100 25732 37156
rect 25788 37212 25844 37268
rect 25228 36204 25284 36260
rect 27244 42082 27300 42084
rect 27244 42030 27246 42082
rect 27246 42030 27298 42082
rect 27298 42030 27300 42082
rect 27244 42028 27300 42030
rect 27132 41916 27188 41972
rect 26460 41132 26516 41188
rect 26124 40962 26180 40964
rect 26124 40910 26126 40962
rect 26126 40910 26178 40962
rect 26178 40910 26180 40962
rect 26124 40908 26180 40910
rect 26012 40684 26068 40740
rect 26460 40402 26516 40404
rect 26460 40350 26462 40402
rect 26462 40350 26514 40402
rect 26514 40350 26516 40402
rect 26460 40348 26516 40350
rect 26236 37884 26292 37940
rect 26124 37490 26180 37492
rect 26124 37438 26126 37490
rect 26126 37438 26178 37490
rect 26178 37438 26180 37490
rect 26124 37436 26180 37438
rect 26348 36540 26404 36596
rect 26460 36652 26516 36708
rect 26460 35980 26516 36036
rect 26012 35922 26068 35924
rect 26012 35870 26014 35922
rect 26014 35870 26066 35922
rect 26066 35870 26068 35922
rect 26012 35868 26068 35870
rect 25228 34412 25284 34468
rect 23660 34130 23716 34132
rect 23660 34078 23662 34130
rect 23662 34078 23714 34130
rect 23714 34078 23716 34130
rect 23660 34076 23716 34078
rect 23212 34018 23268 34020
rect 23212 33966 23214 34018
rect 23214 33966 23266 34018
rect 23266 33966 23268 34018
rect 23212 33964 23268 33966
rect 22876 33292 22932 33348
rect 21980 32620 22036 32676
rect 22540 32674 22596 32676
rect 22540 32622 22542 32674
rect 22542 32622 22594 32674
rect 22594 32622 22596 32674
rect 22540 32620 22596 32622
rect 21308 32172 21364 32228
rect 21532 30828 21588 30884
rect 23100 33068 23156 33124
rect 22764 32172 22820 32228
rect 22540 31500 22596 31556
rect 21756 30156 21812 30212
rect 21868 29820 21924 29876
rect 21756 29596 21812 29652
rect 21084 28140 21140 28196
rect 20748 27356 20804 27412
rect 20636 26124 20692 26180
rect 20860 27186 20916 27188
rect 20860 27134 20862 27186
rect 20862 27134 20914 27186
rect 20914 27134 20916 27186
rect 20860 27132 20916 27134
rect 20972 26066 21028 26068
rect 20972 26014 20974 26066
rect 20974 26014 21026 26066
rect 21026 26014 21028 26066
rect 20972 26012 21028 26014
rect 20748 24444 20804 24500
rect 21308 26962 21364 26964
rect 21308 26910 21310 26962
rect 21310 26910 21362 26962
rect 21362 26910 21364 26962
rect 21308 26908 21364 26910
rect 21868 28642 21924 28644
rect 21868 28590 21870 28642
rect 21870 28590 21922 28642
rect 21922 28590 21924 28642
rect 21868 28588 21924 28590
rect 22316 30210 22372 30212
rect 22316 30158 22318 30210
rect 22318 30158 22370 30210
rect 22370 30158 22372 30210
rect 22316 30156 22372 30158
rect 22204 29932 22260 29988
rect 22092 29036 22148 29092
rect 21980 28364 22036 28420
rect 21532 27916 21588 27972
rect 21644 27580 21700 27636
rect 21980 27468 22036 27524
rect 21532 26348 21588 26404
rect 21644 26290 21700 26292
rect 21644 26238 21646 26290
rect 21646 26238 21698 26290
rect 21698 26238 21700 26290
rect 21644 26236 21700 26238
rect 21644 25564 21700 25620
rect 21532 25228 21588 25284
rect 21420 24668 21476 24724
rect 19836 23546 19892 23548
rect 19836 23494 19838 23546
rect 19838 23494 19890 23546
rect 19890 23494 19892 23546
rect 19836 23492 19892 23494
rect 19940 23546 19996 23548
rect 19940 23494 19942 23546
rect 19942 23494 19994 23546
rect 19994 23494 19996 23546
rect 19940 23492 19996 23494
rect 20044 23546 20100 23548
rect 20044 23494 20046 23546
rect 20046 23494 20098 23546
rect 20098 23494 20100 23546
rect 20300 23548 20356 23604
rect 20044 23492 20100 23494
rect 19068 21756 19124 21812
rect 20300 23100 20356 23156
rect 19628 22764 19684 22820
rect 19516 21644 19572 21700
rect 19836 21978 19892 21980
rect 19836 21926 19838 21978
rect 19838 21926 19890 21978
rect 19890 21926 19892 21978
rect 19836 21924 19892 21926
rect 19940 21978 19996 21980
rect 19940 21926 19942 21978
rect 19942 21926 19994 21978
rect 19994 21926 19996 21978
rect 19940 21924 19996 21926
rect 20044 21978 20100 21980
rect 20044 21926 20046 21978
rect 20046 21926 20098 21978
rect 20098 21926 20100 21978
rect 20044 21924 20100 21926
rect 20524 22764 20580 22820
rect 20636 23548 20692 23604
rect 21644 23436 21700 23492
rect 20972 23266 21028 23268
rect 20972 23214 20974 23266
rect 20974 23214 21026 23266
rect 21026 23214 21028 23266
rect 20972 23212 21028 23214
rect 19292 20188 19348 20244
rect 17948 19292 18004 19348
rect 18620 19852 18676 19908
rect 18060 18338 18116 18340
rect 18060 18286 18062 18338
rect 18062 18286 18114 18338
rect 18114 18286 18116 18338
rect 18060 18284 18116 18286
rect 17724 17724 17780 17780
rect 17948 17836 18004 17892
rect 17500 16828 17556 16884
rect 17276 16268 17332 16324
rect 17836 15260 17892 15316
rect 18060 17666 18116 17668
rect 18060 17614 18062 17666
rect 18062 17614 18114 17666
rect 18114 17614 18116 17666
rect 18060 17612 18116 17614
rect 18284 18284 18340 18340
rect 18284 16828 18340 16884
rect 18620 17388 18676 17444
rect 18620 16210 18676 16212
rect 18620 16158 18622 16210
rect 18622 16158 18674 16210
rect 18674 16158 18676 16210
rect 18620 16156 18676 16158
rect 18508 15260 18564 15316
rect 16380 3388 16436 3444
rect 17724 3388 17780 3444
rect 18956 17836 19012 17892
rect 18956 16268 19012 16324
rect 18956 15596 19012 15652
rect 19068 15484 19124 15540
rect 19292 18284 19348 18340
rect 19292 17612 19348 17668
rect 18396 11452 18452 11508
rect 18732 11394 18788 11396
rect 18732 11342 18734 11394
rect 18734 11342 18786 11394
rect 18786 11342 18788 11394
rect 18732 11340 18788 11342
rect 19292 14252 19348 14308
rect 20412 21420 20468 21476
rect 19836 20410 19892 20412
rect 19836 20358 19838 20410
rect 19838 20358 19890 20410
rect 19890 20358 19892 20410
rect 19836 20356 19892 20358
rect 19940 20410 19996 20412
rect 19940 20358 19942 20410
rect 19942 20358 19994 20410
rect 19994 20358 19996 20410
rect 19940 20356 19996 20358
rect 20044 20410 20100 20412
rect 20044 20358 20046 20410
rect 20046 20358 20098 20410
rect 20098 20358 20100 20410
rect 20044 20356 20100 20358
rect 19628 20076 19684 20132
rect 19516 19964 19572 20020
rect 19964 20018 20020 20020
rect 19964 19966 19966 20018
rect 19966 19966 20018 20018
rect 20018 19966 20020 20018
rect 19964 19964 20020 19966
rect 19852 19346 19908 19348
rect 19852 19294 19854 19346
rect 19854 19294 19906 19346
rect 19906 19294 19908 19346
rect 19852 19292 19908 19294
rect 19836 18842 19892 18844
rect 19836 18790 19838 18842
rect 19838 18790 19890 18842
rect 19890 18790 19892 18842
rect 19836 18788 19892 18790
rect 19940 18842 19996 18844
rect 19940 18790 19942 18842
rect 19942 18790 19994 18842
rect 19994 18790 19996 18842
rect 19940 18788 19996 18790
rect 20044 18842 20100 18844
rect 20044 18790 20046 18842
rect 20046 18790 20098 18842
rect 20098 18790 20100 18842
rect 20044 18788 20100 18790
rect 19740 18396 19796 18452
rect 20076 17778 20132 17780
rect 20076 17726 20078 17778
rect 20078 17726 20130 17778
rect 20130 17726 20132 17778
rect 20076 17724 20132 17726
rect 20188 17612 20244 17668
rect 20188 17388 20244 17444
rect 19836 17274 19892 17276
rect 19836 17222 19838 17274
rect 19838 17222 19890 17274
rect 19890 17222 19892 17274
rect 19836 17220 19892 17222
rect 19940 17274 19996 17276
rect 19940 17222 19942 17274
rect 19942 17222 19994 17274
rect 19994 17222 19996 17274
rect 19940 17220 19996 17222
rect 20044 17274 20100 17276
rect 20044 17222 20046 17274
rect 20046 17222 20098 17274
rect 20098 17222 20100 17274
rect 20044 17220 20100 17222
rect 19516 16156 19572 16212
rect 19836 15706 19892 15708
rect 19628 15596 19684 15652
rect 19836 15654 19838 15706
rect 19838 15654 19890 15706
rect 19890 15654 19892 15706
rect 19836 15652 19892 15654
rect 19940 15706 19996 15708
rect 19940 15654 19942 15706
rect 19942 15654 19994 15706
rect 19994 15654 19996 15706
rect 19940 15652 19996 15654
rect 20044 15706 20100 15708
rect 20044 15654 20046 15706
rect 20046 15654 20098 15706
rect 20098 15654 20100 15706
rect 20044 15652 20100 15654
rect 20412 19964 20468 20020
rect 21868 25116 21924 25172
rect 21868 24556 21924 24612
rect 22540 30210 22596 30212
rect 22540 30158 22542 30210
rect 22542 30158 22594 30210
rect 22594 30158 22596 30210
rect 22540 30156 22596 30158
rect 22876 31276 22932 31332
rect 24444 34130 24500 34132
rect 24444 34078 24446 34130
rect 24446 34078 24498 34130
rect 24498 34078 24500 34130
rect 24444 34076 24500 34078
rect 24668 33964 24724 34020
rect 24780 34076 24836 34132
rect 24220 32732 24276 32788
rect 25452 34130 25508 34132
rect 25452 34078 25454 34130
rect 25454 34078 25506 34130
rect 25506 34078 25508 34130
rect 25452 34076 25508 34078
rect 25676 34130 25732 34132
rect 25676 34078 25678 34130
rect 25678 34078 25730 34130
rect 25730 34078 25732 34130
rect 25676 34076 25732 34078
rect 25228 33740 25284 33796
rect 24892 33180 24948 33236
rect 24444 32562 24500 32564
rect 24444 32510 24446 32562
rect 24446 32510 24498 32562
rect 24498 32510 24500 32562
rect 24444 32508 24500 32510
rect 23436 32172 23492 32228
rect 22988 31052 23044 31108
rect 23100 31890 23156 31892
rect 23100 31838 23102 31890
rect 23102 31838 23154 31890
rect 23154 31838 23156 31890
rect 23100 31836 23156 31838
rect 22540 29820 22596 29876
rect 22652 29148 22708 29204
rect 22204 28364 22260 28420
rect 22092 24892 22148 24948
rect 22540 28082 22596 28084
rect 22540 28030 22542 28082
rect 22542 28030 22594 28082
rect 22594 28030 22596 28082
rect 22540 28028 22596 28030
rect 22204 27132 22260 27188
rect 22428 27746 22484 27748
rect 22428 27694 22430 27746
rect 22430 27694 22482 27746
rect 22482 27694 22484 27746
rect 22428 27692 22484 27694
rect 22540 27580 22596 27636
rect 22428 27468 22484 27524
rect 22652 27186 22708 27188
rect 22652 27134 22654 27186
rect 22654 27134 22706 27186
rect 22706 27134 22708 27186
rect 22652 27132 22708 27134
rect 22316 26236 22372 26292
rect 22428 26796 22484 26852
rect 21868 23324 21924 23380
rect 22204 23378 22260 23380
rect 22204 23326 22206 23378
rect 22206 23326 22258 23378
rect 22258 23326 22260 23378
rect 22204 23324 22260 23326
rect 21420 22316 21476 22372
rect 20860 20076 20916 20132
rect 21868 21644 21924 21700
rect 20748 19122 20804 19124
rect 20748 19070 20750 19122
rect 20750 19070 20802 19122
rect 20802 19070 20804 19122
rect 20748 19068 20804 19070
rect 20748 18396 20804 18452
rect 19836 14138 19892 14140
rect 19836 14086 19838 14138
rect 19838 14086 19890 14138
rect 19890 14086 19892 14138
rect 19836 14084 19892 14086
rect 19940 14138 19996 14140
rect 19940 14086 19942 14138
rect 19942 14086 19994 14138
rect 19994 14086 19996 14138
rect 19940 14084 19996 14086
rect 20044 14138 20100 14140
rect 20044 14086 20046 14138
rect 20046 14086 20098 14138
rect 20098 14086 20100 14138
rect 20044 14084 20100 14086
rect 20748 13074 20804 13076
rect 20748 13022 20750 13074
rect 20750 13022 20802 13074
rect 20802 13022 20804 13074
rect 20748 13020 20804 13022
rect 19836 12570 19892 12572
rect 19836 12518 19838 12570
rect 19838 12518 19890 12570
rect 19890 12518 19892 12570
rect 19836 12516 19892 12518
rect 19940 12570 19996 12572
rect 19940 12518 19942 12570
rect 19942 12518 19994 12570
rect 19994 12518 19996 12570
rect 19940 12516 19996 12518
rect 20044 12570 20100 12572
rect 20044 12518 20046 12570
rect 20046 12518 20098 12570
rect 20098 12518 20100 12570
rect 20044 12516 20100 12518
rect 19964 12402 20020 12404
rect 19964 12350 19966 12402
rect 19966 12350 20018 12402
rect 20018 12350 20020 12402
rect 19964 12348 20020 12350
rect 21420 19964 21476 20020
rect 21084 18450 21140 18452
rect 21084 18398 21086 18450
rect 21086 18398 21138 18450
rect 21138 18398 21140 18450
rect 21084 18396 21140 18398
rect 21868 20018 21924 20020
rect 21868 19966 21870 20018
rect 21870 19966 21922 20018
rect 21922 19966 21924 20018
rect 21868 19964 21924 19966
rect 21756 19292 21812 19348
rect 21868 19180 21924 19236
rect 21532 18060 21588 18116
rect 21868 16156 21924 16212
rect 23212 30882 23268 30884
rect 23212 30830 23214 30882
rect 23214 30830 23266 30882
rect 23266 30830 23268 30882
rect 23212 30828 23268 30830
rect 23212 29932 23268 29988
rect 24220 31948 24276 32004
rect 23996 31836 24052 31892
rect 23548 31276 23604 31332
rect 23996 31276 24052 31332
rect 24556 31388 24612 31444
rect 23772 30940 23828 30996
rect 24444 30994 24500 30996
rect 24444 30942 24446 30994
rect 24446 30942 24498 30994
rect 24498 30942 24500 30994
rect 24444 30940 24500 30942
rect 24108 30156 24164 30212
rect 23772 29932 23828 29988
rect 24892 32620 24948 32676
rect 24668 30492 24724 30548
rect 24556 29932 24612 29988
rect 25788 33964 25844 34020
rect 25116 32786 25172 32788
rect 25116 32734 25118 32786
rect 25118 32734 25170 32786
rect 25170 32734 25172 32786
rect 25116 32732 25172 32734
rect 25788 32732 25844 32788
rect 25452 32562 25508 32564
rect 25452 32510 25454 32562
rect 25454 32510 25506 32562
rect 25506 32510 25508 32562
rect 25452 32508 25508 32510
rect 25340 31948 25396 32004
rect 26012 32450 26068 32452
rect 26012 32398 26014 32450
rect 26014 32398 26066 32450
rect 26066 32398 26068 32450
rect 26012 32396 26068 32398
rect 26012 31948 26068 32004
rect 25676 31724 25732 31780
rect 25900 31724 25956 31780
rect 25228 31276 25284 31332
rect 23436 29036 23492 29092
rect 23100 28476 23156 28532
rect 23212 28700 23268 28756
rect 24444 29148 24500 29204
rect 24108 28700 24164 28756
rect 23996 28642 24052 28644
rect 23996 28590 23998 28642
rect 23998 28590 24050 28642
rect 24050 28590 24052 28642
rect 23996 28588 24052 28590
rect 23436 28530 23492 28532
rect 23436 28478 23438 28530
rect 23438 28478 23490 28530
rect 23490 28478 23492 28530
rect 23436 28476 23492 28478
rect 24780 29426 24836 29428
rect 24780 29374 24782 29426
rect 24782 29374 24834 29426
rect 24834 29374 24836 29426
rect 24780 29372 24836 29374
rect 24668 29260 24724 29316
rect 23324 28082 23380 28084
rect 23324 28030 23326 28082
rect 23326 28030 23378 28082
rect 23378 28030 23380 28082
rect 23324 28028 23380 28030
rect 24668 28082 24724 28084
rect 24668 28030 24670 28082
rect 24670 28030 24722 28082
rect 24722 28030 24724 28082
rect 24668 28028 24724 28030
rect 23548 27916 23604 27972
rect 22988 27858 23044 27860
rect 22988 27806 22990 27858
rect 22990 27806 23042 27858
rect 23042 27806 23044 27858
rect 22988 27804 23044 27806
rect 23212 27634 23268 27636
rect 23212 27582 23214 27634
rect 23214 27582 23266 27634
rect 23266 27582 23268 27634
rect 23212 27580 23268 27582
rect 23324 27356 23380 27412
rect 23436 27244 23492 27300
rect 23548 27020 23604 27076
rect 23996 27244 24052 27300
rect 24220 27244 24276 27300
rect 24108 27132 24164 27188
rect 24220 27074 24276 27076
rect 24220 27022 24222 27074
rect 24222 27022 24274 27074
rect 24274 27022 24276 27074
rect 24220 27020 24276 27022
rect 24108 26908 24164 26964
rect 23324 26348 23380 26404
rect 23436 26460 23492 26516
rect 23660 26460 23716 26516
rect 23100 25788 23156 25844
rect 23884 26850 23940 26852
rect 23884 26798 23886 26850
rect 23886 26798 23938 26850
rect 23938 26798 23940 26850
rect 23884 26796 23940 26798
rect 24556 26962 24612 26964
rect 24556 26910 24558 26962
rect 24558 26910 24610 26962
rect 24610 26910 24612 26962
rect 24556 26908 24612 26910
rect 24220 26290 24276 26292
rect 24220 26238 24222 26290
rect 24222 26238 24274 26290
rect 24274 26238 24276 26290
rect 24220 26236 24276 26238
rect 22764 25116 22820 25172
rect 22652 24444 22708 24500
rect 22652 23266 22708 23268
rect 22652 23214 22654 23266
rect 22654 23214 22706 23266
rect 22706 23214 22708 23266
rect 22652 23212 22708 23214
rect 22540 23100 22596 23156
rect 22988 23996 23044 24052
rect 22988 23324 23044 23380
rect 22764 22316 22820 22372
rect 22876 22988 22932 23044
rect 23212 22652 23268 22708
rect 23100 21810 23156 21812
rect 23100 21758 23102 21810
rect 23102 21758 23154 21810
rect 23154 21758 23156 21810
rect 23100 21756 23156 21758
rect 22316 21474 22372 21476
rect 22316 21422 22318 21474
rect 22318 21422 22370 21474
rect 22370 21422 22372 21474
rect 22316 21420 22372 21422
rect 22540 20860 22596 20916
rect 23660 24050 23716 24052
rect 23660 23998 23662 24050
rect 23662 23998 23714 24050
rect 23714 23998 23716 24050
rect 23660 23996 23716 23998
rect 23548 23154 23604 23156
rect 23548 23102 23550 23154
rect 23550 23102 23602 23154
rect 23602 23102 23604 23154
rect 23548 23100 23604 23102
rect 23884 24834 23940 24836
rect 23884 24782 23886 24834
rect 23886 24782 23938 24834
rect 23938 24782 23940 24834
rect 23884 24780 23940 24782
rect 24444 25788 24500 25844
rect 24332 25564 24388 25620
rect 24556 24946 24612 24948
rect 24556 24894 24558 24946
rect 24558 24894 24610 24946
rect 24610 24894 24612 24946
rect 24556 24892 24612 24894
rect 24780 26460 24836 26516
rect 23884 24444 23940 24500
rect 23772 22988 23828 23044
rect 23324 21644 23380 21700
rect 23436 22428 23492 22484
rect 23548 21586 23604 21588
rect 23548 21534 23550 21586
rect 23550 21534 23602 21586
rect 23602 21534 23604 21586
rect 23548 21532 23604 21534
rect 23324 20860 23380 20916
rect 22204 19068 22260 19124
rect 22092 18956 22148 19012
rect 22428 19122 22484 19124
rect 22428 19070 22430 19122
rect 22430 19070 22482 19122
rect 22482 19070 22484 19122
rect 22428 19068 22484 19070
rect 22876 19010 22932 19012
rect 22876 18958 22878 19010
rect 22878 18958 22930 19010
rect 22930 18958 22932 19010
rect 22876 18956 22932 18958
rect 22540 18508 22596 18564
rect 23100 18508 23156 18564
rect 22764 18284 22820 18340
rect 22204 18060 22260 18116
rect 22204 16716 22260 16772
rect 22652 16156 22708 16212
rect 22652 15596 22708 15652
rect 21308 14306 21364 14308
rect 21308 14254 21310 14306
rect 21310 14254 21362 14306
rect 21362 14254 21364 14306
rect 21308 14252 21364 14254
rect 21420 13634 21476 13636
rect 21420 13582 21422 13634
rect 21422 13582 21474 13634
rect 21474 13582 21476 13634
rect 21420 13580 21476 13582
rect 21532 13132 21588 13188
rect 20860 12348 20916 12404
rect 19404 12124 19460 12180
rect 19516 12236 19572 12292
rect 20300 12178 20356 12180
rect 20300 12126 20302 12178
rect 20302 12126 20354 12178
rect 20354 12126 20356 12178
rect 20300 12124 20356 12126
rect 21756 12908 21812 12964
rect 20972 11788 21028 11844
rect 20300 11340 20356 11396
rect 19852 11116 19908 11172
rect 19836 11002 19892 11004
rect 19836 10950 19838 11002
rect 19838 10950 19890 11002
rect 19890 10950 19892 11002
rect 19836 10948 19892 10950
rect 19940 11002 19996 11004
rect 19940 10950 19942 11002
rect 19942 10950 19994 11002
rect 19994 10950 19996 11002
rect 19940 10948 19996 10950
rect 20044 11002 20100 11004
rect 20044 10950 20046 11002
rect 20046 10950 20098 11002
rect 20098 10950 20100 11002
rect 20044 10948 20100 10950
rect 19836 9434 19892 9436
rect 19836 9382 19838 9434
rect 19838 9382 19890 9434
rect 19890 9382 19892 9434
rect 19836 9380 19892 9382
rect 19940 9434 19996 9436
rect 19940 9382 19942 9434
rect 19942 9382 19994 9434
rect 19994 9382 19996 9434
rect 19940 9380 19996 9382
rect 20044 9434 20100 9436
rect 20044 9382 20046 9434
rect 20046 9382 20098 9434
rect 20098 9382 20100 9434
rect 20044 9380 20100 9382
rect 19628 9100 19684 9156
rect 20524 8876 20580 8932
rect 19836 7866 19892 7868
rect 19836 7814 19838 7866
rect 19838 7814 19890 7866
rect 19890 7814 19892 7866
rect 19836 7812 19892 7814
rect 19940 7866 19996 7868
rect 19940 7814 19942 7866
rect 19942 7814 19994 7866
rect 19994 7814 19996 7866
rect 19940 7812 19996 7814
rect 20044 7866 20100 7868
rect 20044 7814 20046 7866
rect 20046 7814 20098 7866
rect 20098 7814 20100 7866
rect 20044 7812 20100 7814
rect 19836 6298 19892 6300
rect 19836 6246 19838 6298
rect 19838 6246 19890 6298
rect 19890 6246 19892 6298
rect 19836 6244 19892 6246
rect 19940 6298 19996 6300
rect 19940 6246 19942 6298
rect 19942 6246 19994 6298
rect 19994 6246 19996 6298
rect 19940 6244 19996 6246
rect 20044 6298 20100 6300
rect 20044 6246 20046 6298
rect 20046 6246 20098 6298
rect 20098 6246 20100 6298
rect 20044 6244 20100 6246
rect 19836 4730 19892 4732
rect 19836 4678 19838 4730
rect 19838 4678 19890 4730
rect 19890 4678 19892 4730
rect 19836 4676 19892 4678
rect 19940 4730 19996 4732
rect 19940 4678 19942 4730
rect 19942 4678 19994 4730
rect 19994 4678 19996 4730
rect 19940 4676 19996 4678
rect 20044 4730 20100 4732
rect 20044 4678 20046 4730
rect 20046 4678 20098 4730
rect 20098 4678 20100 4730
rect 20044 4676 20100 4678
rect 19180 3442 19236 3444
rect 19180 3390 19182 3442
rect 19182 3390 19234 3442
rect 19234 3390 19236 3442
rect 19180 3388 19236 3390
rect 19852 3442 19908 3444
rect 19852 3390 19854 3442
rect 19854 3390 19906 3442
rect 19906 3390 19908 3442
rect 19852 3388 19908 3390
rect 20188 3442 20244 3444
rect 20188 3390 20190 3442
rect 20190 3390 20242 3442
rect 20242 3390 20244 3442
rect 20188 3388 20244 3390
rect 19836 3162 19892 3164
rect 19836 3110 19838 3162
rect 19838 3110 19890 3162
rect 19890 3110 19892 3162
rect 19836 3108 19892 3110
rect 19940 3162 19996 3164
rect 19940 3110 19942 3162
rect 19942 3110 19994 3162
rect 19994 3110 19996 3162
rect 19940 3108 19996 3110
rect 20044 3162 20100 3164
rect 20044 3110 20046 3162
rect 20046 3110 20098 3162
rect 20098 3110 20100 3162
rect 20044 3108 20100 3110
rect 22092 13132 22148 13188
rect 21644 12124 21700 12180
rect 22540 14252 22596 14308
rect 22652 13580 22708 13636
rect 22316 12796 22372 12852
rect 22540 13020 22596 13076
rect 21980 11788 22036 11844
rect 21868 11228 21924 11284
rect 22988 15538 23044 15540
rect 22988 15486 22990 15538
rect 22990 15486 23042 15538
rect 23042 15486 23044 15538
rect 22988 15484 23044 15486
rect 24444 23826 24500 23828
rect 24444 23774 24446 23826
rect 24446 23774 24498 23826
rect 24498 23774 24500 23826
rect 24444 23772 24500 23774
rect 24556 23212 24612 23268
rect 24556 22540 24612 22596
rect 24332 22428 24388 22484
rect 24892 21868 24948 21924
rect 25452 31554 25508 31556
rect 25452 31502 25454 31554
rect 25454 31502 25506 31554
rect 25506 31502 25508 31554
rect 25452 31500 25508 31502
rect 25676 31554 25732 31556
rect 25676 31502 25678 31554
rect 25678 31502 25730 31554
rect 25730 31502 25732 31554
rect 25676 31500 25732 31502
rect 25340 30604 25396 30660
rect 25788 31276 25844 31332
rect 25788 30380 25844 30436
rect 27020 41074 27076 41076
rect 27020 41022 27022 41074
rect 27022 41022 27074 41074
rect 27074 41022 27076 41074
rect 27020 41020 27076 41022
rect 27244 40402 27300 40404
rect 27244 40350 27246 40402
rect 27246 40350 27298 40402
rect 27298 40350 27300 40402
rect 27244 40348 27300 40350
rect 26236 32674 26292 32676
rect 26236 32622 26238 32674
rect 26238 32622 26290 32674
rect 26290 32622 26292 32674
rect 26236 32620 26292 32622
rect 26572 35196 26628 35252
rect 26460 33740 26516 33796
rect 26796 39618 26852 39620
rect 26796 39566 26798 39618
rect 26798 39566 26850 39618
rect 26850 39566 26852 39618
rect 26796 39564 26852 39566
rect 26908 37772 26964 37828
rect 27132 37436 27188 37492
rect 27244 37660 27300 37716
rect 27020 37324 27076 37380
rect 26908 35922 26964 35924
rect 26908 35870 26910 35922
rect 26910 35870 26962 35922
rect 26962 35870 26964 35922
rect 26908 35868 26964 35870
rect 27020 35980 27076 36036
rect 26908 34914 26964 34916
rect 26908 34862 26910 34914
rect 26910 34862 26962 34914
rect 26962 34862 26964 34914
rect 26908 34860 26964 34862
rect 27244 36428 27300 36484
rect 27580 43484 27636 43540
rect 27916 42866 27972 42868
rect 27916 42814 27918 42866
rect 27918 42814 27970 42866
rect 27970 42814 27972 42866
rect 27916 42812 27972 42814
rect 27580 42252 27636 42308
rect 28252 42476 28308 42532
rect 27692 41970 27748 41972
rect 27692 41918 27694 41970
rect 27694 41918 27746 41970
rect 27746 41918 27748 41970
rect 27692 41916 27748 41918
rect 27468 41298 27524 41300
rect 27468 41246 27470 41298
rect 27470 41246 27522 41298
rect 27522 41246 27524 41298
rect 27468 41244 27524 41246
rect 28028 41298 28084 41300
rect 28028 41246 28030 41298
rect 28030 41246 28082 41298
rect 28082 41246 28084 41298
rect 28028 41244 28084 41246
rect 27580 41132 27636 41188
rect 27468 39394 27524 39396
rect 27468 39342 27470 39394
rect 27470 39342 27522 39394
rect 27522 39342 27524 39394
rect 27468 39340 27524 39342
rect 27468 38722 27524 38724
rect 27468 38670 27470 38722
rect 27470 38670 27522 38722
rect 27522 38670 27524 38722
rect 27468 38668 27524 38670
rect 27916 38162 27972 38164
rect 27916 38110 27918 38162
rect 27918 38110 27970 38162
rect 27970 38110 27972 38162
rect 27916 38108 27972 38110
rect 28476 44044 28532 44100
rect 28700 45106 28756 45108
rect 28700 45054 28702 45106
rect 28702 45054 28754 45106
rect 28754 45054 28756 45106
rect 28700 45052 28756 45054
rect 28476 42028 28532 42084
rect 28700 41356 28756 41412
rect 28700 38668 28756 38724
rect 27468 37436 27524 37492
rect 27468 36988 27524 37044
rect 27468 36594 27524 36596
rect 27468 36542 27470 36594
rect 27470 36542 27522 36594
rect 27522 36542 27524 36594
rect 27468 36540 27524 36542
rect 27356 35980 27412 36036
rect 27356 35084 27412 35140
rect 27244 34690 27300 34692
rect 27244 34638 27246 34690
rect 27246 34638 27298 34690
rect 27298 34638 27300 34690
rect 27244 34636 27300 34638
rect 26908 34130 26964 34132
rect 26908 34078 26910 34130
rect 26910 34078 26962 34130
rect 26962 34078 26964 34130
rect 26908 34076 26964 34078
rect 26348 32508 26404 32564
rect 27132 33234 27188 33236
rect 27132 33182 27134 33234
rect 27134 33182 27186 33234
rect 27186 33182 27188 33234
rect 27132 33180 27188 33182
rect 26572 33122 26628 33124
rect 26572 33070 26574 33122
rect 26574 33070 26626 33122
rect 26626 33070 26628 33122
rect 26572 33068 26628 33070
rect 26908 33068 26964 33124
rect 26236 31554 26292 31556
rect 26236 31502 26238 31554
rect 26238 31502 26290 31554
rect 26290 31502 26292 31554
rect 26236 31500 26292 31502
rect 26348 31388 26404 31444
rect 26348 30828 26404 30884
rect 27020 32396 27076 32452
rect 26684 31948 26740 32004
rect 26572 30828 26628 30884
rect 25900 29484 25956 29540
rect 25788 29426 25844 29428
rect 25788 29374 25790 29426
rect 25790 29374 25842 29426
rect 25842 29374 25844 29426
rect 25788 29372 25844 29374
rect 25676 29314 25732 29316
rect 25676 29262 25678 29314
rect 25678 29262 25730 29314
rect 25730 29262 25732 29314
rect 25676 29260 25732 29262
rect 25452 28476 25508 28532
rect 25228 28028 25284 28084
rect 25228 27468 25284 27524
rect 25116 27244 25172 27300
rect 25116 26514 25172 26516
rect 25116 26462 25118 26514
rect 25118 26462 25170 26514
rect 25170 26462 25172 26514
rect 25116 26460 25172 26462
rect 25900 28028 25956 28084
rect 25564 27858 25620 27860
rect 25564 27806 25566 27858
rect 25566 27806 25618 27858
rect 25618 27806 25620 27858
rect 25564 27804 25620 27806
rect 25452 27132 25508 27188
rect 25900 27244 25956 27300
rect 26012 26514 26068 26516
rect 26012 26462 26014 26514
rect 26014 26462 26066 26514
rect 26066 26462 26068 26514
rect 26012 26460 26068 26462
rect 25452 26402 25508 26404
rect 25452 26350 25454 26402
rect 25454 26350 25506 26402
rect 25506 26350 25508 26402
rect 25452 26348 25508 26350
rect 25788 26348 25844 26404
rect 25452 25004 25508 25060
rect 25116 23996 25172 24052
rect 25564 23826 25620 23828
rect 25564 23774 25566 23826
rect 25566 23774 25618 23826
rect 25618 23774 25620 23826
rect 25564 23772 25620 23774
rect 25340 23154 25396 23156
rect 25340 23102 25342 23154
rect 25342 23102 25394 23154
rect 25394 23102 25396 23154
rect 25340 23100 25396 23102
rect 24444 21644 24500 21700
rect 24332 21586 24388 21588
rect 24332 21534 24334 21586
rect 24334 21534 24386 21586
rect 24386 21534 24388 21586
rect 24332 21532 24388 21534
rect 24108 21420 24164 21476
rect 23996 21196 24052 21252
rect 26908 31666 26964 31668
rect 26908 31614 26910 31666
rect 26910 31614 26962 31666
rect 26962 31614 26964 31666
rect 26908 31612 26964 31614
rect 26796 30380 26852 30436
rect 26572 28588 26628 28644
rect 26684 29148 26740 29204
rect 26124 23996 26180 24052
rect 26236 28364 26292 28420
rect 26348 27244 26404 27300
rect 26348 26908 26404 26964
rect 26572 26012 26628 26068
rect 26348 25900 26404 25956
rect 26572 25004 26628 25060
rect 26460 23436 26516 23492
rect 26348 23324 26404 23380
rect 25228 22370 25284 22372
rect 25228 22318 25230 22370
rect 25230 22318 25282 22370
rect 25282 22318 25284 22370
rect 25228 22316 25284 22318
rect 25676 22316 25732 22372
rect 25004 21644 25060 21700
rect 24556 20188 24612 20244
rect 23548 19122 23604 19124
rect 23548 19070 23550 19122
rect 23550 19070 23602 19122
rect 23602 19070 23604 19122
rect 23548 19068 23604 19070
rect 23324 18396 23380 18452
rect 23212 17948 23268 18004
rect 23660 18732 23716 18788
rect 23772 18508 23828 18564
rect 24108 18338 24164 18340
rect 24108 18286 24110 18338
rect 24110 18286 24162 18338
rect 24162 18286 24164 18338
rect 24108 18284 24164 18286
rect 24332 18450 24388 18452
rect 24332 18398 24334 18450
rect 24334 18398 24386 18450
rect 24386 18398 24388 18450
rect 24332 18396 24388 18398
rect 24220 18172 24276 18228
rect 24780 19964 24836 20020
rect 24780 19180 24836 19236
rect 24668 18732 24724 18788
rect 24556 18674 24612 18676
rect 24556 18622 24558 18674
rect 24558 18622 24610 18674
rect 24610 18622 24612 18674
rect 24556 18620 24612 18622
rect 25452 21698 25508 21700
rect 25452 21646 25454 21698
rect 25454 21646 25506 21698
rect 25506 21646 25508 21698
rect 25452 21644 25508 21646
rect 25564 21420 25620 21476
rect 25340 20188 25396 20244
rect 25676 20018 25732 20020
rect 25676 19966 25678 20018
rect 25678 19966 25730 20018
rect 25730 19966 25732 20018
rect 25676 19964 25732 19966
rect 26124 23042 26180 23044
rect 26124 22990 26126 23042
rect 26126 22990 26178 23042
rect 26178 22990 26180 23042
rect 26124 22988 26180 22990
rect 26012 21644 26068 21700
rect 26348 22428 26404 22484
rect 26572 22652 26628 22708
rect 26460 21532 26516 21588
rect 26796 28082 26852 28084
rect 26796 28030 26798 28082
rect 26798 28030 26850 28082
rect 26850 28030 26852 28082
rect 26796 28028 26852 28030
rect 26796 26460 26852 26516
rect 27468 34300 27524 34356
rect 28252 37660 28308 37716
rect 28140 36428 28196 36484
rect 27580 34860 27636 34916
rect 27468 33570 27524 33572
rect 27468 33518 27470 33570
rect 27470 33518 27522 33570
rect 27522 33518 27524 33570
rect 27468 33516 27524 33518
rect 27916 35980 27972 36036
rect 28140 35644 28196 35700
rect 28028 34802 28084 34804
rect 28028 34750 28030 34802
rect 28030 34750 28082 34802
rect 28082 34750 28084 34802
rect 28028 34748 28084 34750
rect 27692 34354 27748 34356
rect 27692 34302 27694 34354
rect 27694 34302 27746 34354
rect 27746 34302 27748 34354
rect 27692 34300 27748 34302
rect 27580 33292 27636 33348
rect 27916 32844 27972 32900
rect 27692 31836 27748 31892
rect 28588 36092 28644 36148
rect 28476 35084 28532 35140
rect 28476 34300 28532 34356
rect 28364 34188 28420 34244
rect 28588 34018 28644 34020
rect 28588 33966 28590 34018
rect 28590 33966 28642 34018
rect 28642 33966 28644 34018
rect 28588 33964 28644 33966
rect 28476 33516 28532 33572
rect 28476 33122 28532 33124
rect 28476 33070 28478 33122
rect 28478 33070 28530 33122
rect 28530 33070 28532 33122
rect 28476 33068 28532 33070
rect 28364 31836 28420 31892
rect 28140 31724 28196 31780
rect 28588 31666 28644 31668
rect 28588 31614 28590 31666
rect 28590 31614 28642 31666
rect 28642 31614 28644 31666
rect 28588 31612 28644 31614
rect 27132 30940 27188 30996
rect 27356 31388 27412 31444
rect 27244 30882 27300 30884
rect 27244 30830 27246 30882
rect 27246 30830 27298 30882
rect 27298 30830 27300 30882
rect 27244 30828 27300 30830
rect 27244 30098 27300 30100
rect 27244 30046 27246 30098
rect 27246 30046 27298 30098
rect 27298 30046 27300 30098
rect 27244 30044 27300 30046
rect 27804 31554 27860 31556
rect 27804 31502 27806 31554
rect 27806 31502 27858 31554
rect 27858 31502 27860 31554
rect 27804 31500 27860 31502
rect 28140 31388 28196 31444
rect 27692 31276 27748 31332
rect 28700 30940 28756 30996
rect 27468 30210 27524 30212
rect 27468 30158 27470 30210
rect 27470 30158 27522 30210
rect 27522 30158 27524 30210
rect 27468 30156 27524 30158
rect 28588 30156 28644 30212
rect 27692 29986 27748 29988
rect 27692 29934 27694 29986
rect 27694 29934 27746 29986
rect 27746 29934 27748 29986
rect 27692 29932 27748 29934
rect 27132 28028 27188 28084
rect 28364 29932 28420 29988
rect 29036 48972 29092 49028
rect 28924 47516 28980 47572
rect 29036 47180 29092 47236
rect 28924 43650 28980 43652
rect 28924 43598 28926 43650
rect 28926 43598 28978 43650
rect 28978 43598 28980 43650
rect 28924 43596 28980 43598
rect 29708 53564 29764 53620
rect 29596 52556 29652 52612
rect 29484 52444 29540 52500
rect 30828 57874 30884 57876
rect 30828 57822 30830 57874
rect 30830 57822 30882 57874
rect 30882 57822 30884 57874
rect 30828 57820 30884 57822
rect 30940 57650 30996 57652
rect 30940 57598 30942 57650
rect 30942 57598 30994 57650
rect 30994 57598 30996 57650
rect 30940 57596 30996 57598
rect 31276 57484 31332 57540
rect 30380 56924 30436 56980
rect 31052 56812 31108 56868
rect 30380 55356 30436 55412
rect 30156 54626 30212 54628
rect 30156 54574 30158 54626
rect 30158 54574 30210 54626
rect 30210 54574 30212 54626
rect 30156 54572 30212 54574
rect 30044 53618 30100 53620
rect 30044 53566 30046 53618
rect 30046 53566 30098 53618
rect 30098 53566 30100 53618
rect 30044 53564 30100 53566
rect 30268 53676 30324 53732
rect 29932 53452 29988 53508
rect 30044 53170 30100 53172
rect 30044 53118 30046 53170
rect 30046 53118 30098 53170
rect 30098 53118 30100 53170
rect 30044 53116 30100 53118
rect 30492 55244 30548 55300
rect 30492 54460 30548 54516
rect 30716 55074 30772 55076
rect 30716 55022 30718 55074
rect 30718 55022 30770 55074
rect 30770 55022 30772 55074
rect 30716 55020 30772 55022
rect 30828 54684 30884 54740
rect 30156 53004 30212 53060
rect 30380 52668 30436 52724
rect 29932 51938 29988 51940
rect 29932 51886 29934 51938
rect 29934 51886 29986 51938
rect 29986 51886 29988 51938
rect 29932 51884 29988 51886
rect 29484 50764 29540 50820
rect 29260 48802 29316 48804
rect 29260 48750 29262 48802
rect 29262 48750 29314 48802
rect 29314 48750 29316 48802
rect 29260 48748 29316 48750
rect 29372 47068 29428 47124
rect 29260 46844 29316 46900
rect 30380 49922 30436 49924
rect 30380 49870 30382 49922
rect 30382 49870 30434 49922
rect 30434 49870 30436 49922
rect 30380 49868 30436 49870
rect 30156 49810 30212 49812
rect 30156 49758 30158 49810
rect 30158 49758 30210 49810
rect 30210 49758 30212 49810
rect 30156 49756 30212 49758
rect 29820 49026 29876 49028
rect 29820 48974 29822 49026
rect 29822 48974 29874 49026
rect 29874 48974 29876 49026
rect 29820 48972 29876 48974
rect 29932 48188 29988 48244
rect 29820 47458 29876 47460
rect 29820 47406 29822 47458
rect 29822 47406 29874 47458
rect 29874 47406 29876 47458
rect 29820 47404 29876 47406
rect 29596 47346 29652 47348
rect 29596 47294 29598 47346
rect 29598 47294 29650 47346
rect 29650 47294 29652 47346
rect 29596 47292 29652 47294
rect 29708 47068 29764 47124
rect 30156 47068 30212 47124
rect 29260 46172 29316 46228
rect 29148 45106 29204 45108
rect 29148 45054 29150 45106
rect 29150 45054 29202 45106
rect 29202 45054 29204 45106
rect 29148 45052 29204 45054
rect 29372 45218 29428 45220
rect 29372 45166 29374 45218
rect 29374 45166 29426 45218
rect 29426 45166 29428 45218
rect 29372 45164 29428 45166
rect 29596 44994 29652 44996
rect 29596 44942 29598 44994
rect 29598 44942 29650 44994
rect 29650 44942 29652 44994
rect 29596 44940 29652 44942
rect 30940 54514 30996 54516
rect 30940 54462 30942 54514
rect 30942 54462 30994 54514
rect 30994 54462 30996 54514
rect 30940 54460 30996 54462
rect 31612 56642 31668 56644
rect 31612 56590 31614 56642
rect 31614 56590 31666 56642
rect 31666 56590 31668 56642
rect 31612 56588 31668 56590
rect 31276 55020 31332 55076
rect 31500 56140 31556 56196
rect 31164 54796 31220 54852
rect 31052 53676 31108 53732
rect 30828 53170 30884 53172
rect 30828 53118 30830 53170
rect 30830 53118 30882 53170
rect 30882 53118 30884 53170
rect 30828 53116 30884 53118
rect 30940 53228 30996 53284
rect 30716 52722 30772 52724
rect 30716 52670 30718 52722
rect 30718 52670 30770 52722
rect 30770 52670 30772 52722
rect 30716 52668 30772 52670
rect 30940 52050 30996 52052
rect 30940 51998 30942 52050
rect 30942 51998 30994 52050
rect 30994 51998 30996 52050
rect 30940 51996 30996 51998
rect 31052 51884 31108 51940
rect 31388 52946 31444 52948
rect 31388 52894 31390 52946
rect 31390 52894 31442 52946
rect 31442 52894 31444 52946
rect 31388 52892 31444 52894
rect 31388 52668 31444 52724
rect 31612 54348 31668 54404
rect 32732 60956 32788 61012
rect 32060 60898 32116 60900
rect 32060 60846 32062 60898
rect 32062 60846 32114 60898
rect 32114 60846 32116 60898
rect 32060 60844 32116 60846
rect 32508 60786 32564 60788
rect 32508 60734 32510 60786
rect 32510 60734 32562 60786
rect 32562 60734 32564 60786
rect 32508 60732 32564 60734
rect 32284 59948 32340 60004
rect 32396 59836 32452 59892
rect 32172 59612 32228 59668
rect 33180 61404 33236 61460
rect 32844 60620 32900 60676
rect 33068 59948 33124 60004
rect 32396 58380 32452 58436
rect 32620 59276 32676 59332
rect 31948 58210 32004 58212
rect 31948 58158 31950 58210
rect 31950 58158 32002 58210
rect 32002 58158 32004 58210
rect 31948 58156 32004 58158
rect 31836 57596 31892 57652
rect 32844 58828 32900 58884
rect 32732 58604 32788 58660
rect 31836 56140 31892 56196
rect 32060 55468 32116 55524
rect 31612 53452 31668 53508
rect 33516 62466 33572 62468
rect 33516 62414 33518 62466
rect 33518 62414 33570 62466
rect 33570 62414 33572 62466
rect 33516 62412 33572 62414
rect 33964 66050 34020 66052
rect 33964 65998 33966 66050
rect 33966 65998 34018 66050
rect 34018 65998 34020 66050
rect 33964 65996 34020 65998
rect 34188 65602 34244 65604
rect 34188 65550 34190 65602
rect 34190 65550 34242 65602
rect 34242 65550 34244 65602
rect 34188 65548 34244 65550
rect 33964 65324 34020 65380
rect 34076 65212 34132 65268
rect 34076 64540 34132 64596
rect 33964 64204 34020 64260
rect 33852 62354 33908 62356
rect 33852 62302 33854 62354
rect 33854 62302 33906 62354
rect 33906 62302 33908 62354
rect 33852 62300 33908 62302
rect 34188 64034 34244 64036
rect 34188 63982 34190 64034
rect 34190 63982 34242 64034
rect 34242 63982 34244 64034
rect 34188 63980 34244 63982
rect 34412 64428 34468 64484
rect 34972 65436 35028 65492
rect 34524 64204 34580 64260
rect 35532 68908 35588 68964
rect 35756 68572 35812 68628
rect 35980 68460 36036 68516
rect 35196 68234 35252 68236
rect 35196 68182 35198 68234
rect 35198 68182 35250 68234
rect 35250 68182 35252 68234
rect 35196 68180 35252 68182
rect 35300 68234 35356 68236
rect 35300 68182 35302 68234
rect 35302 68182 35354 68234
rect 35354 68182 35356 68234
rect 35300 68180 35356 68182
rect 35404 68234 35460 68236
rect 35404 68182 35406 68234
rect 35406 68182 35458 68234
rect 35458 68182 35460 68234
rect 35404 68180 35460 68182
rect 37212 70476 37268 70532
rect 38444 70588 38500 70644
rect 37212 69580 37268 69636
rect 39564 70476 39620 70532
rect 36988 69356 37044 69412
rect 38556 69356 38612 69412
rect 36316 69298 36372 69300
rect 36316 69246 36318 69298
rect 36318 69246 36370 69298
rect 36370 69246 36372 69298
rect 36316 69244 36372 69246
rect 37548 69298 37604 69300
rect 37548 69246 37550 69298
rect 37550 69246 37602 69298
rect 37602 69246 37604 69298
rect 37548 69244 37604 69246
rect 36428 68572 36484 68628
rect 35868 67618 35924 67620
rect 35868 67566 35870 67618
rect 35870 67566 35922 67618
rect 35922 67566 35924 67618
rect 35868 67564 35924 67566
rect 37100 68460 37156 68516
rect 37436 69186 37492 69188
rect 37436 69134 37438 69186
rect 37438 69134 37490 69186
rect 37490 69134 37492 69186
rect 37436 69132 37492 69134
rect 37324 68850 37380 68852
rect 37324 68798 37326 68850
rect 37326 68798 37378 68850
rect 37378 68798 37380 68850
rect 37324 68796 37380 68798
rect 37324 68572 37380 68628
rect 38108 68850 38164 68852
rect 38108 68798 38110 68850
rect 38110 68798 38162 68850
rect 38162 68798 38164 68850
rect 38108 68796 38164 68798
rect 38332 69186 38388 69188
rect 38332 69134 38334 69186
rect 38334 69134 38386 69186
rect 38386 69134 38388 69186
rect 38332 69132 38388 69134
rect 37884 68460 37940 68516
rect 37660 67788 37716 67844
rect 38444 68908 38500 68964
rect 38108 67452 38164 67508
rect 35532 67004 35588 67060
rect 35196 66666 35252 66668
rect 35196 66614 35198 66666
rect 35198 66614 35250 66666
rect 35250 66614 35252 66666
rect 35196 66612 35252 66614
rect 35300 66666 35356 66668
rect 35300 66614 35302 66666
rect 35302 66614 35354 66666
rect 35354 66614 35356 66666
rect 35300 66612 35356 66614
rect 35404 66666 35460 66668
rect 35404 66614 35406 66666
rect 35406 66614 35458 66666
rect 35458 66614 35460 66666
rect 35404 66612 35460 66614
rect 35420 65996 35476 66052
rect 35196 65436 35252 65492
rect 35196 65098 35252 65100
rect 35196 65046 35198 65098
rect 35198 65046 35250 65098
rect 35250 65046 35252 65098
rect 35196 65044 35252 65046
rect 35300 65098 35356 65100
rect 35300 65046 35302 65098
rect 35302 65046 35354 65098
rect 35354 65046 35356 65098
rect 35300 65044 35356 65046
rect 35404 65098 35460 65100
rect 35404 65046 35406 65098
rect 35406 65046 35458 65098
rect 35458 65046 35460 65098
rect 35404 65044 35460 65046
rect 34972 64540 35028 64596
rect 36204 66162 36260 66164
rect 36204 66110 36206 66162
rect 36206 66110 36258 66162
rect 36258 66110 36260 66162
rect 36204 66108 36260 66110
rect 35756 64706 35812 64708
rect 35756 64654 35758 64706
rect 35758 64654 35810 64706
rect 35810 64654 35812 64706
rect 35756 64652 35812 64654
rect 35980 64316 36036 64372
rect 34636 64092 34692 64148
rect 34524 63810 34580 63812
rect 34524 63758 34526 63810
rect 34526 63758 34578 63810
rect 34578 63758 34580 63810
rect 34524 63756 34580 63758
rect 35196 63530 35252 63532
rect 35196 63478 35198 63530
rect 35198 63478 35250 63530
rect 35250 63478 35252 63530
rect 35196 63476 35252 63478
rect 35300 63530 35356 63532
rect 35300 63478 35302 63530
rect 35302 63478 35354 63530
rect 35354 63478 35356 63530
rect 35300 63476 35356 63478
rect 35404 63530 35460 63532
rect 35404 63478 35406 63530
rect 35406 63478 35458 63530
rect 35458 63478 35460 63530
rect 35404 63476 35460 63478
rect 36316 66050 36372 66052
rect 36316 65998 36318 66050
rect 36318 65998 36370 66050
rect 36370 65998 36372 66050
rect 36316 65996 36372 65998
rect 36428 65212 36484 65268
rect 39340 69298 39396 69300
rect 39340 69246 39342 69298
rect 39342 69246 39394 69298
rect 39394 69246 39396 69298
rect 39340 69244 39396 69246
rect 40236 71596 40292 71652
rect 40908 71650 40964 71652
rect 40908 71598 40910 71650
rect 40910 71598 40962 71650
rect 40962 71598 40964 71650
rect 40908 71596 40964 71598
rect 40348 70588 40404 70644
rect 39900 70252 39956 70308
rect 40908 70252 40964 70308
rect 39340 68908 39396 68964
rect 39116 68796 39172 68852
rect 39228 68738 39284 68740
rect 39228 68686 39230 68738
rect 39230 68686 39282 68738
rect 39282 68686 39284 68738
rect 39228 68684 39284 68686
rect 39004 67788 39060 67844
rect 38780 67452 38836 67508
rect 36988 66162 37044 66164
rect 36988 66110 36990 66162
rect 36990 66110 37042 66162
rect 37042 66110 37044 66162
rect 36988 66108 37044 66110
rect 36652 64316 36708 64372
rect 35756 63196 35812 63252
rect 34300 62860 34356 62916
rect 36092 63308 36148 63364
rect 35196 62914 35252 62916
rect 35196 62862 35198 62914
rect 35198 62862 35250 62914
rect 35250 62862 35252 62914
rect 35196 62860 35252 62862
rect 35644 62914 35700 62916
rect 35644 62862 35646 62914
rect 35646 62862 35698 62914
rect 35698 62862 35700 62914
rect 35644 62860 35700 62862
rect 34748 62524 34804 62580
rect 35644 62636 35700 62692
rect 35196 62354 35252 62356
rect 35196 62302 35198 62354
rect 35198 62302 35250 62354
rect 35250 62302 35252 62354
rect 35196 62300 35252 62302
rect 34188 61964 34244 62020
rect 33628 60732 33684 60788
rect 33740 60844 33796 60900
rect 33292 59500 33348 59556
rect 33180 58828 33236 58884
rect 33516 59330 33572 59332
rect 33516 59278 33518 59330
rect 33518 59278 33570 59330
rect 33570 59278 33572 59330
rect 33516 59276 33572 59278
rect 33516 58828 33572 58884
rect 33180 58380 33236 58436
rect 32284 56476 32340 56532
rect 32508 56588 32564 56644
rect 32396 56028 32452 56084
rect 31836 54738 31892 54740
rect 31836 54686 31838 54738
rect 31838 54686 31890 54738
rect 31890 54686 31892 54738
rect 31836 54684 31892 54686
rect 31724 52668 31780 52724
rect 31836 52108 31892 52164
rect 31164 50316 31220 50372
rect 31388 51212 31444 51268
rect 31164 49868 31220 49924
rect 30604 49308 30660 49364
rect 30716 49756 30772 49812
rect 30492 48914 30548 48916
rect 30492 48862 30494 48914
rect 30494 48862 30546 48914
rect 30546 48862 30548 48914
rect 30492 48860 30548 48862
rect 30492 47458 30548 47460
rect 30492 47406 30494 47458
rect 30494 47406 30546 47458
rect 30546 47406 30548 47458
rect 30492 47404 30548 47406
rect 29260 44098 29316 44100
rect 29260 44046 29262 44098
rect 29262 44046 29314 44098
rect 29314 44046 29316 44098
rect 29260 44044 29316 44046
rect 29596 43596 29652 43652
rect 29596 42754 29652 42756
rect 29596 42702 29598 42754
rect 29598 42702 29650 42754
rect 29650 42702 29652 42754
rect 29596 42700 29652 42702
rect 29596 42476 29652 42532
rect 29708 42028 29764 42084
rect 29148 41356 29204 41412
rect 29372 41858 29428 41860
rect 29372 41806 29374 41858
rect 29374 41806 29426 41858
rect 29426 41806 29428 41858
rect 29372 41804 29428 41806
rect 29484 41580 29540 41636
rect 29260 41186 29316 41188
rect 29260 41134 29262 41186
rect 29262 41134 29314 41186
rect 29314 41134 29316 41186
rect 29260 41132 29316 41134
rect 29596 39564 29652 39620
rect 29372 39340 29428 39396
rect 29596 38946 29652 38948
rect 29596 38894 29598 38946
rect 29598 38894 29650 38946
rect 29650 38894 29652 38946
rect 29596 38892 29652 38894
rect 30380 45724 30436 45780
rect 29932 43538 29988 43540
rect 29932 43486 29934 43538
rect 29934 43486 29986 43538
rect 29986 43486 29988 43538
rect 29932 43484 29988 43486
rect 30156 42476 30212 42532
rect 29932 40796 29988 40852
rect 29820 39506 29876 39508
rect 29820 39454 29822 39506
rect 29822 39454 29874 39506
rect 29874 39454 29876 39506
rect 29820 39452 29876 39454
rect 29708 38556 29764 38612
rect 29372 38108 29428 38164
rect 29372 37436 29428 37492
rect 28924 34300 28980 34356
rect 30044 39452 30100 39508
rect 30156 39228 30212 39284
rect 30380 43426 30436 43428
rect 30380 43374 30382 43426
rect 30382 43374 30434 43426
rect 30434 43374 30436 43426
rect 30380 43372 30436 43374
rect 30492 41970 30548 41972
rect 30492 41918 30494 41970
rect 30494 41918 30546 41970
rect 30546 41918 30548 41970
rect 30492 41916 30548 41918
rect 30380 41074 30436 41076
rect 30380 41022 30382 41074
rect 30382 41022 30434 41074
rect 30434 41022 30436 41074
rect 30380 41020 30436 41022
rect 30380 40796 30436 40852
rect 30716 48188 30772 48244
rect 31388 49810 31444 49812
rect 31388 49758 31390 49810
rect 31390 49758 31442 49810
rect 31442 49758 31444 49810
rect 31388 49756 31444 49758
rect 31388 49308 31444 49364
rect 31388 48300 31444 48356
rect 30716 47516 30772 47572
rect 31276 47068 31332 47124
rect 31836 51266 31892 51268
rect 31836 51214 31838 51266
rect 31838 51214 31890 51266
rect 31890 51214 31892 51266
rect 31836 51212 31892 51214
rect 31836 50204 31892 50260
rect 31612 48972 31668 49028
rect 31612 47292 31668 47348
rect 31836 47458 31892 47460
rect 31836 47406 31838 47458
rect 31838 47406 31890 47458
rect 31890 47406 31892 47458
rect 31836 47404 31892 47406
rect 31276 45218 31332 45220
rect 31276 45166 31278 45218
rect 31278 45166 31330 45218
rect 31330 45166 31332 45218
rect 31276 45164 31332 45166
rect 31052 45052 31108 45108
rect 30940 44994 30996 44996
rect 30940 44942 30942 44994
rect 30942 44942 30994 44994
rect 30994 44942 30996 44994
rect 30940 44940 30996 44942
rect 30940 43372 30996 43428
rect 30716 42754 30772 42756
rect 30716 42702 30718 42754
rect 30718 42702 30770 42754
rect 30770 42702 30772 42754
rect 30716 42700 30772 42702
rect 31612 44940 31668 44996
rect 31500 44828 31556 44884
rect 31500 43708 31556 43764
rect 30828 41804 30884 41860
rect 30604 40514 30660 40516
rect 30604 40462 30606 40514
rect 30606 40462 30658 40514
rect 30658 40462 30660 40514
rect 30604 40460 30660 40462
rect 30492 40124 30548 40180
rect 31612 42700 31668 42756
rect 31388 42476 31444 42532
rect 31276 41020 31332 41076
rect 32172 54514 32228 54516
rect 32172 54462 32174 54514
rect 32174 54462 32226 54514
rect 32226 54462 32228 54514
rect 32172 54460 32228 54462
rect 32284 53170 32340 53172
rect 32284 53118 32286 53170
rect 32286 53118 32338 53170
rect 32338 53118 32340 53170
rect 32284 53116 32340 53118
rect 32396 52892 32452 52948
rect 32620 51938 32676 51940
rect 32620 51886 32622 51938
rect 32622 51886 32674 51938
rect 32674 51886 32676 51938
rect 32620 51884 32676 51886
rect 32732 51660 32788 51716
rect 32620 48860 32676 48916
rect 32060 48242 32116 48244
rect 32060 48190 32062 48242
rect 32062 48190 32114 48242
rect 32114 48190 32116 48242
rect 32060 48188 32116 48190
rect 32508 47628 32564 47684
rect 32732 48188 32788 48244
rect 32956 57932 33012 57988
rect 33404 58546 33460 58548
rect 33404 58494 33406 58546
rect 33406 58494 33458 58546
rect 33458 58494 33460 58546
rect 33404 58492 33460 58494
rect 33740 58492 33796 58548
rect 33516 57650 33572 57652
rect 33516 57598 33518 57650
rect 33518 57598 33570 57650
rect 33570 57598 33572 57650
rect 33516 57596 33572 57598
rect 33180 56642 33236 56644
rect 33180 56590 33182 56642
rect 33182 56590 33234 56642
rect 33234 56590 33236 56642
rect 33180 56588 33236 56590
rect 33068 56476 33124 56532
rect 33516 56082 33572 56084
rect 33516 56030 33518 56082
rect 33518 56030 33570 56082
rect 33570 56030 33572 56082
rect 33516 56028 33572 56030
rect 33292 55356 33348 55412
rect 33292 54402 33348 54404
rect 33292 54350 33294 54402
rect 33294 54350 33346 54402
rect 33346 54350 33348 54402
rect 33292 54348 33348 54350
rect 33180 53564 33236 53620
rect 33068 53170 33124 53172
rect 33068 53118 33070 53170
rect 33070 53118 33122 53170
rect 33122 53118 33124 53170
rect 33068 53116 33124 53118
rect 36540 62578 36596 62580
rect 36540 62526 36542 62578
rect 36542 62526 36594 62578
rect 36594 62526 36596 62578
rect 36540 62524 36596 62526
rect 35196 61962 35252 61964
rect 35196 61910 35198 61962
rect 35198 61910 35250 61962
rect 35250 61910 35252 61962
rect 35196 61908 35252 61910
rect 35300 61962 35356 61964
rect 35300 61910 35302 61962
rect 35302 61910 35354 61962
rect 35354 61910 35356 61962
rect 35300 61908 35356 61910
rect 35404 61962 35460 61964
rect 35404 61910 35406 61962
rect 35406 61910 35458 61962
rect 35458 61910 35460 61962
rect 35404 61908 35460 61910
rect 34748 61740 34804 61796
rect 33964 61292 34020 61348
rect 34188 59724 34244 59780
rect 34860 60674 34916 60676
rect 34860 60622 34862 60674
rect 34862 60622 34914 60674
rect 34914 60622 34916 60674
rect 34860 60620 34916 60622
rect 34636 59948 34692 60004
rect 34188 58716 34244 58772
rect 36092 62412 36148 62468
rect 35308 60508 35364 60564
rect 35196 60394 35252 60396
rect 35196 60342 35198 60394
rect 35198 60342 35250 60394
rect 35250 60342 35252 60394
rect 35196 60340 35252 60342
rect 35300 60394 35356 60396
rect 35300 60342 35302 60394
rect 35302 60342 35354 60394
rect 35354 60342 35356 60394
rect 35300 60340 35356 60342
rect 35404 60394 35460 60396
rect 35404 60342 35406 60394
rect 35406 60342 35458 60394
rect 35458 60342 35460 60394
rect 35404 60340 35460 60342
rect 35420 60172 35476 60228
rect 34860 59612 34916 59668
rect 34860 58940 34916 58996
rect 35084 59612 35140 59668
rect 34748 58828 34804 58884
rect 34636 58716 34692 58772
rect 34076 58380 34132 58436
rect 34188 58492 34244 58548
rect 34524 58268 34580 58324
rect 34076 57538 34132 57540
rect 34076 57486 34078 57538
rect 34078 57486 34130 57538
rect 34130 57486 34132 57538
rect 34076 57484 34132 57486
rect 33964 56978 34020 56980
rect 33964 56926 33966 56978
rect 33966 56926 34018 56978
rect 34018 56926 34020 56978
rect 33964 56924 34020 56926
rect 33964 56082 34020 56084
rect 33964 56030 33966 56082
rect 33966 56030 34018 56082
rect 34018 56030 34020 56082
rect 33964 56028 34020 56030
rect 33964 55356 34020 55412
rect 34300 58210 34356 58212
rect 34300 58158 34302 58210
rect 34302 58158 34354 58210
rect 34354 58158 34356 58210
rect 34300 58156 34356 58158
rect 34412 56588 34468 56644
rect 34300 56194 34356 56196
rect 34300 56142 34302 56194
rect 34302 56142 34354 56194
rect 34354 56142 34356 56194
rect 34300 56140 34356 56142
rect 34412 56028 34468 56084
rect 34076 54796 34132 54852
rect 33404 53058 33460 53060
rect 33404 53006 33406 53058
rect 33406 53006 33458 53058
rect 33458 53006 33460 53058
rect 33404 53004 33460 53006
rect 33292 52274 33348 52276
rect 33292 52222 33294 52274
rect 33294 52222 33346 52274
rect 33346 52222 33348 52274
rect 33292 52220 33348 52222
rect 33404 50594 33460 50596
rect 33404 50542 33406 50594
rect 33406 50542 33458 50594
rect 33458 50542 33460 50594
rect 33404 50540 33460 50542
rect 33516 52220 33572 52276
rect 33068 48354 33124 48356
rect 33068 48302 33070 48354
rect 33070 48302 33122 48354
rect 33122 48302 33124 48354
rect 33068 48300 33124 48302
rect 32508 47404 32564 47460
rect 32732 47458 32788 47460
rect 32732 47406 32734 47458
rect 32734 47406 32786 47458
rect 32786 47406 32788 47458
rect 32732 47404 32788 47406
rect 32508 47234 32564 47236
rect 32508 47182 32510 47234
rect 32510 47182 32562 47234
rect 32562 47182 32564 47234
rect 32508 47180 32564 47182
rect 32060 47068 32116 47124
rect 32284 46898 32340 46900
rect 32284 46846 32286 46898
rect 32286 46846 32338 46898
rect 32338 46846 32340 46898
rect 32284 46844 32340 46846
rect 32060 46396 32116 46452
rect 31948 45612 32004 45668
rect 32396 45276 32452 45332
rect 32844 46956 32900 47012
rect 32284 45106 32340 45108
rect 32284 45054 32286 45106
rect 32286 45054 32338 45106
rect 32338 45054 32340 45106
rect 32284 45052 32340 45054
rect 32396 44156 32452 44212
rect 32284 43708 32340 43764
rect 32620 43596 32676 43652
rect 32508 42866 32564 42868
rect 32508 42814 32510 42866
rect 32510 42814 32562 42866
rect 32562 42814 32564 42866
rect 32508 42812 32564 42814
rect 31948 41804 32004 41860
rect 32060 40348 32116 40404
rect 31388 39618 31444 39620
rect 31388 39566 31390 39618
rect 31390 39566 31442 39618
rect 31442 39566 31444 39618
rect 31388 39564 31444 39566
rect 30380 39340 30436 39396
rect 30156 38108 30212 38164
rect 29820 36482 29876 36484
rect 29820 36430 29822 36482
rect 29822 36430 29874 36482
rect 29874 36430 29876 36482
rect 29820 36428 29876 36430
rect 29148 36258 29204 36260
rect 29148 36206 29150 36258
rect 29150 36206 29202 36258
rect 29202 36206 29204 36258
rect 29148 36204 29204 36206
rect 29260 34748 29316 34804
rect 30716 39228 30772 39284
rect 30604 38556 30660 38612
rect 31836 39506 31892 39508
rect 31836 39454 31838 39506
rect 31838 39454 31890 39506
rect 31890 39454 31892 39506
rect 31836 39452 31892 39454
rect 31724 39058 31780 39060
rect 31724 39006 31726 39058
rect 31726 39006 31778 39058
rect 31778 39006 31780 39058
rect 31724 39004 31780 39006
rect 30828 38108 30884 38164
rect 30156 37436 30212 37492
rect 30492 37378 30548 37380
rect 30492 37326 30494 37378
rect 30494 37326 30546 37378
rect 30546 37326 30548 37378
rect 30492 37324 30548 37326
rect 30156 36092 30212 36148
rect 30380 36428 30436 36484
rect 30380 36258 30436 36260
rect 30380 36206 30382 36258
rect 30382 36206 30434 36258
rect 30434 36206 30436 36258
rect 30380 36204 30436 36206
rect 29596 34636 29652 34692
rect 29484 34242 29540 34244
rect 29484 34190 29486 34242
rect 29486 34190 29538 34242
rect 29538 34190 29540 34242
rect 29484 34188 29540 34190
rect 29820 34300 29876 34356
rect 29260 33628 29316 33684
rect 29372 33234 29428 33236
rect 29372 33182 29374 33234
rect 29374 33182 29426 33234
rect 29426 33182 29428 33234
rect 29372 33180 29428 33182
rect 29148 33122 29204 33124
rect 29148 33070 29150 33122
rect 29150 33070 29202 33122
rect 29202 33070 29204 33122
rect 29148 33068 29204 33070
rect 29708 33964 29764 34020
rect 29596 33122 29652 33124
rect 29596 33070 29598 33122
rect 29598 33070 29650 33122
rect 29650 33070 29652 33122
rect 29596 33068 29652 33070
rect 29148 31500 29204 31556
rect 28812 30492 28868 30548
rect 28588 28364 28644 28420
rect 27916 28082 27972 28084
rect 27916 28030 27918 28082
rect 27918 28030 27970 28082
rect 27970 28030 27972 28082
rect 27916 28028 27972 28030
rect 27580 27692 27636 27748
rect 28476 27746 28532 27748
rect 28476 27694 28478 27746
rect 28478 27694 28530 27746
rect 28530 27694 28532 27746
rect 28476 27692 28532 27694
rect 27132 26460 27188 26516
rect 27692 27020 27748 27076
rect 27244 26178 27300 26180
rect 27244 26126 27246 26178
rect 27246 26126 27298 26178
rect 27298 26126 27300 26178
rect 27244 26124 27300 26126
rect 28028 26572 28084 26628
rect 28140 26908 28196 26964
rect 29036 29820 29092 29876
rect 29372 31948 29428 32004
rect 30268 34972 30324 35028
rect 30044 33346 30100 33348
rect 30044 33294 30046 33346
rect 30046 33294 30098 33346
rect 30098 33294 30100 33346
rect 30044 33292 30100 33294
rect 30156 32732 30212 32788
rect 29484 31836 29540 31892
rect 29372 31778 29428 31780
rect 29372 31726 29374 31778
rect 29374 31726 29426 31778
rect 29426 31726 29428 31778
rect 29372 31724 29428 31726
rect 29372 31500 29428 31556
rect 29260 29372 29316 29428
rect 29148 28530 29204 28532
rect 29148 28478 29150 28530
rect 29150 28478 29202 28530
rect 29202 28478 29204 28530
rect 29148 28476 29204 28478
rect 29260 28418 29316 28420
rect 29260 28366 29262 28418
rect 29262 28366 29314 28418
rect 29314 28366 29316 28418
rect 29260 28364 29316 28366
rect 26908 22988 26964 23044
rect 27132 23154 27188 23156
rect 27132 23102 27134 23154
rect 27134 23102 27186 23154
rect 27186 23102 27188 23154
rect 27132 23100 27188 23102
rect 27468 23436 27524 23492
rect 27580 26348 27636 26404
rect 29036 27858 29092 27860
rect 29036 27806 29038 27858
rect 29038 27806 29090 27858
rect 29090 27806 29092 27858
rect 29036 27804 29092 27806
rect 27356 23324 27412 23380
rect 27692 25452 27748 25508
rect 27692 23212 27748 23268
rect 27244 22988 27300 23044
rect 27804 23100 27860 23156
rect 27132 22764 27188 22820
rect 26796 22428 26852 22484
rect 26684 21420 26740 21476
rect 27692 22370 27748 22372
rect 27692 22318 27694 22370
rect 27694 22318 27746 22370
rect 27746 22318 27748 22370
rect 27692 22316 27748 22318
rect 27020 21644 27076 21700
rect 27244 21868 27300 21924
rect 27804 21868 27860 21924
rect 28140 25788 28196 25844
rect 28140 25506 28196 25508
rect 28140 25454 28142 25506
rect 28142 25454 28194 25506
rect 28194 25454 28196 25506
rect 28140 25452 28196 25454
rect 28364 25394 28420 25396
rect 28364 25342 28366 25394
rect 28366 25342 28418 25394
rect 28418 25342 28420 25394
rect 28364 25340 28420 25342
rect 28252 24050 28308 24052
rect 28252 23998 28254 24050
rect 28254 23998 28306 24050
rect 28306 23998 28308 24050
rect 28252 23996 28308 23998
rect 28588 23772 28644 23828
rect 28252 23436 28308 23492
rect 28140 22482 28196 22484
rect 28140 22430 28142 22482
rect 28142 22430 28194 22482
rect 28194 22430 28196 22482
rect 28140 22428 28196 22430
rect 27020 21420 27076 21476
rect 25228 18620 25284 18676
rect 25676 19292 25732 19348
rect 25452 19122 25508 19124
rect 25452 19070 25454 19122
rect 25454 19070 25506 19122
rect 25506 19070 25508 19122
rect 25452 19068 25508 19070
rect 25676 19010 25732 19012
rect 25676 18958 25678 19010
rect 25678 18958 25730 19010
rect 25730 18958 25732 19010
rect 25676 18956 25732 18958
rect 23884 17724 23940 17780
rect 23548 17164 23604 17220
rect 24108 17164 24164 17220
rect 25004 18172 25060 18228
rect 24444 17164 24500 17220
rect 23660 16716 23716 16772
rect 24780 16604 24836 16660
rect 23660 15484 23716 15540
rect 23324 15260 23380 15316
rect 23212 15090 23268 15092
rect 23212 15038 23214 15090
rect 23214 15038 23266 15090
rect 23266 15038 23268 15090
rect 23212 15036 23268 15038
rect 23772 14924 23828 14980
rect 23884 15484 23940 15540
rect 23548 14700 23604 14756
rect 22988 12962 23044 12964
rect 22988 12910 22990 12962
rect 22990 12910 23042 12962
rect 23042 12910 23044 12962
rect 22988 12908 23044 12910
rect 24668 15484 24724 15540
rect 24108 14700 24164 14756
rect 24332 15036 24388 15092
rect 24444 14924 24500 14980
rect 25340 18172 25396 18228
rect 25340 17778 25396 17780
rect 25340 17726 25342 17778
rect 25342 17726 25394 17778
rect 25394 17726 25396 17778
rect 25340 17724 25396 17726
rect 26012 19404 26068 19460
rect 26460 19292 26516 19348
rect 26124 19010 26180 19012
rect 26124 18958 26126 19010
rect 26126 18958 26178 19010
rect 26178 18958 26180 19010
rect 26124 18956 26180 18958
rect 25788 18172 25844 18228
rect 25900 18620 25956 18676
rect 26460 19010 26516 19012
rect 26460 18958 26462 19010
rect 26462 18958 26514 19010
rect 26514 18958 26516 19010
rect 26460 18956 26516 18958
rect 26236 18508 26292 18564
rect 25340 16658 25396 16660
rect 25340 16606 25342 16658
rect 25342 16606 25394 16658
rect 25394 16606 25396 16658
rect 25340 16604 25396 16606
rect 25452 15932 25508 15988
rect 25228 15314 25284 15316
rect 25228 15262 25230 15314
rect 25230 15262 25282 15314
rect 25282 15262 25284 15314
rect 25228 15260 25284 15262
rect 24444 14364 24500 14420
rect 24220 14306 24276 14308
rect 24220 14254 24222 14306
rect 24222 14254 24274 14306
rect 24274 14254 24276 14306
rect 24220 14252 24276 14254
rect 24668 13692 24724 13748
rect 23100 12236 23156 12292
rect 23436 12796 23492 12852
rect 21644 9602 21700 9604
rect 21644 9550 21646 9602
rect 21646 9550 21698 9602
rect 21698 9550 21700 9602
rect 21644 9548 21700 9550
rect 22988 9714 23044 9716
rect 22988 9662 22990 9714
rect 22990 9662 23042 9714
rect 23042 9662 23044 9714
rect 22988 9660 23044 9662
rect 22988 9154 23044 9156
rect 22988 9102 22990 9154
rect 22990 9102 23042 9154
rect 23042 9102 23044 9154
rect 22988 9100 23044 9102
rect 22988 8876 23044 8932
rect 21868 3442 21924 3444
rect 21868 3390 21870 3442
rect 21870 3390 21922 3442
rect 21922 3390 21924 3442
rect 21868 3388 21924 3390
rect 23436 8876 23492 8932
rect 23996 12908 24052 12964
rect 23772 12236 23828 12292
rect 24108 11788 24164 11844
rect 24668 12124 24724 12180
rect 24668 11452 24724 11508
rect 24444 9660 24500 9716
rect 23884 9042 23940 9044
rect 23884 8990 23886 9042
rect 23886 8990 23938 9042
rect 23938 8990 23940 9042
rect 23884 8988 23940 8990
rect 24220 8876 24276 8932
rect 25228 14700 25284 14756
rect 26460 16770 26516 16772
rect 26460 16718 26462 16770
rect 26462 16718 26514 16770
rect 26514 16718 26516 16770
rect 26460 16716 26516 16718
rect 25676 15036 25732 15092
rect 25116 14418 25172 14420
rect 25116 14366 25118 14418
rect 25118 14366 25170 14418
rect 25170 14366 25172 14418
rect 25116 14364 25172 14366
rect 25788 14364 25844 14420
rect 25340 13692 25396 13748
rect 25340 12962 25396 12964
rect 25340 12910 25342 12962
rect 25342 12910 25394 12962
rect 25394 12910 25396 12962
rect 25340 12908 25396 12910
rect 25004 12236 25060 12292
rect 25004 11116 25060 11172
rect 25228 11788 25284 11844
rect 25116 9996 25172 10052
rect 25452 12178 25508 12180
rect 25452 12126 25454 12178
rect 25454 12126 25506 12178
rect 25506 12126 25508 12178
rect 25452 12124 25508 12126
rect 26236 16658 26292 16660
rect 26236 16606 26238 16658
rect 26238 16606 26290 16658
rect 26290 16606 26292 16658
rect 26236 16604 26292 16606
rect 26236 15932 26292 15988
rect 26572 15932 26628 15988
rect 26572 14418 26628 14420
rect 26572 14366 26574 14418
rect 26574 14366 26626 14418
rect 26626 14366 26628 14418
rect 26572 14364 26628 14366
rect 25900 13746 25956 13748
rect 25900 13694 25902 13746
rect 25902 13694 25954 13746
rect 25954 13694 25956 13746
rect 25900 13692 25956 13694
rect 26348 13692 26404 13748
rect 26124 12066 26180 12068
rect 26124 12014 26126 12066
rect 26126 12014 26178 12066
rect 26178 12014 26180 12066
rect 26124 12012 26180 12014
rect 26796 20412 26852 20468
rect 28364 23266 28420 23268
rect 28364 23214 28366 23266
rect 28366 23214 28418 23266
rect 28418 23214 28420 23266
rect 28364 23212 28420 23214
rect 27804 20578 27860 20580
rect 27804 20526 27806 20578
rect 27806 20526 27858 20578
rect 27858 20526 27860 20578
rect 27804 20524 27860 20526
rect 27244 19852 27300 19908
rect 27244 19458 27300 19460
rect 27244 19406 27246 19458
rect 27246 19406 27298 19458
rect 27298 19406 27300 19458
rect 27244 19404 27300 19406
rect 26908 19122 26964 19124
rect 26908 19070 26910 19122
rect 26910 19070 26962 19122
rect 26962 19070 26964 19122
rect 26908 19068 26964 19070
rect 27692 19906 27748 19908
rect 27692 19854 27694 19906
rect 27694 19854 27746 19906
rect 27746 19854 27748 19906
rect 27692 19852 27748 19854
rect 27692 19404 27748 19460
rect 27356 18620 27412 18676
rect 27468 19234 27524 19236
rect 27468 19182 27470 19234
rect 27470 19182 27522 19234
rect 27522 19182 27524 19234
rect 27468 19180 27524 19182
rect 26908 18508 26964 18564
rect 27804 18956 27860 19012
rect 28252 20802 28308 20804
rect 28252 20750 28254 20802
rect 28254 20750 28306 20802
rect 28306 20750 28308 20802
rect 28252 20748 28308 20750
rect 28252 20412 28308 20468
rect 28140 19234 28196 19236
rect 28140 19182 28142 19234
rect 28142 19182 28194 19234
rect 28194 19182 28196 19234
rect 28140 19180 28196 19182
rect 27804 18620 27860 18676
rect 27468 18508 27524 18564
rect 28140 18508 28196 18564
rect 27020 16716 27076 16772
rect 26796 16604 26852 16660
rect 27692 16604 27748 16660
rect 27916 16716 27972 16772
rect 27804 15932 27860 15988
rect 27692 15820 27748 15876
rect 27244 15314 27300 15316
rect 27244 15262 27246 15314
rect 27246 15262 27298 15314
rect 27298 15262 27300 15314
rect 27244 15260 27300 15262
rect 28364 17724 28420 17780
rect 28588 21756 28644 21812
rect 29484 29484 29540 29540
rect 29484 28028 29540 28084
rect 29932 31948 29988 32004
rect 29932 31500 29988 31556
rect 29820 29932 29876 29988
rect 30380 33122 30436 33124
rect 30380 33070 30382 33122
rect 30382 33070 30434 33122
rect 30434 33070 30436 33122
rect 30380 33068 30436 33070
rect 30268 31724 30324 31780
rect 30380 32508 30436 32564
rect 30268 30210 30324 30212
rect 30268 30158 30270 30210
rect 30270 30158 30322 30210
rect 30322 30158 30324 30210
rect 30268 30156 30324 30158
rect 30044 29426 30100 29428
rect 30044 29374 30046 29426
rect 30046 29374 30098 29426
rect 30098 29374 30100 29426
rect 30044 29372 30100 29374
rect 29932 29260 29988 29316
rect 29820 28700 29876 28756
rect 29708 28028 29764 28084
rect 29820 27970 29876 27972
rect 29820 27918 29822 27970
rect 29822 27918 29874 27970
rect 29874 27918 29876 27970
rect 29820 27916 29876 27918
rect 30156 28418 30212 28420
rect 30156 28366 30158 28418
rect 30158 28366 30210 28418
rect 30210 28366 30212 28418
rect 30156 28364 30212 28366
rect 30156 27916 30212 27972
rect 29260 26348 29316 26404
rect 29036 24556 29092 24612
rect 28924 23042 28980 23044
rect 28924 22990 28926 23042
rect 28926 22990 28978 23042
rect 28978 22990 28980 23042
rect 28924 22988 28980 22990
rect 29596 23826 29652 23828
rect 29596 23774 29598 23826
rect 29598 23774 29650 23826
rect 29650 23774 29652 23826
rect 29596 23772 29652 23774
rect 29148 21980 29204 22036
rect 28588 20748 28644 20804
rect 28700 21308 28756 21364
rect 28812 18732 28868 18788
rect 28924 20636 28980 20692
rect 28588 18172 28644 18228
rect 28140 15036 28196 15092
rect 28140 14642 28196 14644
rect 28140 14590 28142 14642
rect 28142 14590 28194 14642
rect 28194 14590 28196 14642
rect 28140 14588 28196 14590
rect 28700 16716 28756 16772
rect 28364 15314 28420 15316
rect 28364 15262 28366 15314
rect 28366 15262 28418 15314
rect 28418 15262 28420 15314
rect 28364 15260 28420 15262
rect 28588 15036 28644 15092
rect 29036 16156 29092 16212
rect 28924 16044 28980 16100
rect 29036 15874 29092 15876
rect 29036 15822 29038 15874
rect 29038 15822 29090 15874
rect 29090 15822 29092 15874
rect 29036 15820 29092 15822
rect 29260 18172 29316 18228
rect 29260 16044 29316 16100
rect 29148 15484 29204 15540
rect 29260 15260 29316 15316
rect 29372 15484 29428 15540
rect 28700 14588 28756 14644
rect 26684 13244 26740 13300
rect 26908 13356 26964 13412
rect 27356 13580 27412 13636
rect 27132 13356 27188 13412
rect 26460 12124 26516 12180
rect 26908 12012 26964 12068
rect 25340 11282 25396 11284
rect 25340 11230 25342 11282
rect 25342 11230 25394 11282
rect 25394 11230 25396 11282
rect 25340 11228 25396 11230
rect 25452 10556 25508 10612
rect 27020 10610 27076 10612
rect 27020 10558 27022 10610
rect 27022 10558 27074 10610
rect 27074 10558 27076 10610
rect 27020 10556 27076 10558
rect 25564 9996 25620 10052
rect 26572 9996 26628 10052
rect 25004 8988 25060 9044
rect 26236 8988 26292 9044
rect 29036 13634 29092 13636
rect 29036 13582 29038 13634
rect 29038 13582 29090 13634
rect 29090 13582 29092 13634
rect 29036 13580 29092 13582
rect 28588 13468 28644 13524
rect 28252 13074 28308 13076
rect 28252 13022 28254 13074
rect 28254 13022 28306 13074
rect 28306 13022 28308 13074
rect 28252 13020 28308 13022
rect 28700 13244 28756 13300
rect 27244 4284 27300 4340
rect 27132 4060 27188 4116
rect 26236 3612 26292 3668
rect 26796 3442 26852 3444
rect 26796 3390 26798 3442
rect 26798 3390 26850 3442
rect 26850 3390 26852 3442
rect 26796 3388 26852 3390
rect 27244 3554 27300 3556
rect 27244 3502 27246 3554
rect 27246 3502 27298 3554
rect 27298 3502 27300 3554
rect 27244 3500 27300 3502
rect 27580 3388 27636 3444
rect 29372 13074 29428 13076
rect 29372 13022 29374 13074
rect 29374 13022 29426 13074
rect 29426 13022 29428 13074
rect 29372 13020 29428 13022
rect 28140 12066 28196 12068
rect 28140 12014 28142 12066
rect 28142 12014 28194 12066
rect 28194 12014 28196 12066
rect 28140 12012 28196 12014
rect 28028 11340 28084 11396
rect 27916 9884 27972 9940
rect 27804 9042 27860 9044
rect 27804 8990 27806 9042
rect 27806 8990 27858 9042
rect 27858 8990 27860 9042
rect 27804 8988 27860 8990
rect 28140 9996 28196 10052
rect 28812 9996 28868 10052
rect 29372 11394 29428 11396
rect 29372 11342 29374 11394
rect 29374 11342 29426 11394
rect 29426 11342 29428 11394
rect 29372 11340 29428 11342
rect 29260 11228 29316 11284
rect 29260 9884 29316 9940
rect 28364 8988 28420 9044
rect 28700 9772 28756 9828
rect 28140 4114 28196 4116
rect 28140 4062 28142 4114
rect 28142 4062 28194 4114
rect 28194 4062 28196 4114
rect 28140 4060 28196 4062
rect 28364 3554 28420 3556
rect 28364 3502 28366 3554
rect 28366 3502 28418 3554
rect 28418 3502 28420 3554
rect 28364 3500 28420 3502
rect 29932 23714 29988 23716
rect 29932 23662 29934 23714
rect 29934 23662 29986 23714
rect 29986 23662 29988 23714
rect 29932 23660 29988 23662
rect 30268 27804 30324 27860
rect 30828 36428 30884 36484
rect 31164 37548 31220 37604
rect 31164 36988 31220 37044
rect 31612 38220 31668 38276
rect 31388 37378 31444 37380
rect 31388 37326 31390 37378
rect 31390 37326 31442 37378
rect 31442 37326 31444 37378
rect 31388 37324 31444 37326
rect 30716 36204 30772 36260
rect 30604 35026 30660 35028
rect 30604 34974 30606 35026
rect 30606 34974 30658 35026
rect 30658 34974 30660 35026
rect 30604 34972 30660 34974
rect 30940 33516 30996 33572
rect 30828 32620 30884 32676
rect 30716 32450 30772 32452
rect 30716 32398 30718 32450
rect 30718 32398 30770 32450
rect 30770 32398 30772 32450
rect 30716 32396 30772 32398
rect 30492 31276 30548 31332
rect 30940 31106 30996 31108
rect 30940 31054 30942 31106
rect 30942 31054 30994 31106
rect 30994 31054 30996 31106
rect 30940 31052 30996 31054
rect 30940 29596 30996 29652
rect 30492 29484 30548 29540
rect 31164 35308 31220 35364
rect 31276 35196 31332 35252
rect 31276 33404 31332 33460
rect 31164 33292 31220 33348
rect 31164 32844 31220 32900
rect 31276 32732 31332 32788
rect 31612 34802 31668 34804
rect 31612 34750 31614 34802
rect 31614 34750 31666 34802
rect 31666 34750 31668 34802
rect 31612 34748 31668 34750
rect 32396 39788 32452 39844
rect 32172 39564 32228 39620
rect 32396 39452 32452 39508
rect 32172 39058 32228 39060
rect 32172 39006 32174 39058
rect 32174 39006 32226 39058
rect 32226 39006 32228 39058
rect 32172 39004 32228 39006
rect 32508 39228 32564 39284
rect 32172 38556 32228 38612
rect 32732 42588 32788 42644
rect 33068 46956 33124 47012
rect 33404 49026 33460 49028
rect 33404 48974 33406 49026
rect 33406 48974 33458 49026
rect 33458 48974 33460 49026
rect 33404 48972 33460 48974
rect 33292 48242 33348 48244
rect 33292 48190 33294 48242
rect 33294 48190 33346 48242
rect 33346 48190 33348 48242
rect 33292 48188 33348 48190
rect 33516 47852 33572 47908
rect 33516 47068 33572 47124
rect 33180 46396 33236 46452
rect 33180 43260 33236 43316
rect 33180 42812 33236 42868
rect 32620 36988 32676 37044
rect 34076 53452 34132 53508
rect 33964 51772 34020 51828
rect 34076 51660 34132 51716
rect 33852 50764 33908 50820
rect 33740 48914 33796 48916
rect 33740 48862 33742 48914
rect 33742 48862 33794 48914
rect 33794 48862 33796 48914
rect 33740 48860 33796 48862
rect 33852 47852 33908 47908
rect 33740 46508 33796 46564
rect 33740 45948 33796 46004
rect 33628 45836 33684 45892
rect 33404 45724 33460 45780
rect 33516 45500 33572 45556
rect 33740 45276 33796 45332
rect 33404 44434 33460 44436
rect 33404 44382 33406 44434
rect 33406 44382 33458 44434
rect 33458 44382 33460 44434
rect 33404 44380 33460 44382
rect 33740 43538 33796 43540
rect 33740 43486 33742 43538
rect 33742 43486 33794 43538
rect 33794 43486 33796 43538
rect 33740 43484 33796 43486
rect 33628 42754 33684 42756
rect 33628 42702 33630 42754
rect 33630 42702 33682 42754
rect 33682 42702 33684 42754
rect 33628 42700 33684 42702
rect 33964 46956 34020 47012
rect 34412 55132 34468 55188
rect 34412 54796 34468 54852
rect 34636 58380 34692 58436
rect 34636 57484 34692 57540
rect 34860 58044 34916 58100
rect 34860 56812 34916 56868
rect 35532 59948 35588 60004
rect 35532 59778 35588 59780
rect 35532 59726 35534 59778
rect 35534 59726 35586 59778
rect 35586 59726 35588 59778
rect 35532 59724 35588 59726
rect 35196 58826 35252 58828
rect 35196 58774 35198 58826
rect 35198 58774 35250 58826
rect 35250 58774 35252 58826
rect 35196 58772 35252 58774
rect 35300 58826 35356 58828
rect 35300 58774 35302 58826
rect 35302 58774 35354 58826
rect 35354 58774 35356 58826
rect 35300 58772 35356 58774
rect 35404 58826 35460 58828
rect 35404 58774 35406 58826
rect 35406 58774 35458 58826
rect 35458 58774 35460 58826
rect 35404 58772 35460 58774
rect 35196 58492 35252 58548
rect 35756 59052 35812 59108
rect 35980 60284 36036 60340
rect 37660 65996 37716 66052
rect 37324 65436 37380 65492
rect 37212 64652 37268 64708
rect 37324 64092 37380 64148
rect 37996 64146 38052 64148
rect 37996 64094 37998 64146
rect 37998 64094 38050 64146
rect 38050 64094 38052 64146
rect 37996 64092 38052 64094
rect 37100 63756 37156 63812
rect 36876 62914 36932 62916
rect 36876 62862 36878 62914
rect 36878 62862 36930 62914
rect 36930 62862 36932 62914
rect 36876 62860 36932 62862
rect 37100 63420 37156 63476
rect 38892 65436 38948 65492
rect 38332 65212 38388 65268
rect 38332 64204 38388 64260
rect 38220 63756 38276 63812
rect 37884 63308 37940 63364
rect 37212 63138 37268 63140
rect 37212 63086 37214 63138
rect 37214 63086 37266 63138
rect 37266 63086 37268 63138
rect 37212 63084 37268 63086
rect 37884 63138 37940 63140
rect 37884 63086 37886 63138
rect 37886 63086 37938 63138
rect 37938 63086 37940 63138
rect 37884 63084 37940 63086
rect 37100 62636 37156 62692
rect 36204 61346 36260 61348
rect 36204 61294 36206 61346
rect 36206 61294 36258 61346
rect 36258 61294 36260 61346
rect 36204 61292 36260 61294
rect 36092 60172 36148 60228
rect 36428 60674 36484 60676
rect 36428 60622 36430 60674
rect 36430 60622 36482 60674
rect 36482 60622 36484 60674
rect 36428 60620 36484 60622
rect 36092 59612 36148 59668
rect 36988 60396 37044 60452
rect 36988 59276 37044 59332
rect 37100 59724 37156 59780
rect 35868 58940 35924 58996
rect 36316 58828 36372 58884
rect 35532 58268 35588 58324
rect 36092 58322 36148 58324
rect 36092 58270 36094 58322
rect 36094 58270 36146 58322
rect 36146 58270 36148 58322
rect 36092 58268 36148 58270
rect 35196 58156 35252 58212
rect 35644 58044 35700 58100
rect 35196 57258 35252 57260
rect 35196 57206 35198 57258
rect 35198 57206 35250 57258
rect 35250 57206 35252 57258
rect 35196 57204 35252 57206
rect 35300 57258 35356 57260
rect 35300 57206 35302 57258
rect 35302 57206 35354 57258
rect 35354 57206 35356 57258
rect 35300 57204 35356 57206
rect 35404 57258 35460 57260
rect 35404 57206 35406 57258
rect 35406 57206 35458 57258
rect 35458 57206 35460 57258
rect 35404 57204 35460 57206
rect 36428 58604 36484 58660
rect 34860 56642 34916 56644
rect 34860 56590 34862 56642
rect 34862 56590 34914 56642
rect 34914 56590 34916 56642
rect 34860 56588 34916 56590
rect 35196 55690 35252 55692
rect 35196 55638 35198 55690
rect 35198 55638 35250 55690
rect 35250 55638 35252 55690
rect 35196 55636 35252 55638
rect 35300 55690 35356 55692
rect 35300 55638 35302 55690
rect 35302 55638 35354 55690
rect 35354 55638 35356 55690
rect 35300 55636 35356 55638
rect 35404 55690 35460 55692
rect 35404 55638 35406 55690
rect 35406 55638 35458 55690
rect 35458 55638 35460 55690
rect 35404 55636 35460 55638
rect 36316 55468 36372 55524
rect 34972 55244 35028 55300
rect 34860 54684 34916 54740
rect 34636 54460 34692 54516
rect 34412 53564 34468 53620
rect 34748 54236 34804 54292
rect 35644 55020 35700 55076
rect 35868 55074 35924 55076
rect 35868 55022 35870 55074
rect 35870 55022 35922 55074
rect 35922 55022 35924 55074
rect 35868 55020 35924 55022
rect 34972 54348 35028 54404
rect 35084 54236 35140 54292
rect 35420 54290 35476 54292
rect 35420 54238 35422 54290
rect 35422 54238 35474 54290
rect 35474 54238 35476 54290
rect 35420 54236 35476 54238
rect 35196 54122 35252 54124
rect 35196 54070 35198 54122
rect 35198 54070 35250 54122
rect 35250 54070 35252 54122
rect 35196 54068 35252 54070
rect 35300 54122 35356 54124
rect 35300 54070 35302 54122
rect 35302 54070 35354 54122
rect 35354 54070 35356 54122
rect 35300 54068 35356 54070
rect 35404 54122 35460 54124
rect 35404 54070 35406 54122
rect 35406 54070 35458 54122
rect 35458 54070 35460 54122
rect 35404 54068 35460 54070
rect 35084 53788 35140 53844
rect 34860 53506 34916 53508
rect 34860 53454 34862 53506
rect 34862 53454 34914 53506
rect 34914 53454 34916 53506
rect 34860 53452 34916 53454
rect 34748 53228 34804 53284
rect 35196 53170 35252 53172
rect 35196 53118 35198 53170
rect 35198 53118 35250 53170
rect 35250 53118 35252 53170
rect 35196 53116 35252 53118
rect 35420 53228 35476 53284
rect 35756 54236 35812 54292
rect 35756 53900 35812 53956
rect 35980 53788 36036 53844
rect 35644 52892 35700 52948
rect 34972 52780 35028 52836
rect 35868 52780 35924 52836
rect 36428 54514 36484 54516
rect 36428 54462 36430 54514
rect 36430 54462 36482 54514
rect 36482 54462 36484 54514
rect 36428 54460 36484 54462
rect 36204 53788 36260 53844
rect 36204 53452 36260 53508
rect 36428 53900 36484 53956
rect 36092 53004 36148 53060
rect 36204 52780 36260 52836
rect 35196 52554 35252 52556
rect 35196 52502 35198 52554
rect 35198 52502 35250 52554
rect 35250 52502 35252 52554
rect 35196 52500 35252 52502
rect 35300 52554 35356 52556
rect 35300 52502 35302 52554
rect 35302 52502 35354 52554
rect 35354 52502 35356 52554
rect 35300 52500 35356 52502
rect 35404 52554 35460 52556
rect 35404 52502 35406 52554
rect 35406 52502 35458 52554
rect 35458 52502 35460 52554
rect 35404 52500 35460 52502
rect 34412 51884 34468 51940
rect 34748 51772 34804 51828
rect 36540 53676 36596 53732
rect 36540 52780 36596 52836
rect 35644 51436 35700 51492
rect 35196 50986 35252 50988
rect 35196 50934 35198 50986
rect 35198 50934 35250 50986
rect 35250 50934 35252 50986
rect 35196 50932 35252 50934
rect 35300 50986 35356 50988
rect 35300 50934 35302 50986
rect 35302 50934 35354 50986
rect 35354 50934 35356 50986
rect 35300 50932 35356 50934
rect 35404 50986 35460 50988
rect 35404 50934 35406 50986
rect 35406 50934 35458 50986
rect 35458 50934 35460 50986
rect 35404 50932 35460 50934
rect 36092 51266 36148 51268
rect 36092 51214 36094 51266
rect 36094 51214 36146 51266
rect 36146 51214 36148 51266
rect 36092 51212 36148 51214
rect 36876 58940 36932 58996
rect 37100 58828 37156 58884
rect 37100 56642 37156 56644
rect 37100 56590 37102 56642
rect 37102 56590 37154 56642
rect 37154 56590 37156 56642
rect 37100 56588 37156 56590
rect 36988 55468 37044 55524
rect 37100 55020 37156 55076
rect 36764 53564 36820 53620
rect 38108 63196 38164 63252
rect 38220 63084 38276 63140
rect 38444 62636 38500 62692
rect 38892 65100 38948 65156
rect 38892 64146 38948 64148
rect 38892 64094 38894 64146
rect 38894 64094 38946 64146
rect 38946 64094 38948 64146
rect 38892 64092 38948 64094
rect 38780 63810 38836 63812
rect 38780 63758 38782 63810
rect 38782 63758 38834 63810
rect 38834 63758 38836 63810
rect 38780 63756 38836 63758
rect 38892 63644 38948 63700
rect 38892 62860 38948 62916
rect 38556 62524 38612 62580
rect 37548 61292 37604 61348
rect 37324 60396 37380 60452
rect 37436 60732 37492 60788
rect 38220 59724 38276 59780
rect 37660 58604 37716 58660
rect 38220 58380 38276 58436
rect 38220 57932 38276 57988
rect 40348 70194 40404 70196
rect 40348 70142 40350 70194
rect 40350 70142 40402 70194
rect 40402 70142 40404 70194
rect 40348 70140 40404 70142
rect 41916 70700 41972 70756
rect 40460 69298 40516 69300
rect 40460 69246 40462 69298
rect 40462 69246 40514 69298
rect 40514 69246 40516 69298
rect 40460 69244 40516 69246
rect 40124 69132 40180 69188
rect 40124 68460 40180 68516
rect 39676 67564 39732 67620
rect 39676 67282 39732 67284
rect 39676 67230 39678 67282
rect 39678 67230 39730 67282
rect 39730 67230 39732 67282
rect 39676 67228 39732 67230
rect 40236 67618 40292 67620
rect 40236 67566 40238 67618
rect 40238 67566 40290 67618
rect 40290 67566 40292 67618
rect 40236 67564 40292 67566
rect 40908 68908 40964 68964
rect 41244 70140 41300 70196
rect 40460 68684 40516 68740
rect 40796 68460 40852 68516
rect 39116 66780 39172 66836
rect 39116 65212 39172 65268
rect 39340 65324 39396 65380
rect 39228 65100 39284 65156
rect 39340 64092 39396 64148
rect 39900 65996 39956 66052
rect 40572 66780 40628 66836
rect 41468 69468 41524 69524
rect 41356 68850 41412 68852
rect 41356 68798 41358 68850
rect 41358 68798 41410 68850
rect 41410 68798 41412 68850
rect 41356 68796 41412 68798
rect 41244 68738 41300 68740
rect 41244 68686 41246 68738
rect 41246 68686 41298 68738
rect 41298 68686 41300 68738
rect 41244 68684 41300 68686
rect 41132 66892 41188 66948
rect 41356 67116 41412 67172
rect 41468 66780 41524 66836
rect 42700 70754 42756 70756
rect 42700 70702 42702 70754
rect 42702 70702 42754 70754
rect 42754 70702 42756 70754
rect 42700 70700 42756 70702
rect 50556 70586 50612 70588
rect 50556 70534 50558 70586
rect 50558 70534 50610 70586
rect 50610 70534 50612 70586
rect 50556 70532 50612 70534
rect 50660 70586 50716 70588
rect 50660 70534 50662 70586
rect 50662 70534 50714 70586
rect 50714 70534 50716 70586
rect 50660 70532 50716 70534
rect 50764 70586 50820 70588
rect 50764 70534 50766 70586
rect 50766 70534 50818 70586
rect 50818 70534 50820 70586
rect 50764 70532 50820 70534
rect 43820 70140 43876 70196
rect 42588 69522 42644 69524
rect 42588 69470 42590 69522
rect 42590 69470 42642 69522
rect 42642 69470 42644 69522
rect 42588 69468 42644 69470
rect 42924 69186 42980 69188
rect 42924 69134 42926 69186
rect 42926 69134 42978 69186
rect 42978 69134 42980 69186
rect 42924 69132 42980 69134
rect 42364 68908 42420 68964
rect 41916 67564 41972 67620
rect 42028 67228 42084 67284
rect 41244 66274 41300 66276
rect 41244 66222 41246 66274
rect 41246 66222 41298 66274
rect 41298 66222 41300 66274
rect 41244 66220 41300 66222
rect 40348 66050 40404 66052
rect 40348 65998 40350 66050
rect 40350 65998 40402 66050
rect 40402 65998 40404 66050
rect 40348 65996 40404 65998
rect 40236 65490 40292 65492
rect 40236 65438 40238 65490
rect 40238 65438 40290 65490
rect 40290 65438 40292 65490
rect 40236 65436 40292 65438
rect 39900 65324 39956 65380
rect 40124 65212 40180 65268
rect 40124 64540 40180 64596
rect 41132 66050 41188 66052
rect 41132 65998 41134 66050
rect 41134 65998 41186 66050
rect 41186 65998 41188 66050
rect 41132 65996 41188 65998
rect 41916 66162 41972 66164
rect 41916 66110 41918 66162
rect 41918 66110 41970 66162
rect 41970 66110 41972 66162
rect 41916 66108 41972 66110
rect 41692 66050 41748 66052
rect 41692 65998 41694 66050
rect 41694 65998 41746 66050
rect 41746 65998 41748 66050
rect 41692 65996 41748 65998
rect 41692 65660 41748 65716
rect 41020 65378 41076 65380
rect 41020 65326 41022 65378
rect 41022 65326 41074 65378
rect 41074 65326 41076 65378
rect 41020 65324 41076 65326
rect 40460 64482 40516 64484
rect 40460 64430 40462 64482
rect 40462 64430 40514 64482
rect 40514 64430 40516 64482
rect 40460 64428 40516 64430
rect 41244 64876 41300 64932
rect 41020 64428 41076 64484
rect 40684 63868 40740 63924
rect 39788 63420 39844 63476
rect 40348 63644 40404 63700
rect 39116 63196 39172 63252
rect 40236 63250 40292 63252
rect 40236 63198 40238 63250
rect 40238 63198 40290 63250
rect 40290 63198 40292 63250
rect 40236 63196 40292 63198
rect 39452 62466 39508 62468
rect 39452 62414 39454 62466
rect 39454 62414 39506 62466
rect 39506 62414 39508 62466
rect 39452 62412 39508 62414
rect 40124 62636 40180 62692
rect 40012 62524 40068 62580
rect 39788 62300 39844 62356
rect 39900 62242 39956 62244
rect 39900 62190 39902 62242
rect 39902 62190 39954 62242
rect 39954 62190 39956 62242
rect 39900 62188 39956 62190
rect 40012 62076 40068 62132
rect 38444 59948 38500 60004
rect 38556 59890 38612 59892
rect 38556 59838 38558 59890
rect 38558 59838 38610 59890
rect 38610 59838 38612 59890
rect 38556 59836 38612 59838
rect 38444 59330 38500 59332
rect 38444 59278 38446 59330
rect 38446 59278 38498 59330
rect 38498 59278 38500 59330
rect 38444 59276 38500 59278
rect 38668 59218 38724 59220
rect 38668 59166 38670 59218
rect 38670 59166 38722 59218
rect 38722 59166 38724 59218
rect 38668 59164 38724 59166
rect 39116 60786 39172 60788
rect 39116 60734 39118 60786
rect 39118 60734 39170 60786
rect 39170 60734 39172 60786
rect 39116 60732 39172 60734
rect 39004 60674 39060 60676
rect 39004 60622 39006 60674
rect 39006 60622 39058 60674
rect 39058 60622 39060 60674
rect 39004 60620 39060 60622
rect 40460 62748 40516 62804
rect 40572 61682 40628 61684
rect 40572 61630 40574 61682
rect 40574 61630 40626 61682
rect 40626 61630 40628 61682
rect 40572 61628 40628 61630
rect 39340 60620 39396 60676
rect 39004 59948 39060 60004
rect 39564 59778 39620 59780
rect 39564 59726 39566 59778
rect 39566 59726 39618 59778
rect 39618 59726 39620 59778
rect 39564 59724 39620 59726
rect 39452 59612 39508 59668
rect 39340 59442 39396 59444
rect 39340 59390 39342 59442
rect 39342 59390 39394 59442
rect 39394 59390 39396 59442
rect 39340 59388 39396 59390
rect 38780 57932 38836 57988
rect 37660 56588 37716 56644
rect 38332 56642 38388 56644
rect 38332 56590 38334 56642
rect 38334 56590 38386 56642
rect 38386 56590 38388 56642
rect 38332 56588 38388 56590
rect 37996 56476 38052 56532
rect 38780 57484 38836 57540
rect 38668 55356 38724 55412
rect 37884 53900 37940 53956
rect 38220 53730 38276 53732
rect 38220 53678 38222 53730
rect 38222 53678 38274 53730
rect 38274 53678 38276 53730
rect 38220 53676 38276 53678
rect 37324 53506 37380 53508
rect 37324 53454 37326 53506
rect 37326 53454 37378 53506
rect 37378 53454 37380 53506
rect 37324 53452 37380 53454
rect 36764 53170 36820 53172
rect 36764 53118 36766 53170
rect 36766 53118 36818 53170
rect 36818 53118 36820 53170
rect 36764 53116 36820 53118
rect 37100 53004 37156 53060
rect 37212 52946 37268 52948
rect 37212 52894 37214 52946
rect 37214 52894 37266 52946
rect 37266 52894 37268 52946
rect 37212 52892 37268 52894
rect 36764 51212 36820 51268
rect 34300 48860 34356 48916
rect 35308 49810 35364 49812
rect 35308 49758 35310 49810
rect 35310 49758 35362 49810
rect 35362 49758 35364 49810
rect 35308 49756 35364 49758
rect 34636 49026 34692 49028
rect 34636 48974 34638 49026
rect 34638 48974 34690 49026
rect 34690 48974 34692 49026
rect 34636 48972 34692 48974
rect 34748 48748 34804 48804
rect 34412 48524 34468 48580
rect 34300 47628 34356 47684
rect 34188 46956 34244 47012
rect 34412 47180 34468 47236
rect 34076 46786 34132 46788
rect 34076 46734 34078 46786
rect 34078 46734 34130 46786
rect 34130 46734 34132 46786
rect 34076 46732 34132 46734
rect 34188 46674 34244 46676
rect 34188 46622 34190 46674
rect 34190 46622 34242 46674
rect 34242 46622 34244 46674
rect 34188 46620 34244 46622
rect 34076 45836 34132 45892
rect 33964 45388 34020 45444
rect 33964 45218 34020 45220
rect 33964 45166 33966 45218
rect 33966 45166 34018 45218
rect 34018 45166 34020 45218
rect 33964 45164 34020 45166
rect 34188 44716 34244 44772
rect 34412 44492 34468 44548
rect 34076 44380 34132 44436
rect 34748 47964 34804 48020
rect 34972 47404 35028 47460
rect 35196 49418 35252 49420
rect 35196 49366 35198 49418
rect 35198 49366 35250 49418
rect 35250 49366 35252 49418
rect 35196 49364 35252 49366
rect 35300 49418 35356 49420
rect 35300 49366 35302 49418
rect 35302 49366 35354 49418
rect 35354 49366 35356 49418
rect 35300 49364 35356 49366
rect 35404 49418 35460 49420
rect 35404 49366 35406 49418
rect 35406 49366 35458 49418
rect 35458 49366 35460 49418
rect 35404 49364 35460 49366
rect 36540 50034 36596 50036
rect 36540 49982 36542 50034
rect 36542 49982 36594 50034
rect 36594 49982 36596 50034
rect 36540 49980 36596 49982
rect 35756 49026 35812 49028
rect 35756 48974 35758 49026
rect 35758 48974 35810 49026
rect 35810 48974 35812 49026
rect 35756 48972 35812 48974
rect 36988 50764 37044 50820
rect 37212 50764 37268 50820
rect 36204 48972 36260 49028
rect 37100 49756 37156 49812
rect 35196 47850 35252 47852
rect 35196 47798 35198 47850
rect 35198 47798 35250 47850
rect 35250 47798 35252 47850
rect 35196 47796 35252 47798
rect 35300 47850 35356 47852
rect 35300 47798 35302 47850
rect 35302 47798 35354 47850
rect 35354 47798 35356 47850
rect 35300 47796 35356 47798
rect 35404 47850 35460 47852
rect 35404 47798 35406 47850
rect 35406 47798 35458 47850
rect 35458 47798 35460 47850
rect 35404 47796 35460 47798
rect 35756 48076 35812 48132
rect 35980 47628 36036 47684
rect 36204 48524 36260 48580
rect 34972 47234 35028 47236
rect 34972 47182 34974 47234
rect 34974 47182 35026 47234
rect 35026 47182 35028 47234
rect 34972 47180 35028 47182
rect 34636 46508 34692 46564
rect 34636 45890 34692 45892
rect 34636 45838 34638 45890
rect 34638 45838 34690 45890
rect 34690 45838 34692 45890
rect 34636 45836 34692 45838
rect 34636 45388 34692 45444
rect 34748 45276 34804 45332
rect 34972 46786 35028 46788
rect 34972 46734 34974 46786
rect 34974 46734 35026 46786
rect 35026 46734 35028 46786
rect 34972 46732 35028 46734
rect 35196 46674 35252 46676
rect 35196 46622 35198 46674
rect 35198 46622 35250 46674
rect 35250 46622 35252 46674
rect 35196 46620 35252 46622
rect 35196 46282 35252 46284
rect 35196 46230 35198 46282
rect 35198 46230 35250 46282
rect 35250 46230 35252 46282
rect 35196 46228 35252 46230
rect 35300 46282 35356 46284
rect 35300 46230 35302 46282
rect 35302 46230 35354 46282
rect 35354 46230 35356 46282
rect 35300 46228 35356 46230
rect 35404 46282 35460 46284
rect 35404 46230 35406 46282
rect 35406 46230 35458 46282
rect 35458 46230 35460 46282
rect 35404 46228 35460 46230
rect 35420 45948 35476 46004
rect 34972 45778 35028 45780
rect 34972 45726 34974 45778
rect 34974 45726 35026 45778
rect 35026 45726 35028 45778
rect 34972 45724 35028 45726
rect 36204 46844 36260 46900
rect 35308 45666 35364 45668
rect 35308 45614 35310 45666
rect 35310 45614 35362 45666
rect 35362 45614 35364 45666
rect 35308 45612 35364 45614
rect 35532 45500 35588 45556
rect 34972 45164 35028 45220
rect 36204 46284 36260 46340
rect 35868 45836 35924 45892
rect 35196 44714 35252 44716
rect 34524 44434 34580 44436
rect 34524 44382 34526 44434
rect 34526 44382 34578 44434
rect 34578 44382 34580 44434
rect 34524 44380 34580 44382
rect 34972 44604 35028 44660
rect 35196 44662 35198 44714
rect 35198 44662 35250 44714
rect 35250 44662 35252 44714
rect 35196 44660 35252 44662
rect 35300 44714 35356 44716
rect 35300 44662 35302 44714
rect 35302 44662 35354 44714
rect 35354 44662 35356 44714
rect 35300 44660 35356 44662
rect 35404 44714 35460 44716
rect 35404 44662 35406 44714
rect 35406 44662 35458 44714
rect 35458 44662 35460 44714
rect 35404 44660 35460 44662
rect 33964 43820 34020 43876
rect 34076 43148 34132 43204
rect 33404 42642 33460 42644
rect 33404 42590 33406 42642
rect 33406 42590 33458 42642
rect 33458 42590 33460 42642
rect 33404 42588 33460 42590
rect 33292 41916 33348 41972
rect 33404 41468 33460 41524
rect 33404 41132 33460 41188
rect 34188 42588 34244 42644
rect 34636 42754 34692 42756
rect 34636 42702 34638 42754
rect 34638 42702 34690 42754
rect 34690 42702 34692 42754
rect 34636 42700 34692 42702
rect 36204 45500 36260 45556
rect 35868 44434 35924 44436
rect 35868 44382 35870 44434
rect 35870 44382 35922 44434
rect 35922 44382 35924 44434
rect 35868 44380 35924 44382
rect 35308 44322 35364 44324
rect 35308 44270 35310 44322
rect 35310 44270 35362 44322
rect 35362 44270 35364 44322
rect 35308 44268 35364 44270
rect 35084 44210 35140 44212
rect 35084 44158 35086 44210
rect 35086 44158 35138 44210
rect 35138 44158 35140 44210
rect 35084 44156 35140 44158
rect 35308 43820 35364 43876
rect 35980 43650 36036 43652
rect 35980 43598 35982 43650
rect 35982 43598 36034 43650
rect 36034 43598 36036 43650
rect 35980 43596 36036 43598
rect 35196 43426 35252 43428
rect 35196 43374 35198 43426
rect 35198 43374 35250 43426
rect 35250 43374 35252 43426
rect 35196 43372 35252 43374
rect 35196 43146 35252 43148
rect 35196 43094 35198 43146
rect 35198 43094 35250 43146
rect 35250 43094 35252 43146
rect 35196 43092 35252 43094
rect 35300 43146 35356 43148
rect 35300 43094 35302 43146
rect 35302 43094 35354 43146
rect 35354 43094 35356 43146
rect 35300 43092 35356 43094
rect 35404 43146 35460 43148
rect 35404 43094 35406 43146
rect 35406 43094 35458 43146
rect 35458 43094 35460 43146
rect 35404 43092 35460 43094
rect 33964 41468 34020 41524
rect 34188 41132 34244 41188
rect 34860 41970 34916 41972
rect 34860 41918 34862 41970
rect 34862 41918 34914 41970
rect 34914 41918 34916 41970
rect 34860 41916 34916 41918
rect 34300 40908 34356 40964
rect 34748 40962 34804 40964
rect 34748 40910 34750 40962
rect 34750 40910 34802 40962
rect 34802 40910 34804 40962
rect 34748 40908 34804 40910
rect 34748 40572 34804 40628
rect 34188 40514 34244 40516
rect 34188 40462 34190 40514
rect 34190 40462 34242 40514
rect 34242 40462 34244 40514
rect 34188 40460 34244 40462
rect 33964 40402 34020 40404
rect 33964 40350 33966 40402
rect 33966 40350 34018 40402
rect 34018 40350 34020 40402
rect 33964 40348 34020 40350
rect 34412 40402 34468 40404
rect 34412 40350 34414 40402
rect 34414 40350 34466 40402
rect 34466 40350 34468 40402
rect 34412 40348 34468 40350
rect 34748 40348 34804 40404
rect 32508 35420 32564 35476
rect 31948 34802 32004 34804
rect 31948 34750 31950 34802
rect 31950 34750 32002 34802
rect 32002 34750 32004 34802
rect 31948 34748 32004 34750
rect 31500 33404 31556 33460
rect 32620 34188 32676 34244
rect 32060 33964 32116 34020
rect 32396 34018 32452 34020
rect 32396 33966 32398 34018
rect 32398 33966 32450 34018
rect 32450 33966 32452 34018
rect 32396 33964 32452 33966
rect 31836 33516 31892 33572
rect 32620 33458 32676 33460
rect 32620 33406 32622 33458
rect 32622 33406 32674 33458
rect 32674 33406 32676 33458
rect 32620 33404 32676 33406
rect 31388 32396 31444 32452
rect 31724 32844 31780 32900
rect 31612 32396 31668 32452
rect 31500 31724 31556 31780
rect 31500 31218 31556 31220
rect 31500 31166 31502 31218
rect 31502 31166 31554 31218
rect 31554 31166 31556 31218
rect 31500 31164 31556 31166
rect 31276 31052 31332 31108
rect 31164 30994 31220 30996
rect 31164 30942 31166 30994
rect 31166 30942 31218 30994
rect 31218 30942 31220 30994
rect 31164 30940 31220 30942
rect 31164 30156 31220 30212
rect 31052 29372 31108 29428
rect 30604 28642 30660 28644
rect 30604 28590 30606 28642
rect 30606 28590 30658 28642
rect 30658 28590 30660 28642
rect 30604 28588 30660 28590
rect 31612 29708 31668 29764
rect 32172 32732 32228 32788
rect 32284 33292 32340 33348
rect 31836 32620 31892 32676
rect 32172 32562 32228 32564
rect 32172 32510 32174 32562
rect 32174 32510 32226 32562
rect 32226 32510 32228 32562
rect 32172 32508 32228 32510
rect 32060 31948 32116 32004
rect 31836 30268 31892 30324
rect 31724 30044 31780 30100
rect 31500 29538 31556 29540
rect 31500 29486 31502 29538
rect 31502 29486 31554 29538
rect 31554 29486 31556 29538
rect 31500 29484 31556 29486
rect 31388 29314 31444 29316
rect 31388 29262 31390 29314
rect 31390 29262 31442 29314
rect 31442 29262 31444 29314
rect 31388 29260 31444 29262
rect 31164 28754 31220 28756
rect 31164 28702 31166 28754
rect 31166 28702 31218 28754
rect 31218 28702 31220 28754
rect 31164 28700 31220 28702
rect 30940 28476 30996 28532
rect 30604 28082 30660 28084
rect 30604 28030 30606 28082
rect 30606 28030 30658 28082
rect 30658 28030 30660 28082
rect 30604 28028 30660 28030
rect 31164 28364 31220 28420
rect 31948 29372 32004 29428
rect 32284 29650 32340 29652
rect 32284 29598 32286 29650
rect 32286 29598 32338 29650
rect 32338 29598 32340 29650
rect 32284 29596 32340 29598
rect 32172 29426 32228 29428
rect 32172 29374 32174 29426
rect 32174 29374 32226 29426
rect 32226 29374 32228 29426
rect 32172 29372 32228 29374
rect 32620 30380 32676 30436
rect 32508 30268 32564 30324
rect 32284 28588 32340 28644
rect 32172 28140 32228 28196
rect 32284 27970 32340 27972
rect 32284 27918 32286 27970
rect 32286 27918 32338 27970
rect 32338 27918 32340 27970
rect 32284 27916 32340 27918
rect 32956 36370 33012 36372
rect 32956 36318 32958 36370
rect 32958 36318 33010 36370
rect 33010 36318 33012 36370
rect 32956 36316 33012 36318
rect 33292 38556 33348 38612
rect 33852 38274 33908 38276
rect 33852 38222 33854 38274
rect 33854 38222 33906 38274
rect 33906 38222 33908 38274
rect 33852 38220 33908 38222
rect 34636 38220 34692 38276
rect 33516 38162 33572 38164
rect 33516 38110 33518 38162
rect 33518 38110 33570 38162
rect 33570 38110 33572 38162
rect 33516 38108 33572 38110
rect 33964 38162 34020 38164
rect 33964 38110 33966 38162
rect 33966 38110 34018 38162
rect 34018 38110 34020 38162
rect 33964 38108 34020 38110
rect 33852 37996 33908 38052
rect 33516 36316 33572 36372
rect 33628 35980 33684 36036
rect 33740 35922 33796 35924
rect 33740 35870 33742 35922
rect 33742 35870 33794 35922
rect 33794 35870 33796 35922
rect 33740 35868 33796 35870
rect 33180 35420 33236 35476
rect 33964 37884 34020 37940
rect 33180 34802 33236 34804
rect 33180 34750 33182 34802
rect 33182 34750 33234 34802
rect 33234 34750 33236 34802
rect 33180 34748 33236 34750
rect 33292 34690 33348 34692
rect 33292 34638 33294 34690
rect 33294 34638 33346 34690
rect 33346 34638 33348 34690
rect 33292 34636 33348 34638
rect 32844 33180 32900 33236
rect 33068 31500 33124 31556
rect 33068 30268 33124 30324
rect 33292 31948 33348 32004
rect 33404 31164 33460 31220
rect 33404 30210 33460 30212
rect 33404 30158 33406 30210
rect 33406 30158 33458 30210
rect 33458 30158 33460 30210
rect 33404 30156 33460 30158
rect 32732 29708 32788 29764
rect 32732 28588 32788 28644
rect 32844 29596 32900 29652
rect 32620 28252 32676 28308
rect 33068 29820 33124 29876
rect 32508 27186 32564 27188
rect 32508 27134 32510 27186
rect 32510 27134 32562 27186
rect 32562 27134 32564 27186
rect 32508 27132 32564 27134
rect 32620 27804 32676 27860
rect 30492 25340 30548 25396
rect 30268 24722 30324 24724
rect 30268 24670 30270 24722
rect 30270 24670 30322 24722
rect 30322 24670 30324 24722
rect 30268 24668 30324 24670
rect 30156 22988 30212 23044
rect 31052 25004 31108 25060
rect 31724 25394 31780 25396
rect 31724 25342 31726 25394
rect 31726 25342 31778 25394
rect 31778 25342 31780 25394
rect 31724 25340 31780 25342
rect 31724 25004 31780 25060
rect 31500 24780 31556 24836
rect 31164 23660 31220 23716
rect 30268 21980 30324 22036
rect 29708 20188 29764 20244
rect 30044 21474 30100 21476
rect 30044 21422 30046 21474
rect 30046 21422 30098 21474
rect 30098 21422 30100 21474
rect 30044 21420 30100 21422
rect 29596 19010 29652 19012
rect 29596 18958 29598 19010
rect 29598 18958 29650 19010
rect 29650 18958 29652 19010
rect 29596 18956 29652 18958
rect 29708 18508 29764 18564
rect 29932 17724 29988 17780
rect 30828 22988 30884 23044
rect 30716 22428 30772 22484
rect 30492 21532 30548 21588
rect 30604 21420 30660 21476
rect 30492 21362 30548 21364
rect 30492 21310 30494 21362
rect 30494 21310 30546 21362
rect 30546 21310 30548 21362
rect 30492 21308 30548 21310
rect 30380 21196 30436 21252
rect 30828 22316 30884 22372
rect 31164 22652 31220 22708
rect 31164 21756 31220 21812
rect 31500 21532 31556 21588
rect 31948 24668 32004 24724
rect 32172 25340 32228 25396
rect 32396 24610 32452 24612
rect 32396 24558 32398 24610
rect 32398 24558 32450 24610
rect 32450 24558 32452 24610
rect 32396 24556 32452 24558
rect 31836 23212 31892 23268
rect 31836 22092 31892 22148
rect 32284 23772 32340 23828
rect 31500 20524 31556 20580
rect 31276 20188 31332 20244
rect 30380 19964 30436 20020
rect 31164 20018 31220 20020
rect 31164 19966 31166 20018
rect 31166 19966 31218 20018
rect 31218 19966 31220 20018
rect 31164 19964 31220 19966
rect 30492 19010 30548 19012
rect 30492 18958 30494 19010
rect 30494 18958 30546 19010
rect 30546 18958 30548 19010
rect 30492 18956 30548 18958
rect 30380 18508 30436 18564
rect 29820 17500 29876 17556
rect 30268 18396 30324 18452
rect 30268 17164 30324 17220
rect 30604 16828 30660 16884
rect 30044 16604 30100 16660
rect 29596 15708 29652 15764
rect 30604 16210 30660 16212
rect 30604 16158 30606 16210
rect 30606 16158 30658 16210
rect 30658 16158 30660 16210
rect 30604 16156 30660 16158
rect 30044 15596 30100 15652
rect 31724 20076 31780 20132
rect 31388 19852 31444 19908
rect 30828 17778 30884 17780
rect 30828 17726 30830 17778
rect 30830 17726 30882 17778
rect 30882 17726 30884 17778
rect 30828 17724 30884 17726
rect 31388 17612 31444 17668
rect 31500 18396 31556 18452
rect 31388 17442 31444 17444
rect 31388 17390 31390 17442
rect 31390 17390 31442 17442
rect 31442 17390 31444 17442
rect 31388 17388 31444 17390
rect 31388 17164 31444 17220
rect 30828 17106 30884 17108
rect 30828 17054 30830 17106
rect 30830 17054 30882 17106
rect 30882 17054 30884 17106
rect 30828 17052 30884 17054
rect 32396 22370 32452 22372
rect 32396 22318 32398 22370
rect 32398 22318 32450 22370
rect 32450 22318 32452 22370
rect 32396 22316 32452 22318
rect 32396 22092 32452 22148
rect 31948 19906 32004 19908
rect 31948 19854 31950 19906
rect 31950 19854 32002 19906
rect 32002 19854 32004 19906
rect 31948 19852 32004 19854
rect 31836 19068 31892 19124
rect 31612 17554 31668 17556
rect 31612 17502 31614 17554
rect 31614 17502 31666 17554
rect 31666 17502 31668 17554
rect 31612 17500 31668 17502
rect 29932 14530 29988 14532
rect 29932 14478 29934 14530
rect 29934 14478 29986 14530
rect 29986 14478 29988 14530
rect 29932 14476 29988 14478
rect 29708 14364 29764 14420
rect 29596 13580 29652 13636
rect 30828 15372 30884 15428
rect 30268 14812 30324 14868
rect 30268 13468 30324 13524
rect 31500 15148 31556 15204
rect 30604 14530 30660 14532
rect 30604 14478 30606 14530
rect 30606 14478 30658 14530
rect 30658 14478 30660 14530
rect 30604 14476 30660 14478
rect 30828 14418 30884 14420
rect 30828 14366 30830 14418
rect 30830 14366 30882 14418
rect 30882 14366 30884 14418
rect 30828 14364 30884 14366
rect 31164 14364 31220 14420
rect 31276 14476 31332 14532
rect 31388 13468 31444 13524
rect 29708 12178 29764 12180
rect 29708 12126 29710 12178
rect 29710 12126 29762 12178
rect 29762 12126 29764 12178
rect 29708 12124 29764 12126
rect 29708 9602 29764 9604
rect 29708 9550 29710 9602
rect 29710 9550 29762 9602
rect 29762 9550 29764 9602
rect 29708 9548 29764 9550
rect 30828 12178 30884 12180
rect 30828 12126 30830 12178
rect 30830 12126 30882 12178
rect 30882 12126 30884 12178
rect 30828 12124 30884 12126
rect 30716 11340 30772 11396
rect 30716 10668 30772 10724
rect 30380 9548 30436 9604
rect 29372 3666 29428 3668
rect 29372 3614 29374 3666
rect 29374 3614 29426 3666
rect 29426 3614 29428 3666
rect 29372 3612 29428 3614
rect 30828 10108 30884 10164
rect 30828 8876 30884 8932
rect 31276 12290 31332 12292
rect 31276 12238 31278 12290
rect 31278 12238 31330 12290
rect 31330 12238 31332 12290
rect 31276 12236 31332 12238
rect 31052 11394 31108 11396
rect 31052 11342 31054 11394
rect 31054 11342 31106 11394
rect 31106 11342 31108 11394
rect 31052 11340 31108 11342
rect 31500 12962 31556 12964
rect 31500 12910 31502 12962
rect 31502 12910 31554 12962
rect 31554 12910 31556 12962
rect 31500 12908 31556 12910
rect 32284 18450 32340 18452
rect 32284 18398 32286 18450
rect 32286 18398 32338 18450
rect 32338 18398 32340 18450
rect 32284 18396 32340 18398
rect 31948 17052 32004 17108
rect 32060 17164 32116 17220
rect 32284 17612 32340 17668
rect 31948 16882 32004 16884
rect 31948 16830 31950 16882
rect 31950 16830 32002 16882
rect 32002 16830 32004 16882
rect 31948 16828 32004 16830
rect 31724 16604 31780 16660
rect 31724 15932 31780 15988
rect 32172 15708 32228 15764
rect 32060 15596 32116 15652
rect 32732 24050 32788 24052
rect 32732 23998 32734 24050
rect 32734 23998 32786 24050
rect 32786 23998 32788 24050
rect 32732 23996 32788 23998
rect 33068 24668 33124 24724
rect 33292 27356 33348 27412
rect 33292 27074 33348 27076
rect 33292 27022 33294 27074
rect 33294 27022 33346 27074
rect 33346 27022 33348 27074
rect 33292 27020 33348 27022
rect 33628 33292 33684 33348
rect 33852 34690 33908 34692
rect 33852 34638 33854 34690
rect 33854 34638 33906 34690
rect 33906 34638 33908 34690
rect 33852 34636 33908 34638
rect 33852 34412 33908 34468
rect 33740 31500 33796 31556
rect 33852 31106 33908 31108
rect 33852 31054 33854 31106
rect 33854 31054 33906 31106
rect 33906 31054 33908 31106
rect 33852 31052 33908 31054
rect 33628 30268 33684 30324
rect 33628 29820 33684 29876
rect 34524 37826 34580 37828
rect 34524 37774 34526 37826
rect 34526 37774 34578 37826
rect 34578 37774 34580 37826
rect 34524 37772 34580 37774
rect 34412 35980 34468 36036
rect 34524 35810 34580 35812
rect 34524 35758 34526 35810
rect 34526 35758 34578 35810
rect 34578 35758 34580 35810
rect 34524 35756 34580 35758
rect 34300 35644 34356 35700
rect 35084 42588 35140 42644
rect 35644 41692 35700 41748
rect 35196 41578 35252 41580
rect 35196 41526 35198 41578
rect 35198 41526 35250 41578
rect 35250 41526 35252 41578
rect 35196 41524 35252 41526
rect 35300 41578 35356 41580
rect 35300 41526 35302 41578
rect 35302 41526 35354 41578
rect 35354 41526 35356 41578
rect 35300 41524 35356 41526
rect 35404 41578 35460 41580
rect 35404 41526 35406 41578
rect 35406 41526 35458 41578
rect 35458 41526 35460 41578
rect 35404 41524 35460 41526
rect 35196 41186 35252 41188
rect 35196 41134 35198 41186
rect 35198 41134 35250 41186
rect 35250 41134 35252 41186
rect 35196 41132 35252 41134
rect 36428 48802 36484 48804
rect 36428 48750 36430 48802
rect 36430 48750 36482 48802
rect 36482 48750 36484 48802
rect 36428 48748 36484 48750
rect 37100 48636 37156 48692
rect 36876 48076 36932 48132
rect 36764 46562 36820 46564
rect 36764 46510 36766 46562
rect 36766 46510 36818 46562
rect 36818 46510 36820 46562
rect 36764 46508 36820 46510
rect 36988 47458 37044 47460
rect 36988 47406 36990 47458
rect 36990 47406 37042 47458
rect 37042 47406 37044 47458
rect 36988 47404 37044 47406
rect 37212 48802 37268 48804
rect 37212 48750 37214 48802
rect 37214 48750 37266 48802
rect 37266 48750 37268 48802
rect 37212 48748 37268 48750
rect 37212 47628 37268 47684
rect 37436 53170 37492 53172
rect 37436 53118 37438 53170
rect 37438 53118 37490 53170
rect 37490 53118 37492 53170
rect 37436 53116 37492 53118
rect 37996 53116 38052 53172
rect 37548 52946 37604 52948
rect 37548 52894 37550 52946
rect 37550 52894 37602 52946
rect 37602 52894 37604 52946
rect 37548 52892 37604 52894
rect 39116 59164 39172 59220
rect 39564 59442 39620 59444
rect 39564 59390 39566 59442
rect 39566 59390 39618 59442
rect 39618 59390 39620 59442
rect 39564 59388 39620 59390
rect 39788 60002 39844 60004
rect 39788 59950 39790 60002
rect 39790 59950 39842 60002
rect 39842 59950 39844 60002
rect 39788 59948 39844 59950
rect 40012 60396 40068 60452
rect 40348 60674 40404 60676
rect 40348 60622 40350 60674
rect 40350 60622 40402 60674
rect 40402 60622 40404 60674
rect 40348 60620 40404 60622
rect 40012 60172 40068 60228
rect 40012 59724 40068 59780
rect 40012 59218 40068 59220
rect 40012 59166 40014 59218
rect 40014 59166 40066 59218
rect 40066 59166 40068 59218
rect 40012 59164 40068 59166
rect 39900 59052 39956 59108
rect 39004 57372 39060 57428
rect 39116 57148 39172 57204
rect 39116 56140 39172 56196
rect 39564 58546 39620 58548
rect 39564 58494 39566 58546
rect 39566 58494 39618 58546
rect 39618 58494 39620 58546
rect 39564 58492 39620 58494
rect 39340 56978 39396 56980
rect 39340 56926 39342 56978
rect 39342 56926 39394 56978
rect 39394 56926 39396 56978
rect 39340 56924 39396 56926
rect 39452 57372 39508 57428
rect 38668 52220 38724 52276
rect 38108 52108 38164 52164
rect 37996 51490 38052 51492
rect 37996 51438 37998 51490
rect 37998 51438 38050 51490
rect 38050 51438 38052 51490
rect 37996 51436 38052 51438
rect 37884 51378 37940 51380
rect 37884 51326 37886 51378
rect 37886 51326 37938 51378
rect 37938 51326 37940 51378
rect 37884 51324 37940 51326
rect 37996 51154 38052 51156
rect 37996 51102 37998 51154
rect 37998 51102 38050 51154
rect 38050 51102 38052 51154
rect 37996 51100 38052 51102
rect 38444 52162 38500 52164
rect 38444 52110 38446 52162
rect 38446 52110 38498 52162
rect 38498 52110 38500 52162
rect 38444 52108 38500 52110
rect 38892 52274 38948 52276
rect 38892 52222 38894 52274
rect 38894 52222 38946 52274
rect 38946 52222 38948 52274
rect 38892 52220 38948 52222
rect 38780 51660 38836 51716
rect 39004 51602 39060 51604
rect 39004 51550 39006 51602
rect 39006 51550 39058 51602
rect 39058 51550 39060 51602
rect 39004 51548 39060 51550
rect 38108 50428 38164 50484
rect 37548 49980 37604 50036
rect 37436 48636 37492 48692
rect 37548 48412 37604 48468
rect 37996 49980 38052 50036
rect 38220 49922 38276 49924
rect 38220 49870 38222 49922
rect 38222 49870 38274 49922
rect 38274 49870 38276 49922
rect 38220 49868 38276 49870
rect 38108 49026 38164 49028
rect 38108 48974 38110 49026
rect 38110 48974 38162 49026
rect 38162 48974 38164 49026
rect 38108 48972 38164 48974
rect 37884 48748 37940 48804
rect 37772 47964 37828 48020
rect 37324 47852 37380 47908
rect 38220 48636 38276 48692
rect 38332 48412 38388 48468
rect 38108 47682 38164 47684
rect 38108 47630 38110 47682
rect 38110 47630 38162 47682
rect 38162 47630 38164 47682
rect 38108 47628 38164 47630
rect 37996 47234 38052 47236
rect 37996 47182 37998 47234
rect 37998 47182 38050 47234
rect 38050 47182 38052 47234
rect 37996 47180 38052 47182
rect 38444 48354 38500 48356
rect 38444 48302 38446 48354
rect 38446 48302 38498 48354
rect 38498 48302 38500 48354
rect 38444 48300 38500 48302
rect 38444 47404 38500 47460
rect 38332 47180 38388 47236
rect 37212 46620 37268 46676
rect 36988 46396 37044 46452
rect 36428 46002 36484 46004
rect 36428 45950 36430 46002
rect 36430 45950 36482 46002
rect 36482 45950 36484 46002
rect 36428 45948 36484 45950
rect 37212 45388 37268 45444
rect 37772 45948 37828 46004
rect 37100 45276 37156 45332
rect 37100 44156 37156 44212
rect 37436 45164 37492 45220
rect 36428 42642 36484 42644
rect 36428 42590 36430 42642
rect 36430 42590 36482 42642
rect 36482 42590 36484 42642
rect 36428 42588 36484 42590
rect 36764 42364 36820 42420
rect 35868 40908 35924 40964
rect 35532 40796 35588 40852
rect 35308 40626 35364 40628
rect 35308 40574 35310 40626
rect 35310 40574 35362 40626
rect 35362 40574 35364 40626
rect 35308 40572 35364 40574
rect 35196 40402 35252 40404
rect 35196 40350 35198 40402
rect 35198 40350 35250 40402
rect 35250 40350 35252 40402
rect 35196 40348 35252 40350
rect 34748 35868 34804 35924
rect 34748 35532 34804 35588
rect 35196 40010 35252 40012
rect 35196 39958 35198 40010
rect 35198 39958 35250 40010
rect 35250 39958 35252 40010
rect 35196 39956 35252 39958
rect 35300 40010 35356 40012
rect 35300 39958 35302 40010
rect 35302 39958 35354 40010
rect 35354 39958 35356 40010
rect 35300 39956 35356 39958
rect 35404 40010 35460 40012
rect 35404 39958 35406 40010
rect 35406 39958 35458 40010
rect 35458 39958 35460 40010
rect 35404 39956 35460 39958
rect 36316 40572 36372 40628
rect 35756 40514 35812 40516
rect 35756 40462 35758 40514
rect 35758 40462 35810 40514
rect 35810 40462 35812 40514
rect 35756 40460 35812 40462
rect 36204 40402 36260 40404
rect 36204 40350 36206 40402
rect 36206 40350 36258 40402
rect 36258 40350 36260 40402
rect 36204 40348 36260 40350
rect 36092 39452 36148 39508
rect 35532 38556 35588 38612
rect 35196 38442 35252 38444
rect 35196 38390 35198 38442
rect 35198 38390 35250 38442
rect 35250 38390 35252 38442
rect 35196 38388 35252 38390
rect 35300 38442 35356 38444
rect 35300 38390 35302 38442
rect 35302 38390 35354 38442
rect 35354 38390 35356 38442
rect 35300 38388 35356 38390
rect 35404 38442 35460 38444
rect 35404 38390 35406 38442
rect 35406 38390 35458 38442
rect 35458 38390 35460 38442
rect 35404 38388 35460 38390
rect 35420 37826 35476 37828
rect 35420 37774 35422 37826
rect 35422 37774 35474 37826
rect 35474 37774 35476 37826
rect 35420 37772 35476 37774
rect 35196 36874 35252 36876
rect 35196 36822 35198 36874
rect 35198 36822 35250 36874
rect 35250 36822 35252 36874
rect 35196 36820 35252 36822
rect 35300 36874 35356 36876
rect 35300 36822 35302 36874
rect 35302 36822 35354 36874
rect 35354 36822 35356 36874
rect 35300 36820 35356 36822
rect 35404 36874 35460 36876
rect 35404 36822 35406 36874
rect 35406 36822 35458 36874
rect 35458 36822 35460 36874
rect 35404 36820 35460 36822
rect 37324 42700 37380 42756
rect 37324 42476 37380 42532
rect 36764 41970 36820 41972
rect 36764 41918 36766 41970
rect 36766 41918 36818 41970
rect 36818 41918 36820 41970
rect 36764 41916 36820 41918
rect 36876 39452 36932 39508
rect 35644 35868 35700 35924
rect 35084 35756 35140 35812
rect 35532 35644 35588 35700
rect 35196 35306 35252 35308
rect 35196 35254 35198 35306
rect 35198 35254 35250 35306
rect 35250 35254 35252 35306
rect 35196 35252 35252 35254
rect 35300 35306 35356 35308
rect 35300 35254 35302 35306
rect 35302 35254 35354 35306
rect 35354 35254 35356 35306
rect 35300 35252 35356 35254
rect 35404 35306 35460 35308
rect 35404 35254 35406 35306
rect 35406 35254 35458 35306
rect 35458 35254 35460 35306
rect 35404 35252 35460 35254
rect 34188 34412 34244 34468
rect 35420 34802 35476 34804
rect 35420 34750 35422 34802
rect 35422 34750 35474 34802
rect 35474 34750 35476 34802
rect 35420 34748 35476 34750
rect 35308 34690 35364 34692
rect 35308 34638 35310 34690
rect 35310 34638 35362 34690
rect 35362 34638 35364 34690
rect 35308 34636 35364 34638
rect 34412 34300 34468 34356
rect 34076 33292 34132 33348
rect 34188 33122 34244 33124
rect 34188 33070 34190 33122
rect 34190 33070 34242 33122
rect 34242 33070 34244 33122
rect 34188 33068 34244 33070
rect 35084 33964 35140 34020
rect 35868 35084 35924 35140
rect 36540 35756 36596 35812
rect 35756 34802 35812 34804
rect 35756 34750 35758 34802
rect 35758 34750 35810 34802
rect 35810 34750 35812 34802
rect 35756 34748 35812 34750
rect 35196 33738 35252 33740
rect 35196 33686 35198 33738
rect 35198 33686 35250 33738
rect 35250 33686 35252 33738
rect 35196 33684 35252 33686
rect 35300 33738 35356 33740
rect 35300 33686 35302 33738
rect 35302 33686 35354 33738
rect 35354 33686 35356 33738
rect 35300 33684 35356 33686
rect 35404 33738 35460 33740
rect 35404 33686 35406 33738
rect 35406 33686 35458 33738
rect 35458 33686 35460 33738
rect 35404 33684 35460 33686
rect 35532 33516 35588 33572
rect 36428 34636 36484 34692
rect 35868 33404 35924 33460
rect 35084 33346 35140 33348
rect 35084 33294 35086 33346
rect 35086 33294 35138 33346
rect 35138 33294 35140 33346
rect 35084 33292 35140 33294
rect 34188 32786 34244 32788
rect 34188 32734 34190 32786
rect 34190 32734 34242 32786
rect 34242 32734 34244 32786
rect 34188 32732 34244 32734
rect 35532 33122 35588 33124
rect 35532 33070 35534 33122
rect 35534 33070 35586 33122
rect 35586 33070 35588 33122
rect 35532 33068 35588 33070
rect 34412 32786 34468 32788
rect 34412 32734 34414 32786
rect 34414 32734 34466 32786
rect 34466 32734 34468 32786
rect 34412 32732 34468 32734
rect 34300 32508 34356 32564
rect 34076 30210 34132 30212
rect 34076 30158 34078 30210
rect 34078 30158 34130 30210
rect 34130 30158 34132 30210
rect 34076 30156 34132 30158
rect 34076 29820 34132 29876
rect 33516 27804 33572 27860
rect 33292 26236 33348 26292
rect 33404 26124 33460 26180
rect 33292 24780 33348 24836
rect 33292 23996 33348 24052
rect 33404 24556 33460 24612
rect 33180 22428 33236 22484
rect 33068 21810 33124 21812
rect 33068 21758 33070 21810
rect 33070 21758 33122 21810
rect 33122 21758 33124 21810
rect 33068 21756 33124 21758
rect 32844 18396 32900 18452
rect 33068 18620 33124 18676
rect 32844 17612 32900 17668
rect 32620 16156 32676 16212
rect 32508 15314 32564 15316
rect 32508 15262 32510 15314
rect 32510 15262 32562 15314
rect 32562 15262 32564 15314
rect 32508 15260 32564 15262
rect 33180 17724 33236 17780
rect 33180 17164 33236 17220
rect 33068 15820 33124 15876
rect 33516 20524 33572 20580
rect 33740 28418 33796 28420
rect 33740 28366 33742 28418
rect 33742 28366 33794 28418
rect 33794 28366 33796 28418
rect 33740 28364 33796 28366
rect 33740 27244 33796 27300
rect 34412 29538 34468 29540
rect 34412 29486 34414 29538
rect 34414 29486 34466 29538
rect 34466 29486 34468 29538
rect 34412 29484 34468 29486
rect 35196 32844 35252 32900
rect 35980 33068 36036 33124
rect 34748 32284 34804 32340
rect 35196 32170 35252 32172
rect 35196 32118 35198 32170
rect 35198 32118 35250 32170
rect 35250 32118 35252 32170
rect 35196 32116 35252 32118
rect 35300 32170 35356 32172
rect 35300 32118 35302 32170
rect 35302 32118 35354 32170
rect 35354 32118 35356 32170
rect 35300 32116 35356 32118
rect 35404 32170 35460 32172
rect 35404 32118 35406 32170
rect 35406 32118 35458 32170
rect 35458 32118 35460 32170
rect 35404 32116 35460 32118
rect 35420 31948 35476 32004
rect 34748 30268 34804 30324
rect 34188 28364 34244 28420
rect 34188 27020 34244 27076
rect 34524 28642 34580 28644
rect 34524 28590 34526 28642
rect 34526 28590 34578 28642
rect 34578 28590 34580 28642
rect 34524 28588 34580 28590
rect 34412 27356 34468 27412
rect 34524 27074 34580 27076
rect 34524 27022 34526 27074
rect 34526 27022 34578 27074
rect 34578 27022 34580 27074
rect 34524 27020 34580 27022
rect 35644 32562 35700 32564
rect 35644 32510 35646 32562
rect 35646 32510 35698 32562
rect 35698 32510 35700 32562
rect 35644 32508 35700 32510
rect 37324 41970 37380 41972
rect 37324 41918 37326 41970
rect 37326 41918 37378 41970
rect 37378 41918 37380 41970
rect 37324 41916 37380 41918
rect 37212 40626 37268 40628
rect 37212 40574 37214 40626
rect 37214 40574 37266 40626
rect 37266 40574 37268 40626
rect 37212 40572 37268 40574
rect 37772 45388 37828 45444
rect 38108 45276 38164 45332
rect 38892 51378 38948 51380
rect 38892 51326 38894 51378
rect 38894 51326 38946 51378
rect 38946 51326 38948 51378
rect 38892 51324 38948 51326
rect 40460 59388 40516 59444
rect 39788 57148 39844 57204
rect 40460 58156 40516 58212
rect 40572 57820 40628 57876
rect 40348 57538 40404 57540
rect 40348 57486 40350 57538
rect 40350 57486 40402 57538
rect 40402 57486 40404 57538
rect 40348 57484 40404 57486
rect 40124 56924 40180 56980
rect 40236 57036 40292 57092
rect 40236 56588 40292 56644
rect 39900 54460 39956 54516
rect 40124 53730 40180 53732
rect 40124 53678 40126 53730
rect 40126 53678 40178 53730
rect 40178 53678 40180 53730
rect 40124 53676 40180 53678
rect 39564 52892 39620 52948
rect 39228 51996 39284 52052
rect 39564 51660 39620 51716
rect 39228 51548 39284 51604
rect 38668 49868 38724 49924
rect 39452 51378 39508 51380
rect 39452 51326 39454 51378
rect 39454 51326 39506 51378
rect 39506 51326 39508 51378
rect 39452 51324 39508 51326
rect 38668 49644 38724 49700
rect 38668 48748 38724 48804
rect 38668 47404 38724 47460
rect 38556 45948 38612 46004
rect 39228 50988 39284 51044
rect 38892 50876 38948 50932
rect 39340 50204 39396 50260
rect 39228 49922 39284 49924
rect 39228 49870 39230 49922
rect 39230 49870 39282 49922
rect 39282 49870 39284 49922
rect 39228 49868 39284 49870
rect 39900 51378 39956 51380
rect 39900 51326 39902 51378
rect 39902 51326 39954 51378
rect 39954 51326 39956 51378
rect 39900 51324 39956 51326
rect 40012 51212 40068 51268
rect 39564 50876 39620 50932
rect 39676 51100 39732 51156
rect 39340 49644 39396 49700
rect 39564 49084 39620 49140
rect 39116 48802 39172 48804
rect 39116 48750 39118 48802
rect 39118 48750 39170 48802
rect 39170 48750 39172 48802
rect 39116 48748 39172 48750
rect 39116 48466 39172 48468
rect 39116 48414 39118 48466
rect 39118 48414 39170 48466
rect 39170 48414 39172 48466
rect 39116 48412 39172 48414
rect 39340 48242 39396 48244
rect 39340 48190 39342 48242
rect 39342 48190 39394 48242
rect 39394 48190 39396 48242
rect 39340 48188 39396 48190
rect 39228 48130 39284 48132
rect 39228 48078 39230 48130
rect 39230 48078 39282 48130
rect 39282 48078 39284 48130
rect 39228 48076 39284 48078
rect 38892 47570 38948 47572
rect 38892 47518 38894 47570
rect 38894 47518 38946 47570
rect 38946 47518 38948 47570
rect 38892 47516 38948 47518
rect 37660 42754 37716 42756
rect 37660 42702 37662 42754
rect 37662 42702 37714 42754
rect 37714 42702 37716 42754
rect 37660 42700 37716 42702
rect 37548 41970 37604 41972
rect 37548 41918 37550 41970
rect 37550 41918 37602 41970
rect 37602 41918 37604 41970
rect 37548 41916 37604 41918
rect 37996 43148 38052 43204
rect 37884 42812 37940 42868
rect 38668 44210 38724 44212
rect 38668 44158 38670 44210
rect 38670 44158 38722 44210
rect 38722 44158 38724 44210
rect 38668 44156 38724 44158
rect 38332 43484 38388 43540
rect 38780 43372 38836 43428
rect 38668 43148 38724 43204
rect 38332 42754 38388 42756
rect 38332 42702 38334 42754
rect 38334 42702 38386 42754
rect 38386 42702 38388 42754
rect 38332 42700 38388 42702
rect 40572 57372 40628 57428
rect 40348 55970 40404 55972
rect 40348 55918 40350 55970
rect 40350 55918 40402 55970
rect 40402 55918 40404 55970
rect 40348 55916 40404 55918
rect 40460 53116 40516 53172
rect 41244 64316 41300 64372
rect 41356 63922 41412 63924
rect 41356 63870 41358 63922
rect 41358 63870 41410 63922
rect 41410 63870 41412 63922
rect 41356 63868 41412 63870
rect 40796 63756 40852 63812
rect 42252 66892 42308 66948
rect 42476 66780 42532 66836
rect 42588 67116 42644 67172
rect 42476 66220 42532 66276
rect 43260 67170 43316 67172
rect 43260 67118 43262 67170
rect 43262 67118 43314 67170
rect 43314 67118 43316 67170
rect 43260 67116 43316 67118
rect 44156 69186 44212 69188
rect 44156 69134 44158 69186
rect 44158 69134 44210 69186
rect 44210 69134 44212 69186
rect 44156 69132 44212 69134
rect 44156 68908 44212 68964
rect 45164 68908 45220 68964
rect 43484 67170 43540 67172
rect 43484 67118 43486 67170
rect 43486 67118 43538 67170
rect 43538 67118 43540 67170
rect 43484 67116 43540 67118
rect 42812 67004 42868 67060
rect 42700 66108 42756 66164
rect 42812 65996 42868 66052
rect 43036 66050 43092 66052
rect 43036 65998 43038 66050
rect 43038 65998 43090 66050
rect 43090 65998 43092 66050
rect 43036 65996 43092 65998
rect 44492 67170 44548 67172
rect 44492 67118 44494 67170
rect 44494 67118 44546 67170
rect 44546 67118 44548 67170
rect 44492 67116 44548 67118
rect 43260 66780 43316 66836
rect 43372 66498 43428 66500
rect 43372 66446 43374 66498
rect 43374 66446 43426 66498
rect 43426 66446 43428 66498
rect 43372 66444 43428 66446
rect 44044 66444 44100 66500
rect 44492 66332 44548 66388
rect 43596 66162 43652 66164
rect 43596 66110 43598 66162
rect 43598 66110 43650 66162
rect 43650 66110 43652 66162
rect 43596 66108 43652 66110
rect 43708 65996 43764 66052
rect 42588 65548 42644 65604
rect 43372 65548 43428 65604
rect 43036 65436 43092 65492
rect 42028 65100 42084 65156
rect 41692 64930 41748 64932
rect 41692 64878 41694 64930
rect 41694 64878 41746 64930
rect 41746 64878 41748 64930
rect 41692 64876 41748 64878
rect 42252 64594 42308 64596
rect 42252 64542 42254 64594
rect 42254 64542 42306 64594
rect 42306 64542 42308 64594
rect 42252 64540 42308 64542
rect 42140 64428 42196 64484
rect 42700 65324 42756 65380
rect 43260 65100 43316 65156
rect 43036 64594 43092 64596
rect 43036 64542 43038 64594
rect 43038 64542 43090 64594
rect 43090 64542 43092 64594
rect 43036 64540 43092 64542
rect 42252 64204 42308 64260
rect 42588 64204 42644 64260
rect 42476 64146 42532 64148
rect 42476 64094 42478 64146
rect 42478 64094 42530 64146
rect 42530 64094 42532 64146
rect 42476 64092 42532 64094
rect 41468 63756 41524 63812
rect 41692 63196 41748 63252
rect 41916 63698 41972 63700
rect 41916 63646 41918 63698
rect 41918 63646 41970 63698
rect 41970 63646 41972 63698
rect 41916 63644 41972 63646
rect 41020 62748 41076 62804
rect 41692 62636 41748 62692
rect 41132 62578 41188 62580
rect 41132 62526 41134 62578
rect 41134 62526 41186 62578
rect 41186 62526 41188 62578
rect 41132 62524 41188 62526
rect 40908 62354 40964 62356
rect 40908 62302 40910 62354
rect 40910 62302 40962 62354
rect 40962 62302 40964 62354
rect 40908 62300 40964 62302
rect 40796 62188 40852 62244
rect 41356 62466 41412 62468
rect 41356 62414 41358 62466
rect 41358 62414 41410 62466
rect 41410 62414 41412 62466
rect 41356 62412 41412 62414
rect 41244 62300 41300 62356
rect 40908 61964 40964 62020
rect 41356 61628 41412 61684
rect 42700 63308 42756 63364
rect 43148 62972 43204 63028
rect 42924 62860 42980 62916
rect 41916 61740 41972 61796
rect 42140 61794 42196 61796
rect 42140 61742 42142 61794
rect 42142 61742 42194 61794
rect 42194 61742 42196 61794
rect 42140 61740 42196 61742
rect 42812 62354 42868 62356
rect 42812 62302 42814 62354
rect 42814 62302 42866 62354
rect 42866 62302 42868 62354
rect 42812 62300 42868 62302
rect 43260 62578 43316 62580
rect 43260 62526 43262 62578
rect 43262 62526 43314 62578
rect 43314 62526 43316 62578
rect 43260 62524 43316 62526
rect 43372 62412 43428 62468
rect 42364 61740 42420 61796
rect 41692 61628 41748 61684
rect 42252 61628 42308 61684
rect 40908 61180 40964 61236
rect 41020 60508 41076 60564
rect 41020 60172 41076 60228
rect 41020 59778 41076 59780
rect 41020 59726 41022 59778
rect 41022 59726 41074 59778
rect 41074 59726 41076 59778
rect 41020 59724 41076 59726
rect 41804 61404 41860 61460
rect 41580 61180 41636 61236
rect 42252 61180 42308 61236
rect 42140 61068 42196 61124
rect 41580 59836 41636 59892
rect 41468 59778 41524 59780
rect 41468 59726 41470 59778
rect 41470 59726 41522 59778
rect 41522 59726 41524 59778
rect 41468 59724 41524 59726
rect 41244 58772 41300 58828
rect 41468 58546 41524 58548
rect 41468 58494 41470 58546
rect 41470 58494 41522 58546
rect 41522 58494 41524 58546
rect 41468 58492 41524 58494
rect 41244 58156 41300 58212
rect 41132 58044 41188 58100
rect 41356 57650 41412 57652
rect 41356 57598 41358 57650
rect 41358 57598 41410 57650
rect 41410 57598 41412 57650
rect 41356 57596 41412 57598
rect 41580 58044 41636 58100
rect 42028 58044 42084 58100
rect 41916 57874 41972 57876
rect 41916 57822 41918 57874
rect 41918 57822 41970 57874
rect 41970 57822 41972 57874
rect 41916 57820 41972 57822
rect 41020 56588 41076 56644
rect 43484 64204 43540 64260
rect 42700 61458 42756 61460
rect 42700 61406 42702 61458
rect 42702 61406 42754 61458
rect 42754 61406 42756 61458
rect 42700 61404 42756 61406
rect 42252 60396 42308 60452
rect 42588 59836 42644 59892
rect 42252 59724 42308 59780
rect 42364 59612 42420 59668
rect 42252 57596 42308 57652
rect 43148 61180 43204 61236
rect 42588 59442 42644 59444
rect 42588 59390 42590 59442
rect 42590 59390 42642 59442
rect 42642 59390 42644 59442
rect 42588 59388 42644 59390
rect 43596 63868 43652 63924
rect 43820 65714 43876 65716
rect 43820 65662 43822 65714
rect 43822 65662 43874 65714
rect 43874 65662 43876 65714
rect 43820 65660 43876 65662
rect 44268 66108 44324 66164
rect 43932 65436 43988 65492
rect 44044 64428 44100 64484
rect 43596 62860 43652 62916
rect 44044 62914 44100 62916
rect 44044 62862 44046 62914
rect 44046 62862 44098 62914
rect 44098 62862 44100 62914
rect 44044 62860 44100 62862
rect 44380 65714 44436 65716
rect 44380 65662 44382 65714
rect 44382 65662 44434 65714
rect 44434 65662 44436 65714
rect 44380 65660 44436 65662
rect 44604 65996 44660 66052
rect 45052 67116 45108 67172
rect 44940 67058 44996 67060
rect 44940 67006 44942 67058
rect 44942 67006 44994 67058
rect 44994 67006 44996 67058
rect 44940 67004 44996 67006
rect 44828 66332 44884 66388
rect 44716 64316 44772 64372
rect 44268 62914 44324 62916
rect 44268 62862 44270 62914
rect 44270 62862 44322 62914
rect 44322 62862 44324 62914
rect 44268 62860 44324 62862
rect 44604 62578 44660 62580
rect 44604 62526 44606 62578
rect 44606 62526 44658 62578
rect 44658 62526 44660 62578
rect 44604 62524 44660 62526
rect 44156 62466 44212 62468
rect 44156 62414 44158 62466
rect 44158 62414 44210 62466
rect 44210 62414 44212 62466
rect 44156 62412 44212 62414
rect 43596 61740 43652 61796
rect 44380 61346 44436 61348
rect 44380 61294 44382 61346
rect 44382 61294 44434 61346
rect 44434 61294 44436 61346
rect 44380 61292 44436 61294
rect 43596 60396 43652 60452
rect 43148 59612 43204 59668
rect 42924 59388 42980 59444
rect 42588 59052 42644 59108
rect 42588 58828 42644 58884
rect 42252 57036 42308 57092
rect 40796 53730 40852 53732
rect 40796 53678 40798 53730
rect 40798 53678 40850 53730
rect 40850 53678 40852 53730
rect 40796 53676 40852 53678
rect 42364 55356 42420 55412
rect 42476 55916 42532 55972
rect 41580 55298 41636 55300
rect 41580 55246 41582 55298
rect 41582 55246 41634 55298
rect 41634 55246 41636 55298
rect 41580 55244 41636 55246
rect 41020 55186 41076 55188
rect 41020 55134 41022 55186
rect 41022 55134 41074 55186
rect 41074 55134 41076 55186
rect 41020 55132 41076 55134
rect 42252 55186 42308 55188
rect 42252 55134 42254 55186
rect 42254 55134 42306 55186
rect 42306 55134 42308 55186
rect 42252 55132 42308 55134
rect 41804 55074 41860 55076
rect 41804 55022 41806 55074
rect 41806 55022 41858 55074
rect 41858 55022 41860 55074
rect 41804 55020 41860 55022
rect 41020 54514 41076 54516
rect 41020 54462 41022 54514
rect 41022 54462 41074 54514
rect 41074 54462 41076 54514
rect 41020 54460 41076 54462
rect 42140 54348 42196 54404
rect 42364 55074 42420 55076
rect 42364 55022 42366 55074
rect 42366 55022 42418 55074
rect 42418 55022 42420 55074
rect 42364 55020 42420 55022
rect 42700 56194 42756 56196
rect 42700 56142 42702 56194
rect 42702 56142 42754 56194
rect 42754 56142 42756 56194
rect 42700 56140 42756 56142
rect 42588 55244 42644 55300
rect 41244 53116 41300 53172
rect 41356 53452 41412 53508
rect 41020 53004 41076 53060
rect 40908 52108 40964 52164
rect 40236 50204 40292 50260
rect 41132 50428 41188 50484
rect 41356 51212 41412 51268
rect 41356 50706 41412 50708
rect 41356 50654 41358 50706
rect 41358 50654 41410 50706
rect 41410 50654 41412 50706
rect 41356 50652 41412 50654
rect 40012 49810 40068 49812
rect 40012 49758 40014 49810
rect 40014 49758 40066 49810
rect 40066 49758 40068 49810
rect 40012 49756 40068 49758
rect 39900 48972 39956 49028
rect 39788 48914 39844 48916
rect 39788 48862 39790 48914
rect 39790 48862 39842 48914
rect 39842 48862 39844 48914
rect 39788 48860 39844 48862
rect 39676 48636 39732 48692
rect 39564 47570 39620 47572
rect 39564 47518 39566 47570
rect 39566 47518 39618 47570
rect 39618 47518 39620 47570
rect 39564 47516 39620 47518
rect 39452 46956 39508 47012
rect 38892 43596 38948 43652
rect 39788 47346 39844 47348
rect 39788 47294 39790 47346
rect 39790 47294 39842 47346
rect 39842 47294 39844 47346
rect 39788 47292 39844 47294
rect 38780 42588 38836 42644
rect 37660 41692 37716 41748
rect 38108 41298 38164 41300
rect 38108 41246 38110 41298
rect 38110 41246 38162 41298
rect 38162 41246 38164 41298
rect 38108 41244 38164 41246
rect 39564 43650 39620 43652
rect 39564 43598 39566 43650
rect 39566 43598 39618 43650
rect 39618 43598 39620 43650
rect 39564 43596 39620 43598
rect 39116 42812 39172 42868
rect 39676 42754 39732 42756
rect 39676 42702 39678 42754
rect 39678 42702 39730 42754
rect 39730 42702 39732 42754
rect 39676 42700 39732 42702
rect 39228 42642 39284 42644
rect 39228 42590 39230 42642
rect 39230 42590 39282 42642
rect 39282 42590 39284 42642
rect 39228 42588 39284 42590
rect 38556 41244 38612 41300
rect 37884 40236 37940 40292
rect 38220 39004 38276 39060
rect 38332 38668 38388 38724
rect 38220 35868 38276 35924
rect 38444 36316 38500 36372
rect 38444 36092 38500 36148
rect 37212 35644 37268 35700
rect 37100 35138 37156 35140
rect 37100 35086 37102 35138
rect 37102 35086 37154 35138
rect 37154 35086 37156 35138
rect 37100 35084 37156 35086
rect 36988 34188 37044 34244
rect 37212 33964 37268 34020
rect 37436 33516 37492 33572
rect 36092 32172 36148 32228
rect 35644 31724 35700 31780
rect 36540 32396 36596 32452
rect 36428 31948 36484 32004
rect 36316 31724 36372 31780
rect 37548 33404 37604 33460
rect 37660 33346 37716 33348
rect 37660 33294 37662 33346
rect 37662 33294 37714 33346
rect 37714 33294 37716 33346
rect 37660 33292 37716 33294
rect 38780 40290 38836 40292
rect 38780 40238 38782 40290
rect 38782 40238 38834 40290
rect 38834 40238 38836 40290
rect 38780 40236 38836 40238
rect 39004 40402 39060 40404
rect 39004 40350 39006 40402
rect 39006 40350 39058 40402
rect 39058 40350 39060 40402
rect 39004 40348 39060 40350
rect 39676 41970 39732 41972
rect 39676 41918 39678 41970
rect 39678 41918 39730 41970
rect 39730 41918 39732 41970
rect 39676 41916 39732 41918
rect 39676 41244 39732 41300
rect 40236 49980 40292 50036
rect 40236 49138 40292 49140
rect 40236 49086 40238 49138
rect 40238 49086 40290 49138
rect 40290 49086 40292 49138
rect 40236 49084 40292 49086
rect 40012 48466 40068 48468
rect 40012 48414 40014 48466
rect 40014 48414 40066 48466
rect 40066 48414 40068 48466
rect 40012 48412 40068 48414
rect 40236 48242 40292 48244
rect 40236 48190 40238 48242
rect 40238 48190 40290 48242
rect 40290 48190 40292 48242
rect 40236 48188 40292 48190
rect 40460 48300 40516 48356
rect 40460 48076 40516 48132
rect 41132 48972 41188 49028
rect 41020 48748 41076 48804
rect 40796 48188 40852 48244
rect 40572 47570 40628 47572
rect 40572 47518 40574 47570
rect 40574 47518 40626 47570
rect 40626 47518 40628 47570
rect 40572 47516 40628 47518
rect 40908 48130 40964 48132
rect 40908 48078 40910 48130
rect 40910 48078 40962 48130
rect 40962 48078 40964 48130
rect 40908 48076 40964 48078
rect 41020 47404 41076 47460
rect 41132 47346 41188 47348
rect 41132 47294 41134 47346
rect 41134 47294 41186 47346
rect 41186 47294 41188 47346
rect 41132 47292 41188 47294
rect 41132 46956 41188 47012
rect 41468 48914 41524 48916
rect 41468 48862 41470 48914
rect 41470 48862 41522 48914
rect 41522 48862 41524 48914
rect 41468 48860 41524 48862
rect 41804 53116 41860 53172
rect 42252 53506 42308 53508
rect 42252 53454 42254 53506
rect 42254 53454 42306 53506
rect 42306 53454 42308 53506
rect 42252 53452 42308 53454
rect 42364 53116 42420 53172
rect 42476 53452 42532 53508
rect 42700 53618 42756 53620
rect 42700 53566 42702 53618
rect 42702 53566 42754 53618
rect 42754 53566 42756 53618
rect 42700 53564 42756 53566
rect 42588 53058 42644 53060
rect 42588 53006 42590 53058
rect 42590 53006 42642 53058
rect 42642 53006 42644 53058
rect 42588 53004 42644 53006
rect 43260 59164 43316 59220
rect 43148 59106 43204 59108
rect 43148 59054 43150 59106
rect 43150 59054 43202 59106
rect 43202 59054 43204 59106
rect 43148 59052 43204 59054
rect 43484 59724 43540 59780
rect 43596 59836 43652 59892
rect 43484 59052 43540 59108
rect 44940 65436 44996 65492
rect 50556 69018 50612 69020
rect 50556 68966 50558 69018
rect 50558 68966 50610 69018
rect 50610 68966 50612 69018
rect 50556 68964 50612 68966
rect 50660 69018 50716 69020
rect 50660 68966 50662 69018
rect 50662 68966 50714 69018
rect 50714 68966 50716 69018
rect 50660 68964 50716 68966
rect 50764 69018 50820 69020
rect 50764 68966 50766 69018
rect 50766 68966 50818 69018
rect 50818 68966 50820 69018
rect 50764 68964 50820 68966
rect 45836 67564 45892 67620
rect 45388 67058 45444 67060
rect 45388 67006 45390 67058
rect 45390 67006 45442 67058
rect 45442 67006 45444 67058
rect 45388 67004 45444 67006
rect 45612 66332 45668 66388
rect 45164 65996 45220 66052
rect 45276 64482 45332 64484
rect 45276 64430 45278 64482
rect 45278 64430 45330 64482
rect 45330 64430 45332 64482
rect 45276 64428 45332 64430
rect 45500 64092 45556 64148
rect 45276 63980 45332 64036
rect 45388 63026 45444 63028
rect 45388 62974 45390 63026
rect 45390 62974 45442 63026
rect 45442 62974 45444 63026
rect 45388 62972 45444 62974
rect 44940 61516 44996 61572
rect 45388 61346 45444 61348
rect 45388 61294 45390 61346
rect 45390 61294 45442 61346
rect 45442 61294 45444 61346
rect 45388 61292 45444 61294
rect 45052 60396 45108 60452
rect 43708 59164 43764 59220
rect 43484 58492 43540 58548
rect 43820 58716 43876 58772
rect 43932 58940 43988 58996
rect 43708 58268 43764 58324
rect 44268 59218 44324 59220
rect 44268 59166 44270 59218
rect 44270 59166 44322 59218
rect 44322 59166 44324 59218
rect 44268 59164 44324 59166
rect 44044 58604 44100 58660
rect 43484 57874 43540 57876
rect 43484 57822 43486 57874
rect 43486 57822 43538 57874
rect 43538 57822 43540 57874
rect 43484 57820 43540 57822
rect 43820 56252 43876 56308
rect 42924 56082 42980 56084
rect 42924 56030 42926 56082
rect 42926 56030 42978 56082
rect 42978 56030 42980 56082
rect 42924 56028 42980 56030
rect 43036 55074 43092 55076
rect 43036 55022 43038 55074
rect 43038 55022 43090 55074
rect 43090 55022 43092 55074
rect 43036 55020 43092 55022
rect 42924 54908 42980 54964
rect 46844 64092 46900 64148
rect 47180 64146 47236 64148
rect 47180 64094 47182 64146
rect 47182 64094 47234 64146
rect 47234 64094 47236 64146
rect 47180 64092 47236 64094
rect 47068 63980 47124 64036
rect 47292 63980 47348 64036
rect 45724 63308 45780 63364
rect 45500 59890 45556 59892
rect 45500 59838 45502 59890
rect 45502 59838 45554 59890
rect 45554 59838 45556 59890
rect 45500 59836 45556 59838
rect 45612 59612 45668 59668
rect 44492 58156 44548 58212
rect 44268 56476 44324 56532
rect 44044 56140 44100 56196
rect 43932 56082 43988 56084
rect 43932 56030 43934 56082
rect 43934 56030 43986 56082
rect 43986 56030 43988 56082
rect 43932 56028 43988 56030
rect 43372 55356 43428 55412
rect 43820 55468 43876 55524
rect 43932 55074 43988 55076
rect 43932 55022 43934 55074
rect 43934 55022 43986 55074
rect 43986 55022 43988 55074
rect 43932 55020 43988 55022
rect 43820 54402 43876 54404
rect 43820 54350 43822 54402
rect 43822 54350 43874 54402
rect 43874 54350 43876 54402
rect 43820 54348 43876 54350
rect 44156 54514 44212 54516
rect 44156 54462 44158 54514
rect 44158 54462 44210 54514
rect 44210 54462 44212 54514
rect 44156 54460 44212 54462
rect 43820 53618 43876 53620
rect 43820 53566 43822 53618
rect 43822 53566 43874 53618
rect 43874 53566 43876 53618
rect 43820 53564 43876 53566
rect 43372 53228 43428 53284
rect 43708 53228 43764 53284
rect 42812 52892 42868 52948
rect 42588 52108 42644 52164
rect 41804 51436 41860 51492
rect 41916 50876 41972 50932
rect 41580 48802 41636 48804
rect 41580 48750 41582 48802
rect 41582 48750 41634 48802
rect 41634 48750 41636 48802
rect 41580 48748 41636 48750
rect 41692 50652 41748 50708
rect 41468 48242 41524 48244
rect 41468 48190 41470 48242
rect 41470 48190 41522 48242
rect 41522 48190 41524 48242
rect 41468 48188 41524 48190
rect 42364 50706 42420 50708
rect 42364 50654 42366 50706
rect 42366 50654 42418 50706
rect 42418 50654 42420 50706
rect 42364 50652 42420 50654
rect 42140 49532 42196 49588
rect 42028 49026 42084 49028
rect 42028 48974 42030 49026
rect 42030 48974 42082 49026
rect 42082 48974 42084 49026
rect 42028 48972 42084 48974
rect 41356 46844 41412 46900
rect 41804 48524 41860 48580
rect 40908 45948 40964 46004
rect 40684 44156 40740 44212
rect 41356 44492 41412 44548
rect 40572 42754 40628 42756
rect 40572 42702 40574 42754
rect 40574 42702 40626 42754
rect 40626 42702 40628 42754
rect 40572 42700 40628 42702
rect 40908 43372 40964 43428
rect 40236 42588 40292 42644
rect 39788 40796 39844 40852
rect 39564 40402 39620 40404
rect 39564 40350 39566 40402
rect 39566 40350 39618 40402
rect 39618 40350 39620 40402
rect 39564 40348 39620 40350
rect 39452 38946 39508 38948
rect 39452 38894 39454 38946
rect 39454 38894 39506 38946
rect 39506 38894 39508 38946
rect 39452 38892 39508 38894
rect 39788 39004 39844 39060
rect 39676 38780 39732 38836
rect 38892 38722 38948 38724
rect 38892 38670 38894 38722
rect 38894 38670 38946 38722
rect 38946 38670 38948 38722
rect 38892 38668 38948 38670
rect 41020 42642 41076 42644
rect 41020 42590 41022 42642
rect 41022 42590 41074 42642
rect 41074 42590 41076 42642
rect 41020 42588 41076 42590
rect 40796 42476 40852 42532
rect 41020 41804 41076 41860
rect 41356 42754 41412 42756
rect 41356 42702 41358 42754
rect 41358 42702 41410 42754
rect 41410 42702 41412 42754
rect 41356 42700 41412 42702
rect 41580 47180 41636 47236
rect 41916 48188 41972 48244
rect 41916 47068 41972 47124
rect 42252 48914 42308 48916
rect 42252 48862 42254 48914
rect 42254 48862 42306 48914
rect 42306 48862 42308 48914
rect 42252 48860 42308 48862
rect 42364 48412 42420 48468
rect 42476 48300 42532 48356
rect 42700 50204 42756 50260
rect 43148 53116 43204 53172
rect 44268 52162 44324 52164
rect 44268 52110 44270 52162
rect 44270 52110 44322 52162
rect 44322 52110 44324 52162
rect 44268 52108 44324 52110
rect 44156 51996 44212 52052
rect 43820 51212 43876 51268
rect 43484 50594 43540 50596
rect 43484 50542 43486 50594
rect 43486 50542 43538 50594
rect 43538 50542 43540 50594
rect 43484 50540 43540 50542
rect 43148 49980 43204 50036
rect 43820 49980 43876 50036
rect 42924 49532 42980 49588
rect 43484 49810 43540 49812
rect 43484 49758 43486 49810
rect 43486 49758 43538 49810
rect 43538 49758 43540 49810
rect 43484 49756 43540 49758
rect 44268 49810 44324 49812
rect 44268 49758 44270 49810
rect 44270 49758 44322 49810
rect 44322 49758 44324 49810
rect 44268 49756 44324 49758
rect 42924 48802 42980 48804
rect 42924 48750 42926 48802
rect 42926 48750 42978 48802
rect 42978 48750 42980 48802
rect 42924 48748 42980 48750
rect 43148 48802 43204 48804
rect 43148 48750 43150 48802
rect 43150 48750 43202 48802
rect 43202 48750 43204 48802
rect 43148 48748 43204 48750
rect 43260 48354 43316 48356
rect 43260 48302 43262 48354
rect 43262 48302 43314 48354
rect 43314 48302 43316 48354
rect 43260 48300 43316 48302
rect 42924 47852 42980 47908
rect 42924 47346 42980 47348
rect 42924 47294 42926 47346
rect 42926 47294 42978 47346
rect 42978 47294 42980 47346
rect 42924 47292 42980 47294
rect 42364 46956 42420 47012
rect 43260 47234 43316 47236
rect 43260 47182 43262 47234
rect 43262 47182 43314 47234
rect 43314 47182 43316 47234
rect 43260 47180 43316 47182
rect 43260 46956 43316 47012
rect 42588 46732 42644 46788
rect 42924 46674 42980 46676
rect 42924 46622 42926 46674
rect 42926 46622 42978 46674
rect 42978 46622 42980 46674
rect 42924 46620 42980 46622
rect 42812 46508 42868 46564
rect 41804 45388 41860 45444
rect 41580 44210 41636 44212
rect 41580 44158 41582 44210
rect 41582 44158 41634 44210
rect 41634 44158 41636 44210
rect 41580 44156 41636 44158
rect 42140 44156 42196 44212
rect 42812 44380 42868 44436
rect 42924 45164 42980 45220
rect 43596 48914 43652 48916
rect 43596 48862 43598 48914
rect 43598 48862 43650 48914
rect 43650 48862 43652 48914
rect 43596 48860 43652 48862
rect 44716 58044 44772 58100
rect 44940 58828 44996 58884
rect 45500 59106 45556 59108
rect 45500 59054 45502 59106
rect 45502 59054 45554 59106
rect 45554 59054 45556 59106
rect 45500 59052 45556 59054
rect 45276 58994 45332 58996
rect 45276 58942 45278 58994
rect 45278 58942 45330 58994
rect 45330 58942 45332 58994
rect 45276 58940 45332 58942
rect 45724 59052 45780 59108
rect 45164 58716 45220 58772
rect 44940 58210 44996 58212
rect 44940 58158 44942 58210
rect 44942 58158 44994 58210
rect 44994 58158 44996 58210
rect 44940 58156 44996 58158
rect 50556 67450 50612 67452
rect 50556 67398 50558 67450
rect 50558 67398 50610 67450
rect 50610 67398 50612 67450
rect 50556 67396 50612 67398
rect 50660 67450 50716 67452
rect 50660 67398 50662 67450
rect 50662 67398 50714 67450
rect 50714 67398 50716 67450
rect 50660 67396 50716 67398
rect 50764 67450 50820 67452
rect 50764 67398 50766 67450
rect 50766 67398 50818 67450
rect 50818 67398 50820 67450
rect 50764 67396 50820 67398
rect 47404 62188 47460 62244
rect 47516 65436 47572 65492
rect 50556 65882 50612 65884
rect 50556 65830 50558 65882
rect 50558 65830 50610 65882
rect 50610 65830 50612 65882
rect 50556 65828 50612 65830
rect 50660 65882 50716 65884
rect 50660 65830 50662 65882
rect 50662 65830 50714 65882
rect 50714 65830 50716 65882
rect 50660 65828 50716 65830
rect 50764 65882 50820 65884
rect 50764 65830 50766 65882
rect 50766 65830 50818 65882
rect 50818 65830 50820 65882
rect 50764 65828 50820 65830
rect 47628 64034 47684 64036
rect 47628 63982 47630 64034
rect 47630 63982 47682 64034
rect 47682 63982 47684 64034
rect 47628 63980 47684 63982
rect 50556 64314 50612 64316
rect 50556 64262 50558 64314
rect 50558 64262 50610 64314
rect 50610 64262 50612 64314
rect 50556 64260 50612 64262
rect 50660 64314 50716 64316
rect 50660 64262 50662 64314
rect 50662 64262 50714 64314
rect 50714 64262 50716 64314
rect 50660 64260 50716 64262
rect 50764 64314 50820 64316
rect 50764 64262 50766 64314
rect 50766 64262 50818 64314
rect 50818 64262 50820 64314
rect 50764 64260 50820 64262
rect 48188 63980 48244 64036
rect 48076 63420 48132 63476
rect 47852 62972 47908 63028
rect 48972 64034 49028 64036
rect 48972 63982 48974 64034
rect 48974 63982 49026 64034
rect 49026 63982 49028 64034
rect 48972 63980 49028 63982
rect 48748 63868 48804 63924
rect 49420 63922 49476 63924
rect 49420 63870 49422 63922
rect 49422 63870 49474 63922
rect 49474 63870 49476 63922
rect 49420 63868 49476 63870
rect 48860 63420 48916 63476
rect 46396 61570 46452 61572
rect 46396 61518 46398 61570
rect 46398 61518 46450 61570
rect 46450 61518 46452 61570
rect 46396 61516 46452 61518
rect 46172 61458 46228 61460
rect 46172 61406 46174 61458
rect 46174 61406 46226 61458
rect 46226 61406 46228 61458
rect 46172 61404 46228 61406
rect 46172 60786 46228 60788
rect 46172 60734 46174 60786
rect 46174 60734 46226 60786
rect 46226 60734 46228 60786
rect 46172 60732 46228 60734
rect 45948 60284 46004 60340
rect 45276 58604 45332 58660
rect 45164 58210 45220 58212
rect 45164 58158 45166 58210
rect 45166 58158 45218 58210
rect 45218 58158 45220 58210
rect 45164 58156 45220 58158
rect 45276 58044 45332 58100
rect 45388 57932 45444 57988
rect 44828 57708 44884 57764
rect 45276 57708 45332 57764
rect 44940 57148 44996 57204
rect 44716 56082 44772 56084
rect 44716 56030 44718 56082
rect 44718 56030 44770 56082
rect 44770 56030 44772 56082
rect 44716 56028 44772 56030
rect 46396 60508 46452 60564
rect 46844 60508 46900 60564
rect 46732 60002 46788 60004
rect 46732 59950 46734 60002
rect 46734 59950 46786 60002
rect 46786 59950 46788 60002
rect 46732 59948 46788 59950
rect 46060 59612 46116 59668
rect 47516 61516 47572 61572
rect 47180 60732 47236 60788
rect 46956 59890 47012 59892
rect 46956 59838 46958 59890
rect 46958 59838 47010 59890
rect 47010 59838 47012 59890
rect 46956 59836 47012 59838
rect 45948 58604 46004 58660
rect 46060 59052 46116 59108
rect 45836 58210 45892 58212
rect 45836 58158 45838 58210
rect 45838 58158 45890 58210
rect 45890 58158 45892 58210
rect 45836 58156 45892 58158
rect 46172 58828 46228 58884
rect 46060 58044 46116 58100
rect 46956 59218 47012 59220
rect 46956 59166 46958 59218
rect 46958 59166 47010 59218
rect 47010 59166 47012 59218
rect 46956 59164 47012 59166
rect 46732 58322 46788 58324
rect 46732 58270 46734 58322
rect 46734 58270 46786 58322
rect 46786 58270 46788 58322
rect 46732 58268 46788 58270
rect 46172 57650 46228 57652
rect 46172 57598 46174 57650
rect 46174 57598 46226 57650
rect 46226 57598 46228 57650
rect 46172 57596 46228 57598
rect 45612 57484 45668 57540
rect 46060 57484 46116 57540
rect 46508 57372 46564 57428
rect 45500 56364 45556 56420
rect 45388 56306 45444 56308
rect 45388 56254 45390 56306
rect 45390 56254 45442 56306
rect 45442 56254 45444 56306
rect 45388 56252 45444 56254
rect 46396 56364 46452 56420
rect 45164 54460 45220 54516
rect 44828 53618 44884 53620
rect 44828 53566 44830 53618
rect 44830 53566 44882 53618
rect 44882 53566 44884 53618
rect 44828 53564 44884 53566
rect 45052 53228 45108 53284
rect 45052 52780 45108 52836
rect 46732 57036 46788 57092
rect 46732 56642 46788 56644
rect 46732 56590 46734 56642
rect 46734 56590 46786 56642
rect 46786 56590 46788 56642
rect 46732 56588 46788 56590
rect 45836 55468 45892 55524
rect 45388 53058 45444 53060
rect 45388 53006 45390 53058
rect 45390 53006 45442 53058
rect 45442 53006 45444 53058
rect 45388 53004 45444 53006
rect 45500 54460 45556 54516
rect 45948 53228 46004 53284
rect 46732 53788 46788 53844
rect 46620 53506 46676 53508
rect 46620 53454 46622 53506
rect 46622 53454 46674 53506
rect 46674 53454 46676 53506
rect 46620 53452 46676 53454
rect 46508 53116 46564 53172
rect 45500 51996 45556 52052
rect 45388 51490 45444 51492
rect 45388 51438 45390 51490
rect 45390 51438 45442 51490
rect 45442 51438 45444 51490
rect 45388 51436 45444 51438
rect 44716 50540 44772 50596
rect 43932 48748 43988 48804
rect 43820 48466 43876 48468
rect 43820 48414 43822 48466
rect 43822 48414 43874 48466
rect 43874 48414 43876 48466
rect 43820 48412 43876 48414
rect 44156 48802 44212 48804
rect 44156 48750 44158 48802
rect 44158 48750 44210 48802
rect 44210 48750 44212 48802
rect 44156 48748 44212 48750
rect 43932 48130 43988 48132
rect 43932 48078 43934 48130
rect 43934 48078 43986 48130
rect 43986 48078 43988 48130
rect 43932 48076 43988 48078
rect 43596 47964 43652 48020
rect 45276 48748 45332 48804
rect 45388 48524 45444 48580
rect 44828 48466 44884 48468
rect 44828 48414 44830 48466
rect 44830 48414 44882 48466
rect 44882 48414 44884 48466
rect 44828 48412 44884 48414
rect 44044 47516 44100 47572
rect 44380 47964 44436 48020
rect 43932 47234 43988 47236
rect 43932 47182 43934 47234
rect 43934 47182 43986 47234
rect 43986 47182 43988 47234
rect 43932 47180 43988 47182
rect 43484 46674 43540 46676
rect 43484 46622 43486 46674
rect 43486 46622 43538 46674
rect 43538 46622 43540 46674
rect 43484 46620 43540 46622
rect 43708 46956 43764 47012
rect 43708 46450 43764 46452
rect 43708 46398 43710 46450
rect 43710 46398 43762 46450
rect 43762 46398 43764 46450
rect 43708 46396 43764 46398
rect 43820 46844 43876 46900
rect 43484 45836 43540 45892
rect 44268 46956 44324 47012
rect 45164 47516 45220 47572
rect 46508 52892 46564 52948
rect 45724 51436 45780 51492
rect 46732 51490 46788 51492
rect 46732 51438 46734 51490
rect 46734 51438 46786 51490
rect 46786 51438 46788 51490
rect 46732 51436 46788 51438
rect 46396 51266 46452 51268
rect 46396 51214 46398 51266
rect 46398 51214 46450 51266
rect 46450 51214 46452 51266
rect 46396 51212 46452 51214
rect 46732 50706 46788 50708
rect 46732 50654 46734 50706
rect 46734 50654 46786 50706
rect 46786 50654 46788 50706
rect 46732 50652 46788 50654
rect 45948 49980 46004 50036
rect 46172 48188 46228 48244
rect 45724 47458 45780 47460
rect 45724 47406 45726 47458
rect 45726 47406 45778 47458
rect 45778 47406 45780 47458
rect 45724 47404 45780 47406
rect 44492 47292 44548 47348
rect 45052 46956 45108 47012
rect 44604 46844 44660 46900
rect 45948 47292 46004 47348
rect 43708 45164 43764 45220
rect 44156 45330 44212 45332
rect 44156 45278 44158 45330
rect 44158 45278 44210 45330
rect 44210 45278 44212 45330
rect 44156 45276 44212 45278
rect 44828 46396 44884 46452
rect 45052 45890 45108 45892
rect 45052 45838 45054 45890
rect 45054 45838 45106 45890
rect 45106 45838 45108 45890
rect 45052 45836 45108 45838
rect 44940 45276 44996 45332
rect 45276 45836 45332 45892
rect 45388 46284 45444 46340
rect 45948 47068 46004 47124
rect 46508 48914 46564 48916
rect 46508 48862 46510 48914
rect 46510 48862 46562 48914
rect 46562 48862 46564 48914
rect 46508 48860 46564 48862
rect 46620 48802 46676 48804
rect 46620 48750 46622 48802
rect 46622 48750 46674 48802
rect 46674 48750 46676 48802
rect 46620 48748 46676 48750
rect 46396 48524 46452 48580
rect 46396 48300 46452 48356
rect 46620 47458 46676 47460
rect 46620 47406 46622 47458
rect 46622 47406 46674 47458
rect 46674 47406 46676 47458
rect 46620 47404 46676 47406
rect 47404 61292 47460 61348
rect 47404 60674 47460 60676
rect 47404 60622 47406 60674
rect 47406 60622 47458 60674
rect 47458 60622 47460 60674
rect 47404 60620 47460 60622
rect 48076 60396 48132 60452
rect 47516 60002 47572 60004
rect 47516 59950 47518 60002
rect 47518 59950 47570 60002
rect 47570 59950 47572 60002
rect 47516 59948 47572 59950
rect 47404 59890 47460 59892
rect 47404 59838 47406 59890
rect 47406 59838 47458 59890
rect 47458 59838 47460 59890
rect 47404 59836 47460 59838
rect 47292 59218 47348 59220
rect 47292 59166 47294 59218
rect 47294 59166 47346 59218
rect 47346 59166 47348 59218
rect 47292 59164 47348 59166
rect 47292 58156 47348 58212
rect 47516 58268 47572 58324
rect 48972 62972 49028 63028
rect 48860 60674 48916 60676
rect 48860 60622 48862 60674
rect 48862 60622 48914 60674
rect 48914 60622 48916 60674
rect 48860 60620 48916 60622
rect 50556 62746 50612 62748
rect 50556 62694 50558 62746
rect 50558 62694 50610 62746
rect 50610 62694 50612 62746
rect 50556 62692 50612 62694
rect 50660 62746 50716 62748
rect 50660 62694 50662 62746
rect 50662 62694 50714 62746
rect 50714 62694 50716 62746
rect 50660 62692 50716 62694
rect 50764 62746 50820 62748
rect 50764 62694 50766 62746
rect 50766 62694 50818 62746
rect 50818 62694 50820 62746
rect 50764 62692 50820 62694
rect 50764 62242 50820 62244
rect 50764 62190 50766 62242
rect 50766 62190 50818 62242
rect 50818 62190 50820 62242
rect 50764 62188 50820 62190
rect 49084 61516 49140 61572
rect 49196 61292 49252 61348
rect 49196 60620 49252 60676
rect 49084 60396 49140 60452
rect 50204 61516 50260 61572
rect 50876 61570 50932 61572
rect 50876 61518 50878 61570
rect 50878 61518 50930 61570
rect 50930 61518 50932 61570
rect 50876 61516 50932 61518
rect 50316 61292 50372 61348
rect 47964 59276 48020 59332
rect 48748 59276 48804 59332
rect 47852 59164 47908 59220
rect 47628 58156 47684 58212
rect 47740 58268 47796 58324
rect 47404 58044 47460 58100
rect 47292 57820 47348 57876
rect 47180 57260 47236 57316
rect 47516 57148 47572 57204
rect 48076 57260 48132 57316
rect 48188 57484 48244 57540
rect 47292 56306 47348 56308
rect 47292 56254 47294 56306
rect 47294 56254 47346 56306
rect 47346 56254 47348 56306
rect 47292 56252 47348 56254
rect 46956 56028 47012 56084
rect 46956 53170 47012 53172
rect 46956 53118 46958 53170
rect 46958 53118 47010 53170
rect 47010 53118 47012 53170
rect 46956 53116 47012 53118
rect 46956 52220 47012 52276
rect 47180 53228 47236 53284
rect 47852 56194 47908 56196
rect 47852 56142 47854 56194
rect 47854 56142 47906 56194
rect 47906 56142 47908 56194
rect 47852 56140 47908 56142
rect 47628 56082 47684 56084
rect 47628 56030 47630 56082
rect 47630 56030 47682 56082
rect 47682 56030 47684 56082
rect 47628 56028 47684 56030
rect 48076 56028 48132 56084
rect 48972 59218 49028 59220
rect 48972 59166 48974 59218
rect 48974 59166 49026 59218
rect 49026 59166 49028 59218
rect 48972 59164 49028 59166
rect 48860 57538 48916 57540
rect 48860 57486 48862 57538
rect 48862 57486 48914 57538
rect 48914 57486 48916 57538
rect 48860 57484 48916 57486
rect 49308 57538 49364 57540
rect 49308 57486 49310 57538
rect 49310 57486 49362 57538
rect 49362 57486 49364 57538
rect 49308 57484 49364 57486
rect 49420 57036 49476 57092
rect 47628 53900 47684 53956
rect 48636 56252 48692 56308
rect 48972 56194 49028 56196
rect 48972 56142 48974 56194
rect 48974 56142 49026 56194
rect 49026 56142 49028 56194
rect 48972 56140 49028 56142
rect 48860 56082 48916 56084
rect 48860 56030 48862 56082
rect 48862 56030 48914 56082
rect 48914 56030 48916 56082
rect 48860 56028 48916 56030
rect 47964 54738 48020 54740
rect 47964 54686 47966 54738
rect 47966 54686 48018 54738
rect 48018 54686 48020 54738
rect 47964 54684 48020 54686
rect 47852 53842 47908 53844
rect 47852 53790 47854 53842
rect 47854 53790 47906 53842
rect 47906 53790 47908 53842
rect 47852 53788 47908 53790
rect 48524 54460 48580 54516
rect 47516 53452 47572 53508
rect 47180 52946 47236 52948
rect 47180 52894 47182 52946
rect 47182 52894 47234 52946
rect 47234 52894 47236 52946
rect 47180 52892 47236 52894
rect 47292 52834 47348 52836
rect 47292 52782 47294 52834
rect 47294 52782 47346 52834
rect 47346 52782 47348 52834
rect 47292 52780 47348 52782
rect 47068 51548 47124 51604
rect 47068 51324 47124 51380
rect 47404 51378 47460 51380
rect 47404 51326 47406 51378
rect 47406 51326 47458 51378
rect 47458 51326 47460 51378
rect 47404 51324 47460 51326
rect 48524 53900 48580 53956
rect 48636 53842 48692 53844
rect 48636 53790 48638 53842
rect 48638 53790 48690 53842
rect 48690 53790 48692 53842
rect 48636 53788 48692 53790
rect 48748 54402 48804 54404
rect 48748 54350 48750 54402
rect 48750 54350 48802 54402
rect 48802 54350 48804 54402
rect 48748 54348 48804 54350
rect 48076 53058 48132 53060
rect 48076 53006 48078 53058
rect 48078 53006 48130 53058
rect 48130 53006 48132 53058
rect 48076 53004 48132 53006
rect 48076 51154 48132 51156
rect 48076 51102 48078 51154
rect 48078 51102 48130 51154
rect 48130 51102 48132 51154
rect 48076 51100 48132 51102
rect 47180 50316 47236 50372
rect 47180 47404 47236 47460
rect 46396 47068 46452 47124
rect 46284 46844 46340 46900
rect 46060 46674 46116 46676
rect 46060 46622 46062 46674
rect 46062 46622 46114 46674
rect 46114 46622 46116 46674
rect 46060 46620 46116 46622
rect 46956 47180 47012 47236
rect 46396 45836 46452 45892
rect 45164 45276 45220 45332
rect 44044 45164 44100 45220
rect 44828 45106 44884 45108
rect 44828 45054 44830 45106
rect 44830 45054 44882 45106
rect 44882 45054 44884 45106
rect 44828 45052 44884 45054
rect 45948 45276 46004 45332
rect 43372 44940 43428 44996
rect 43820 44994 43876 44996
rect 43820 44942 43822 44994
rect 43822 44942 43874 44994
rect 43874 44942 43876 44994
rect 43820 44940 43876 44942
rect 41580 43148 41636 43204
rect 41916 42642 41972 42644
rect 41916 42590 41918 42642
rect 41918 42590 41970 42642
rect 41970 42590 41972 42642
rect 41916 42588 41972 42590
rect 40908 40348 40964 40404
rect 40908 39340 40964 39396
rect 40684 39228 40740 39284
rect 40012 38892 40068 38948
rect 40908 39004 40964 39060
rect 41132 41356 41188 41412
rect 41468 41970 41524 41972
rect 41468 41918 41470 41970
rect 41470 41918 41522 41970
rect 41522 41918 41524 41970
rect 41468 41916 41524 41918
rect 41580 41804 41636 41860
rect 41580 40348 41636 40404
rect 41468 39676 41524 39732
rect 42924 43484 42980 43540
rect 42588 43148 42644 43204
rect 42700 43036 42756 43092
rect 42252 42476 42308 42532
rect 42028 40402 42084 40404
rect 42028 40350 42030 40402
rect 42030 40350 42082 40402
rect 42082 40350 42084 40402
rect 42028 40348 42084 40350
rect 41356 39394 41412 39396
rect 41356 39342 41358 39394
rect 41358 39342 41410 39394
rect 41410 39342 41412 39394
rect 41356 39340 41412 39342
rect 38780 36316 38836 36372
rect 38780 34972 38836 35028
rect 38220 34690 38276 34692
rect 38220 34638 38222 34690
rect 38222 34638 38274 34690
rect 38274 34638 38276 34690
rect 38220 34636 38276 34638
rect 38780 34636 38836 34692
rect 41132 38780 41188 38836
rect 40348 36876 40404 36932
rect 41132 36876 41188 36932
rect 39340 34690 39396 34692
rect 39340 34638 39342 34690
rect 39342 34638 39394 34690
rect 39394 34638 39396 34690
rect 39340 34636 39396 34638
rect 41020 35980 41076 36036
rect 39788 35922 39844 35924
rect 39788 35870 39790 35922
rect 39790 35870 39842 35922
rect 39842 35870 39844 35922
rect 39788 35868 39844 35870
rect 40124 35868 40180 35924
rect 39676 34802 39732 34804
rect 39676 34750 39678 34802
rect 39678 34750 39730 34802
rect 39730 34750 39732 34802
rect 39676 34748 39732 34750
rect 39900 35698 39956 35700
rect 39900 35646 39902 35698
rect 39902 35646 39954 35698
rect 39954 35646 39956 35698
rect 39900 35644 39956 35646
rect 41468 37772 41524 37828
rect 41468 37490 41524 37492
rect 41468 37438 41470 37490
rect 41470 37438 41522 37490
rect 41522 37438 41524 37490
rect 41468 37436 41524 37438
rect 41356 37212 41412 37268
rect 40908 35698 40964 35700
rect 40908 35646 40910 35698
rect 40910 35646 40962 35698
rect 40962 35646 40964 35698
rect 40908 35644 40964 35646
rect 42028 38668 42084 38724
rect 41916 37266 41972 37268
rect 41916 37214 41918 37266
rect 41918 37214 41970 37266
rect 41970 37214 41972 37266
rect 41916 37212 41972 37214
rect 41692 36988 41748 37044
rect 42924 41916 42980 41972
rect 43036 41356 43092 41412
rect 45612 45106 45668 45108
rect 45612 45054 45614 45106
rect 45614 45054 45666 45106
rect 45666 45054 45668 45106
rect 45612 45052 45668 45054
rect 44940 44322 44996 44324
rect 44940 44270 44942 44322
rect 44942 44270 44994 44322
rect 44994 44270 44996 44322
rect 44940 44268 44996 44270
rect 45612 43148 45668 43204
rect 45052 42924 45108 42980
rect 44828 42642 44884 42644
rect 44828 42590 44830 42642
rect 44830 42590 44882 42642
rect 44882 42590 44884 42642
rect 44828 42588 44884 42590
rect 43372 41132 43428 41188
rect 43036 40348 43092 40404
rect 43484 40012 43540 40068
rect 43372 39730 43428 39732
rect 43372 39678 43374 39730
rect 43374 39678 43426 39730
rect 43426 39678 43428 39730
rect 43372 39676 43428 39678
rect 43036 39618 43092 39620
rect 43036 39566 43038 39618
rect 43038 39566 43090 39618
rect 43090 39566 43092 39618
rect 43036 39564 43092 39566
rect 45388 42588 45444 42644
rect 45164 42530 45220 42532
rect 45164 42478 45166 42530
rect 45166 42478 45218 42530
rect 45218 42478 45220 42530
rect 45164 42476 45220 42478
rect 46060 43708 46116 43764
rect 46732 46844 46788 46900
rect 47068 46786 47124 46788
rect 47068 46734 47070 46786
rect 47070 46734 47122 46786
rect 47122 46734 47124 46786
rect 47068 46732 47124 46734
rect 46844 44268 46900 44324
rect 46844 43708 46900 43764
rect 47516 50652 47572 50708
rect 49308 54348 49364 54404
rect 49532 54684 49588 54740
rect 49084 53228 49140 53284
rect 49420 53842 49476 53844
rect 49420 53790 49422 53842
rect 49422 53790 49474 53842
rect 49474 53790 49476 53842
rect 49420 53788 49476 53790
rect 49756 59276 49812 59332
rect 49868 59442 49924 59444
rect 49868 59390 49870 59442
rect 49870 59390 49922 59442
rect 49922 59390 49924 59442
rect 49868 59388 49924 59390
rect 49868 59164 49924 59220
rect 49756 57260 49812 57316
rect 50556 61178 50612 61180
rect 50556 61126 50558 61178
rect 50558 61126 50610 61178
rect 50610 61126 50612 61178
rect 50556 61124 50612 61126
rect 50660 61178 50716 61180
rect 50660 61126 50662 61178
rect 50662 61126 50714 61178
rect 50714 61126 50716 61178
rect 50660 61124 50716 61126
rect 50764 61178 50820 61180
rect 50764 61126 50766 61178
rect 50766 61126 50818 61178
rect 50818 61126 50820 61178
rect 50764 61124 50820 61126
rect 52108 59724 52164 59780
rect 50556 59610 50612 59612
rect 50556 59558 50558 59610
rect 50558 59558 50610 59610
rect 50610 59558 50612 59610
rect 50556 59556 50612 59558
rect 50660 59610 50716 59612
rect 50660 59558 50662 59610
rect 50662 59558 50714 59610
rect 50714 59558 50716 59610
rect 50660 59556 50716 59558
rect 50764 59610 50820 59612
rect 50764 59558 50766 59610
rect 50766 59558 50818 59610
rect 50818 59558 50820 59610
rect 50764 59556 50820 59558
rect 50316 59388 50372 59444
rect 50092 57484 50148 57540
rect 49980 56252 50036 56308
rect 49980 55074 50036 55076
rect 49980 55022 49982 55074
rect 49982 55022 50034 55074
rect 50034 55022 50036 55074
rect 49980 55020 50036 55022
rect 49868 54460 49924 54516
rect 49756 53954 49812 53956
rect 49756 53902 49758 53954
rect 49758 53902 49810 53954
rect 49810 53902 49812 53954
rect 49756 53900 49812 53902
rect 50556 58042 50612 58044
rect 50556 57990 50558 58042
rect 50558 57990 50610 58042
rect 50610 57990 50612 58042
rect 50556 57988 50612 57990
rect 50660 58042 50716 58044
rect 50660 57990 50662 58042
rect 50662 57990 50714 58042
rect 50714 57990 50716 58042
rect 50660 57988 50716 57990
rect 50764 58042 50820 58044
rect 50764 57990 50766 58042
rect 50766 57990 50818 58042
rect 50818 57990 50820 58042
rect 50764 57988 50820 57990
rect 50556 56474 50612 56476
rect 50556 56422 50558 56474
rect 50558 56422 50610 56474
rect 50610 56422 50612 56474
rect 50556 56420 50612 56422
rect 50660 56474 50716 56476
rect 50660 56422 50662 56474
rect 50662 56422 50714 56474
rect 50714 56422 50716 56474
rect 50660 56420 50716 56422
rect 50764 56474 50820 56476
rect 50764 56422 50766 56474
rect 50766 56422 50818 56474
rect 50818 56422 50820 56474
rect 50764 56420 50820 56422
rect 49644 53564 49700 53620
rect 49084 52668 49140 52724
rect 48636 52220 48692 52276
rect 48860 51602 48916 51604
rect 48860 51550 48862 51602
rect 48862 51550 48914 51602
rect 48914 51550 48916 51602
rect 48860 51548 48916 51550
rect 48972 51436 49028 51492
rect 47852 48914 47908 48916
rect 47852 48862 47854 48914
rect 47854 48862 47906 48914
rect 47906 48862 47908 48914
rect 47852 48860 47908 48862
rect 47740 47404 47796 47460
rect 47628 46786 47684 46788
rect 47628 46734 47630 46786
rect 47630 46734 47682 46786
rect 47682 46734 47684 46786
rect 47628 46732 47684 46734
rect 47404 46674 47460 46676
rect 47404 46622 47406 46674
rect 47406 46622 47458 46674
rect 47458 46622 47460 46674
rect 47404 46620 47460 46622
rect 47516 46562 47572 46564
rect 47516 46510 47518 46562
rect 47518 46510 47570 46562
rect 47570 46510 47572 46562
rect 47516 46508 47572 46510
rect 47628 46284 47684 46340
rect 47964 45836 48020 45892
rect 47516 44156 47572 44212
rect 48748 48748 48804 48804
rect 48188 48130 48244 48132
rect 48188 48078 48190 48130
rect 48190 48078 48242 48130
rect 48242 48078 48244 48130
rect 48188 48076 48244 48078
rect 48300 47570 48356 47572
rect 48300 47518 48302 47570
rect 48302 47518 48354 47570
rect 48354 47518 48356 47570
rect 48300 47516 48356 47518
rect 48748 47570 48804 47572
rect 48748 47518 48750 47570
rect 48750 47518 48802 47570
rect 48802 47518 48804 47570
rect 48748 47516 48804 47518
rect 48300 46508 48356 46564
rect 48412 44322 48468 44324
rect 48412 44270 48414 44322
rect 48414 44270 48466 44322
rect 48466 44270 48468 44322
rect 48412 44268 48468 44270
rect 49308 51548 49364 51604
rect 49420 52162 49476 52164
rect 49420 52110 49422 52162
rect 49422 52110 49474 52162
rect 49474 52110 49476 52162
rect 49420 52108 49476 52110
rect 49196 51100 49252 51156
rect 49308 50316 49364 50372
rect 50876 55020 50932 55076
rect 50556 54906 50612 54908
rect 50556 54854 50558 54906
rect 50558 54854 50610 54906
rect 50610 54854 50612 54906
rect 50556 54852 50612 54854
rect 50660 54906 50716 54908
rect 50660 54854 50662 54906
rect 50662 54854 50714 54906
rect 50714 54854 50716 54906
rect 50660 54852 50716 54854
rect 50764 54906 50820 54908
rect 50764 54854 50766 54906
rect 50766 54854 50818 54906
rect 50818 54854 50820 54906
rect 50764 54852 50820 54854
rect 49756 51602 49812 51604
rect 49756 51550 49758 51602
rect 49758 51550 49810 51602
rect 49810 51550 49812 51602
rect 49756 51548 49812 51550
rect 49756 47516 49812 47572
rect 49644 44322 49700 44324
rect 49644 44270 49646 44322
rect 49646 44270 49698 44322
rect 49698 44270 49700 44322
rect 49644 44268 49700 44270
rect 48860 44210 48916 44212
rect 48860 44158 48862 44210
rect 48862 44158 48914 44210
rect 48914 44158 48916 44210
rect 48860 44156 48916 44158
rect 46284 43148 46340 43204
rect 45164 41186 45220 41188
rect 45164 41134 45166 41186
rect 45166 41134 45218 41186
rect 45218 41134 45220 41186
rect 45164 41132 45220 41134
rect 45052 40684 45108 40740
rect 45276 40572 45332 40628
rect 44940 40402 44996 40404
rect 44940 40350 44942 40402
rect 44942 40350 44994 40402
rect 44994 40350 44996 40402
rect 44940 40348 44996 40350
rect 44156 40012 44212 40068
rect 43932 39564 43988 39620
rect 45164 39452 45220 39508
rect 43260 38668 43316 38724
rect 45388 39228 45444 39284
rect 45276 39004 45332 39060
rect 46172 42476 46228 42532
rect 46956 42754 47012 42756
rect 46956 42702 46958 42754
rect 46958 42702 47010 42754
rect 47010 42702 47012 42754
rect 46956 42700 47012 42702
rect 47292 43148 47348 43204
rect 46172 40124 46228 40180
rect 46508 41916 46564 41972
rect 47068 42252 47124 42308
rect 47628 42812 47684 42868
rect 47180 42140 47236 42196
rect 47628 42364 47684 42420
rect 46732 41356 46788 41412
rect 46956 40124 47012 40180
rect 45612 39004 45668 39060
rect 46396 39394 46452 39396
rect 46396 39342 46398 39394
rect 46398 39342 46450 39394
rect 46450 39342 46452 39394
rect 46396 39340 46452 39342
rect 46620 39004 46676 39060
rect 45164 37996 45220 38052
rect 42588 37826 42644 37828
rect 42588 37774 42590 37826
rect 42590 37774 42642 37826
rect 42642 37774 42644 37826
rect 42588 37772 42644 37774
rect 42364 36876 42420 36932
rect 40460 34860 40516 34916
rect 40124 34748 40180 34804
rect 40124 34412 40180 34468
rect 39340 34242 39396 34244
rect 39340 34190 39342 34242
rect 39342 34190 39394 34242
rect 39394 34190 39396 34242
rect 39340 34188 39396 34190
rect 38332 34018 38388 34020
rect 38332 33966 38334 34018
rect 38334 33966 38386 34018
rect 38386 33966 38388 34018
rect 38332 33964 38388 33966
rect 38108 32620 38164 32676
rect 38444 33068 38500 33124
rect 37100 32284 37156 32340
rect 37324 32396 37380 32452
rect 36988 32172 37044 32228
rect 38220 31836 38276 31892
rect 37548 31778 37604 31780
rect 37548 31726 37550 31778
rect 37550 31726 37602 31778
rect 37602 31726 37604 31778
rect 37548 31724 37604 31726
rect 35532 31554 35588 31556
rect 35532 31502 35534 31554
rect 35534 31502 35586 31554
rect 35586 31502 35588 31554
rect 35532 31500 35588 31502
rect 35420 31052 35476 31108
rect 36316 31554 36372 31556
rect 36316 31502 36318 31554
rect 36318 31502 36370 31554
rect 36370 31502 36372 31554
rect 36316 31500 36372 31502
rect 35756 30716 35812 30772
rect 36428 31106 36484 31108
rect 36428 31054 36430 31106
rect 36430 31054 36482 31106
rect 36482 31054 36484 31106
rect 36428 31052 36484 31054
rect 35196 30602 35252 30604
rect 35196 30550 35198 30602
rect 35198 30550 35250 30602
rect 35250 30550 35252 30602
rect 35196 30548 35252 30550
rect 35300 30602 35356 30604
rect 35300 30550 35302 30602
rect 35302 30550 35354 30602
rect 35354 30550 35356 30602
rect 35300 30548 35356 30550
rect 35404 30602 35460 30604
rect 35404 30550 35406 30602
rect 35406 30550 35458 30602
rect 35458 30550 35460 30602
rect 35404 30548 35460 30550
rect 35756 30492 35812 30548
rect 34972 29426 35028 29428
rect 34972 29374 34974 29426
rect 34974 29374 35026 29426
rect 35026 29374 35028 29426
rect 34972 29372 35028 29374
rect 34972 28642 35028 28644
rect 34972 28590 34974 28642
rect 34974 28590 35026 28642
rect 35026 28590 35028 28642
rect 34972 28588 35028 28590
rect 34748 27356 34804 27412
rect 34972 28140 35028 28196
rect 34860 27074 34916 27076
rect 34860 27022 34862 27074
rect 34862 27022 34914 27074
rect 34914 27022 34916 27074
rect 34860 27020 34916 27022
rect 34300 26290 34356 26292
rect 34300 26238 34302 26290
rect 34302 26238 34354 26290
rect 34354 26238 34356 26290
rect 34300 26236 34356 26238
rect 34748 26962 34804 26964
rect 34748 26910 34750 26962
rect 34750 26910 34802 26962
rect 34802 26910 34804 26962
rect 34748 26908 34804 26910
rect 34748 26124 34804 26180
rect 34972 26124 35028 26180
rect 33740 23772 33796 23828
rect 33852 25228 33908 25284
rect 33964 25004 34020 25060
rect 34076 24892 34132 24948
rect 33964 24834 34020 24836
rect 33964 24782 33966 24834
rect 33966 24782 34018 24834
rect 34018 24782 34020 24834
rect 33964 24780 34020 24782
rect 33628 20300 33684 20356
rect 34748 25004 34804 25060
rect 34860 24780 34916 24836
rect 34636 24610 34692 24612
rect 34636 24558 34638 24610
rect 34638 24558 34690 24610
rect 34690 24558 34692 24610
rect 34636 24556 34692 24558
rect 34636 24108 34692 24164
rect 34524 23660 34580 23716
rect 34412 21868 34468 21924
rect 34300 20690 34356 20692
rect 34300 20638 34302 20690
rect 34302 20638 34354 20690
rect 34354 20638 34356 20690
rect 34300 20636 34356 20638
rect 34076 20076 34132 20132
rect 34300 20188 34356 20244
rect 33516 19852 33572 19908
rect 33404 18172 33460 18228
rect 34412 18844 34468 18900
rect 34524 18732 34580 18788
rect 33740 18450 33796 18452
rect 33740 18398 33742 18450
rect 33742 18398 33794 18450
rect 33794 18398 33796 18450
rect 33740 18396 33796 18398
rect 33852 18060 33908 18116
rect 33964 18396 34020 18452
rect 33628 17778 33684 17780
rect 33628 17726 33630 17778
rect 33630 17726 33682 17778
rect 33682 17726 33684 17778
rect 33628 17724 33684 17726
rect 33516 17164 33572 17220
rect 34188 18284 34244 18340
rect 34076 17612 34132 17668
rect 34412 18060 34468 18116
rect 34524 18172 34580 18228
rect 34524 17500 34580 17556
rect 34188 17106 34244 17108
rect 34188 17054 34190 17106
rect 34190 17054 34242 17106
rect 34242 17054 34244 17106
rect 34188 17052 34244 17054
rect 34188 16716 34244 16772
rect 36204 30716 36260 30772
rect 35644 29372 35700 29428
rect 35196 29034 35252 29036
rect 35196 28982 35198 29034
rect 35198 28982 35250 29034
rect 35250 28982 35252 29034
rect 35196 28980 35252 28982
rect 35300 29034 35356 29036
rect 35300 28982 35302 29034
rect 35302 28982 35354 29034
rect 35354 28982 35356 29034
rect 35300 28980 35356 28982
rect 35404 29034 35460 29036
rect 35404 28982 35406 29034
rect 35406 28982 35458 29034
rect 35458 28982 35460 29034
rect 35404 28980 35460 28982
rect 36092 29426 36148 29428
rect 36092 29374 36094 29426
rect 36094 29374 36146 29426
rect 36146 29374 36148 29426
rect 36092 29372 36148 29374
rect 36316 28812 36372 28868
rect 35532 28642 35588 28644
rect 35532 28590 35534 28642
rect 35534 28590 35586 28642
rect 35586 28590 35588 28642
rect 35532 28588 35588 28590
rect 35868 28642 35924 28644
rect 35868 28590 35870 28642
rect 35870 28590 35922 28642
rect 35922 28590 35924 28642
rect 35868 28588 35924 28590
rect 35196 28140 35252 28196
rect 36428 28700 36484 28756
rect 35196 27466 35252 27468
rect 35196 27414 35198 27466
rect 35198 27414 35250 27466
rect 35250 27414 35252 27466
rect 35196 27412 35252 27414
rect 35300 27466 35356 27468
rect 35300 27414 35302 27466
rect 35302 27414 35354 27466
rect 35354 27414 35356 27466
rect 35300 27412 35356 27414
rect 35404 27466 35460 27468
rect 35404 27414 35406 27466
rect 35406 27414 35458 27466
rect 35458 27414 35460 27466
rect 35404 27412 35460 27414
rect 35196 27298 35252 27300
rect 35196 27246 35198 27298
rect 35198 27246 35250 27298
rect 35250 27246 35252 27298
rect 35196 27244 35252 27246
rect 35756 27074 35812 27076
rect 35756 27022 35758 27074
rect 35758 27022 35810 27074
rect 35810 27022 35812 27074
rect 35756 27020 35812 27022
rect 35308 26962 35364 26964
rect 35308 26910 35310 26962
rect 35310 26910 35362 26962
rect 35362 26910 35364 26962
rect 35308 26908 35364 26910
rect 35532 26962 35588 26964
rect 35532 26910 35534 26962
rect 35534 26910 35586 26962
rect 35586 26910 35588 26962
rect 35532 26908 35588 26910
rect 36316 26962 36372 26964
rect 36316 26910 36318 26962
rect 36318 26910 36370 26962
rect 36370 26910 36372 26962
rect 36316 26908 36372 26910
rect 35196 26348 35252 26404
rect 36092 26290 36148 26292
rect 36092 26238 36094 26290
rect 36094 26238 36146 26290
rect 36146 26238 36148 26290
rect 36092 26236 36148 26238
rect 35868 26124 35924 26180
rect 35196 25898 35252 25900
rect 35196 25846 35198 25898
rect 35198 25846 35250 25898
rect 35250 25846 35252 25898
rect 35196 25844 35252 25846
rect 35300 25898 35356 25900
rect 35300 25846 35302 25898
rect 35302 25846 35354 25898
rect 35354 25846 35356 25898
rect 35300 25844 35356 25846
rect 35404 25898 35460 25900
rect 35404 25846 35406 25898
rect 35406 25846 35458 25898
rect 35458 25846 35460 25898
rect 35404 25844 35460 25846
rect 36204 25452 36260 25508
rect 35868 25282 35924 25284
rect 35868 25230 35870 25282
rect 35870 25230 35922 25282
rect 35922 25230 35924 25282
rect 35868 25228 35924 25230
rect 35196 25004 35252 25060
rect 35196 24330 35252 24332
rect 35196 24278 35198 24330
rect 35198 24278 35250 24330
rect 35250 24278 35252 24330
rect 35196 24276 35252 24278
rect 35300 24330 35356 24332
rect 35300 24278 35302 24330
rect 35302 24278 35354 24330
rect 35354 24278 35356 24330
rect 35300 24276 35356 24278
rect 35404 24330 35460 24332
rect 35404 24278 35406 24330
rect 35406 24278 35458 24330
rect 35458 24278 35460 24330
rect 35404 24276 35460 24278
rect 35084 24108 35140 24164
rect 35196 23714 35252 23716
rect 35196 23662 35198 23714
rect 35198 23662 35250 23714
rect 35250 23662 35252 23714
rect 35196 23660 35252 23662
rect 35756 23548 35812 23604
rect 35644 23266 35700 23268
rect 35644 23214 35646 23266
rect 35646 23214 35698 23266
rect 35698 23214 35700 23266
rect 35644 23212 35700 23214
rect 35196 22762 35252 22764
rect 35196 22710 35198 22762
rect 35198 22710 35250 22762
rect 35250 22710 35252 22762
rect 35196 22708 35252 22710
rect 35300 22762 35356 22764
rect 35300 22710 35302 22762
rect 35302 22710 35354 22762
rect 35354 22710 35356 22762
rect 35300 22708 35356 22710
rect 35404 22762 35460 22764
rect 35404 22710 35406 22762
rect 35406 22710 35458 22762
rect 35458 22710 35460 22762
rect 35404 22708 35460 22710
rect 34972 21756 35028 21812
rect 35196 21586 35252 21588
rect 35196 21534 35198 21586
rect 35198 21534 35250 21586
rect 35250 21534 35252 21586
rect 35196 21532 35252 21534
rect 35644 22482 35700 22484
rect 35644 22430 35646 22482
rect 35646 22430 35698 22482
rect 35698 22430 35700 22482
rect 35644 22428 35700 22430
rect 35868 21756 35924 21812
rect 35196 21194 35252 21196
rect 35196 21142 35198 21194
rect 35198 21142 35250 21194
rect 35250 21142 35252 21194
rect 35196 21140 35252 21142
rect 35300 21194 35356 21196
rect 35300 21142 35302 21194
rect 35302 21142 35354 21194
rect 35354 21142 35356 21194
rect 35300 21140 35356 21142
rect 35404 21194 35460 21196
rect 35404 21142 35406 21194
rect 35406 21142 35458 21194
rect 35458 21142 35460 21194
rect 35404 21140 35460 21142
rect 34860 20188 34916 20244
rect 34860 20018 34916 20020
rect 34860 19966 34862 20018
rect 34862 19966 34914 20018
rect 34914 19966 34916 20018
rect 34860 19964 34916 19966
rect 34748 19740 34804 19796
rect 35084 20188 35140 20244
rect 34972 19346 35028 19348
rect 34972 19294 34974 19346
rect 34974 19294 35026 19346
rect 35026 19294 35028 19346
rect 34972 19292 35028 19294
rect 35196 19626 35252 19628
rect 35196 19574 35198 19626
rect 35198 19574 35250 19626
rect 35250 19574 35252 19626
rect 35196 19572 35252 19574
rect 35300 19626 35356 19628
rect 35300 19574 35302 19626
rect 35302 19574 35354 19626
rect 35354 19574 35356 19626
rect 35300 19572 35356 19574
rect 35404 19626 35460 19628
rect 35404 19574 35406 19626
rect 35406 19574 35458 19626
rect 35458 19574 35460 19626
rect 35404 19572 35460 19574
rect 35308 19458 35364 19460
rect 35308 19406 35310 19458
rect 35310 19406 35362 19458
rect 35362 19406 35364 19458
rect 35308 19404 35364 19406
rect 35420 19292 35476 19348
rect 35084 18844 35140 18900
rect 35420 18508 35476 18564
rect 35084 18338 35140 18340
rect 35084 18286 35086 18338
rect 35086 18286 35138 18338
rect 35138 18286 35140 18338
rect 35084 18284 35140 18286
rect 34972 18172 35028 18228
rect 35756 20578 35812 20580
rect 35756 20526 35758 20578
rect 35758 20526 35810 20578
rect 35810 20526 35812 20578
rect 35756 20524 35812 20526
rect 36316 23212 36372 23268
rect 36428 22764 36484 22820
rect 36316 22370 36372 22372
rect 36316 22318 36318 22370
rect 36318 22318 36370 22370
rect 36370 22318 36372 22370
rect 36316 22316 36372 22318
rect 36428 21698 36484 21700
rect 36428 21646 36430 21698
rect 36430 21646 36482 21698
rect 36482 21646 36484 21698
rect 36428 21644 36484 21646
rect 35644 20300 35700 20356
rect 36092 20300 36148 20356
rect 35644 19404 35700 19460
rect 36204 19404 36260 19460
rect 35756 19234 35812 19236
rect 35756 19182 35758 19234
rect 35758 19182 35810 19234
rect 35810 19182 35812 19234
rect 35756 19180 35812 19182
rect 36092 19292 36148 19348
rect 35644 18620 35700 18676
rect 35196 18058 35252 18060
rect 35196 18006 35198 18058
rect 35198 18006 35250 18058
rect 35250 18006 35252 18058
rect 35196 18004 35252 18006
rect 35300 18058 35356 18060
rect 35300 18006 35302 18058
rect 35302 18006 35354 18058
rect 35354 18006 35356 18058
rect 35300 18004 35356 18006
rect 35404 18058 35460 18060
rect 35404 18006 35406 18058
rect 35406 18006 35458 18058
rect 35458 18006 35460 18058
rect 35404 18004 35460 18006
rect 35196 17612 35252 17668
rect 34748 17554 34804 17556
rect 34748 17502 34750 17554
rect 34750 17502 34802 17554
rect 34802 17502 34804 17554
rect 34748 17500 34804 17502
rect 35756 18284 35812 18340
rect 36988 31052 37044 31108
rect 38108 30994 38164 30996
rect 38108 30942 38110 30994
rect 38110 30942 38162 30994
rect 38162 30942 38164 30994
rect 38108 30940 38164 30942
rect 38332 30828 38388 30884
rect 36988 30716 37044 30772
rect 36652 29596 36708 29652
rect 38332 30044 38388 30100
rect 37100 29986 37156 29988
rect 37100 29934 37102 29986
rect 37102 29934 37154 29986
rect 37154 29934 37156 29986
rect 37100 29932 37156 29934
rect 39452 31948 39508 32004
rect 40796 34860 40852 34916
rect 40684 34076 40740 34132
rect 40908 34748 40964 34804
rect 41132 34524 41188 34580
rect 40908 34242 40964 34244
rect 40908 34190 40910 34242
rect 40910 34190 40962 34242
rect 40962 34190 40964 34242
rect 40908 34188 40964 34190
rect 41020 34076 41076 34132
rect 41580 36204 41636 36260
rect 41468 34524 41524 34580
rect 41804 34524 41860 34580
rect 42252 35532 42308 35588
rect 43708 37826 43764 37828
rect 43708 37774 43710 37826
rect 43710 37774 43762 37826
rect 43762 37774 43764 37826
rect 43708 37772 43764 37774
rect 42812 37436 42868 37492
rect 42812 36482 42868 36484
rect 42812 36430 42814 36482
rect 42814 36430 42866 36482
rect 42866 36430 42868 36482
rect 42812 36428 42868 36430
rect 43260 36988 43316 37044
rect 42700 35868 42756 35924
rect 42588 35420 42644 35476
rect 45164 37266 45220 37268
rect 45164 37214 45166 37266
rect 45166 37214 45218 37266
rect 45218 37214 45220 37266
rect 45164 37212 45220 37214
rect 43820 36988 43876 37044
rect 44716 36988 44772 37044
rect 44940 36876 44996 36932
rect 43484 36594 43540 36596
rect 43484 36542 43486 36594
rect 43486 36542 43538 36594
rect 43538 36542 43540 36594
rect 43484 36540 43540 36542
rect 44380 36540 44436 36596
rect 43372 36258 43428 36260
rect 43372 36206 43374 36258
rect 43374 36206 43426 36258
rect 43426 36206 43428 36258
rect 43372 36204 43428 36206
rect 44268 35644 44324 35700
rect 44156 35420 44212 35476
rect 42364 34690 42420 34692
rect 42364 34638 42366 34690
rect 42366 34638 42418 34690
rect 42418 34638 42420 34690
rect 42364 34636 42420 34638
rect 43148 34802 43204 34804
rect 43148 34750 43150 34802
rect 43150 34750 43202 34802
rect 43202 34750 43204 34802
rect 43148 34748 43204 34750
rect 43932 34802 43988 34804
rect 43932 34750 43934 34802
rect 43934 34750 43986 34802
rect 43986 34750 43988 34802
rect 43932 34748 43988 34750
rect 42700 34524 42756 34580
rect 40684 33122 40740 33124
rect 40684 33070 40686 33122
rect 40686 33070 40738 33122
rect 40738 33070 40740 33122
rect 40684 33068 40740 33070
rect 41020 33122 41076 33124
rect 41020 33070 41022 33122
rect 41022 33070 41074 33122
rect 41074 33070 41076 33122
rect 41020 33068 41076 33070
rect 39900 32284 39956 32340
rect 39004 31890 39060 31892
rect 39004 31838 39006 31890
rect 39006 31838 39058 31890
rect 39058 31838 39060 31890
rect 39004 31836 39060 31838
rect 38892 31554 38948 31556
rect 38892 31502 38894 31554
rect 38894 31502 38946 31554
rect 38946 31502 38948 31554
rect 38892 31500 38948 31502
rect 38556 29932 38612 29988
rect 37436 29484 37492 29540
rect 37212 29426 37268 29428
rect 37212 29374 37214 29426
rect 37214 29374 37266 29426
rect 37266 29374 37268 29426
rect 37212 29372 37268 29374
rect 36988 28642 37044 28644
rect 36988 28590 36990 28642
rect 36990 28590 37042 28642
rect 37042 28590 37044 28642
rect 36988 28588 37044 28590
rect 37100 28476 37156 28532
rect 36652 28140 36708 28196
rect 36988 28140 37044 28196
rect 36652 27916 36708 27972
rect 36876 26178 36932 26180
rect 36876 26126 36878 26178
rect 36878 26126 36930 26178
rect 36930 26126 36932 26178
rect 36876 26124 36932 26126
rect 37548 29372 37604 29428
rect 38108 29314 38164 29316
rect 38108 29262 38110 29314
rect 38110 29262 38162 29314
rect 38162 29262 38164 29314
rect 38108 29260 38164 29262
rect 37548 28812 37604 28868
rect 36764 22428 36820 22484
rect 38108 28418 38164 28420
rect 38108 28366 38110 28418
rect 38110 28366 38162 28418
rect 38162 28366 38164 28418
rect 38108 28364 38164 28366
rect 38332 29426 38388 29428
rect 38332 29374 38334 29426
rect 38334 29374 38386 29426
rect 38386 29374 38388 29426
rect 38332 29372 38388 29374
rect 38332 28700 38388 28756
rect 37772 27074 37828 27076
rect 37772 27022 37774 27074
rect 37774 27022 37826 27074
rect 37826 27022 37828 27074
rect 37772 27020 37828 27022
rect 37324 26962 37380 26964
rect 37324 26910 37326 26962
rect 37326 26910 37378 26962
rect 37378 26910 37380 26962
rect 37324 26908 37380 26910
rect 37548 26962 37604 26964
rect 37548 26910 37550 26962
rect 37550 26910 37602 26962
rect 37602 26910 37604 26962
rect 37548 26908 37604 26910
rect 37996 26850 38052 26852
rect 37996 26798 37998 26850
rect 37998 26798 38050 26850
rect 38050 26798 38052 26850
rect 37996 26796 38052 26798
rect 37212 26572 37268 26628
rect 37100 24108 37156 24164
rect 36988 23826 37044 23828
rect 36988 23774 36990 23826
rect 36990 23774 37042 23826
rect 37042 23774 37044 23826
rect 36988 23772 37044 23774
rect 37884 26290 37940 26292
rect 37884 26238 37886 26290
rect 37886 26238 37938 26290
rect 37938 26238 37940 26290
rect 37884 26236 37940 26238
rect 37436 23938 37492 23940
rect 37436 23886 37438 23938
rect 37438 23886 37490 23938
rect 37490 23886 37492 23938
rect 37436 23884 37492 23886
rect 37996 23938 38052 23940
rect 37996 23886 37998 23938
rect 37998 23886 38050 23938
rect 38050 23886 38052 23938
rect 37996 23884 38052 23886
rect 37324 23772 37380 23828
rect 36876 21868 36932 21924
rect 37100 22764 37156 22820
rect 37548 22370 37604 22372
rect 37548 22318 37550 22370
rect 37550 22318 37602 22370
rect 37602 22318 37604 22370
rect 37548 22316 37604 22318
rect 37996 21756 38052 21812
rect 38780 30940 38836 30996
rect 39340 30994 39396 30996
rect 39340 30942 39342 30994
rect 39342 30942 39394 30994
rect 39394 30942 39396 30994
rect 39340 30940 39396 30942
rect 39452 30828 39508 30884
rect 39228 30210 39284 30212
rect 39228 30158 39230 30210
rect 39230 30158 39282 30210
rect 39282 30158 39284 30210
rect 39228 30156 39284 30158
rect 39564 30604 39620 30660
rect 39340 29986 39396 29988
rect 39340 29934 39342 29986
rect 39342 29934 39394 29986
rect 39394 29934 39396 29986
rect 39340 29932 39396 29934
rect 38780 29820 38836 29876
rect 39004 29820 39060 29876
rect 38668 28754 38724 28756
rect 38668 28702 38670 28754
rect 38670 28702 38722 28754
rect 38722 28702 38724 28754
rect 38668 28700 38724 28702
rect 38556 27020 38612 27076
rect 38332 26572 38388 26628
rect 38780 24108 38836 24164
rect 38668 23772 38724 23828
rect 38332 21756 38388 21812
rect 38556 21586 38612 21588
rect 38556 21534 38558 21586
rect 38558 21534 38610 21586
rect 38610 21534 38612 21586
rect 38556 21532 38612 21534
rect 38108 21420 38164 21476
rect 39788 29820 39844 29876
rect 39900 31164 39956 31220
rect 43036 32786 43092 32788
rect 43036 32734 43038 32786
rect 43038 32734 43090 32786
rect 43090 32734 43092 32786
rect 43036 32732 43092 32734
rect 43596 34690 43652 34692
rect 43596 34638 43598 34690
rect 43598 34638 43650 34690
rect 43650 34638 43652 34690
rect 43596 34636 43652 34638
rect 44716 35586 44772 35588
rect 44716 35534 44718 35586
rect 44718 35534 44770 35586
rect 44770 35534 44772 35586
rect 44716 35532 44772 35534
rect 45164 36428 45220 36484
rect 45164 35922 45220 35924
rect 45164 35870 45166 35922
rect 45166 35870 45218 35922
rect 45218 35870 45220 35922
rect 45164 35868 45220 35870
rect 45836 37154 45892 37156
rect 45836 37102 45838 37154
rect 45838 37102 45890 37154
rect 45890 37102 45892 37154
rect 45836 37100 45892 37102
rect 45500 35922 45556 35924
rect 45500 35870 45502 35922
rect 45502 35870 45554 35922
rect 45554 35870 45556 35922
rect 45500 35868 45556 35870
rect 45836 35922 45892 35924
rect 45836 35870 45838 35922
rect 45838 35870 45890 35922
rect 45890 35870 45892 35922
rect 45836 35868 45892 35870
rect 45388 35420 45444 35476
rect 44828 34802 44884 34804
rect 44828 34750 44830 34802
rect 44830 34750 44882 34802
rect 44882 34750 44884 34802
rect 44828 34748 44884 34750
rect 45948 34690 46004 34692
rect 45948 34638 45950 34690
rect 45950 34638 46002 34690
rect 46002 34638 46004 34690
rect 45948 34636 46004 34638
rect 45724 34412 45780 34468
rect 45612 34242 45668 34244
rect 45612 34190 45614 34242
rect 45614 34190 45666 34242
rect 45666 34190 45668 34242
rect 45612 34188 45668 34190
rect 44380 33852 44436 33908
rect 44156 33068 44212 33124
rect 43148 31836 43204 31892
rect 42812 31724 42868 31780
rect 40572 30210 40628 30212
rect 40572 30158 40574 30210
rect 40574 30158 40626 30210
rect 40626 30158 40628 30210
rect 40572 30156 40628 30158
rect 40012 30044 40068 30100
rect 40796 30044 40852 30100
rect 40460 29986 40516 29988
rect 40460 29934 40462 29986
rect 40462 29934 40514 29986
rect 40514 29934 40516 29986
rect 40460 29932 40516 29934
rect 39452 29148 39508 29204
rect 40012 29148 40068 29204
rect 39116 28530 39172 28532
rect 39116 28478 39118 28530
rect 39118 28478 39170 28530
rect 39170 28478 39172 28530
rect 39116 28476 39172 28478
rect 39788 27916 39844 27972
rect 41244 31218 41300 31220
rect 41244 31166 41246 31218
rect 41246 31166 41298 31218
rect 41298 31166 41300 31218
rect 41244 31164 41300 31166
rect 42812 31164 42868 31220
rect 41356 30994 41412 30996
rect 41356 30942 41358 30994
rect 41358 30942 41410 30994
rect 41410 30942 41412 30994
rect 41356 30940 41412 30942
rect 42252 30716 42308 30772
rect 41132 29538 41188 29540
rect 41132 29486 41134 29538
rect 41134 29486 41186 29538
rect 41186 29486 41188 29538
rect 41132 29484 41188 29486
rect 42140 30044 42196 30100
rect 41468 29932 41524 29988
rect 41356 29820 41412 29876
rect 40460 29372 40516 29428
rect 42476 30940 42532 30996
rect 40236 28588 40292 28644
rect 40012 28028 40068 28084
rect 39116 26908 39172 26964
rect 39004 26796 39060 26852
rect 37100 20578 37156 20580
rect 37100 20526 37102 20578
rect 37102 20526 37154 20578
rect 37154 20526 37156 20578
rect 37100 20524 37156 20526
rect 37212 19628 37268 19684
rect 37660 20524 37716 20580
rect 36652 19292 36708 19348
rect 36540 18956 36596 19012
rect 36316 18732 36372 18788
rect 35980 18172 36036 18228
rect 36092 18508 36148 18564
rect 35868 18060 35924 18116
rect 35644 17276 35700 17332
rect 34748 16882 34804 16884
rect 34748 16830 34750 16882
rect 34750 16830 34802 16882
rect 34802 16830 34804 16882
rect 34748 16828 34804 16830
rect 34748 16044 34804 16100
rect 35756 17106 35812 17108
rect 35756 17054 35758 17106
rect 35758 17054 35810 17106
rect 35810 17054 35812 17106
rect 35756 17052 35812 17054
rect 35644 16828 35700 16884
rect 32844 15708 32900 15764
rect 35420 16604 35476 16660
rect 33404 15596 33460 15652
rect 31612 12124 31668 12180
rect 32508 12908 32564 12964
rect 32508 12348 32564 12404
rect 32284 12236 32340 12292
rect 31948 11676 32004 11732
rect 32620 11900 32676 11956
rect 33292 15538 33348 15540
rect 33292 15486 33294 15538
rect 33294 15486 33346 15538
rect 33346 15486 33348 15538
rect 33292 15484 33348 15486
rect 33068 15372 33124 15428
rect 33516 15260 33572 15316
rect 33180 15202 33236 15204
rect 33180 15150 33182 15202
rect 33182 15150 33234 15202
rect 33234 15150 33236 15202
rect 33180 15148 33236 15150
rect 33964 15314 34020 15316
rect 33964 15262 33966 15314
rect 33966 15262 34018 15314
rect 34018 15262 34020 15314
rect 33964 15260 34020 15262
rect 33628 14924 33684 14980
rect 33404 13858 33460 13860
rect 33404 13806 33406 13858
rect 33406 13806 33458 13858
rect 33458 13806 33460 13858
rect 33404 13804 33460 13806
rect 34748 14812 34804 14868
rect 35196 16490 35252 16492
rect 35196 16438 35198 16490
rect 35198 16438 35250 16490
rect 35250 16438 35252 16490
rect 35196 16436 35252 16438
rect 35300 16490 35356 16492
rect 35300 16438 35302 16490
rect 35302 16438 35354 16490
rect 35354 16438 35356 16490
rect 35300 16436 35356 16438
rect 35404 16490 35460 16492
rect 35404 16438 35406 16490
rect 35406 16438 35458 16490
rect 35458 16438 35460 16490
rect 35404 16436 35460 16438
rect 35644 16098 35700 16100
rect 35644 16046 35646 16098
rect 35646 16046 35698 16098
rect 35698 16046 35700 16098
rect 35644 16044 35700 16046
rect 35196 15596 35252 15652
rect 35308 15314 35364 15316
rect 35308 15262 35310 15314
rect 35310 15262 35362 15314
rect 35362 15262 35364 15314
rect 35308 15260 35364 15262
rect 35420 15036 35476 15092
rect 36204 17388 36260 17444
rect 36204 17052 36260 17108
rect 36652 18396 36708 18452
rect 36652 17724 36708 17780
rect 36540 17612 36596 17668
rect 36540 17164 36596 17220
rect 36652 17052 36708 17108
rect 36540 16828 36596 16884
rect 35980 15820 36036 15876
rect 36316 15820 36372 15876
rect 35980 15596 36036 15652
rect 35644 15148 35700 15204
rect 35196 14922 35252 14924
rect 35196 14870 35198 14922
rect 35198 14870 35250 14922
rect 35250 14870 35252 14922
rect 35196 14868 35252 14870
rect 35300 14922 35356 14924
rect 35300 14870 35302 14922
rect 35302 14870 35354 14922
rect 35354 14870 35356 14922
rect 35300 14868 35356 14870
rect 35404 14922 35460 14924
rect 35404 14870 35406 14922
rect 35406 14870 35458 14922
rect 35458 14870 35460 14922
rect 35404 14868 35460 14870
rect 35084 14700 35140 14756
rect 35980 15036 36036 15092
rect 34300 13804 34356 13860
rect 35756 14476 35812 14532
rect 35532 14364 35588 14420
rect 34972 13804 35028 13860
rect 34076 13580 34132 13636
rect 33964 12796 34020 12852
rect 33292 12402 33348 12404
rect 33292 12350 33294 12402
rect 33294 12350 33346 12402
rect 33346 12350 33348 12402
rect 33292 12348 33348 12350
rect 35084 14252 35140 14308
rect 35196 13858 35252 13860
rect 35196 13806 35198 13858
rect 35198 13806 35250 13858
rect 35250 13806 35252 13858
rect 35196 13804 35252 13806
rect 35084 13692 35140 13748
rect 35196 13354 35252 13356
rect 35196 13302 35198 13354
rect 35198 13302 35250 13354
rect 35250 13302 35252 13354
rect 35196 13300 35252 13302
rect 35300 13354 35356 13356
rect 35300 13302 35302 13354
rect 35302 13302 35354 13354
rect 35354 13302 35356 13354
rect 35300 13300 35356 13302
rect 35404 13354 35460 13356
rect 35404 13302 35406 13354
rect 35406 13302 35458 13354
rect 35458 13302 35460 13354
rect 35404 13300 35460 13302
rect 34188 12850 34244 12852
rect 34188 12798 34190 12850
rect 34190 12798 34242 12850
rect 34242 12798 34244 12850
rect 34188 12796 34244 12798
rect 31948 11228 32004 11284
rect 31276 9826 31332 9828
rect 31276 9774 31278 9826
rect 31278 9774 31330 9826
rect 31330 9774 31332 9826
rect 31276 9772 31332 9774
rect 33180 11900 33236 11956
rect 32396 10108 32452 10164
rect 32508 9826 32564 9828
rect 32508 9774 32510 9826
rect 32510 9774 32562 9826
rect 32562 9774 32564 9826
rect 32508 9772 32564 9774
rect 33068 10722 33124 10724
rect 33068 10670 33070 10722
rect 33070 10670 33122 10722
rect 33122 10670 33124 10722
rect 33068 10668 33124 10670
rect 33180 9884 33236 9940
rect 31612 8876 31668 8932
rect 33740 11340 33796 11396
rect 33740 10444 33796 10500
rect 34748 11900 34804 11956
rect 33516 9884 33572 9940
rect 33628 9772 33684 9828
rect 33180 8876 33236 8932
rect 34748 10444 34804 10500
rect 35308 12066 35364 12068
rect 35308 12014 35310 12066
rect 35310 12014 35362 12066
rect 35362 12014 35364 12066
rect 35308 12012 35364 12014
rect 35196 11786 35252 11788
rect 35196 11734 35198 11786
rect 35198 11734 35250 11786
rect 35250 11734 35252 11786
rect 35196 11732 35252 11734
rect 35300 11786 35356 11788
rect 35300 11734 35302 11786
rect 35302 11734 35354 11786
rect 35354 11734 35356 11786
rect 35300 11732 35356 11734
rect 35404 11786 35460 11788
rect 35404 11734 35406 11786
rect 35406 11734 35458 11786
rect 35458 11734 35460 11786
rect 35404 11732 35460 11734
rect 36316 15260 36372 15316
rect 37100 19458 37156 19460
rect 37100 19406 37102 19458
rect 37102 19406 37154 19458
rect 37154 19406 37156 19458
rect 37100 19404 37156 19406
rect 37100 19122 37156 19124
rect 37100 19070 37102 19122
rect 37102 19070 37154 19122
rect 37154 19070 37156 19122
rect 37100 19068 37156 19070
rect 37324 18562 37380 18564
rect 37324 18510 37326 18562
rect 37326 18510 37378 18562
rect 37378 18510 37380 18562
rect 37324 18508 37380 18510
rect 36988 18060 37044 18116
rect 37212 18338 37268 18340
rect 37212 18286 37214 18338
rect 37214 18286 37266 18338
rect 37266 18286 37268 18338
rect 37212 18284 37268 18286
rect 37660 19346 37716 19348
rect 37660 19294 37662 19346
rect 37662 19294 37714 19346
rect 37714 19294 37716 19346
rect 37660 19292 37716 19294
rect 39340 26852 39396 26908
rect 40348 27804 40404 27860
rect 40348 27074 40404 27076
rect 40348 27022 40350 27074
rect 40350 27022 40402 27074
rect 40402 27022 40404 27074
rect 40348 27020 40404 27022
rect 40012 26796 40068 26852
rect 39340 26348 39396 26404
rect 40236 25228 40292 25284
rect 39116 24050 39172 24052
rect 39116 23998 39118 24050
rect 39118 23998 39170 24050
rect 39170 23998 39172 24050
rect 39116 23996 39172 23998
rect 39228 23884 39284 23940
rect 39004 22428 39060 22484
rect 38108 20188 38164 20244
rect 38892 21420 38948 21476
rect 38108 19180 38164 19236
rect 37660 18284 37716 18340
rect 36988 17500 37044 17556
rect 36988 17052 37044 17108
rect 37212 16940 37268 16996
rect 37324 17500 37380 17556
rect 37100 16828 37156 16884
rect 37324 15820 37380 15876
rect 36988 14418 37044 14420
rect 36988 14366 36990 14418
rect 36990 14366 37042 14418
rect 37042 14366 37044 14418
rect 36988 14364 37044 14366
rect 35868 13074 35924 13076
rect 35868 13022 35870 13074
rect 35870 13022 35922 13074
rect 35922 13022 35924 13074
rect 35868 13020 35924 13022
rect 37324 14364 37380 14420
rect 37212 14306 37268 14308
rect 37212 14254 37214 14306
rect 37214 14254 37266 14306
rect 37266 14254 37268 14306
rect 37212 14252 37268 14254
rect 36764 13858 36820 13860
rect 36764 13806 36766 13858
rect 36766 13806 36818 13858
rect 36818 13806 36820 13858
rect 36764 13804 36820 13806
rect 35756 12066 35812 12068
rect 35756 12014 35758 12066
rect 35758 12014 35810 12066
rect 35810 12014 35812 12066
rect 35756 12012 35812 12014
rect 35756 10722 35812 10724
rect 35756 10670 35758 10722
rect 35758 10670 35810 10722
rect 35810 10670 35812 10722
rect 35756 10668 35812 10670
rect 35644 10556 35700 10612
rect 34972 10332 35028 10388
rect 35196 10218 35252 10220
rect 35196 10166 35198 10218
rect 35198 10166 35250 10218
rect 35250 10166 35252 10218
rect 35196 10164 35252 10166
rect 35300 10218 35356 10220
rect 35300 10166 35302 10218
rect 35302 10166 35354 10218
rect 35354 10166 35356 10218
rect 35300 10164 35356 10166
rect 35404 10218 35460 10220
rect 35404 10166 35406 10218
rect 35406 10166 35458 10218
rect 35458 10166 35460 10218
rect 35404 10164 35460 10166
rect 34188 9772 34244 9828
rect 36316 12796 36372 12852
rect 36204 12012 36260 12068
rect 36204 10386 36260 10388
rect 36204 10334 36206 10386
rect 36206 10334 36258 10386
rect 36258 10334 36260 10386
rect 36204 10332 36260 10334
rect 36764 13020 36820 13076
rect 36428 9938 36484 9940
rect 36428 9886 36430 9938
rect 36430 9886 36482 9938
rect 36482 9886 36484 9938
rect 36428 9884 36484 9886
rect 36204 9212 36260 9268
rect 36316 8930 36372 8932
rect 36316 8878 36318 8930
rect 36318 8878 36370 8930
rect 36370 8878 36372 8930
rect 36316 8876 36372 8878
rect 37436 13692 37492 13748
rect 37324 13468 37380 13524
rect 37324 12796 37380 12852
rect 37324 12348 37380 12404
rect 37436 12124 37492 12180
rect 37212 11676 37268 11732
rect 37324 11452 37380 11508
rect 36764 10668 36820 10724
rect 37100 11116 37156 11172
rect 36988 9884 37044 9940
rect 35196 8650 35252 8652
rect 35196 8598 35198 8650
rect 35198 8598 35250 8650
rect 35250 8598 35252 8650
rect 35196 8596 35252 8598
rect 35300 8650 35356 8652
rect 35300 8598 35302 8650
rect 35302 8598 35354 8650
rect 35354 8598 35356 8650
rect 35300 8596 35356 8598
rect 35404 8650 35460 8652
rect 35404 8598 35406 8650
rect 35406 8598 35458 8650
rect 35458 8598 35460 8650
rect 35404 8596 35460 8598
rect 36988 8876 37044 8932
rect 36428 8146 36484 8148
rect 36428 8094 36430 8146
rect 36430 8094 36482 8146
rect 36482 8094 36484 8146
rect 36428 8092 36484 8094
rect 37212 10610 37268 10612
rect 37212 10558 37214 10610
rect 37214 10558 37266 10610
rect 37266 10558 37268 10610
rect 37212 10556 37268 10558
rect 35196 7082 35252 7084
rect 35196 7030 35198 7082
rect 35198 7030 35250 7082
rect 35250 7030 35252 7082
rect 35196 7028 35252 7030
rect 35300 7082 35356 7084
rect 35300 7030 35302 7082
rect 35302 7030 35354 7082
rect 35354 7030 35356 7082
rect 35300 7028 35356 7030
rect 35404 7082 35460 7084
rect 35404 7030 35406 7082
rect 35406 7030 35458 7082
rect 35458 7030 35460 7082
rect 35404 7028 35460 7030
rect 35196 5514 35252 5516
rect 35196 5462 35198 5514
rect 35198 5462 35250 5514
rect 35250 5462 35252 5514
rect 35196 5460 35252 5462
rect 35300 5514 35356 5516
rect 35300 5462 35302 5514
rect 35302 5462 35354 5514
rect 35354 5462 35356 5514
rect 35300 5460 35356 5462
rect 35404 5514 35460 5516
rect 35404 5462 35406 5514
rect 35406 5462 35458 5514
rect 35458 5462 35460 5514
rect 35404 5460 35460 5462
rect 34860 4956 34916 5012
rect 34188 3442 34244 3444
rect 34188 3390 34190 3442
rect 34190 3390 34242 3442
rect 34242 3390 34244 3442
rect 34188 3388 34244 3390
rect 35196 3946 35252 3948
rect 35196 3894 35198 3946
rect 35198 3894 35250 3946
rect 35250 3894 35252 3946
rect 35196 3892 35252 3894
rect 35300 3946 35356 3948
rect 35300 3894 35302 3946
rect 35302 3894 35354 3946
rect 35354 3894 35356 3946
rect 35300 3892 35356 3894
rect 35404 3946 35460 3948
rect 35404 3894 35406 3946
rect 35406 3894 35458 3946
rect 35458 3894 35460 3946
rect 35404 3892 35460 3894
rect 36316 3442 36372 3444
rect 36316 3390 36318 3442
rect 36318 3390 36370 3442
rect 36370 3390 36372 3442
rect 36316 3388 36372 3390
rect 37212 3388 37268 3444
rect 37884 17948 37940 18004
rect 37660 17052 37716 17108
rect 38556 19122 38612 19124
rect 38556 19070 38558 19122
rect 38558 19070 38610 19122
rect 38610 19070 38612 19122
rect 38556 19068 38612 19070
rect 38332 18060 38388 18116
rect 41132 28700 41188 28756
rect 41020 28588 41076 28644
rect 40908 28082 40964 28084
rect 40908 28030 40910 28082
rect 40910 28030 40962 28082
rect 40962 28030 40964 28082
rect 40908 28028 40964 28030
rect 40460 24108 40516 24164
rect 40348 23996 40404 24052
rect 40236 23884 40292 23940
rect 39788 23212 39844 23268
rect 41244 27858 41300 27860
rect 41244 27806 41246 27858
rect 41246 27806 41298 27858
rect 41298 27806 41300 27858
rect 41244 27804 41300 27806
rect 41692 27804 41748 27860
rect 41244 27580 41300 27636
rect 41580 27186 41636 27188
rect 41580 27134 41582 27186
rect 41582 27134 41634 27186
rect 41634 27134 41636 27186
rect 41580 27132 41636 27134
rect 42700 29932 42756 29988
rect 43260 31724 43316 31780
rect 43708 32732 43764 32788
rect 44044 31890 44100 31892
rect 44044 31838 44046 31890
rect 44046 31838 44098 31890
rect 44098 31838 44100 31890
rect 44044 31836 44100 31838
rect 42924 30716 42980 30772
rect 42812 29820 42868 29876
rect 42476 28140 42532 28196
rect 42700 28588 42756 28644
rect 42140 27074 42196 27076
rect 42140 27022 42142 27074
rect 42142 27022 42194 27074
rect 42194 27022 42196 27074
rect 42140 27020 42196 27022
rect 42476 27132 42532 27188
rect 43148 30994 43204 30996
rect 43148 30942 43150 30994
rect 43150 30942 43202 30994
rect 43202 30942 43204 30994
rect 43148 30940 43204 30942
rect 43148 30604 43204 30660
rect 43260 30716 43316 30772
rect 43260 30210 43316 30212
rect 43260 30158 43262 30210
rect 43262 30158 43314 30210
rect 43314 30158 43316 30210
rect 43260 30156 43316 30158
rect 42028 26850 42084 26852
rect 42028 26798 42030 26850
rect 42030 26798 42082 26850
rect 42082 26798 42084 26850
rect 42028 26796 42084 26798
rect 44380 29596 44436 29652
rect 44268 29148 44324 29204
rect 43484 28364 43540 28420
rect 43484 28140 43540 28196
rect 43484 27244 43540 27300
rect 43260 27074 43316 27076
rect 43260 27022 43262 27074
rect 43262 27022 43314 27074
rect 43314 27022 43316 27074
rect 43260 27020 43316 27022
rect 44044 28418 44100 28420
rect 44044 28366 44046 28418
rect 44046 28366 44098 28418
rect 44098 28366 44100 28418
rect 44044 28364 44100 28366
rect 43932 27244 43988 27300
rect 41020 25282 41076 25284
rect 41020 25230 41022 25282
rect 41022 25230 41074 25282
rect 41074 25230 41076 25282
rect 41020 25228 41076 25230
rect 40908 22876 40964 22932
rect 40124 21810 40180 21812
rect 40124 21758 40126 21810
rect 40126 21758 40178 21810
rect 40178 21758 40180 21810
rect 40124 21756 40180 21758
rect 40012 21532 40068 21588
rect 40460 21532 40516 21588
rect 40348 20748 40404 20804
rect 39452 20130 39508 20132
rect 39452 20078 39454 20130
rect 39454 20078 39506 20130
rect 39506 20078 39508 20130
rect 39452 20076 39508 20078
rect 39900 19740 39956 19796
rect 39116 18450 39172 18452
rect 39116 18398 39118 18450
rect 39118 18398 39170 18450
rect 39170 18398 39172 18450
rect 39116 18396 39172 18398
rect 39340 18396 39396 18452
rect 38668 17724 38724 17780
rect 38556 16828 38612 16884
rect 37884 15260 37940 15316
rect 38892 17948 38948 18004
rect 38556 15932 38612 15988
rect 38444 15874 38500 15876
rect 38444 15822 38446 15874
rect 38446 15822 38498 15874
rect 38498 15822 38500 15874
rect 38444 15820 38500 15822
rect 37884 14924 37940 14980
rect 38332 14530 38388 14532
rect 38332 14478 38334 14530
rect 38334 14478 38386 14530
rect 38386 14478 38388 14530
rect 38332 14476 38388 14478
rect 37996 14364 38052 14420
rect 38220 13916 38276 13972
rect 38444 13746 38500 13748
rect 38444 13694 38446 13746
rect 38446 13694 38498 13746
rect 38498 13694 38500 13746
rect 38444 13692 38500 13694
rect 37996 13580 38052 13636
rect 37660 13356 37716 13412
rect 38108 13522 38164 13524
rect 38108 13470 38110 13522
rect 38110 13470 38162 13522
rect 38162 13470 38164 13522
rect 38108 13468 38164 13470
rect 37660 12012 37716 12068
rect 37772 12796 37828 12852
rect 37660 10498 37716 10500
rect 37660 10446 37662 10498
rect 37662 10446 37714 10498
rect 37714 10446 37716 10498
rect 37660 10444 37716 10446
rect 37772 9436 37828 9492
rect 37772 8146 37828 8148
rect 37772 8094 37774 8146
rect 37774 8094 37826 8146
rect 37826 8094 37828 8146
rect 37772 8092 37828 8094
rect 38108 12012 38164 12068
rect 37996 11452 38052 11508
rect 38108 11004 38164 11060
rect 39228 18060 39284 18116
rect 39228 17052 39284 17108
rect 39116 16994 39172 16996
rect 39116 16942 39118 16994
rect 39118 16942 39170 16994
rect 39170 16942 39172 16994
rect 39116 16940 39172 16942
rect 40236 19740 40292 19796
rect 40236 18732 40292 18788
rect 40348 18674 40404 18676
rect 40348 18622 40350 18674
rect 40350 18622 40402 18674
rect 40402 18622 40404 18674
rect 40348 18620 40404 18622
rect 40236 18508 40292 18564
rect 40012 18284 40068 18340
rect 39564 17724 39620 17780
rect 40796 22540 40852 22596
rect 40796 21868 40852 21924
rect 40684 20578 40740 20580
rect 40684 20526 40686 20578
rect 40686 20526 40738 20578
rect 40738 20526 40740 20578
rect 40684 20524 40740 20526
rect 41020 21868 41076 21924
rect 41244 23826 41300 23828
rect 41244 23774 41246 23826
rect 41246 23774 41298 23826
rect 41298 23774 41300 23826
rect 41244 23772 41300 23774
rect 41244 22876 41300 22932
rect 41580 23212 41636 23268
rect 41692 23996 41748 24052
rect 41468 23100 41524 23156
rect 42028 23548 42084 23604
rect 42140 23154 42196 23156
rect 42140 23102 42142 23154
rect 42142 23102 42194 23154
rect 42194 23102 42196 23154
rect 42140 23100 42196 23102
rect 42140 22482 42196 22484
rect 42140 22430 42142 22482
rect 42142 22430 42194 22482
rect 42194 22430 42196 22482
rect 42140 22428 42196 22430
rect 42364 26236 42420 26292
rect 43148 26290 43204 26292
rect 43148 26238 43150 26290
rect 43150 26238 43202 26290
rect 43202 26238 43204 26290
rect 43148 26236 43204 26238
rect 42700 26124 42756 26180
rect 41916 21868 41972 21924
rect 41468 21810 41524 21812
rect 41468 21758 41470 21810
rect 41470 21758 41522 21810
rect 41522 21758 41524 21810
rect 41468 21756 41524 21758
rect 42140 21756 42196 21812
rect 41356 20860 41412 20916
rect 41132 20524 41188 20580
rect 41244 20636 41300 20692
rect 40796 19180 40852 19236
rect 40684 18732 40740 18788
rect 40796 18620 40852 18676
rect 40908 18562 40964 18564
rect 40908 18510 40910 18562
rect 40910 18510 40962 18562
rect 40962 18510 40964 18562
rect 40908 18508 40964 18510
rect 41020 18338 41076 18340
rect 41020 18286 41022 18338
rect 41022 18286 41074 18338
rect 41074 18286 41076 18338
rect 41020 18284 41076 18286
rect 41580 20802 41636 20804
rect 41580 20750 41582 20802
rect 41582 20750 41634 20802
rect 41634 20750 41636 20802
rect 41580 20748 41636 20750
rect 41468 20690 41524 20692
rect 41468 20638 41470 20690
rect 41470 20638 41522 20690
rect 41522 20638 41524 20690
rect 41468 20636 41524 20638
rect 41692 20018 41748 20020
rect 41692 19966 41694 20018
rect 41694 19966 41746 20018
rect 41746 19966 41748 20018
rect 41692 19964 41748 19966
rect 41580 19292 41636 19348
rect 43932 26124 43988 26180
rect 42924 25900 42980 25956
rect 42588 23154 42644 23156
rect 42588 23102 42590 23154
rect 42590 23102 42642 23154
rect 42642 23102 42644 23154
rect 42588 23100 42644 23102
rect 42812 23660 42868 23716
rect 43372 24892 43428 24948
rect 43036 24498 43092 24500
rect 43036 24446 43038 24498
rect 43038 24446 43090 24498
rect 43090 24446 43092 24498
rect 43036 24444 43092 24446
rect 43596 25228 43652 25284
rect 44492 27244 44548 27300
rect 43708 24556 43764 24612
rect 43596 24444 43652 24500
rect 43036 23324 43092 23380
rect 42924 23212 42980 23268
rect 43372 23548 43428 23604
rect 43148 23100 43204 23156
rect 43260 23436 43316 23492
rect 42812 22428 42868 22484
rect 42588 21868 42644 21924
rect 42252 21698 42308 21700
rect 42252 21646 42254 21698
rect 42254 21646 42306 21698
rect 42306 21646 42308 21698
rect 42252 21644 42308 21646
rect 42364 20690 42420 20692
rect 42364 20638 42366 20690
rect 42366 20638 42418 20690
rect 42418 20638 42420 20690
rect 42364 20636 42420 20638
rect 42476 20242 42532 20244
rect 42476 20190 42478 20242
rect 42478 20190 42530 20242
rect 42530 20190 42532 20242
rect 42476 20188 42532 20190
rect 41804 19068 41860 19124
rect 42588 19740 42644 19796
rect 42924 20802 42980 20804
rect 42924 20750 42926 20802
rect 42926 20750 42978 20802
rect 42978 20750 42980 20802
rect 42924 20748 42980 20750
rect 42252 18956 42308 19012
rect 42700 19346 42756 19348
rect 42700 19294 42702 19346
rect 42702 19294 42754 19346
rect 42754 19294 42756 19346
rect 42700 19292 42756 19294
rect 42588 19234 42644 19236
rect 42588 19182 42590 19234
rect 42590 19182 42642 19234
rect 42642 19182 42644 19234
rect 42588 19180 42644 19182
rect 43484 22876 43540 22932
rect 44156 24780 44212 24836
rect 43932 23826 43988 23828
rect 43932 23774 43934 23826
rect 43934 23774 43986 23826
rect 43986 23774 43988 23826
rect 43932 23772 43988 23774
rect 44044 23660 44100 23716
rect 44156 23548 44212 23604
rect 44380 25116 44436 25172
rect 43596 21868 43652 21924
rect 43596 20300 43652 20356
rect 43372 20076 43428 20132
rect 43932 22930 43988 22932
rect 43932 22878 43934 22930
rect 43934 22878 43986 22930
rect 43986 22878 43988 22930
rect 43932 22876 43988 22878
rect 44044 20914 44100 20916
rect 44044 20862 44046 20914
rect 44046 20862 44098 20914
rect 44098 20862 44100 20914
rect 44044 20860 44100 20862
rect 43708 19628 43764 19684
rect 42924 19122 42980 19124
rect 42924 19070 42926 19122
rect 42926 19070 42978 19122
rect 42978 19070 42980 19122
rect 42924 19068 42980 19070
rect 42812 18844 42868 18900
rect 42588 18620 42644 18676
rect 39676 17164 39732 17220
rect 39452 16940 39508 16996
rect 39340 16828 39396 16884
rect 39228 15986 39284 15988
rect 39228 15934 39230 15986
rect 39230 15934 39282 15986
rect 39282 15934 39284 15986
rect 39228 15932 39284 15934
rect 38668 14530 38724 14532
rect 38668 14478 38670 14530
rect 38670 14478 38722 14530
rect 38722 14478 38724 14530
rect 38668 14476 38724 14478
rect 38780 14418 38836 14420
rect 38780 14366 38782 14418
rect 38782 14366 38834 14418
rect 38834 14366 38836 14418
rect 38780 14364 38836 14366
rect 39788 15372 39844 15428
rect 39004 14252 39060 14308
rect 38780 13970 38836 13972
rect 38780 13918 38782 13970
rect 38782 13918 38834 13970
rect 38834 13918 38836 13970
rect 38780 13916 38836 13918
rect 39564 14924 39620 14980
rect 39004 13746 39060 13748
rect 39004 13694 39006 13746
rect 39006 13694 39058 13746
rect 39058 13694 39060 13746
rect 39004 13692 39060 13694
rect 40124 17106 40180 17108
rect 40124 17054 40126 17106
rect 40126 17054 40178 17106
rect 40178 17054 40180 17106
rect 40124 17052 40180 17054
rect 40796 17388 40852 17444
rect 40348 16828 40404 16884
rect 40236 16044 40292 16100
rect 40012 15314 40068 15316
rect 40012 15262 40014 15314
rect 40014 15262 40066 15314
rect 40066 15262 40068 15314
rect 40012 15260 40068 15262
rect 42140 18450 42196 18452
rect 42140 18398 42142 18450
rect 42142 18398 42194 18450
rect 42194 18398 42196 18450
rect 42140 18396 42196 18398
rect 40908 16604 40964 16660
rect 40684 15820 40740 15876
rect 40460 15260 40516 15316
rect 39900 14924 39956 14980
rect 40236 14812 40292 14868
rect 39900 14252 39956 14308
rect 38892 13634 38948 13636
rect 38892 13582 38894 13634
rect 38894 13582 38946 13634
rect 38946 13582 38948 13634
rect 38892 13580 38948 13582
rect 38668 13468 38724 13524
rect 40908 15932 40964 15988
rect 41020 15820 41076 15876
rect 41580 17948 41636 18004
rect 41356 17106 41412 17108
rect 41356 17054 41358 17106
rect 41358 17054 41410 17106
rect 41410 17054 41412 17106
rect 41356 17052 41412 17054
rect 41804 17724 41860 17780
rect 41580 17052 41636 17108
rect 41692 16940 41748 16996
rect 41580 15372 41636 15428
rect 42924 18508 42980 18564
rect 43148 18956 43204 19012
rect 42028 16882 42084 16884
rect 42028 16830 42030 16882
rect 42030 16830 42082 16882
rect 42082 16830 42084 16882
rect 42028 16828 42084 16830
rect 41804 16044 41860 16100
rect 41916 15932 41972 15988
rect 42028 16604 42084 16660
rect 40796 13804 40852 13860
rect 38892 12178 38948 12180
rect 38892 12126 38894 12178
rect 38894 12126 38946 12178
rect 38946 12126 38948 12178
rect 38892 12124 38948 12126
rect 40236 12402 40292 12404
rect 40236 12350 40238 12402
rect 40238 12350 40290 12402
rect 40290 12350 40292 12402
rect 40236 12348 40292 12350
rect 39564 12178 39620 12180
rect 39564 12126 39566 12178
rect 39566 12126 39618 12178
rect 39618 12126 39620 12178
rect 39564 12124 39620 12126
rect 38556 11676 38612 11732
rect 39340 11676 39396 11732
rect 38332 11228 38388 11284
rect 37884 3388 37940 3444
rect 38108 9436 38164 9492
rect 38332 9212 38388 9268
rect 38780 11228 38836 11284
rect 38556 10108 38612 10164
rect 38780 10108 38836 10164
rect 38892 9548 38948 9604
rect 38444 9100 38500 9156
rect 38220 4956 38276 5012
rect 40348 11564 40404 11620
rect 39900 11452 39956 11508
rect 39676 11282 39732 11284
rect 39676 11230 39678 11282
rect 39678 11230 39730 11282
rect 39730 11230 39732 11282
rect 39676 11228 39732 11230
rect 40012 11004 40068 11060
rect 39228 9266 39284 9268
rect 39228 9214 39230 9266
rect 39230 9214 39282 9266
rect 39282 9214 39284 9266
rect 39228 9212 39284 9214
rect 39676 9154 39732 9156
rect 39676 9102 39678 9154
rect 39678 9102 39730 9154
rect 39730 9102 39732 9154
rect 39676 9100 39732 9102
rect 40572 12124 40628 12180
rect 40908 11282 40964 11284
rect 40908 11230 40910 11282
rect 40910 11230 40962 11282
rect 40962 11230 40964 11282
rect 40908 11228 40964 11230
rect 40796 11116 40852 11172
rect 40908 9548 40964 9604
rect 40236 8988 40292 9044
rect 40348 8316 40404 8372
rect 41692 15036 41748 15092
rect 41916 15260 41972 15316
rect 41580 14812 41636 14868
rect 41468 13916 41524 13972
rect 41132 13804 41188 13860
rect 42364 15036 42420 15092
rect 42476 13916 42532 13972
rect 41244 12124 41300 12180
rect 41468 11618 41524 11620
rect 41468 11566 41470 11618
rect 41470 11566 41522 11618
rect 41522 11566 41524 11618
rect 41468 11564 41524 11566
rect 42140 11116 42196 11172
rect 42812 17388 42868 17444
rect 42812 16604 42868 16660
rect 42700 15148 42756 15204
rect 43036 17778 43092 17780
rect 43036 17726 43038 17778
rect 43038 17726 43090 17778
rect 43090 17726 43092 17778
rect 43036 17724 43092 17726
rect 43372 18844 43428 18900
rect 43596 18508 43652 18564
rect 43372 18396 43428 18452
rect 46284 35922 46340 35924
rect 46284 35870 46286 35922
rect 46286 35870 46338 35922
rect 46338 35870 46340 35922
rect 46284 35868 46340 35870
rect 46508 37100 46564 37156
rect 46844 37100 46900 37156
rect 47852 42754 47908 42756
rect 47852 42702 47854 42754
rect 47854 42702 47906 42754
rect 47906 42702 47908 42754
rect 47852 42700 47908 42702
rect 48188 42754 48244 42756
rect 48188 42702 48190 42754
rect 48190 42702 48242 42754
rect 48242 42702 48244 42754
rect 48188 42700 48244 42702
rect 48748 43148 48804 43204
rect 47740 40290 47796 40292
rect 47740 40238 47742 40290
rect 47742 40238 47794 40290
rect 47794 40238 47796 40290
rect 47740 40236 47796 40238
rect 47628 39394 47684 39396
rect 47628 39342 47630 39394
rect 47630 39342 47682 39394
rect 47682 39342 47684 39394
rect 47628 39340 47684 39342
rect 46172 35532 46228 35588
rect 46396 35420 46452 35476
rect 46844 34636 46900 34692
rect 46284 33404 46340 33460
rect 46732 34242 46788 34244
rect 46732 34190 46734 34242
rect 46734 34190 46786 34242
rect 46786 34190 46788 34242
rect 46732 34188 46788 34190
rect 44940 33068 44996 33124
rect 46284 33122 46340 33124
rect 46284 33070 46286 33122
rect 46286 33070 46338 33122
rect 46338 33070 46340 33122
rect 46284 33068 46340 33070
rect 45164 31612 45220 31668
rect 45164 30994 45220 30996
rect 45164 30942 45166 30994
rect 45166 30942 45218 30994
rect 45218 30942 45220 30994
rect 45164 30940 45220 30942
rect 45052 30268 45108 30324
rect 45164 30716 45220 30772
rect 44940 30210 44996 30212
rect 44940 30158 44942 30210
rect 44942 30158 44994 30210
rect 44994 30158 44996 30210
rect 44940 30156 44996 30158
rect 46508 31612 46564 31668
rect 47628 37826 47684 37828
rect 47628 37774 47630 37826
rect 47630 37774 47682 37826
rect 47682 37774 47684 37826
rect 47628 37772 47684 37774
rect 47740 37436 47796 37492
rect 48524 40460 48580 40516
rect 48636 40348 48692 40404
rect 48860 40460 48916 40516
rect 48412 37826 48468 37828
rect 48412 37774 48414 37826
rect 48414 37774 48466 37826
rect 48466 37774 48468 37826
rect 48412 37772 48468 37774
rect 48076 37436 48132 37492
rect 47964 37154 48020 37156
rect 47964 37102 47966 37154
rect 47966 37102 48018 37154
rect 48018 37102 48020 37154
rect 47964 37100 48020 37102
rect 47964 36204 48020 36260
rect 48524 37212 48580 37268
rect 49532 42530 49588 42532
rect 49532 42478 49534 42530
rect 49534 42478 49586 42530
rect 49586 42478 49588 42530
rect 49532 42476 49588 42478
rect 49308 42082 49364 42084
rect 49308 42030 49310 42082
rect 49310 42030 49362 42082
rect 49362 42030 49364 42082
rect 49308 42028 49364 42030
rect 49084 41970 49140 41972
rect 49084 41918 49086 41970
rect 49086 41918 49138 41970
rect 49138 41918 49140 41970
rect 49084 41916 49140 41918
rect 49196 41186 49252 41188
rect 49196 41134 49198 41186
rect 49198 41134 49250 41186
rect 49250 41134 49252 41186
rect 49196 41132 49252 41134
rect 49196 40908 49252 40964
rect 49084 39058 49140 39060
rect 49084 39006 49086 39058
rect 49086 39006 49138 39058
rect 49138 39006 49140 39058
rect 49084 39004 49140 39006
rect 49532 41356 49588 41412
rect 50316 53618 50372 53620
rect 50316 53566 50318 53618
rect 50318 53566 50370 53618
rect 50370 53566 50372 53618
rect 50316 53564 50372 53566
rect 50876 53618 50932 53620
rect 50876 53566 50878 53618
rect 50878 53566 50930 53618
rect 50930 53566 50932 53618
rect 50876 53564 50932 53566
rect 50204 53228 50260 53284
rect 50556 53338 50612 53340
rect 50556 53286 50558 53338
rect 50558 53286 50610 53338
rect 50610 53286 50612 53338
rect 50556 53284 50612 53286
rect 50660 53338 50716 53340
rect 50660 53286 50662 53338
rect 50662 53286 50714 53338
rect 50714 53286 50716 53338
rect 50660 53284 50716 53286
rect 50764 53338 50820 53340
rect 50764 53286 50766 53338
rect 50766 53286 50818 53338
rect 50818 53286 50820 53338
rect 50764 53284 50820 53286
rect 50092 52668 50148 52724
rect 50556 51770 50612 51772
rect 50556 51718 50558 51770
rect 50558 51718 50610 51770
rect 50610 51718 50612 51770
rect 50556 51716 50612 51718
rect 50660 51770 50716 51772
rect 50660 51718 50662 51770
rect 50662 51718 50714 51770
rect 50714 51718 50716 51770
rect 50660 51716 50716 51718
rect 50764 51770 50820 51772
rect 50764 51718 50766 51770
rect 50766 51718 50818 51770
rect 50818 51718 50820 51770
rect 50764 51716 50820 51718
rect 49980 50316 50036 50372
rect 51660 50316 51716 50372
rect 50556 50202 50612 50204
rect 50556 50150 50558 50202
rect 50558 50150 50610 50202
rect 50610 50150 50612 50202
rect 50556 50148 50612 50150
rect 50660 50202 50716 50204
rect 50660 50150 50662 50202
rect 50662 50150 50714 50202
rect 50714 50150 50716 50202
rect 50660 50148 50716 50150
rect 50764 50202 50820 50204
rect 50764 50150 50766 50202
rect 50766 50150 50818 50202
rect 50818 50150 50820 50202
rect 50764 50148 50820 50150
rect 50316 48802 50372 48804
rect 50316 48750 50318 48802
rect 50318 48750 50370 48802
rect 50370 48750 50372 48802
rect 50316 48748 50372 48750
rect 50556 48634 50612 48636
rect 50556 48582 50558 48634
rect 50558 48582 50610 48634
rect 50610 48582 50612 48634
rect 50556 48580 50612 48582
rect 50660 48634 50716 48636
rect 50660 48582 50662 48634
rect 50662 48582 50714 48634
rect 50714 48582 50716 48634
rect 50660 48580 50716 48582
rect 50764 48634 50820 48636
rect 50764 48582 50766 48634
rect 50766 48582 50818 48634
rect 50818 48582 50820 48634
rect 50764 48580 50820 48582
rect 50556 47066 50612 47068
rect 50556 47014 50558 47066
rect 50558 47014 50610 47066
rect 50610 47014 50612 47066
rect 50556 47012 50612 47014
rect 50660 47066 50716 47068
rect 50660 47014 50662 47066
rect 50662 47014 50714 47066
rect 50714 47014 50716 47066
rect 50660 47012 50716 47014
rect 50764 47066 50820 47068
rect 50764 47014 50766 47066
rect 50766 47014 50818 47066
rect 50818 47014 50820 47066
rect 50764 47012 50820 47014
rect 51100 45836 51156 45892
rect 50556 45498 50612 45500
rect 50556 45446 50558 45498
rect 50558 45446 50610 45498
rect 50610 45446 50612 45498
rect 50556 45444 50612 45446
rect 50660 45498 50716 45500
rect 50660 45446 50662 45498
rect 50662 45446 50714 45498
rect 50714 45446 50716 45498
rect 50660 45444 50716 45446
rect 50764 45498 50820 45500
rect 50764 45446 50766 45498
rect 50766 45446 50818 45498
rect 50818 45446 50820 45498
rect 50764 45444 50820 45446
rect 50556 43930 50612 43932
rect 50556 43878 50558 43930
rect 50558 43878 50610 43930
rect 50610 43878 50612 43930
rect 50556 43876 50612 43878
rect 50660 43930 50716 43932
rect 50660 43878 50662 43930
rect 50662 43878 50714 43930
rect 50714 43878 50716 43930
rect 50660 43876 50716 43878
rect 50764 43930 50820 43932
rect 50764 43878 50766 43930
rect 50766 43878 50818 43930
rect 50818 43878 50820 43930
rect 50764 43876 50820 43878
rect 50652 43708 50708 43764
rect 49868 42812 49924 42868
rect 50204 42866 50260 42868
rect 50204 42814 50206 42866
rect 50206 42814 50258 42866
rect 50258 42814 50260 42866
rect 50204 42812 50260 42814
rect 50540 42530 50596 42532
rect 50540 42478 50542 42530
rect 50542 42478 50594 42530
rect 50594 42478 50596 42530
rect 50540 42476 50596 42478
rect 50556 42362 50612 42364
rect 50556 42310 50558 42362
rect 50558 42310 50610 42362
rect 50610 42310 50612 42362
rect 50556 42308 50612 42310
rect 50660 42362 50716 42364
rect 50660 42310 50662 42362
rect 50662 42310 50714 42362
rect 50714 42310 50716 42362
rect 50660 42308 50716 42310
rect 50764 42362 50820 42364
rect 50764 42310 50766 42362
rect 50766 42310 50818 42362
rect 50818 42310 50820 42362
rect 50764 42308 50820 42310
rect 50316 42028 50372 42084
rect 49756 39004 49812 39060
rect 49308 37490 49364 37492
rect 49308 37438 49310 37490
rect 49310 37438 49362 37490
rect 49362 37438 49364 37490
rect 49308 37436 49364 37438
rect 48076 35922 48132 35924
rect 48076 35870 48078 35922
rect 48078 35870 48130 35922
rect 48130 35870 48132 35922
rect 48076 35868 48132 35870
rect 48188 35980 48244 36036
rect 47740 34860 47796 34916
rect 47516 34636 47572 34692
rect 47628 34354 47684 34356
rect 47628 34302 47630 34354
rect 47630 34302 47682 34354
rect 47682 34302 47684 34354
rect 47628 34300 47684 34302
rect 48748 35420 48804 35476
rect 49196 36652 49252 36708
rect 49308 37212 49364 37268
rect 49084 35868 49140 35924
rect 49420 35868 49476 35924
rect 48188 34636 48244 34692
rect 47964 34188 48020 34244
rect 48188 34300 48244 34356
rect 47068 33628 47124 33684
rect 48188 34018 48244 34020
rect 48188 33966 48190 34018
rect 48190 33966 48242 34018
rect 48242 33966 48244 34018
rect 48188 33964 48244 33966
rect 48188 33740 48244 33796
rect 48860 34860 48916 34916
rect 48636 33740 48692 33796
rect 48748 33628 48804 33684
rect 49532 34242 49588 34244
rect 49532 34190 49534 34242
rect 49534 34190 49586 34242
rect 49586 34190 49588 34242
rect 49532 34188 49588 34190
rect 49532 33404 49588 33460
rect 47964 33346 48020 33348
rect 47964 33294 47966 33346
rect 47966 33294 48018 33346
rect 48018 33294 48020 33346
rect 47964 33292 48020 33294
rect 48748 33346 48804 33348
rect 48748 33294 48750 33346
rect 48750 33294 48802 33346
rect 48802 33294 48804 33346
rect 48748 33292 48804 33294
rect 50988 41410 51044 41412
rect 50988 41358 50990 41410
rect 50990 41358 51042 41410
rect 51042 41358 51044 41410
rect 50988 41356 51044 41358
rect 51660 44268 51716 44324
rect 51660 43708 51716 43764
rect 52332 58940 52388 58996
rect 52220 56924 52276 56980
rect 52332 48300 52388 48356
rect 52220 44492 52276 44548
rect 52108 43260 52164 43316
rect 51660 42028 51716 42084
rect 50556 40794 50612 40796
rect 50556 40742 50558 40794
rect 50558 40742 50610 40794
rect 50610 40742 50612 40794
rect 50556 40740 50612 40742
rect 50660 40794 50716 40796
rect 50660 40742 50662 40794
rect 50662 40742 50714 40794
rect 50714 40742 50716 40794
rect 50660 40740 50716 40742
rect 50764 40794 50820 40796
rect 50764 40742 50766 40794
rect 50766 40742 50818 40794
rect 50818 40742 50820 40794
rect 50764 40740 50820 40742
rect 55356 46450 55412 46452
rect 55356 46398 55358 46450
rect 55358 46398 55410 46450
rect 55410 46398 55412 46450
rect 55356 46396 55412 46398
rect 55020 45724 55076 45780
rect 53228 42924 53284 42980
rect 52668 42028 52724 42084
rect 53788 42700 53844 42756
rect 52108 41916 52164 41972
rect 51436 40962 51492 40964
rect 51436 40910 51438 40962
rect 51438 40910 51490 40962
rect 51490 40910 51492 40962
rect 51436 40908 51492 40910
rect 53228 41468 53284 41524
rect 52108 40236 52164 40292
rect 50556 39226 50612 39228
rect 50556 39174 50558 39226
rect 50558 39174 50610 39226
rect 50610 39174 50612 39226
rect 50556 39172 50612 39174
rect 50660 39226 50716 39228
rect 50660 39174 50662 39226
rect 50662 39174 50714 39226
rect 50714 39174 50716 39226
rect 50660 39172 50716 39174
rect 50764 39226 50820 39228
rect 50764 39174 50766 39226
rect 50766 39174 50818 39226
rect 50818 39174 50820 39226
rect 50764 39172 50820 39174
rect 53452 40402 53508 40404
rect 53452 40350 53454 40402
rect 53454 40350 53506 40402
rect 53506 40350 53508 40402
rect 53452 40348 53508 40350
rect 55580 45890 55636 45892
rect 55580 45838 55582 45890
rect 55582 45838 55634 45890
rect 55634 45838 55636 45890
rect 55580 45836 55636 45838
rect 57932 45052 57988 45108
rect 57820 44380 57876 44436
rect 55580 44322 55636 44324
rect 55580 44270 55582 44322
rect 55582 44270 55634 44322
rect 55634 44270 55636 44322
rect 55580 44268 55636 44270
rect 57932 43708 57988 43764
rect 57932 43036 57988 43092
rect 55580 42754 55636 42756
rect 55580 42702 55582 42754
rect 55582 42702 55634 42754
rect 55634 42702 55636 42754
rect 55580 42700 55636 42702
rect 55468 41916 55524 41972
rect 57932 42364 57988 42420
rect 55356 41746 55412 41748
rect 55356 41694 55358 41746
rect 55358 41694 55410 41746
rect 55410 41694 55412 41746
rect 55356 41692 55412 41694
rect 55020 40348 55076 40404
rect 53788 40124 53844 40180
rect 55356 39676 55412 39732
rect 55468 39788 55524 39844
rect 57932 41020 57988 41076
rect 55580 39618 55636 39620
rect 55580 39566 55582 39618
rect 55582 39566 55634 39618
rect 55634 39566 55636 39618
rect 55580 39564 55636 39566
rect 52668 38892 52724 38948
rect 57932 39004 57988 39060
rect 55356 38610 55412 38612
rect 55356 38558 55358 38610
rect 55358 38558 55410 38610
rect 55410 38558 55412 38610
rect 55356 38556 55412 38558
rect 53228 38108 53284 38164
rect 55356 38050 55412 38052
rect 55356 37998 55358 38050
rect 55358 37998 55410 38050
rect 55410 37998 55412 38050
rect 55356 37996 55412 37998
rect 50556 37658 50612 37660
rect 50556 37606 50558 37658
rect 50558 37606 50610 37658
rect 50610 37606 50612 37658
rect 50556 37604 50612 37606
rect 50660 37658 50716 37660
rect 50660 37606 50662 37658
rect 50662 37606 50714 37658
rect 50714 37606 50716 37658
rect 50660 37604 50716 37606
rect 50764 37658 50820 37660
rect 50764 37606 50766 37658
rect 50766 37606 50818 37658
rect 50818 37606 50820 37658
rect 50764 37604 50820 37606
rect 57932 37660 57988 37716
rect 53452 37266 53508 37268
rect 53452 37214 53454 37266
rect 53454 37214 53506 37266
rect 53506 37214 53508 37266
rect 53452 37212 53508 37214
rect 52668 37100 52724 37156
rect 49868 35644 49924 35700
rect 50428 36706 50484 36708
rect 50428 36654 50430 36706
rect 50430 36654 50482 36706
rect 50482 36654 50484 36706
rect 50428 36652 50484 36654
rect 52108 36428 52164 36484
rect 50876 36258 50932 36260
rect 50876 36206 50878 36258
rect 50878 36206 50930 36258
rect 50930 36206 50932 36258
rect 50876 36204 50932 36206
rect 50556 36090 50612 36092
rect 50556 36038 50558 36090
rect 50558 36038 50610 36090
rect 50610 36038 50612 36090
rect 50556 36036 50612 36038
rect 50660 36090 50716 36092
rect 50660 36038 50662 36090
rect 50662 36038 50714 36090
rect 50714 36038 50716 36090
rect 50660 36036 50716 36038
rect 50764 36090 50820 36092
rect 50764 36038 50766 36090
rect 50766 36038 50818 36090
rect 50818 36038 50820 36090
rect 50764 36036 50820 36038
rect 50540 35532 50596 35588
rect 49868 35308 49924 35364
rect 50556 34522 50612 34524
rect 50556 34470 50558 34522
rect 50558 34470 50610 34522
rect 50610 34470 50612 34522
rect 50556 34468 50612 34470
rect 50660 34522 50716 34524
rect 50660 34470 50662 34522
rect 50662 34470 50714 34522
rect 50714 34470 50716 34522
rect 50660 34468 50716 34470
rect 50764 34522 50820 34524
rect 50764 34470 50766 34522
rect 50766 34470 50818 34522
rect 50818 34470 50820 34522
rect 50764 34468 50820 34470
rect 52108 35756 52164 35812
rect 51660 35586 51716 35588
rect 51660 35534 51662 35586
rect 51662 35534 51714 35586
rect 51714 35534 51716 35586
rect 51660 35532 51716 35534
rect 50988 33964 51044 34020
rect 51660 34018 51716 34020
rect 51660 33966 51662 34018
rect 51662 33966 51714 34018
rect 51714 33966 51716 34018
rect 51660 33964 51716 33966
rect 50092 33404 50148 33460
rect 50652 33404 50708 33460
rect 46284 31164 46340 31220
rect 45836 30828 45892 30884
rect 46508 30882 46564 30884
rect 46508 30830 46510 30882
rect 46510 30830 46562 30882
rect 46562 30830 46564 30882
rect 46508 30828 46564 30830
rect 45612 30492 45668 30548
rect 45948 30492 46004 30548
rect 46620 30492 46676 30548
rect 45276 29986 45332 29988
rect 45276 29934 45278 29986
rect 45278 29934 45330 29986
rect 45330 29934 45332 29986
rect 45276 29932 45332 29934
rect 45164 28028 45220 28084
rect 45388 29596 45444 29652
rect 46060 30268 46116 30324
rect 45836 29148 45892 29204
rect 45948 29932 46004 29988
rect 46172 30044 46228 30100
rect 46172 29426 46228 29428
rect 46172 29374 46174 29426
rect 46174 29374 46226 29426
rect 46226 29374 46228 29426
rect 46172 29372 46228 29374
rect 46060 29148 46116 29204
rect 46508 29650 46564 29652
rect 46508 29598 46510 29650
rect 46510 29598 46562 29650
rect 46562 29598 46564 29650
rect 46508 29596 46564 29598
rect 46844 30210 46900 30212
rect 46844 30158 46846 30210
rect 46846 30158 46898 30210
rect 46898 30158 46900 30210
rect 46844 30156 46900 30158
rect 46732 30098 46788 30100
rect 46732 30046 46734 30098
rect 46734 30046 46786 30098
rect 46786 30046 46788 30098
rect 46732 30044 46788 30046
rect 46844 29820 46900 29876
rect 47180 30380 47236 30436
rect 48860 32396 48916 32452
rect 49196 32450 49252 32452
rect 49196 32398 49198 32450
rect 49198 32398 49250 32450
rect 49250 32398 49252 32450
rect 49196 32396 49252 32398
rect 49420 31836 49476 31892
rect 48076 31164 48132 31220
rect 48636 31164 48692 31220
rect 47628 31052 47684 31108
rect 47404 30994 47460 30996
rect 47404 30942 47406 30994
rect 47406 30942 47458 30994
rect 47458 30942 47460 30994
rect 47404 30940 47460 30942
rect 47628 30716 47684 30772
rect 47292 30044 47348 30100
rect 47740 29820 47796 29876
rect 47964 30156 48020 30212
rect 47852 30044 47908 30100
rect 47404 29538 47460 29540
rect 47404 29486 47406 29538
rect 47406 29486 47458 29538
rect 47458 29486 47460 29538
rect 47404 29484 47460 29486
rect 45724 28082 45780 28084
rect 45724 28030 45726 28082
rect 45726 28030 45778 28082
rect 45778 28030 45780 28082
rect 45724 28028 45780 28030
rect 45388 27916 45444 27972
rect 45052 27580 45108 27636
rect 44940 26850 44996 26852
rect 44940 26798 44942 26850
rect 44942 26798 44994 26850
rect 44994 26798 44996 26850
rect 44940 26796 44996 26798
rect 45612 26796 45668 26852
rect 44828 24780 44884 24836
rect 45276 26012 45332 26068
rect 46172 27132 46228 27188
rect 46060 27074 46116 27076
rect 46060 27022 46062 27074
rect 46062 27022 46114 27074
rect 46114 27022 46116 27074
rect 46060 27020 46116 27022
rect 45836 26796 45892 26852
rect 44940 25228 44996 25284
rect 44716 24610 44772 24612
rect 44716 24558 44718 24610
rect 44718 24558 44770 24610
rect 44770 24558 44772 24610
rect 44716 24556 44772 24558
rect 44604 23324 44660 23380
rect 44604 21868 44660 21924
rect 44492 20018 44548 20020
rect 44492 19966 44494 20018
rect 44494 19966 44546 20018
rect 44546 19966 44548 20018
rect 44492 19964 44548 19966
rect 44380 19852 44436 19908
rect 45836 25116 45892 25172
rect 44940 23436 44996 23492
rect 45836 23436 45892 23492
rect 45276 23212 45332 23268
rect 44940 23154 44996 23156
rect 44940 23102 44942 23154
rect 44942 23102 44994 23154
rect 44994 23102 44996 23154
rect 44940 23100 44996 23102
rect 44828 22370 44884 22372
rect 44828 22318 44830 22370
rect 44830 22318 44882 22370
rect 44882 22318 44884 22370
rect 44828 22316 44884 22318
rect 45052 21980 45108 22036
rect 45836 23100 45892 23156
rect 45276 22146 45332 22148
rect 45276 22094 45278 22146
rect 45278 22094 45330 22146
rect 45330 22094 45332 22146
rect 45276 22092 45332 22094
rect 45948 22092 46004 22148
rect 45948 20972 46004 21028
rect 44044 19068 44100 19124
rect 43932 19010 43988 19012
rect 43932 18958 43934 19010
rect 43934 18958 43986 19010
rect 43986 18958 43988 19010
rect 43932 18956 43988 18958
rect 43820 18620 43876 18676
rect 44716 19010 44772 19012
rect 44716 18958 44718 19010
rect 44718 18958 44770 19010
rect 44770 18958 44772 19010
rect 44716 18956 44772 18958
rect 44604 17948 44660 18004
rect 43932 17778 43988 17780
rect 43932 17726 43934 17778
rect 43934 17726 43986 17778
rect 43986 17726 43988 17778
rect 43932 17724 43988 17726
rect 43372 17500 43428 17556
rect 43708 16994 43764 16996
rect 43708 16942 43710 16994
rect 43710 16942 43762 16994
rect 43762 16942 43764 16994
rect 43708 16940 43764 16942
rect 43484 16044 43540 16100
rect 43036 14812 43092 14868
rect 44940 19122 44996 19124
rect 44940 19070 44942 19122
rect 44942 19070 44994 19122
rect 44994 19070 44996 19122
rect 44940 19068 44996 19070
rect 45388 20524 45444 20580
rect 45500 20300 45556 20356
rect 45500 19234 45556 19236
rect 45500 19182 45502 19234
rect 45502 19182 45554 19234
rect 45554 19182 45556 19234
rect 45500 19180 45556 19182
rect 45500 18508 45556 18564
rect 45276 18396 45332 18452
rect 45052 17276 45108 17332
rect 44940 17052 44996 17108
rect 44828 16828 44884 16884
rect 45388 17442 45444 17444
rect 45388 17390 45390 17442
rect 45390 17390 45442 17442
rect 45442 17390 45444 17442
rect 45388 17388 45444 17390
rect 45276 16940 45332 16996
rect 45164 16770 45220 16772
rect 45164 16718 45166 16770
rect 45166 16718 45218 16770
rect 45218 16718 45220 16770
rect 45164 16716 45220 16718
rect 45052 16098 45108 16100
rect 45052 16046 45054 16098
rect 45054 16046 45106 16098
rect 45106 16046 45108 16098
rect 45052 16044 45108 16046
rect 46508 29148 46564 29204
rect 46172 22988 46228 23044
rect 46172 22370 46228 22372
rect 46172 22318 46174 22370
rect 46174 22318 46226 22370
rect 46226 22318 46228 22370
rect 46172 22316 46228 22318
rect 46172 21532 46228 21588
rect 46508 26796 46564 26852
rect 46844 27692 46900 27748
rect 46732 27132 46788 27188
rect 46620 25900 46676 25956
rect 46844 25116 46900 25172
rect 48076 29596 48132 29652
rect 48412 30268 48468 30324
rect 48412 29596 48468 29652
rect 47964 29484 48020 29540
rect 47852 28754 47908 28756
rect 47852 28702 47854 28754
rect 47854 28702 47906 28754
rect 47906 28702 47908 28754
rect 47852 28700 47908 28702
rect 48076 27858 48132 27860
rect 48076 27806 48078 27858
rect 48078 27806 48130 27858
rect 48130 27806 48132 27858
rect 48076 27804 48132 27806
rect 47964 27746 48020 27748
rect 47964 27694 47966 27746
rect 47966 27694 48018 27746
rect 48018 27694 48020 27746
rect 47964 27692 48020 27694
rect 47404 27020 47460 27076
rect 47740 27132 47796 27188
rect 48524 27186 48580 27188
rect 48524 27134 48526 27186
rect 48526 27134 48578 27186
rect 48578 27134 48580 27186
rect 48524 27132 48580 27134
rect 48188 26962 48244 26964
rect 48188 26910 48190 26962
rect 48190 26910 48242 26962
rect 48242 26910 48244 26962
rect 48188 26908 48244 26910
rect 47068 26236 47124 26292
rect 47740 26236 47796 26292
rect 48076 26514 48132 26516
rect 48076 26462 48078 26514
rect 48078 26462 48130 26514
rect 48130 26462 48132 26514
rect 48076 26460 48132 26462
rect 48412 26348 48468 26404
rect 48076 26236 48132 26292
rect 46956 25004 47012 25060
rect 47292 23884 47348 23940
rect 46844 23772 46900 23828
rect 46396 23324 46452 23380
rect 48076 25900 48132 25956
rect 48188 24834 48244 24836
rect 48188 24782 48190 24834
rect 48190 24782 48242 24834
rect 48242 24782 48244 24834
rect 48188 24780 48244 24782
rect 47852 23772 47908 23828
rect 47068 23548 47124 23604
rect 47852 23266 47908 23268
rect 47852 23214 47854 23266
rect 47854 23214 47906 23266
rect 47906 23214 47908 23266
rect 47852 23212 47908 23214
rect 47292 23154 47348 23156
rect 47292 23102 47294 23154
rect 47294 23102 47346 23154
rect 47346 23102 47348 23154
rect 47292 23100 47348 23102
rect 46508 22092 46564 22148
rect 46620 21980 46676 22036
rect 46844 21586 46900 21588
rect 46844 21534 46846 21586
rect 46846 21534 46898 21586
rect 46898 21534 46900 21586
rect 46844 21532 46900 21534
rect 46284 20972 46340 21028
rect 46284 19964 46340 20020
rect 46060 19906 46116 19908
rect 46060 19854 46062 19906
rect 46062 19854 46114 19906
rect 46114 19854 46116 19906
rect 46060 19852 46116 19854
rect 45724 18172 45780 18228
rect 45724 17554 45780 17556
rect 45724 17502 45726 17554
rect 45726 17502 45778 17554
rect 45778 17502 45780 17554
rect 45724 17500 45780 17502
rect 46844 20578 46900 20580
rect 46844 20526 46846 20578
rect 46846 20526 46898 20578
rect 46898 20526 46900 20578
rect 46844 20524 46900 20526
rect 46508 20188 46564 20244
rect 46396 18956 46452 19012
rect 47516 22316 47572 22372
rect 47292 21532 47348 21588
rect 47180 20524 47236 20580
rect 47852 20802 47908 20804
rect 47852 20750 47854 20802
rect 47854 20750 47906 20802
rect 47906 20750 47908 20802
rect 47852 20748 47908 20750
rect 47292 19852 47348 19908
rect 47628 19628 47684 19684
rect 47740 19292 47796 19348
rect 46284 18284 46340 18340
rect 46844 18562 46900 18564
rect 46844 18510 46846 18562
rect 46846 18510 46898 18562
rect 46898 18510 46900 18562
rect 46844 18508 46900 18510
rect 47068 18620 47124 18676
rect 47516 18284 47572 18340
rect 46620 17836 46676 17892
rect 46956 17948 47012 18004
rect 46396 17778 46452 17780
rect 46396 17726 46398 17778
rect 46398 17726 46450 17778
rect 46450 17726 46452 17778
rect 46396 17724 46452 17726
rect 45612 16716 45668 16772
rect 45612 16044 45668 16100
rect 43932 15372 43988 15428
rect 43036 14642 43092 14644
rect 43036 14590 43038 14642
rect 43038 14590 43090 14642
rect 43090 14590 43092 14642
rect 43036 14588 43092 14590
rect 43036 13970 43092 13972
rect 43036 13918 43038 13970
rect 43038 13918 43090 13970
rect 43090 13918 43092 13970
rect 43036 13916 43092 13918
rect 42588 12402 42644 12404
rect 42588 12350 42590 12402
rect 42590 12350 42642 12402
rect 42642 12350 42644 12402
rect 42588 12348 42644 12350
rect 42812 12012 42868 12068
rect 42588 11394 42644 11396
rect 42588 11342 42590 11394
rect 42590 11342 42642 11394
rect 42642 11342 42644 11394
rect 42588 11340 42644 11342
rect 41580 10444 41636 10500
rect 41916 10556 41972 10612
rect 42364 10220 42420 10276
rect 41916 9212 41972 9268
rect 41356 8988 41412 9044
rect 42364 9042 42420 9044
rect 42364 8990 42366 9042
rect 42366 8990 42418 9042
rect 42418 8990 42420 9042
rect 42364 8988 42420 8990
rect 42812 10220 42868 10276
rect 43484 14306 43540 14308
rect 43484 14254 43486 14306
rect 43486 14254 43538 14306
rect 43538 14254 43540 14306
rect 43484 14252 43540 14254
rect 43484 13970 43540 13972
rect 43484 13918 43486 13970
rect 43486 13918 43538 13970
rect 43538 13918 43540 13970
rect 43484 13916 43540 13918
rect 44940 15372 44996 15428
rect 45164 15148 45220 15204
rect 46060 17052 46116 17108
rect 46284 17388 46340 17444
rect 46396 17164 46452 17220
rect 46732 17276 46788 17332
rect 46620 16882 46676 16884
rect 46620 16830 46622 16882
rect 46622 16830 46674 16882
rect 46674 16830 46676 16882
rect 46620 16828 46676 16830
rect 44828 14588 44884 14644
rect 46060 15820 46116 15876
rect 45500 14642 45556 14644
rect 45500 14590 45502 14642
rect 45502 14590 45554 14642
rect 45554 14590 45556 14642
rect 45500 14588 45556 14590
rect 43260 12066 43316 12068
rect 43260 12014 43262 12066
rect 43262 12014 43314 12066
rect 43314 12014 43316 12066
rect 43260 12012 43316 12014
rect 43036 10220 43092 10276
rect 43596 10108 43652 10164
rect 41468 8204 41524 8260
rect 42364 8258 42420 8260
rect 42364 8206 42366 8258
rect 42366 8206 42418 8258
rect 42418 8206 42420 8258
rect 42364 8204 42420 8206
rect 43372 8092 43428 8148
rect 43596 8204 43652 8260
rect 42140 7196 42196 7252
rect 42588 6130 42644 6132
rect 42588 6078 42590 6130
rect 42590 6078 42642 6130
rect 42642 6078 42644 6130
rect 42588 6076 42644 6078
rect 45612 13746 45668 13748
rect 45612 13694 45614 13746
rect 45614 13694 45666 13746
rect 45666 13694 45668 13746
rect 45612 13692 45668 13694
rect 46732 16156 46788 16212
rect 46620 16098 46676 16100
rect 46620 16046 46622 16098
rect 46622 16046 46674 16098
rect 46674 16046 46676 16098
rect 46620 16044 46676 16046
rect 46508 15202 46564 15204
rect 46508 15150 46510 15202
rect 46510 15150 46562 15202
rect 46562 15150 46564 15202
rect 46508 15148 46564 15150
rect 44604 13020 44660 13076
rect 43932 12796 43988 12852
rect 45500 13074 45556 13076
rect 45500 13022 45502 13074
rect 45502 13022 45554 13074
rect 45554 13022 45556 13074
rect 45500 13020 45556 13022
rect 44380 12012 44436 12068
rect 44156 11564 44212 11620
rect 44380 11340 44436 11396
rect 44156 10108 44212 10164
rect 44828 11394 44884 11396
rect 44828 11342 44830 11394
rect 44830 11342 44882 11394
rect 44882 11342 44884 11394
rect 44828 11340 44884 11342
rect 45724 12348 45780 12404
rect 45276 11564 45332 11620
rect 43148 7250 43204 7252
rect 43148 7198 43150 7250
rect 43150 7198 43202 7250
rect 43202 7198 43204 7250
rect 43148 7196 43204 7198
rect 43036 3388 43092 3444
rect 43372 3388 43428 3444
rect 43708 7644 43764 7700
rect 44828 10498 44884 10500
rect 44828 10446 44830 10498
rect 44830 10446 44882 10498
rect 44882 10446 44884 10498
rect 44828 10444 44884 10446
rect 44828 8988 44884 9044
rect 45500 11282 45556 11284
rect 45500 11230 45502 11282
rect 45502 11230 45554 11282
rect 45554 11230 45556 11282
rect 45500 11228 45556 11230
rect 45388 11170 45444 11172
rect 45388 11118 45390 11170
rect 45390 11118 45442 11170
rect 45442 11118 45444 11170
rect 45388 11116 45444 11118
rect 45948 12348 46004 12404
rect 48076 19292 48132 19348
rect 48412 21196 48468 21252
rect 48524 26124 48580 26180
rect 47628 17836 47684 17892
rect 47404 17554 47460 17556
rect 47404 17502 47406 17554
rect 47406 17502 47458 17554
rect 47458 17502 47460 17554
rect 47404 17500 47460 17502
rect 47740 17612 47796 17668
rect 47628 17442 47684 17444
rect 47628 17390 47630 17442
rect 47630 17390 47682 17442
rect 47682 17390 47684 17442
rect 47628 17388 47684 17390
rect 48076 18620 48132 18676
rect 48300 18284 48356 18340
rect 48412 17836 48468 17892
rect 48188 17666 48244 17668
rect 48188 17614 48190 17666
rect 48190 17614 48242 17666
rect 48242 17614 48244 17666
rect 48188 17612 48244 17614
rect 47292 16210 47348 16212
rect 47292 16158 47294 16210
rect 47294 16158 47346 16210
rect 47346 16158 47348 16210
rect 47292 16156 47348 16158
rect 47740 16156 47796 16212
rect 47628 15708 47684 15764
rect 47404 15372 47460 15428
rect 47852 15484 47908 15540
rect 48076 17500 48132 17556
rect 48300 17052 48356 17108
rect 48412 16604 48468 16660
rect 48412 16098 48468 16100
rect 48412 16046 48414 16098
rect 48414 16046 48466 16098
rect 48466 16046 48468 16098
rect 48412 16044 48468 16046
rect 48076 15932 48132 15988
rect 48076 15426 48132 15428
rect 48076 15374 48078 15426
rect 48078 15374 48130 15426
rect 48130 15374 48132 15426
rect 48076 15372 48132 15374
rect 47068 14530 47124 14532
rect 47068 14478 47070 14530
rect 47070 14478 47122 14530
rect 47122 14478 47124 14530
rect 47068 14476 47124 14478
rect 47964 15036 48020 15092
rect 46732 13858 46788 13860
rect 46732 13806 46734 13858
rect 46734 13806 46786 13858
rect 46786 13806 46788 13858
rect 46732 13804 46788 13806
rect 45836 11116 45892 11172
rect 46284 13468 46340 13524
rect 46732 13634 46788 13636
rect 46732 13582 46734 13634
rect 46734 13582 46786 13634
rect 46786 13582 46788 13634
rect 46732 13580 46788 13582
rect 47068 13580 47124 13636
rect 46844 13468 46900 13524
rect 47180 12850 47236 12852
rect 47180 12798 47182 12850
rect 47182 12798 47234 12850
rect 47234 12798 47236 12850
rect 47180 12796 47236 12798
rect 46508 12348 46564 12404
rect 47852 13970 47908 13972
rect 47852 13918 47854 13970
rect 47854 13918 47906 13970
rect 47906 13918 47908 13970
rect 47852 13916 47908 13918
rect 47628 13858 47684 13860
rect 47628 13806 47630 13858
rect 47630 13806 47682 13858
rect 47682 13806 47684 13858
rect 47628 13804 47684 13806
rect 47404 13580 47460 13636
rect 47740 12850 47796 12852
rect 47740 12798 47742 12850
rect 47742 12798 47794 12850
rect 47794 12798 47796 12850
rect 47740 12796 47796 12798
rect 46060 11282 46116 11284
rect 46060 11230 46062 11282
rect 46062 11230 46114 11282
rect 46114 11230 46116 11282
rect 46060 11228 46116 11230
rect 44268 8146 44324 8148
rect 44268 8094 44270 8146
rect 44270 8094 44322 8146
rect 44322 8094 44324 8146
rect 44268 8092 44324 8094
rect 44268 7308 44324 7364
rect 43708 6076 43764 6132
rect 43932 3442 43988 3444
rect 43932 3390 43934 3442
rect 43934 3390 43986 3442
rect 43986 3390 43988 3442
rect 43932 3388 43988 3390
rect 45612 7644 45668 7700
rect 45276 7532 45332 7588
rect 45164 7362 45220 7364
rect 45164 7310 45166 7362
rect 45166 7310 45218 7362
rect 45218 7310 45220 7362
rect 45164 7308 45220 7310
rect 45164 6972 45220 7028
rect 45612 7308 45668 7364
rect 46508 10610 46564 10612
rect 46508 10558 46510 10610
rect 46510 10558 46562 10610
rect 46562 10558 46564 10610
rect 46508 10556 46564 10558
rect 47404 12066 47460 12068
rect 47404 12014 47406 12066
rect 47406 12014 47458 12066
rect 47458 12014 47460 12066
rect 47404 12012 47460 12014
rect 47852 12348 47908 12404
rect 48748 30210 48804 30212
rect 48748 30158 48750 30210
rect 48750 30158 48802 30210
rect 48802 30158 48804 30210
rect 48748 30156 48804 30158
rect 48972 29986 49028 29988
rect 48972 29934 48974 29986
rect 48974 29934 49026 29986
rect 49026 29934 49028 29986
rect 48972 29932 49028 29934
rect 48860 29372 48916 29428
rect 49868 30322 49924 30324
rect 49868 30270 49870 30322
rect 49870 30270 49922 30322
rect 49922 30270 49924 30322
rect 49868 30268 49924 30270
rect 49420 30210 49476 30212
rect 49420 30158 49422 30210
rect 49422 30158 49474 30210
rect 49474 30158 49476 30210
rect 49420 30156 49476 30158
rect 49644 29820 49700 29876
rect 48748 27858 48804 27860
rect 48748 27806 48750 27858
rect 48750 27806 48802 27858
rect 48802 27806 48804 27858
rect 48748 27804 48804 27806
rect 48748 26236 48804 26292
rect 48972 26908 49028 26964
rect 50556 32954 50612 32956
rect 50556 32902 50558 32954
rect 50558 32902 50610 32954
rect 50610 32902 50612 32954
rect 50556 32900 50612 32902
rect 50660 32954 50716 32956
rect 50660 32902 50662 32954
rect 50662 32902 50714 32954
rect 50714 32902 50716 32954
rect 50660 32900 50716 32902
rect 50764 32954 50820 32956
rect 50764 32902 50766 32954
rect 50766 32902 50818 32954
rect 50818 32902 50820 32954
rect 50764 32900 50820 32902
rect 50540 31890 50596 31892
rect 50540 31838 50542 31890
rect 50542 31838 50594 31890
rect 50594 31838 50596 31890
rect 50540 31836 50596 31838
rect 55356 37042 55412 37044
rect 55356 36990 55358 37042
rect 55358 36990 55410 37042
rect 55410 36990 55412 37042
rect 55356 36988 55412 36990
rect 55580 36876 55636 36932
rect 52780 36482 52836 36484
rect 52780 36430 52782 36482
rect 52782 36430 52834 36482
rect 52834 36430 52836 36482
rect 52780 36428 52836 36430
rect 55020 35644 55076 35700
rect 55244 36316 55300 36372
rect 53228 35420 53284 35476
rect 55468 35532 55524 35588
rect 55244 35084 55300 35140
rect 55356 34972 55412 35028
rect 55244 34636 55300 34692
rect 53452 33964 53508 34020
rect 53452 33628 53508 33684
rect 53228 32732 53284 32788
rect 50556 31386 50612 31388
rect 50556 31334 50558 31386
rect 50558 31334 50610 31386
rect 50610 31334 50612 31386
rect 50556 31332 50612 31334
rect 50660 31386 50716 31388
rect 50660 31334 50662 31386
rect 50662 31334 50714 31386
rect 50714 31334 50716 31386
rect 50660 31332 50716 31334
rect 50764 31386 50820 31388
rect 50764 31334 50766 31386
rect 50766 31334 50818 31386
rect 50818 31334 50820 31386
rect 50764 31332 50820 31334
rect 50764 31106 50820 31108
rect 50764 31054 50766 31106
rect 50766 31054 50818 31106
rect 50818 31054 50820 31106
rect 50764 31052 50820 31054
rect 50428 30210 50484 30212
rect 50428 30158 50430 30210
rect 50430 30158 50482 30210
rect 50482 30158 50484 30210
rect 50428 30156 50484 30158
rect 50764 30098 50820 30100
rect 50764 30046 50766 30098
rect 50766 30046 50818 30098
rect 50818 30046 50820 30098
rect 50764 30044 50820 30046
rect 51324 31052 51380 31108
rect 50204 29986 50260 29988
rect 50204 29934 50206 29986
rect 50206 29934 50258 29986
rect 50258 29934 50260 29986
rect 50204 29932 50260 29934
rect 50652 29986 50708 29988
rect 50652 29934 50654 29986
rect 50654 29934 50706 29986
rect 50706 29934 50708 29986
rect 50652 29932 50708 29934
rect 50316 29820 50372 29876
rect 49756 26908 49812 26964
rect 49644 26514 49700 26516
rect 49644 26462 49646 26514
rect 49646 26462 49698 26514
rect 49698 26462 49700 26514
rect 49644 26460 49700 26462
rect 49532 26236 49588 26292
rect 50556 29818 50612 29820
rect 50556 29766 50558 29818
rect 50558 29766 50610 29818
rect 50610 29766 50612 29818
rect 50556 29764 50612 29766
rect 50660 29818 50716 29820
rect 50660 29766 50662 29818
rect 50662 29766 50714 29818
rect 50714 29766 50716 29818
rect 50660 29764 50716 29766
rect 50764 29818 50820 29820
rect 50764 29766 50766 29818
rect 50766 29766 50818 29818
rect 50818 29766 50820 29818
rect 50764 29764 50820 29766
rect 50556 28250 50612 28252
rect 50556 28198 50558 28250
rect 50558 28198 50610 28250
rect 50610 28198 50612 28250
rect 50556 28196 50612 28198
rect 50660 28250 50716 28252
rect 50660 28198 50662 28250
rect 50662 28198 50714 28250
rect 50714 28198 50716 28250
rect 50660 28196 50716 28198
rect 50764 28250 50820 28252
rect 50764 28198 50766 28250
rect 50766 28198 50818 28250
rect 50818 28198 50820 28250
rect 50764 28196 50820 28198
rect 50428 27132 50484 27188
rect 55020 30940 55076 30996
rect 55356 33906 55412 33908
rect 55356 33854 55358 33906
rect 55358 33854 55410 33906
rect 55410 33854 55412 33906
rect 55356 33852 55412 33854
rect 55356 33234 55412 33236
rect 55356 33182 55358 33234
rect 55358 33182 55410 33234
rect 55410 33182 55412 33234
rect 55356 33180 55412 33182
rect 55356 32338 55412 32340
rect 55356 32286 55358 32338
rect 55358 32286 55410 32338
rect 55410 32286 55412 32338
rect 55356 32284 55412 32286
rect 56588 35138 56644 35140
rect 56588 35086 56590 35138
rect 56590 35086 56642 35138
rect 56642 35086 56644 35138
rect 56588 35084 56644 35086
rect 55580 34914 55636 34916
rect 55580 34862 55582 34914
rect 55582 34862 55634 34914
rect 55634 34862 55636 34914
rect 55580 34860 55636 34862
rect 57932 34300 57988 34356
rect 55580 33346 55636 33348
rect 55580 33294 55582 33346
rect 55582 33294 55634 33346
rect 55634 33294 55636 33346
rect 55580 33292 55636 33294
rect 57932 32956 57988 33012
rect 57932 31612 57988 31668
rect 55356 30322 55412 30324
rect 55356 30270 55358 30322
rect 55358 30270 55410 30322
rect 55410 30270 55412 30322
rect 55356 30268 55412 30270
rect 50652 26962 50708 26964
rect 50652 26910 50654 26962
rect 50654 26910 50706 26962
rect 50706 26910 50708 26962
rect 50652 26908 50708 26910
rect 50556 26682 50612 26684
rect 50556 26630 50558 26682
rect 50558 26630 50610 26682
rect 50610 26630 50612 26682
rect 50556 26628 50612 26630
rect 50660 26682 50716 26684
rect 50660 26630 50662 26682
rect 50662 26630 50714 26682
rect 50714 26630 50716 26682
rect 50660 26628 50716 26630
rect 50764 26682 50820 26684
rect 50764 26630 50766 26682
rect 50766 26630 50818 26682
rect 50818 26630 50820 26682
rect 50764 26628 50820 26630
rect 50316 25900 50372 25956
rect 57036 26012 57092 26068
rect 50556 25114 50612 25116
rect 50556 25062 50558 25114
rect 50558 25062 50610 25114
rect 50610 25062 50612 25114
rect 50556 25060 50612 25062
rect 50660 25114 50716 25116
rect 50660 25062 50662 25114
rect 50662 25062 50714 25114
rect 50714 25062 50716 25114
rect 50660 25060 50716 25062
rect 50764 25114 50820 25116
rect 50764 25062 50766 25114
rect 50766 25062 50818 25114
rect 50818 25062 50820 25114
rect 50764 25060 50820 25062
rect 57596 25394 57652 25396
rect 57596 25342 57598 25394
rect 57598 25342 57650 25394
rect 57650 25342 57652 25394
rect 57596 25340 57652 25342
rect 58156 25394 58212 25396
rect 58156 25342 58158 25394
rect 58158 25342 58210 25394
rect 58210 25342 58212 25394
rect 58156 25340 58212 25342
rect 57820 25282 57876 25284
rect 57820 25230 57822 25282
rect 57822 25230 57874 25282
rect 57874 25230 57876 25282
rect 57820 25228 57876 25230
rect 57036 24892 57092 24948
rect 57820 24946 57876 24948
rect 57820 24894 57822 24946
rect 57822 24894 57874 24946
rect 57874 24894 57876 24946
rect 57820 24892 57876 24894
rect 58156 24892 58212 24948
rect 49868 24780 49924 24836
rect 49420 24722 49476 24724
rect 49420 24670 49422 24722
rect 49422 24670 49474 24722
rect 49474 24670 49476 24722
rect 49420 24668 49476 24670
rect 48860 23884 48916 23940
rect 48748 23042 48804 23044
rect 48748 22990 48750 23042
rect 48750 22990 48802 23042
rect 48802 22990 48804 23042
rect 48748 22988 48804 22990
rect 49420 23772 49476 23828
rect 49868 23772 49924 23828
rect 49644 23548 49700 23604
rect 49868 23436 49924 23492
rect 50540 24722 50596 24724
rect 50540 24670 50542 24722
rect 50542 24670 50594 24722
rect 50594 24670 50596 24722
rect 50540 24668 50596 24670
rect 50092 23938 50148 23940
rect 50092 23886 50094 23938
rect 50094 23886 50146 23938
rect 50146 23886 50148 23938
rect 50092 23884 50148 23886
rect 50204 23660 50260 23716
rect 58156 24220 58212 24276
rect 50428 23826 50484 23828
rect 50428 23774 50430 23826
rect 50430 23774 50482 23826
rect 50482 23774 50484 23826
rect 50428 23772 50484 23774
rect 50652 23660 50708 23716
rect 50988 23884 51044 23940
rect 50316 23548 50372 23604
rect 50204 23436 50260 23492
rect 50556 23546 50612 23548
rect 50556 23494 50558 23546
rect 50558 23494 50610 23546
rect 50610 23494 50612 23546
rect 50556 23492 50612 23494
rect 50660 23546 50716 23548
rect 50660 23494 50662 23546
rect 50662 23494 50714 23546
rect 50714 23494 50716 23546
rect 50660 23492 50716 23494
rect 50764 23546 50820 23548
rect 50764 23494 50766 23546
rect 50766 23494 50818 23546
rect 50818 23494 50820 23546
rect 50764 23492 50820 23494
rect 48972 22316 49028 22372
rect 49644 21196 49700 21252
rect 48860 19628 48916 19684
rect 48748 18338 48804 18340
rect 48748 18286 48750 18338
rect 48750 18286 48802 18338
rect 48802 18286 48804 18338
rect 48748 18284 48804 18286
rect 48972 17890 49028 17892
rect 48972 17838 48974 17890
rect 48974 17838 49026 17890
rect 49026 17838 49028 17890
rect 48972 17836 49028 17838
rect 48748 17666 48804 17668
rect 48748 17614 48750 17666
rect 48750 17614 48802 17666
rect 48802 17614 48804 17666
rect 48748 17612 48804 17614
rect 48860 17388 48916 17444
rect 49308 17106 49364 17108
rect 49308 17054 49310 17106
rect 49310 17054 49362 17106
rect 49362 17054 49364 17106
rect 49308 17052 49364 17054
rect 50556 21978 50612 21980
rect 50556 21926 50558 21978
rect 50558 21926 50610 21978
rect 50610 21926 50612 21978
rect 50556 21924 50612 21926
rect 50660 21978 50716 21980
rect 50660 21926 50662 21978
rect 50662 21926 50714 21978
rect 50714 21926 50716 21978
rect 50660 21924 50716 21926
rect 50764 21978 50820 21980
rect 50764 21926 50766 21978
rect 50766 21926 50818 21978
rect 50818 21926 50820 21978
rect 50764 21924 50820 21926
rect 50092 20748 50148 20804
rect 50556 20410 50612 20412
rect 50556 20358 50558 20410
rect 50558 20358 50610 20410
rect 50610 20358 50612 20410
rect 50556 20356 50612 20358
rect 50660 20410 50716 20412
rect 50660 20358 50662 20410
rect 50662 20358 50714 20410
rect 50714 20358 50716 20410
rect 50660 20356 50716 20358
rect 50764 20410 50820 20412
rect 50764 20358 50766 20410
rect 50766 20358 50818 20410
rect 50818 20358 50820 20410
rect 50764 20356 50820 20358
rect 50556 18842 50612 18844
rect 50556 18790 50558 18842
rect 50558 18790 50610 18842
rect 50610 18790 50612 18842
rect 50556 18788 50612 18790
rect 50660 18842 50716 18844
rect 50660 18790 50662 18842
rect 50662 18790 50714 18842
rect 50714 18790 50716 18842
rect 50660 18788 50716 18790
rect 50764 18842 50820 18844
rect 50764 18790 50766 18842
rect 50766 18790 50818 18842
rect 50818 18790 50820 18842
rect 50764 18788 50820 18790
rect 49756 18284 49812 18340
rect 50556 17274 50612 17276
rect 50556 17222 50558 17274
rect 50558 17222 50610 17274
rect 50610 17222 50612 17274
rect 50556 17220 50612 17222
rect 50660 17274 50716 17276
rect 50660 17222 50662 17274
rect 50662 17222 50714 17274
rect 50714 17222 50716 17274
rect 50660 17220 50716 17222
rect 50764 17274 50820 17276
rect 50764 17222 50766 17274
rect 50766 17222 50818 17274
rect 50818 17222 50820 17274
rect 50764 17220 50820 17222
rect 49196 16994 49252 16996
rect 49196 16942 49198 16994
rect 49198 16942 49250 16994
rect 49250 16942 49252 16994
rect 49196 16940 49252 16942
rect 48748 15874 48804 15876
rect 48748 15822 48750 15874
rect 48750 15822 48802 15874
rect 48802 15822 48804 15874
rect 48748 15820 48804 15822
rect 48748 15538 48804 15540
rect 48748 15486 48750 15538
rect 48750 15486 48802 15538
rect 48802 15486 48804 15538
rect 48748 15484 48804 15486
rect 48412 13580 48468 13636
rect 48524 13244 48580 13300
rect 48972 15874 49028 15876
rect 48972 15822 48974 15874
rect 48974 15822 49026 15874
rect 49026 15822 49028 15874
rect 48972 15820 49028 15822
rect 48972 15148 49028 15204
rect 50876 16940 50932 16996
rect 49980 16210 50036 16212
rect 49980 16158 49982 16210
rect 49982 16158 50034 16210
rect 50034 16158 50036 16210
rect 49980 16156 50036 16158
rect 49756 16044 49812 16100
rect 49420 15986 49476 15988
rect 49420 15934 49422 15986
rect 49422 15934 49474 15986
rect 49474 15934 49476 15986
rect 49420 15932 49476 15934
rect 49532 15820 49588 15876
rect 50428 16098 50484 16100
rect 50428 16046 50430 16098
rect 50430 16046 50482 16098
rect 50482 16046 50484 16098
rect 50428 16044 50484 16046
rect 50556 15706 50612 15708
rect 50556 15654 50558 15706
rect 50558 15654 50610 15706
rect 50610 15654 50612 15706
rect 50556 15652 50612 15654
rect 50660 15706 50716 15708
rect 50660 15654 50662 15706
rect 50662 15654 50714 15706
rect 50714 15654 50716 15706
rect 50660 15652 50716 15654
rect 50764 15706 50820 15708
rect 50764 15654 50766 15706
rect 50766 15654 50818 15706
rect 50818 15654 50820 15706
rect 50764 15652 50820 15654
rect 57820 23714 57876 23716
rect 57820 23662 57822 23714
rect 57822 23662 57874 23714
rect 57874 23662 57876 23714
rect 57820 23660 57876 23662
rect 57596 23548 57652 23604
rect 58156 23548 58212 23604
rect 57596 22258 57652 22260
rect 57596 22206 57598 22258
rect 57598 22206 57650 22258
rect 57650 22206 57652 22258
rect 57596 22204 57652 22206
rect 58156 22258 58212 22260
rect 58156 22206 58158 22258
rect 58158 22206 58210 22258
rect 58210 22206 58212 22258
rect 58156 22204 58212 22206
rect 57820 22146 57876 22148
rect 57820 22094 57822 22146
rect 57822 22094 57874 22146
rect 57874 22094 57876 22146
rect 57820 22092 57876 22094
rect 53788 21868 53844 21924
rect 58156 21532 58212 21588
rect 53788 20076 53844 20132
rect 48972 13746 49028 13748
rect 48972 13694 48974 13746
rect 48974 13694 49026 13746
rect 49026 13694 49028 13746
rect 48972 13692 49028 13694
rect 49420 15036 49476 15092
rect 48860 13634 48916 13636
rect 48860 13582 48862 13634
rect 48862 13582 48914 13634
rect 48914 13582 48916 13634
rect 48860 13580 48916 13582
rect 48860 13244 48916 13300
rect 49196 13970 49252 13972
rect 49196 13918 49198 13970
rect 49198 13918 49250 13970
rect 49250 13918 49252 13970
rect 49196 13916 49252 13918
rect 51660 15036 51716 15092
rect 52780 15036 52836 15092
rect 49868 14476 49924 14532
rect 50556 14138 50612 14140
rect 50556 14086 50558 14138
rect 50558 14086 50610 14138
rect 50610 14086 50612 14138
rect 50556 14084 50612 14086
rect 50660 14138 50716 14140
rect 50660 14086 50662 14138
rect 50662 14086 50714 14138
rect 50714 14086 50716 14138
rect 50660 14084 50716 14086
rect 50764 14138 50820 14140
rect 50764 14086 50766 14138
rect 50766 14086 50818 14138
rect 50818 14086 50820 14138
rect 50764 14084 50820 14086
rect 48860 12402 48916 12404
rect 48860 12350 48862 12402
rect 48862 12350 48914 12402
rect 48914 12350 48916 12402
rect 48860 12348 48916 12350
rect 49420 13244 49476 13300
rect 50556 12570 50612 12572
rect 50556 12518 50558 12570
rect 50558 12518 50610 12570
rect 50610 12518 50612 12570
rect 50556 12516 50612 12518
rect 50660 12570 50716 12572
rect 50660 12518 50662 12570
rect 50662 12518 50714 12570
rect 50714 12518 50716 12570
rect 50660 12516 50716 12518
rect 50764 12570 50820 12572
rect 50764 12518 50766 12570
rect 50766 12518 50818 12570
rect 50818 12518 50820 12570
rect 50764 12516 50820 12518
rect 50556 11002 50612 11004
rect 50556 10950 50558 11002
rect 50558 10950 50610 11002
rect 50610 10950 50612 11002
rect 50556 10948 50612 10950
rect 50660 11002 50716 11004
rect 50660 10950 50662 11002
rect 50662 10950 50714 11002
rect 50714 10950 50716 11002
rect 50660 10948 50716 10950
rect 50764 11002 50820 11004
rect 50764 10950 50766 11002
rect 50766 10950 50818 11002
rect 50818 10950 50820 11002
rect 50764 10948 50820 10950
rect 50556 9434 50612 9436
rect 50556 9382 50558 9434
rect 50558 9382 50610 9434
rect 50610 9382 50612 9434
rect 50556 9380 50612 9382
rect 50660 9434 50716 9436
rect 50660 9382 50662 9434
rect 50662 9382 50714 9434
rect 50714 9382 50716 9434
rect 50660 9380 50716 9382
rect 50764 9434 50820 9436
rect 50764 9382 50766 9434
rect 50766 9382 50818 9434
rect 50818 9382 50820 9434
rect 50764 9380 50820 9382
rect 46172 8316 46228 8372
rect 47852 8370 47908 8372
rect 47852 8318 47854 8370
rect 47854 8318 47906 8370
rect 47906 8318 47908 8370
rect 47852 8316 47908 8318
rect 50556 7866 50612 7868
rect 50556 7814 50558 7866
rect 50558 7814 50610 7866
rect 50610 7814 50612 7866
rect 50556 7812 50612 7814
rect 50660 7866 50716 7868
rect 50660 7814 50662 7866
rect 50662 7814 50714 7866
rect 50714 7814 50716 7866
rect 50660 7812 50716 7814
rect 50764 7866 50820 7868
rect 50764 7814 50766 7866
rect 50766 7814 50818 7866
rect 50818 7814 50820 7866
rect 50764 7812 50820 7814
rect 46172 7532 46228 7588
rect 46060 6972 46116 7028
rect 50556 6298 50612 6300
rect 50556 6246 50558 6298
rect 50558 6246 50610 6298
rect 50610 6246 50612 6298
rect 50556 6244 50612 6246
rect 50660 6298 50716 6300
rect 50660 6246 50662 6298
rect 50662 6246 50714 6298
rect 50714 6246 50716 6298
rect 50660 6244 50716 6246
rect 50764 6298 50820 6300
rect 50764 6246 50766 6298
rect 50766 6246 50818 6298
rect 50818 6246 50820 6298
rect 50764 6244 50820 6246
rect 50556 4730 50612 4732
rect 50556 4678 50558 4730
rect 50558 4678 50610 4730
rect 50610 4678 50612 4730
rect 50556 4676 50612 4678
rect 50660 4730 50716 4732
rect 50660 4678 50662 4730
rect 50662 4678 50714 4730
rect 50714 4678 50716 4730
rect 50660 4676 50716 4678
rect 50764 4730 50820 4732
rect 50764 4678 50766 4730
rect 50766 4678 50818 4730
rect 50818 4678 50820 4730
rect 50764 4676 50820 4678
rect 50556 3162 50612 3164
rect 50556 3110 50558 3162
rect 50558 3110 50610 3162
rect 50610 3110 50612 3162
rect 50556 3108 50612 3110
rect 50660 3162 50716 3164
rect 50660 3110 50662 3162
rect 50662 3110 50714 3162
rect 50714 3110 50716 3162
rect 50660 3108 50716 3110
rect 50764 3162 50820 3164
rect 50764 3110 50766 3162
rect 50766 3110 50818 3162
rect 50818 3110 50820 3162
rect 50764 3108 50820 3110
<< metal3 >>
rect 19826 76804 19836 76860
rect 19892 76804 19940 76860
rect 19996 76804 20044 76860
rect 20100 76804 20110 76860
rect 50546 76804 50556 76860
rect 50612 76804 50660 76860
rect 50716 76804 50764 76860
rect 50820 76804 50830 76860
rect 4466 76020 4476 76076
rect 4532 76020 4580 76076
rect 4636 76020 4684 76076
rect 4740 76020 4750 76076
rect 35186 76020 35196 76076
rect 35252 76020 35300 76076
rect 35356 76020 35404 76076
rect 35460 76020 35470 76076
rect 19826 75236 19836 75292
rect 19892 75236 19940 75292
rect 19996 75236 20044 75292
rect 20100 75236 20110 75292
rect 50546 75236 50556 75292
rect 50612 75236 50660 75292
rect 50716 75236 50764 75292
rect 50820 75236 50830 75292
rect 4466 74452 4476 74508
rect 4532 74452 4580 74508
rect 4636 74452 4684 74508
rect 4740 74452 4750 74508
rect 35186 74452 35196 74508
rect 35252 74452 35300 74508
rect 35356 74452 35404 74508
rect 35460 74452 35470 74508
rect 19826 73668 19836 73724
rect 19892 73668 19940 73724
rect 19996 73668 20044 73724
rect 20100 73668 20110 73724
rect 50546 73668 50556 73724
rect 50612 73668 50660 73724
rect 50716 73668 50764 73724
rect 50820 73668 50830 73724
rect 4466 72884 4476 72940
rect 4532 72884 4580 72940
rect 4636 72884 4684 72940
rect 4740 72884 4750 72940
rect 35186 72884 35196 72940
rect 35252 72884 35300 72940
rect 35356 72884 35404 72940
rect 35460 72884 35470 72940
rect 19826 72100 19836 72156
rect 19892 72100 19940 72156
rect 19996 72100 20044 72156
rect 20100 72100 20110 72156
rect 50546 72100 50556 72156
rect 50612 72100 50660 72156
rect 50716 72100 50764 72156
rect 50820 72100 50830 72156
rect 40226 71596 40236 71652
rect 40292 71596 40908 71652
rect 40964 71596 40974 71652
rect 4466 71316 4476 71372
rect 4532 71316 4580 71372
rect 4636 71316 4684 71372
rect 4740 71316 4750 71372
rect 35186 71316 35196 71372
rect 35252 71316 35300 71372
rect 35356 71316 35404 71372
rect 35460 71316 35470 71372
rect 41906 70700 41916 70756
rect 41972 70700 42700 70756
rect 42756 70700 42766 70756
rect 0 70644 800 70672
rect 0 70588 4172 70644
rect 4228 70588 4238 70644
rect 38434 70588 38444 70644
rect 38500 70588 40348 70644
rect 40404 70588 40414 70644
rect 0 70560 800 70588
rect 19826 70532 19836 70588
rect 19892 70532 19940 70588
rect 19996 70532 20044 70588
rect 20100 70532 20110 70588
rect 50546 70532 50556 70588
rect 50612 70532 50660 70588
rect 50716 70532 50764 70588
rect 50820 70532 50830 70588
rect 31602 70476 31612 70532
rect 31668 70476 33180 70532
rect 33236 70476 36428 70532
rect 36484 70476 37212 70532
rect 37268 70476 39564 70532
rect 39620 70476 39630 70532
rect 39890 70252 39900 70308
rect 39956 70252 40908 70308
rect 40964 70252 40974 70308
rect 40338 70140 40348 70196
rect 40404 70140 41244 70196
rect 41300 70140 43820 70196
rect 43876 70140 43886 70196
rect 29698 70028 29708 70084
rect 29764 70028 30716 70084
rect 30772 70028 30782 70084
rect 22866 69916 22876 69972
rect 22932 69916 23884 69972
rect 23940 69916 23950 69972
rect 4466 69748 4476 69804
rect 4532 69748 4580 69804
rect 4636 69748 4684 69804
rect 4740 69748 4750 69804
rect 35186 69748 35196 69804
rect 35252 69748 35300 69804
rect 35356 69748 35404 69804
rect 35460 69748 35470 69804
rect 30370 69580 30380 69636
rect 30436 69580 31276 69636
rect 31332 69580 31342 69636
rect 36418 69580 36428 69636
rect 36484 69580 37212 69636
rect 37268 69580 37278 69636
rect 41458 69468 41468 69524
rect 41524 69468 42588 69524
rect 42644 69468 42654 69524
rect 25330 69356 25340 69412
rect 25396 69356 27804 69412
rect 27860 69356 27870 69412
rect 34402 69356 34412 69412
rect 34468 69356 36092 69412
rect 36148 69356 36158 69412
rect 36978 69356 36988 69412
rect 37044 69356 38556 69412
rect 38612 69356 38622 69412
rect 29026 69244 29036 69300
rect 29092 69244 31836 69300
rect 31892 69244 31902 69300
rect 33282 69244 33292 69300
rect 33348 69244 34972 69300
rect 35028 69244 35038 69300
rect 36306 69244 36316 69300
rect 36372 69244 37548 69300
rect 37604 69244 37614 69300
rect 39330 69244 39340 69300
rect 39396 69244 40460 69300
rect 40516 69244 40526 69300
rect 33292 69188 33348 69244
rect 29222 69132 29260 69188
rect 29316 69132 29326 69188
rect 30818 69132 30828 69188
rect 30884 69132 31276 69188
rect 31332 69132 31612 69188
rect 31668 69132 33348 69188
rect 33954 69132 33964 69188
rect 34020 69132 34636 69188
rect 34692 69132 34702 69188
rect 37426 69132 37436 69188
rect 37492 69132 38332 69188
rect 38388 69132 40124 69188
rect 40180 69132 40190 69188
rect 42130 69132 42140 69188
rect 42196 69132 42924 69188
rect 42980 69132 44156 69188
rect 44212 69132 44222 69188
rect 29922 69020 29932 69076
rect 29988 69020 33068 69076
rect 33124 69020 34188 69076
rect 34244 69020 34254 69076
rect 19826 68964 19836 69020
rect 19892 68964 19940 69020
rect 19996 68964 20044 69020
rect 20100 68964 20110 69020
rect 50546 68964 50556 69020
rect 50612 68964 50660 69020
rect 50716 68964 50764 69020
rect 50820 68964 50830 69020
rect 22194 68908 22204 68964
rect 22260 68908 22988 68964
rect 23044 68908 25340 68964
rect 25396 68908 25406 68964
rect 29698 68908 29708 68964
rect 29764 68908 30828 68964
rect 30884 68908 30894 68964
rect 32834 68908 32844 68964
rect 32900 68908 35084 68964
rect 35140 68908 35532 68964
rect 35588 68908 35598 68964
rect 38434 68908 38444 68964
rect 38500 68908 39340 68964
rect 39396 68908 39406 68964
rect 40898 68908 40908 68964
rect 40964 68908 42364 68964
rect 42420 68908 44156 68964
rect 44212 68908 45164 68964
rect 45220 68908 45230 68964
rect 29362 68796 29372 68852
rect 29428 68796 30044 68852
rect 30100 68796 30110 68852
rect 33506 68796 33516 68852
rect 33572 68796 34972 68852
rect 35028 68796 37324 68852
rect 37380 68796 38108 68852
rect 38164 68796 38174 68852
rect 39106 68796 39116 68852
rect 39172 68796 41356 68852
rect 41412 68796 41422 68852
rect 34412 68740 34468 68796
rect 34402 68684 34412 68740
rect 34468 68684 34478 68740
rect 39218 68684 39228 68740
rect 39284 68684 39294 68740
rect 40450 68684 40460 68740
rect 40516 68684 41244 68740
rect 41300 68684 41310 68740
rect 39228 68628 39284 68684
rect 31042 68572 31052 68628
rect 31108 68572 32956 68628
rect 33012 68572 33022 68628
rect 35746 68572 35756 68628
rect 35812 68572 36428 68628
rect 36484 68572 37324 68628
rect 37380 68572 39284 68628
rect 35970 68460 35980 68516
rect 36036 68460 37100 68516
rect 37156 68460 37884 68516
rect 37940 68460 40124 68516
rect 40180 68460 40796 68516
rect 40852 68460 40862 68516
rect 4466 68180 4476 68236
rect 4532 68180 4580 68236
rect 4636 68180 4684 68236
rect 4740 68180 4750 68236
rect 35186 68180 35196 68236
rect 35252 68180 35300 68236
rect 35356 68180 35404 68236
rect 35460 68180 35470 68236
rect 20738 68124 20748 68180
rect 20804 68124 21308 68180
rect 21364 68124 22876 68180
rect 22932 68124 31500 68180
rect 31556 68124 31566 68180
rect 23426 68012 23436 68068
rect 23492 68012 26628 68068
rect 26572 67844 26628 68012
rect 19842 67788 19852 67844
rect 19908 67788 21868 67844
rect 21924 67788 22428 67844
rect 22484 67788 22494 67844
rect 24658 67788 24668 67844
rect 24724 67788 25452 67844
rect 25508 67788 26124 67844
rect 26180 67788 26190 67844
rect 26572 67788 28028 67844
rect 28084 67788 28094 67844
rect 37650 67788 37660 67844
rect 37716 67788 39004 67844
rect 39060 67788 39070 67844
rect 21298 67676 21308 67732
rect 21364 67676 21980 67732
rect 22036 67676 22046 67732
rect 24882 67676 24892 67732
rect 24948 67676 26348 67732
rect 26404 67676 26414 67732
rect 22082 67564 22092 67620
rect 22148 67564 23772 67620
rect 23828 67564 24332 67620
rect 24388 67564 25564 67620
rect 25620 67564 25630 67620
rect 25778 67564 25788 67620
rect 25844 67564 28364 67620
rect 28420 67564 28430 67620
rect 35858 67564 35868 67620
rect 35924 67564 39676 67620
rect 39732 67564 39742 67620
rect 40226 67564 40236 67620
rect 40292 67564 41916 67620
rect 41972 67564 45836 67620
rect 45892 67564 45902 67620
rect 23986 67452 23996 67508
rect 24052 67452 24444 67508
rect 24500 67452 29708 67508
rect 29764 67452 31164 67508
rect 31220 67452 31230 67508
rect 38098 67452 38108 67508
rect 38164 67452 38780 67508
rect 38836 67452 42140 67508
rect 42196 67452 42206 67508
rect 19826 67396 19836 67452
rect 19892 67396 19940 67452
rect 19996 67396 20044 67452
rect 20100 67396 20110 67452
rect 50546 67396 50556 67452
rect 50612 67396 50660 67452
rect 50716 67396 50764 67452
rect 50820 67396 50830 67452
rect 22194 67340 22204 67396
rect 22260 67340 22876 67396
rect 22932 67340 23100 67396
rect 23156 67340 23548 67396
rect 23604 67340 24668 67396
rect 24724 67340 24734 67396
rect 30034 67340 30044 67396
rect 30100 67340 30380 67396
rect 30436 67340 33068 67396
rect 33124 67340 33134 67396
rect 20514 67228 20524 67284
rect 20580 67228 26236 67284
rect 26292 67228 29260 67284
rect 29316 67228 29326 67284
rect 29474 67228 29484 67284
rect 29540 67228 30604 67284
rect 30660 67228 30670 67284
rect 39666 67228 39676 67284
rect 39732 67228 42028 67284
rect 42084 67228 42094 67284
rect 23314 67116 23324 67172
rect 23380 67116 23996 67172
rect 24052 67116 24062 67172
rect 28354 67116 28364 67172
rect 28420 67116 29148 67172
rect 29204 67116 29214 67172
rect 32498 67116 32508 67172
rect 32564 67116 33404 67172
rect 33460 67116 33470 67172
rect 41346 67116 41356 67172
rect 41412 67116 42588 67172
rect 42644 67116 43260 67172
rect 43316 67116 43326 67172
rect 43474 67116 43484 67172
rect 43540 67116 44492 67172
rect 44548 67116 45052 67172
rect 45108 67116 45220 67172
rect 45164 67060 45220 67116
rect 21074 67004 21084 67060
rect 21140 67004 23100 67060
rect 23156 67004 23166 67060
rect 28578 67004 28588 67060
rect 28644 67004 30156 67060
rect 30212 67004 30604 67060
rect 30660 67004 30670 67060
rect 32050 67004 32060 67060
rect 32116 67004 35532 67060
rect 35588 67004 35598 67060
rect 42802 67004 42812 67060
rect 42868 67004 44940 67060
rect 44996 67004 45006 67060
rect 45164 67004 45388 67060
rect 45444 67004 45454 67060
rect 20514 66892 20524 66948
rect 20580 66892 21308 66948
rect 21364 66892 24220 66948
rect 24276 66892 24286 66948
rect 30034 66892 30044 66948
rect 30100 66892 30716 66948
rect 30772 66892 34748 66948
rect 34804 66892 41132 66948
rect 41188 66892 42252 66948
rect 42308 66892 42318 66948
rect 14242 66780 14252 66836
rect 14308 66780 15260 66836
rect 15316 66780 15326 66836
rect 22418 66780 22428 66836
rect 22484 66780 22876 66836
rect 22932 66780 24332 66836
rect 24388 66780 24398 66836
rect 39106 66780 39116 66836
rect 39172 66780 39452 66836
rect 39508 66780 39518 66836
rect 40562 66780 40572 66836
rect 40628 66780 41468 66836
rect 41524 66780 42476 66836
rect 42532 66780 43260 66836
rect 43316 66780 43326 66836
rect 4466 66612 4476 66668
rect 4532 66612 4580 66668
rect 4636 66612 4684 66668
rect 4740 66612 4750 66668
rect 35186 66612 35196 66668
rect 35252 66612 35300 66668
rect 35356 66612 35404 66668
rect 35460 66612 35470 66668
rect 26236 66444 27020 66500
rect 27076 66444 34188 66500
rect 34244 66444 34524 66500
rect 34580 66444 34590 66500
rect 43362 66444 43372 66500
rect 43428 66444 44044 66500
rect 44100 66444 44110 66500
rect 21410 66332 21420 66388
rect 21476 66332 21868 66388
rect 21924 66332 21934 66388
rect 26236 66276 26292 66444
rect 44482 66332 44492 66388
rect 44548 66332 44828 66388
rect 44884 66332 45612 66388
rect 45668 66332 45678 66388
rect 26226 66220 26236 66276
rect 26292 66220 26302 66276
rect 27794 66220 27804 66276
rect 27860 66220 28252 66276
rect 28308 66220 28700 66276
rect 28756 66220 28766 66276
rect 29250 66220 29260 66276
rect 29316 66220 31052 66276
rect 31108 66220 31118 66276
rect 41206 66220 41244 66276
rect 41300 66220 41310 66276
rect 42466 66220 42476 66276
rect 42532 66220 43652 66276
rect 43596 66164 43652 66220
rect 25414 66108 25452 66164
rect 25508 66108 26124 66164
rect 26180 66108 26190 66164
rect 36194 66108 36204 66164
rect 36260 66108 36988 66164
rect 37044 66108 37054 66164
rect 41906 66108 41916 66164
rect 41972 66108 42700 66164
rect 42756 66108 42766 66164
rect 43586 66108 43596 66164
rect 43652 66108 44268 66164
rect 44324 66108 44334 66164
rect 20178 65996 20188 66052
rect 20244 65996 20524 66052
rect 20580 65996 21420 66052
rect 21476 65996 21486 66052
rect 24770 65996 24780 66052
rect 24836 65996 25564 66052
rect 25620 65996 25630 66052
rect 26898 65996 26908 66052
rect 26964 65996 27244 66052
rect 27300 65996 27310 66052
rect 29250 65996 29260 66052
rect 29316 65996 30044 66052
rect 30100 65996 30110 66052
rect 31602 65996 31612 66052
rect 31668 65996 33292 66052
rect 33348 65996 33358 66052
rect 33506 65996 33516 66052
rect 33572 65996 33964 66052
rect 34020 65996 34030 66052
rect 35410 65996 35420 66052
rect 35476 65996 36316 66052
rect 36372 65996 37660 66052
rect 37716 65996 37726 66052
rect 39890 65996 39900 66052
rect 39956 65996 40348 66052
rect 40404 65996 40414 66052
rect 41122 65996 41132 66052
rect 41188 65996 41692 66052
rect 41748 65996 41758 66052
rect 42802 65996 42812 66052
rect 42868 65996 43036 66052
rect 43092 65996 43708 66052
rect 43764 65996 43774 66052
rect 44594 65996 44604 66052
rect 44660 65996 45164 66052
rect 45220 65996 45230 66052
rect 33394 65884 33404 65940
rect 33460 65884 33740 65940
rect 33796 65884 33806 65940
rect 19826 65828 19836 65884
rect 19892 65828 19940 65884
rect 19996 65828 20044 65884
rect 20100 65828 20110 65884
rect 50546 65828 50556 65884
rect 50612 65828 50660 65884
rect 50716 65828 50764 65884
rect 50820 65828 50830 65884
rect 25218 65772 25228 65828
rect 25284 65772 25676 65828
rect 25732 65772 26180 65828
rect 26124 65716 26180 65772
rect 14018 65660 14028 65716
rect 14084 65660 14924 65716
rect 14980 65660 16380 65716
rect 16436 65660 16446 65716
rect 24434 65660 24444 65716
rect 24500 65660 24510 65716
rect 24994 65660 25004 65716
rect 25060 65660 25788 65716
rect 25844 65660 25854 65716
rect 26114 65660 26124 65716
rect 26180 65660 26190 65716
rect 33394 65660 33404 65716
rect 33460 65660 34244 65716
rect 41682 65660 41692 65716
rect 41748 65660 43820 65716
rect 43876 65660 44380 65716
rect 44436 65660 44446 65716
rect 24444 65604 24500 65660
rect 34188 65604 34244 65660
rect 16482 65548 16492 65604
rect 16548 65548 17500 65604
rect 17556 65548 18508 65604
rect 18564 65548 18574 65604
rect 24444 65548 25340 65604
rect 25396 65548 25900 65604
rect 25956 65548 25966 65604
rect 32610 65548 32620 65604
rect 32676 65548 33516 65604
rect 33572 65548 33582 65604
rect 34178 65548 34188 65604
rect 34244 65548 34254 65604
rect 42578 65548 42588 65604
rect 42644 65548 43372 65604
rect 43428 65548 43438 65604
rect 15250 65436 15260 65492
rect 15316 65436 17724 65492
rect 17780 65436 17790 65492
rect 23090 65436 23100 65492
rect 23156 65436 26572 65492
rect 26628 65436 26638 65492
rect 27458 65436 27468 65492
rect 27524 65436 30156 65492
rect 30212 65436 30222 65492
rect 31938 65436 31948 65492
rect 32004 65436 32284 65492
rect 32340 65436 32350 65492
rect 32498 65436 32508 65492
rect 32564 65436 34972 65492
rect 35028 65436 35038 65492
rect 35186 65436 35196 65492
rect 35252 65436 37324 65492
rect 37380 65436 37390 65492
rect 38882 65436 38892 65492
rect 38948 65436 40236 65492
rect 40292 65436 43036 65492
rect 43092 65436 43102 65492
rect 43922 65436 43932 65492
rect 43988 65436 44940 65492
rect 44996 65436 47516 65492
rect 47572 65436 47582 65492
rect 12674 65324 12684 65380
rect 12740 65324 13916 65380
rect 13972 65324 13982 65380
rect 21746 65324 21756 65380
rect 21812 65324 23212 65380
rect 23268 65324 23278 65380
rect 25218 65324 25228 65380
rect 25284 65324 26012 65380
rect 26068 65324 26908 65380
rect 28354 65324 28364 65380
rect 28420 65324 29372 65380
rect 29428 65324 29438 65380
rect 32834 65324 32844 65380
rect 32900 65324 32910 65380
rect 33618 65324 33628 65380
rect 33684 65324 33964 65380
rect 34020 65324 34030 65380
rect 26852 65268 26908 65324
rect 32844 65268 32900 65324
rect 35196 65268 35252 65436
rect 39330 65324 39340 65380
rect 39396 65324 39900 65380
rect 39956 65324 41020 65380
rect 41076 65324 42700 65380
rect 42756 65324 42766 65380
rect 22866 65212 22876 65268
rect 22932 65212 23436 65268
rect 23492 65212 23502 65268
rect 26852 65212 32900 65268
rect 34066 65212 34076 65268
rect 34132 65212 35252 65268
rect 36418 65212 36428 65268
rect 36484 65212 38332 65268
rect 38388 65212 38398 65268
rect 39106 65212 39116 65268
rect 39172 65212 40124 65268
rect 40180 65212 40190 65268
rect 38882 65100 38892 65156
rect 38948 65100 39228 65156
rect 39284 65100 39294 65156
rect 42018 65100 42028 65156
rect 42084 65100 43260 65156
rect 43316 65100 43326 65156
rect 4466 65044 4476 65100
rect 4532 65044 4580 65100
rect 4636 65044 4684 65100
rect 4740 65044 4750 65100
rect 35186 65044 35196 65100
rect 35252 65044 35300 65100
rect 35356 65044 35404 65100
rect 35460 65044 35470 65100
rect 16370 64876 16380 64932
rect 16436 64876 17836 64932
rect 17892 64876 17902 64932
rect 41234 64876 41244 64932
rect 41300 64876 41692 64932
rect 41748 64876 41758 64932
rect 10098 64764 10108 64820
rect 10164 64764 13132 64820
rect 13188 64764 14364 64820
rect 14420 64764 14430 64820
rect 17938 64764 17948 64820
rect 18004 64764 19964 64820
rect 20020 64764 20030 64820
rect 14812 64652 26908 64708
rect 27458 64652 27468 64708
rect 27524 64652 29372 64708
rect 29428 64652 30268 64708
rect 30324 64652 30334 64708
rect 35746 64652 35756 64708
rect 35812 64652 37212 64708
rect 37268 64652 37278 64708
rect 14812 64596 14868 64652
rect 26852 64596 26908 64652
rect 14466 64540 14476 64596
rect 14532 64540 14868 64596
rect 15026 64540 15036 64596
rect 15092 64540 17388 64596
rect 17444 64540 17454 64596
rect 26852 64540 27356 64596
rect 27412 64540 27804 64596
rect 27860 64540 27870 64596
rect 34066 64540 34076 64596
rect 34132 64540 34972 64596
rect 35028 64540 35038 64596
rect 40114 64540 40124 64596
rect 40180 64540 42252 64596
rect 42308 64540 42318 64596
rect 43026 64540 43036 64596
rect 43092 64540 43204 64596
rect 14018 64428 14028 64484
rect 14084 64428 15148 64484
rect 15204 64428 16380 64484
rect 16436 64428 16446 64484
rect 23538 64428 23548 64484
rect 23604 64428 26460 64484
rect 26516 64428 26526 64484
rect 26852 64428 32172 64484
rect 32228 64428 32238 64484
rect 32386 64428 32396 64484
rect 32452 64428 34412 64484
rect 34468 64428 34478 64484
rect 40450 64428 40460 64484
rect 40516 64428 41020 64484
rect 41076 64428 42140 64484
rect 42196 64428 42206 64484
rect 26852 64372 26908 64428
rect 43148 64372 43204 64540
rect 44034 64428 44044 64484
rect 44100 64428 45276 64484
rect 45332 64428 45342 64484
rect 15092 64316 16156 64372
rect 16212 64316 17612 64372
rect 17668 64316 17678 64372
rect 26338 64316 26348 64372
rect 26404 64316 26908 64372
rect 27234 64316 27244 64372
rect 27300 64316 28588 64372
rect 28644 64316 29820 64372
rect 29876 64316 29886 64372
rect 30706 64316 30716 64372
rect 30772 64316 35812 64372
rect 35970 64316 35980 64372
rect 36036 64316 36652 64372
rect 36708 64316 41244 64372
rect 41300 64316 44716 64372
rect 44772 64316 44782 64372
rect 15092 64260 15148 64316
rect 19826 64260 19836 64316
rect 19892 64260 19940 64316
rect 19996 64260 20044 64316
rect 20100 64260 20110 64316
rect 35756 64260 35812 64316
rect 50546 64260 50556 64316
rect 50612 64260 50660 64316
rect 50716 64260 50764 64316
rect 50820 64260 50830 64316
rect 13794 64204 13804 64260
rect 13860 64204 15148 64260
rect 15586 64204 15596 64260
rect 15652 64204 16604 64260
rect 16660 64204 17948 64260
rect 18004 64204 18014 64260
rect 24546 64204 24556 64260
rect 24612 64204 26460 64260
rect 26516 64204 26526 64260
rect 27346 64204 27356 64260
rect 27412 64204 28924 64260
rect 28980 64204 29484 64260
rect 29540 64204 30156 64260
rect 30212 64204 30222 64260
rect 31714 64204 31724 64260
rect 31780 64204 33964 64260
rect 34020 64204 34524 64260
rect 34580 64204 34590 64260
rect 35756 64204 38332 64260
rect 38388 64204 38398 64260
rect 38612 64204 42252 64260
rect 42308 64204 42588 64260
rect 42644 64204 43484 64260
rect 43540 64204 43550 64260
rect 15362 64092 15372 64148
rect 15428 64092 16268 64148
rect 16324 64092 16334 64148
rect 22978 64092 22988 64148
rect 23044 64092 24444 64148
rect 24500 64092 24510 64148
rect 27010 64092 27020 64148
rect 27076 64092 28588 64148
rect 28644 64092 28654 64148
rect 33506 64092 33516 64148
rect 33572 64092 34636 64148
rect 34692 64092 34702 64148
rect 37314 64092 37324 64148
rect 37380 64092 37996 64148
rect 38052 64092 38062 64148
rect 38612 64036 38668 64204
rect 38882 64092 38892 64148
rect 38948 64092 39340 64148
rect 39396 64092 39406 64148
rect 41234 64092 41244 64148
rect 41300 64092 42476 64148
rect 42532 64092 42542 64148
rect 45490 64092 45500 64148
rect 45556 64092 46844 64148
rect 46900 64092 47180 64148
rect 47236 64092 47246 64148
rect 12450 63980 12460 64036
rect 12516 63980 13916 64036
rect 13972 63980 13982 64036
rect 14914 63980 14924 64036
rect 14980 63980 15932 64036
rect 15988 63980 15998 64036
rect 29362 63980 29372 64036
rect 29428 63980 30380 64036
rect 30436 63980 31388 64036
rect 31444 63980 31454 64036
rect 31938 63980 31948 64036
rect 32004 63980 33628 64036
rect 33684 63980 33694 64036
rect 34150 63980 34188 64036
rect 34244 63980 38668 64036
rect 45266 63980 45276 64036
rect 45332 63980 47068 64036
rect 47124 63980 47134 64036
rect 47282 63980 47292 64036
rect 47348 63980 47628 64036
rect 47684 63980 47694 64036
rect 48178 63980 48188 64036
rect 48244 63980 48972 64036
rect 49028 63980 49038 64036
rect 11554 63868 11564 63924
rect 11620 63868 11900 63924
rect 11956 63868 12572 63924
rect 12628 63868 12638 63924
rect 13010 63868 13020 63924
rect 13076 63868 13692 63924
rect 13748 63868 13758 63924
rect 16594 63868 16604 63924
rect 16660 63868 17388 63924
rect 17444 63868 17454 63924
rect 26002 63868 26012 63924
rect 26068 63868 27468 63924
rect 27524 63868 27534 63924
rect 31826 63868 31836 63924
rect 31892 63868 33068 63924
rect 33124 63868 33292 63924
rect 33348 63868 33358 63924
rect 40674 63868 40684 63924
rect 40740 63868 41356 63924
rect 41412 63868 41422 63924
rect 43586 63868 43596 63924
rect 43652 63868 48748 63924
rect 48804 63868 49420 63924
rect 49476 63868 49486 63924
rect 10546 63756 10556 63812
rect 10612 63756 12460 63812
rect 12516 63756 12526 63812
rect 13458 63756 13468 63812
rect 13524 63756 14700 63812
rect 14756 63756 15260 63812
rect 15316 63756 15326 63812
rect 22642 63756 22652 63812
rect 22708 63756 24332 63812
rect 24388 63756 24398 63812
rect 25554 63756 25564 63812
rect 25620 63756 25900 63812
rect 25956 63756 25966 63812
rect 28130 63756 28140 63812
rect 28196 63756 29484 63812
rect 29540 63756 29550 63812
rect 34514 63756 34524 63812
rect 34580 63756 37100 63812
rect 37156 63756 37166 63812
rect 38210 63756 38220 63812
rect 38276 63756 38780 63812
rect 38836 63756 38846 63812
rect 39004 63756 40796 63812
rect 40852 63756 41468 63812
rect 41524 63756 41534 63812
rect 39004 63700 39060 63756
rect 23314 63644 23324 63700
rect 23380 63644 25116 63700
rect 25172 63644 25182 63700
rect 38882 63644 38892 63700
rect 38948 63644 39060 63700
rect 40338 63644 40348 63700
rect 40404 63644 41916 63700
rect 41972 63644 41982 63700
rect 4466 63476 4476 63532
rect 4532 63476 4580 63532
rect 4636 63476 4684 63532
rect 4740 63476 4750 63532
rect 35186 63476 35196 63532
rect 35252 63476 35300 63532
rect 35356 63476 35404 63532
rect 35460 63476 35470 63532
rect 22418 63420 22428 63476
rect 22484 63420 22764 63476
rect 22820 63420 22830 63476
rect 37090 63420 37100 63476
rect 37156 63420 39788 63476
rect 39844 63420 40012 63476
rect 40068 63420 40078 63476
rect 48066 63420 48076 63476
rect 48132 63420 48860 63476
rect 48916 63420 48926 63476
rect 11442 63308 11452 63364
rect 11508 63308 12572 63364
rect 12628 63308 12638 63364
rect 22194 63308 22204 63364
rect 22260 63308 22876 63364
rect 22932 63308 22942 63364
rect 25218 63308 25228 63364
rect 25284 63308 25564 63364
rect 25620 63308 25630 63364
rect 36082 63308 36092 63364
rect 36148 63308 37884 63364
rect 37940 63308 37950 63364
rect 42690 63308 42700 63364
rect 42756 63308 45724 63364
rect 45780 63308 45790 63364
rect 28802 63196 28812 63252
rect 28868 63196 31164 63252
rect 31220 63196 31230 63252
rect 35746 63196 35756 63252
rect 35812 63196 38108 63252
rect 38164 63196 38174 63252
rect 39106 63196 39116 63252
rect 39172 63196 40236 63252
rect 40292 63196 41692 63252
rect 41748 63196 41758 63252
rect 17490 63084 17500 63140
rect 17556 63084 18732 63140
rect 18788 63084 18798 63140
rect 19730 63084 19740 63140
rect 19796 63084 21308 63140
rect 21364 63084 23380 63140
rect 23538 63084 23548 63140
rect 23604 63084 24332 63140
rect 24388 63084 24398 63140
rect 37202 63084 37212 63140
rect 37268 63084 37884 63140
rect 37940 63084 38220 63140
rect 38276 63084 38286 63140
rect 23324 63028 23380 63084
rect 21634 62972 21644 63028
rect 21700 62972 23100 63028
rect 23156 62972 23166 63028
rect 23324 62972 27132 63028
rect 27188 62972 27198 63028
rect 30034 62972 30044 63028
rect 30100 62972 32396 63028
rect 32452 62972 32462 63028
rect 43138 62972 43148 63028
rect 43204 62972 45388 63028
rect 45444 62972 45454 63028
rect 47842 62972 47852 63028
rect 47908 62972 48972 63028
rect 49028 62972 49038 63028
rect 20178 62860 20188 62916
rect 20244 62860 21308 62916
rect 21364 62860 21374 62916
rect 22306 62860 22316 62916
rect 22372 62860 24220 62916
rect 24276 62860 24286 62916
rect 24770 62860 24780 62916
rect 24836 62860 26012 62916
rect 26068 62860 26078 62916
rect 34290 62860 34300 62916
rect 34356 62860 35196 62916
rect 35252 62860 35262 62916
rect 35634 62860 35644 62916
rect 35700 62860 36876 62916
rect 36932 62860 36942 62916
rect 38612 62860 38892 62916
rect 38948 62860 38958 62916
rect 42914 62860 42924 62916
rect 42980 62860 43596 62916
rect 43652 62860 44044 62916
rect 44100 62860 44110 62916
rect 44258 62860 44268 62916
rect 44324 62860 44362 62916
rect 22082 62748 22092 62804
rect 22148 62748 22764 62804
rect 22820 62748 22830 62804
rect 19826 62692 19836 62748
rect 19892 62692 19940 62748
rect 19996 62692 20044 62748
rect 20100 62692 20110 62748
rect 38612 62692 38668 62860
rect 40450 62748 40460 62804
rect 40516 62748 41020 62804
rect 41076 62748 41086 62804
rect 50546 62692 50556 62748
rect 50612 62692 50660 62748
rect 50716 62692 50764 62748
rect 50820 62692 50830 62748
rect 33058 62636 33068 62692
rect 33124 62636 35644 62692
rect 35700 62636 35710 62692
rect 37090 62636 37100 62692
rect 37156 62636 38444 62692
rect 38500 62636 38668 62692
rect 40114 62636 40124 62692
rect 40180 62636 41692 62692
rect 41748 62636 41758 62692
rect 11442 62524 11452 62580
rect 11508 62524 11676 62580
rect 11732 62524 12908 62580
rect 12964 62524 12974 62580
rect 17938 62524 17948 62580
rect 18004 62524 18508 62580
rect 18564 62524 23660 62580
rect 23716 62524 23726 62580
rect 34738 62524 34748 62580
rect 34804 62524 36540 62580
rect 36596 62524 38556 62580
rect 38612 62524 38622 62580
rect 40002 62524 40012 62580
rect 40068 62524 41132 62580
rect 41188 62524 41198 62580
rect 43222 62524 43260 62580
rect 43316 62524 44604 62580
rect 44660 62524 44670 62580
rect 33506 62412 33516 62468
rect 33572 62412 36092 62468
rect 36148 62412 36158 62468
rect 38612 62412 39452 62468
rect 39508 62412 41356 62468
rect 41412 62412 41422 62468
rect 43362 62412 43372 62468
rect 43428 62412 44156 62468
rect 44212 62412 44222 62468
rect 23090 62300 23100 62356
rect 23156 62300 26908 62356
rect 28466 62300 28476 62356
rect 28532 62300 29484 62356
rect 29540 62300 29550 62356
rect 31154 62300 31164 62356
rect 31220 62300 32564 62356
rect 33170 62300 33180 62356
rect 33236 62300 33852 62356
rect 33908 62300 35196 62356
rect 35252 62300 35262 62356
rect 26852 62244 26908 62300
rect 32508 62244 32564 62300
rect 38612 62244 38668 62412
rect 39778 62300 39788 62356
rect 39844 62300 40908 62356
rect 40964 62300 40974 62356
rect 41234 62300 41244 62356
rect 41300 62300 42812 62356
rect 42868 62300 42878 62356
rect 9986 62188 9996 62244
rect 10052 62188 12460 62244
rect 12516 62188 13020 62244
rect 13076 62188 13086 62244
rect 15026 62188 15036 62244
rect 15092 62188 15932 62244
rect 15988 62188 15998 62244
rect 26852 62188 30044 62244
rect 30100 62188 30110 62244
rect 31042 62188 31052 62244
rect 31108 62188 31612 62244
rect 31668 62188 32284 62244
rect 32340 62188 32350 62244
rect 32508 62188 32844 62244
rect 32900 62188 38668 62244
rect 39890 62188 39900 62244
rect 39956 62188 40796 62244
rect 40852 62188 40862 62244
rect 47394 62188 47404 62244
rect 47460 62188 50764 62244
rect 50820 62188 50830 62244
rect 11890 62076 11900 62132
rect 11956 62076 11966 62132
rect 26562 62076 26572 62132
rect 26628 62076 28700 62132
rect 28756 62076 28766 62132
rect 29708 62076 30716 62132
rect 30772 62076 30940 62132
rect 30996 62076 31006 62132
rect 32498 62076 32508 62132
rect 32564 62076 38668 62132
rect 39974 62076 40012 62132
rect 40068 62076 40078 62132
rect 4466 61908 4476 61964
rect 4532 61908 4580 61964
rect 4636 61908 4684 61964
rect 4740 61908 4750 61964
rect 11900 61572 11956 62076
rect 26002 61964 26012 62020
rect 26068 61964 27468 62020
rect 27524 61964 27534 62020
rect 27906 61964 27916 62020
rect 27972 61964 29260 62020
rect 29316 61964 29326 62020
rect 29708 61908 29764 62076
rect 38612 62020 38668 62076
rect 29922 61964 29932 62020
rect 29988 61964 30268 62020
rect 30324 61964 30828 62020
rect 30884 61964 30894 62020
rect 34150 61964 34188 62020
rect 34244 61964 34254 62020
rect 38612 61964 40908 62020
rect 40964 61964 40974 62020
rect 35186 61908 35196 61964
rect 35252 61908 35300 61964
rect 35356 61908 35404 61964
rect 35460 61908 35470 61964
rect 27570 61852 27580 61908
rect 27636 61852 29764 61908
rect 24210 61740 24220 61796
rect 24276 61740 25340 61796
rect 25396 61740 25406 61796
rect 28242 61740 28252 61796
rect 28308 61740 29036 61796
rect 29092 61740 29102 61796
rect 32722 61740 32732 61796
rect 32788 61740 34748 61796
rect 34804 61740 34814 61796
rect 41906 61740 41916 61796
rect 41972 61740 42140 61796
rect 42196 61740 42206 61796
rect 42354 61740 42364 61796
rect 42420 61740 43596 61796
rect 43652 61740 43662 61796
rect 40562 61628 40572 61684
rect 40628 61628 41356 61684
rect 41412 61628 41422 61684
rect 41682 61628 41692 61684
rect 41748 61628 42252 61684
rect 42308 61628 42318 61684
rect 44716 61628 49364 61684
rect 44716 61572 44772 61628
rect 10658 61516 10668 61572
rect 10724 61516 11900 61572
rect 11956 61516 12572 61572
rect 12628 61516 12638 61572
rect 17714 61516 17724 61572
rect 17780 61516 21308 61572
rect 21364 61516 21374 61572
rect 22418 61516 22428 61572
rect 22484 61516 30604 61572
rect 30660 61516 30670 61572
rect 31378 61516 31388 61572
rect 31444 61516 32172 61572
rect 32228 61516 32238 61572
rect 37548 61516 44772 61572
rect 44930 61516 44940 61572
rect 44996 61516 46396 61572
rect 46452 61516 47516 61572
rect 47572 61516 49084 61572
rect 49140 61516 49150 61572
rect 22194 61404 22204 61460
rect 22260 61404 29260 61460
rect 29316 61404 29326 61460
rect 29586 61404 29596 61460
rect 29652 61404 31500 61460
rect 31556 61404 32508 61460
rect 32564 61404 33180 61460
rect 33236 61404 33246 61460
rect 37548 61348 37604 61516
rect 41794 61404 41804 61460
rect 41860 61404 42700 61460
rect 42756 61404 42766 61460
rect 44380 61404 46172 61460
rect 46228 61404 46238 61460
rect 44380 61348 44436 61404
rect 49308 61348 49364 61628
rect 50194 61516 50204 61572
rect 50260 61516 50876 61572
rect 50932 61516 50942 61572
rect 10322 61292 10332 61348
rect 10388 61292 11788 61348
rect 11844 61292 11854 61348
rect 12898 61292 12908 61348
rect 12964 61292 14476 61348
rect 14532 61292 14542 61348
rect 18274 61292 18284 61348
rect 18340 61292 18844 61348
rect 18900 61292 18910 61348
rect 26898 61292 26908 61348
rect 26964 61292 28252 61348
rect 28308 61292 28318 61348
rect 28466 61292 28476 61348
rect 28532 61292 28570 61348
rect 33954 61292 33964 61348
rect 34020 61292 36204 61348
rect 36260 61292 37548 61348
rect 37604 61292 37614 61348
rect 38612 61292 44380 61348
rect 44436 61292 44446 61348
rect 45378 61292 45388 61348
rect 45444 61292 47404 61348
rect 47460 61292 47470 61348
rect 49186 61292 49196 61348
rect 49252 61292 50316 61348
rect 50372 61292 50382 61348
rect 38612 61236 38668 61292
rect 18946 61180 18956 61236
rect 19012 61180 19022 61236
rect 31714 61180 31724 61236
rect 31780 61180 38668 61236
rect 40898 61180 40908 61236
rect 40964 61180 41580 61236
rect 41636 61180 41646 61236
rect 42242 61180 42252 61236
rect 42308 61180 42588 61236
rect 42644 61180 43148 61236
rect 43204 61180 43214 61236
rect 18956 61012 19012 61180
rect 19826 61124 19836 61180
rect 19892 61124 19940 61180
rect 19996 61124 20044 61180
rect 20100 61124 20110 61180
rect 50546 61124 50556 61180
rect 50612 61124 50660 61180
rect 50716 61124 50764 61180
rect 50820 61124 50830 61180
rect 22978 61068 22988 61124
rect 23044 61068 23884 61124
rect 23940 61068 25676 61124
rect 25732 61068 26348 61124
rect 26404 61068 26414 61124
rect 31500 61068 33964 61124
rect 34020 61068 34030 61124
rect 42102 61068 42140 61124
rect 42196 61068 42206 61124
rect 31500 61012 31556 61068
rect 10882 60956 10892 61012
rect 10948 60956 11676 61012
rect 11732 60956 12796 61012
rect 12852 60956 12862 61012
rect 18956 60956 19740 61012
rect 19796 60956 19806 61012
rect 20850 60956 20860 61012
rect 20916 60956 21756 61012
rect 21812 60956 21822 61012
rect 23090 60956 23100 61012
rect 23156 60956 23772 61012
rect 23828 60956 23838 61012
rect 26562 60956 26572 61012
rect 26628 60956 28924 61012
rect 28980 60956 28990 61012
rect 30594 60956 30604 61012
rect 30660 60956 31500 61012
rect 31556 60956 31566 61012
rect 31836 60956 32732 61012
rect 32788 60956 32798 61012
rect 31836 60900 31892 60956
rect 16146 60844 16156 60900
rect 16212 60844 17388 60900
rect 17444 60844 17454 60900
rect 22642 60844 22652 60900
rect 22708 60844 23044 60900
rect 23202 60844 23212 60900
rect 23268 60844 23996 60900
rect 24052 60844 25340 60900
rect 25396 60844 25406 60900
rect 25564 60844 31892 60900
rect 32050 60844 32060 60900
rect 32116 60844 33740 60900
rect 33796 60844 33806 60900
rect 22988 60788 23044 60844
rect 25564 60788 25620 60844
rect 13122 60732 13132 60788
rect 13188 60732 13580 60788
rect 13636 60732 13916 60788
rect 13972 60732 13982 60788
rect 16034 60732 16044 60788
rect 16100 60732 16110 60788
rect 16594 60732 16604 60788
rect 16660 60732 17948 60788
rect 18004 60732 18014 60788
rect 19506 60732 19516 60788
rect 19572 60732 19964 60788
rect 20020 60732 20030 60788
rect 20132 60732 20300 60788
rect 20356 60732 20366 60788
rect 22082 60732 22092 60788
rect 22148 60732 22764 60788
rect 22820 60732 22830 60788
rect 22988 60732 23100 60788
rect 23156 60732 25620 60788
rect 26562 60732 26572 60788
rect 26628 60732 28700 60788
rect 28756 60732 28766 60788
rect 29362 60732 29372 60788
rect 29428 60732 29820 60788
rect 29876 60732 30156 60788
rect 30212 60732 31052 60788
rect 31108 60732 31118 60788
rect 32498 60732 32508 60788
rect 32564 60732 33628 60788
rect 33684 60732 33694 60788
rect 37426 60732 37436 60788
rect 37492 60732 39116 60788
rect 39172 60732 39182 60788
rect 46162 60732 46172 60788
rect 46228 60732 47180 60788
rect 47236 60732 47246 60788
rect 16044 60676 16100 60732
rect 20132 60676 20188 60732
rect 29596 60676 29652 60732
rect 16044 60620 16828 60676
rect 16884 60620 17836 60676
rect 17892 60620 17902 60676
rect 19394 60620 19404 60676
rect 19460 60620 20188 60676
rect 27346 60620 27356 60676
rect 27412 60620 28588 60676
rect 28644 60620 28654 60676
rect 29586 60620 29596 60676
rect 29652 60620 29662 60676
rect 32834 60620 32844 60676
rect 32900 60620 34860 60676
rect 34916 60620 34926 60676
rect 36418 60620 36428 60676
rect 36484 60620 39004 60676
rect 39060 60620 39070 60676
rect 39330 60620 39340 60676
rect 39396 60620 40348 60676
rect 40404 60620 40414 60676
rect 47394 60620 47404 60676
rect 47460 60620 48860 60676
rect 48916 60620 49196 60676
rect 49252 60620 49262 60676
rect 15698 60508 15708 60564
rect 15764 60508 17388 60564
rect 17444 60508 17454 60564
rect 25218 60508 25228 60564
rect 25284 60508 26236 60564
rect 26292 60508 26908 60564
rect 26964 60508 26974 60564
rect 28242 60508 28252 60564
rect 28308 60508 29036 60564
rect 29092 60508 29102 60564
rect 35298 60508 35308 60564
rect 35364 60508 35588 60564
rect 41010 60508 41020 60564
rect 41076 60508 46396 60564
rect 46452 60508 46844 60564
rect 46900 60508 46910 60564
rect 20626 60396 20636 60452
rect 20692 60396 21532 60452
rect 21588 60396 21598 60452
rect 4466 60340 4476 60396
rect 4532 60340 4580 60396
rect 4636 60340 4684 60396
rect 4740 60340 4750 60396
rect 35186 60340 35196 60396
rect 35252 60340 35300 60396
rect 35356 60340 35404 60396
rect 35460 60340 35470 60396
rect 26002 60284 26012 60340
rect 26068 60284 27020 60340
rect 27076 60284 27086 60340
rect 35532 60228 35588 60508
rect 36978 60396 36988 60452
rect 37044 60396 37324 60452
rect 37380 60396 37390 60452
rect 39330 60396 39340 60452
rect 39396 60396 40012 60452
rect 40068 60396 40078 60452
rect 42242 60396 42252 60452
rect 42308 60396 43596 60452
rect 43652 60396 43662 60452
rect 45042 60396 45052 60452
rect 45108 60396 48076 60452
rect 48132 60396 49084 60452
rect 49140 60396 49150 60452
rect 35970 60284 35980 60340
rect 36036 60284 45948 60340
rect 46004 60284 46014 60340
rect 26226 60172 26236 60228
rect 26292 60172 26796 60228
rect 26852 60172 28028 60228
rect 28084 60172 28094 60228
rect 35410 60172 35420 60228
rect 35476 60172 35588 60228
rect 36082 60172 36092 60228
rect 36148 60172 40012 60228
rect 40068 60172 41020 60228
rect 41076 60172 41086 60228
rect 21522 60060 21532 60116
rect 21588 60060 22204 60116
rect 22260 60060 22270 60116
rect 31042 60060 31052 60116
rect 31108 60060 42084 60116
rect 42028 60004 42084 60060
rect 19618 59948 19628 60004
rect 19684 59948 20524 60004
rect 20580 59948 21644 60004
rect 21700 59948 21710 60004
rect 23874 59948 23884 60004
rect 23940 59948 24892 60004
rect 24948 59948 29148 60004
rect 29204 59948 29214 60004
rect 32274 59948 32284 60004
rect 32340 59948 33068 60004
rect 33124 59948 33134 60004
rect 34626 59948 34636 60004
rect 34692 59948 35532 60004
rect 35588 59948 35598 60004
rect 38434 59948 38444 60004
rect 38500 59948 39004 60004
rect 39060 59948 39788 60004
rect 39844 59948 39854 60004
rect 42028 59948 45780 60004
rect 46722 59948 46732 60004
rect 46788 59948 47516 60004
rect 47572 59948 47582 60004
rect 16482 59836 16492 59892
rect 16548 59836 16828 59892
rect 16884 59836 16894 59892
rect 19170 59836 19180 59892
rect 19236 59836 20748 59892
rect 20804 59836 20814 59892
rect 21410 59836 21420 59892
rect 21476 59836 26012 59892
rect 26068 59836 26078 59892
rect 32386 59836 32396 59892
rect 32452 59836 32462 59892
rect 38546 59836 38556 59892
rect 38612 59836 41580 59892
rect 41636 59836 41646 59892
rect 42028 59836 42588 59892
rect 42644 59836 42654 59892
rect 43586 59836 43596 59892
rect 43652 59836 45500 59892
rect 45556 59836 45566 59892
rect 32396 59780 32452 59836
rect 14690 59724 14700 59780
rect 14756 59724 15708 59780
rect 15764 59724 15774 59780
rect 19842 59724 19852 59780
rect 19908 59724 20244 59780
rect 22642 59724 22652 59780
rect 22708 59724 23996 59780
rect 24052 59724 24332 59780
rect 24388 59724 24398 59780
rect 32396 59724 34188 59780
rect 34244 59724 34254 59780
rect 35522 59724 35532 59780
rect 35588 59724 37100 59780
rect 37156 59724 38220 59780
rect 38276 59724 38286 59780
rect 39554 59724 39564 59780
rect 39620 59724 40012 59780
rect 40068 59724 41020 59780
rect 41076 59724 41468 59780
rect 41524 59724 41534 59780
rect 19826 59556 19836 59612
rect 19892 59556 19940 59612
rect 19996 59556 20044 59612
rect 20100 59556 20110 59612
rect 20188 59332 20244 59724
rect 42028 59668 42084 59836
rect 45724 59780 45780 59948
rect 46946 59836 46956 59892
rect 47012 59836 47404 59892
rect 47460 59836 47470 59892
rect 42242 59724 42252 59780
rect 42308 59724 43484 59780
rect 43540 59724 43550 59780
rect 45724 59724 52108 59780
rect 52164 59724 52174 59780
rect 32162 59612 32172 59668
rect 32228 59612 34860 59668
rect 34916 59612 34926 59668
rect 35074 59612 35084 59668
rect 35140 59612 36092 59668
rect 36148 59612 36158 59668
rect 39414 59612 39452 59668
rect 39508 59612 39518 59668
rect 42028 59612 42364 59668
rect 42420 59612 42430 59668
rect 43138 59612 43148 59668
rect 43204 59612 45612 59668
rect 45668 59612 46060 59668
rect 46116 59612 46126 59668
rect 50546 59556 50556 59612
rect 50612 59556 50660 59612
rect 50716 59556 50764 59612
rect 50820 59556 50830 59612
rect 21494 59500 21532 59556
rect 21588 59500 21598 59556
rect 22418 59500 22428 59556
rect 22484 59500 22988 59556
rect 23044 59500 23054 59556
rect 23772 59500 25452 59556
rect 25508 59500 33292 59556
rect 33348 59500 33358 59556
rect 23772 59332 23828 59500
rect 23986 59388 23996 59444
rect 24052 59388 24556 59444
rect 24612 59388 26460 59444
rect 26516 59388 26526 59444
rect 27122 59388 27132 59444
rect 27188 59388 27692 59444
rect 27748 59388 27758 59444
rect 39302 59388 39340 59444
rect 39396 59388 39406 59444
rect 39554 59388 39564 59444
rect 39620 59388 40460 59444
rect 40516 59388 40526 59444
rect 42578 59388 42588 59444
rect 42644 59388 42924 59444
rect 42980 59388 42990 59444
rect 49858 59388 49868 59444
rect 49924 59388 50316 59444
rect 50372 59388 50382 59444
rect 19730 59276 19740 59332
rect 19796 59276 23828 59332
rect 25778 59276 25788 59332
rect 25844 59276 26236 59332
rect 26292 59276 26908 59332
rect 26964 59276 26974 59332
rect 27794 59276 27804 59332
rect 27860 59276 28476 59332
rect 28532 59276 28542 59332
rect 32610 59276 32620 59332
rect 32676 59276 33516 59332
rect 33572 59276 36988 59332
rect 37044 59276 38444 59332
rect 38500 59276 47964 59332
rect 48020 59276 48748 59332
rect 48804 59276 49756 59332
rect 49812 59276 49822 59332
rect 20066 59164 20076 59220
rect 20132 59164 20748 59220
rect 20804 59164 21756 59220
rect 21812 59164 21822 59220
rect 22754 59164 22764 59220
rect 22820 59164 24444 59220
rect 24500 59164 24510 59220
rect 26002 59164 26012 59220
rect 26068 59164 27132 59220
rect 27188 59164 27198 59220
rect 38658 59164 38668 59220
rect 38724 59164 39116 59220
rect 39172 59164 40012 59220
rect 40068 59164 40078 59220
rect 43250 59164 43260 59220
rect 43316 59164 43708 59220
rect 43764 59164 44268 59220
rect 44324 59164 44334 59220
rect 46946 59164 46956 59220
rect 47012 59164 47292 59220
rect 47348 59164 47358 59220
rect 47842 59164 47852 59220
rect 47908 59164 48972 59220
rect 49028 59164 49868 59220
rect 49924 59164 49934 59220
rect 16818 59052 16828 59108
rect 16884 59052 17164 59108
rect 17220 59052 17230 59108
rect 22978 59052 22988 59108
rect 23044 59052 26236 59108
rect 26292 59052 26302 59108
rect 30258 59052 30268 59108
rect 30324 59052 35756 59108
rect 35812 59052 35822 59108
rect 39890 59052 39900 59108
rect 39956 59052 39966 59108
rect 42578 59052 42588 59108
rect 42644 59052 43148 59108
rect 43204 59052 43214 59108
rect 43474 59052 43484 59108
rect 43540 59052 45500 59108
rect 45556 59052 45566 59108
rect 45714 59052 45724 59108
rect 45780 59052 46060 59108
rect 46116 59052 46126 59108
rect 23314 58940 23324 58996
rect 23380 58940 24556 58996
rect 24612 58940 24622 58996
rect 34850 58940 34860 58996
rect 34916 58940 35868 58996
rect 35924 58940 36876 58996
rect 36932 58940 36942 58996
rect 18722 58828 18732 58884
rect 18788 58828 19180 58884
rect 19236 58828 19246 58884
rect 22866 58828 22876 58884
rect 22932 58828 25228 58884
rect 25284 58828 25294 58884
rect 32834 58828 32844 58884
rect 32900 58828 33180 58884
rect 33236 58828 33246 58884
rect 33506 58828 33516 58884
rect 33572 58828 34748 58884
rect 34804 58828 34814 58884
rect 36306 58828 36316 58884
rect 36372 58828 37100 58884
rect 37156 58828 37166 58884
rect 4466 58772 4476 58828
rect 4532 58772 4580 58828
rect 4636 58772 4684 58828
rect 4740 58772 4750 58828
rect 35186 58772 35196 58828
rect 35252 58772 35300 58828
rect 35356 58772 35404 58828
rect 35460 58772 35470 58828
rect 23762 58716 23772 58772
rect 23828 58716 24220 58772
rect 24276 58716 24668 58772
rect 24724 58716 26684 58772
rect 26740 58716 26750 58772
rect 27234 58716 27244 58772
rect 27300 58716 27916 58772
rect 27972 58716 27982 58772
rect 34178 58716 34188 58772
rect 34244 58716 34636 58772
rect 34692 58716 34702 58772
rect 39900 58660 39956 59052
rect 41244 58940 43260 58996
rect 43316 58940 43326 58996
rect 43922 58940 43932 58996
rect 43988 58940 44268 58996
rect 44324 58940 44334 58996
rect 45266 58940 45276 58996
rect 45332 58940 52332 58996
rect 52388 58940 52398 58996
rect 41244 58828 41300 58940
rect 42550 58828 42588 58884
rect 42644 58828 42654 58884
rect 44930 58828 44940 58884
rect 44996 58828 46172 58884
rect 46228 58828 46238 58884
rect 41234 58772 41244 58828
rect 41300 58772 41310 58828
rect 43810 58716 43820 58772
rect 43876 58716 45164 58772
rect 45220 58716 45230 58772
rect 32722 58604 32732 58660
rect 32788 58604 33796 58660
rect 36418 58604 36428 58660
rect 36484 58604 37660 58660
rect 37716 58604 37726 58660
rect 38612 58604 39956 58660
rect 44034 58604 44044 58660
rect 44100 58604 45276 58660
rect 45332 58604 45342 58660
rect 45910 58604 45948 58660
rect 46004 58604 46014 58660
rect 33740 58548 33796 58604
rect 38612 58548 38668 58604
rect 6178 58492 6188 58548
rect 6244 58492 9660 58548
rect 9716 58492 9726 58548
rect 13010 58492 13020 58548
rect 13076 58492 14924 58548
rect 14980 58492 14990 58548
rect 21522 58492 21532 58548
rect 21588 58492 21980 58548
rect 22036 58492 30940 58548
rect 30996 58492 31006 58548
rect 32396 58492 33404 58548
rect 33460 58492 33470 58548
rect 33730 58492 33740 58548
rect 33796 58492 34188 58548
rect 34244 58492 34254 58548
rect 35186 58492 35196 58548
rect 35252 58492 38668 58548
rect 39554 58492 39564 58548
rect 39620 58492 41468 58548
rect 41524 58492 41534 58548
rect 43474 58492 43484 58548
rect 43540 58492 43764 58548
rect 32396 58436 32452 58492
rect 13794 58380 13804 58436
rect 13860 58380 14812 58436
rect 14868 58380 14878 58436
rect 15474 58380 15484 58436
rect 15540 58380 17612 58436
rect 17668 58380 17678 58436
rect 19842 58380 19852 58436
rect 19908 58380 20636 58436
rect 20692 58380 20702 58436
rect 24658 58380 24668 58436
rect 24724 58380 26908 58436
rect 26964 58380 26974 58436
rect 28018 58380 28028 58436
rect 28084 58380 28812 58436
rect 28868 58380 29820 58436
rect 29876 58380 29886 58436
rect 30146 58380 30156 58436
rect 30212 58380 32396 58436
rect 32452 58380 32462 58436
rect 33170 58380 33180 58436
rect 33236 58380 34076 58436
rect 34132 58380 34142 58436
rect 34626 58380 34636 58436
rect 34692 58380 38220 58436
rect 38276 58380 38286 58436
rect 43708 58324 43764 58492
rect 16482 58268 16492 58324
rect 16548 58268 17500 58324
rect 17556 58268 17566 58324
rect 20738 58268 20748 58324
rect 20804 58268 21532 58324
rect 21588 58268 21598 58324
rect 28130 58268 28140 58324
rect 28196 58268 29932 58324
rect 29988 58268 29998 58324
rect 34514 58268 34524 58324
rect 34580 58268 35532 58324
rect 35588 58268 36092 58324
rect 36148 58268 36158 58324
rect 43698 58268 43708 58324
rect 43764 58268 43774 58324
rect 46722 58268 46732 58324
rect 46788 58268 47516 58324
rect 47572 58268 47740 58324
rect 47796 58268 47806 58324
rect 14354 58156 14364 58212
rect 14420 58156 15148 58212
rect 17266 58156 17276 58212
rect 17332 58156 17836 58212
rect 17892 58156 17902 58212
rect 19170 58156 19180 58212
rect 19236 58156 20300 58212
rect 20356 58156 20366 58212
rect 26450 58156 26460 58212
rect 26516 58156 28252 58212
rect 28308 58156 28318 58212
rect 31490 58156 31500 58212
rect 31556 58156 31948 58212
rect 32004 58156 32014 58212
rect 34290 58156 34300 58212
rect 34356 58156 35196 58212
rect 35252 58156 35262 58212
rect 40450 58156 40460 58212
rect 40516 58156 41244 58212
rect 41300 58156 41310 58212
rect 44482 58156 44492 58212
rect 44548 58156 44940 58212
rect 44996 58156 45006 58212
rect 45154 58156 45164 58212
rect 45220 58156 45836 58212
rect 45892 58156 45902 58212
rect 47282 58156 47292 58212
rect 47348 58156 47628 58212
rect 47684 58156 47694 58212
rect 15092 58100 15148 58156
rect 44716 58100 44772 58156
rect 15092 58044 15260 58100
rect 15316 58044 16044 58100
rect 16100 58044 16110 58100
rect 20178 58044 20188 58100
rect 20244 58044 21420 58100
rect 21476 58044 21486 58100
rect 34850 58044 34860 58100
rect 34916 58044 35644 58100
rect 35700 58044 35710 58100
rect 41122 58044 41132 58100
rect 41188 58044 41580 58100
rect 41636 58044 42028 58100
rect 42084 58044 42094 58100
rect 44706 58044 44716 58100
rect 44772 58044 44782 58100
rect 44930 58044 44940 58100
rect 44996 58044 45276 58100
rect 45332 58044 45342 58100
rect 46050 58044 46060 58100
rect 46116 58044 46126 58100
rect 47292 58044 47404 58100
rect 47460 58044 47470 58100
rect 19826 57988 19836 58044
rect 19892 57988 19940 58044
rect 19996 57988 20044 58044
rect 20100 57988 20110 58044
rect 46060 57988 46116 58044
rect 18610 57932 18620 57988
rect 18676 57932 19404 57988
rect 19460 57932 19470 57988
rect 23202 57932 23212 57988
rect 23268 57932 25340 57988
rect 25396 57932 25676 57988
rect 25732 57932 26908 57988
rect 27906 57932 27916 57988
rect 27972 57932 32956 57988
rect 33012 57932 33022 57988
rect 38210 57932 38220 57988
rect 38276 57932 38780 57988
rect 38836 57932 45388 57988
rect 45444 57932 46116 57988
rect 26852 57876 26908 57932
rect 47292 57876 47348 58044
rect 50546 57988 50556 58044
rect 50612 57988 50660 58044
rect 50716 57988 50764 58044
rect 50820 57988 50830 58044
rect 9538 57820 9548 57876
rect 9604 57820 12236 57876
rect 12292 57820 13468 57876
rect 13524 57820 14924 57876
rect 14980 57820 14990 57876
rect 23762 57820 23772 57876
rect 23828 57820 24556 57876
rect 24612 57820 25788 57876
rect 25844 57820 25854 57876
rect 26852 57820 28364 57876
rect 28420 57820 30828 57876
rect 30884 57820 30894 57876
rect 40562 57820 40572 57876
rect 40628 57820 41916 57876
rect 41972 57820 41982 57876
rect 43474 57820 43484 57876
rect 43540 57820 44940 57876
rect 44996 57820 45006 57876
rect 47282 57820 47292 57876
rect 47348 57820 47358 57876
rect 21074 57708 21084 57764
rect 21140 57708 22428 57764
rect 22484 57708 23996 57764
rect 24052 57708 24062 57764
rect 44818 57708 44828 57764
rect 44884 57708 45276 57764
rect 45332 57708 46228 57764
rect 46172 57652 46228 57708
rect 10434 57596 10444 57652
rect 10500 57596 11340 57652
rect 11396 57596 11406 57652
rect 12786 57596 12796 57652
rect 12852 57596 16940 57652
rect 16996 57596 17006 57652
rect 23426 57596 23436 57652
rect 23492 57596 24108 57652
rect 24164 57596 25228 57652
rect 25284 57596 25294 57652
rect 28578 57596 28588 57652
rect 28644 57596 30940 57652
rect 30996 57596 31006 57652
rect 31826 57596 31836 57652
rect 31892 57596 33516 57652
rect 33572 57596 33582 57652
rect 41346 57596 41356 57652
rect 41412 57596 42252 57652
rect 42308 57596 42318 57652
rect 46162 57596 46172 57652
rect 46228 57596 46238 57652
rect 23100 57484 24892 57540
rect 24948 57484 24958 57540
rect 26852 57484 27244 57540
rect 27300 57484 27310 57540
rect 29810 57484 29820 57540
rect 29876 57484 31276 57540
rect 31332 57484 31342 57540
rect 34066 57484 34076 57540
rect 34132 57484 34636 57540
rect 34692 57484 34702 57540
rect 38770 57484 38780 57540
rect 38836 57484 40348 57540
rect 40404 57484 40414 57540
rect 45602 57484 45612 57540
rect 45668 57484 46060 57540
rect 46116 57484 48188 57540
rect 48244 57484 48860 57540
rect 48916 57484 49308 57540
rect 49364 57484 50092 57540
rect 50148 57484 50158 57540
rect 23100 57428 23156 57484
rect 22978 57372 22988 57428
rect 23044 57372 23156 57428
rect 23650 57372 23660 57428
rect 23716 57372 26124 57428
rect 26180 57372 26190 57428
rect 23538 57260 23548 57316
rect 23604 57260 24892 57316
rect 24948 57260 25452 57316
rect 25508 57260 25518 57316
rect 4466 57204 4476 57260
rect 4532 57204 4580 57260
rect 4636 57204 4684 57260
rect 4740 57204 4750 57260
rect 26852 57204 26908 57484
rect 38994 57372 39004 57428
rect 39060 57372 39452 57428
rect 39508 57372 40572 57428
rect 40628 57372 46508 57428
rect 46564 57372 46574 57428
rect 47170 57260 47180 57316
rect 47236 57260 48076 57316
rect 48132 57260 49756 57316
rect 49812 57260 49822 57316
rect 35186 57204 35196 57260
rect 35252 57204 35300 57260
rect 35356 57204 35404 57260
rect 35460 57204 35470 57260
rect 21858 57148 21868 57204
rect 21924 57148 25676 57204
rect 25732 57148 26572 57204
rect 26628 57148 26908 57204
rect 39106 57148 39116 57204
rect 39172 57148 39788 57204
rect 39844 57148 44940 57204
rect 44996 57148 45006 57204
rect 47506 57148 47516 57204
rect 47572 57148 47582 57204
rect 47516 57092 47572 57148
rect 18498 57036 18508 57092
rect 18564 57036 19628 57092
rect 19684 57036 20300 57092
rect 20356 57036 20366 57092
rect 20626 57036 20636 57092
rect 20692 57036 21644 57092
rect 21700 57036 22428 57092
rect 22484 57036 22494 57092
rect 23874 57036 23884 57092
rect 23940 57036 24668 57092
rect 24724 57036 30156 57092
rect 30212 57036 30222 57092
rect 40226 57036 40236 57092
rect 40292 57036 42252 57092
rect 42308 57036 42318 57092
rect 46722 57036 46732 57092
rect 46788 57036 49420 57092
rect 49476 57036 49486 57092
rect 6850 56924 6860 56980
rect 6916 56924 8988 56980
rect 9044 56924 9054 56980
rect 19058 56924 19068 56980
rect 19124 56924 29148 56980
rect 29204 56924 30380 56980
rect 30436 56924 30446 56980
rect 33926 56924 33964 56980
rect 34020 56924 34030 56980
rect 39330 56924 39340 56980
rect 39396 56924 40124 56980
rect 40180 56924 52220 56980
rect 52276 56924 52286 56980
rect 19506 56812 19516 56868
rect 19572 56812 21308 56868
rect 21364 56812 21374 56868
rect 21634 56812 21644 56868
rect 21700 56812 22092 56868
rect 22148 56812 22876 56868
rect 22932 56812 24220 56868
rect 24276 56812 24286 56868
rect 31042 56812 31052 56868
rect 31108 56812 34860 56868
rect 34916 56812 34926 56868
rect 9090 56700 9100 56756
rect 9156 56700 10444 56756
rect 10500 56700 10510 56756
rect 13682 56700 13692 56756
rect 13748 56700 15148 56756
rect 15204 56700 15214 56756
rect 18386 56700 18396 56756
rect 18452 56700 19404 56756
rect 19460 56700 19470 56756
rect 21410 56700 21420 56756
rect 21476 56700 21756 56756
rect 21812 56700 21822 56756
rect 22642 56700 22652 56756
rect 22708 56700 23100 56756
rect 23156 56700 24332 56756
rect 24388 56700 24398 56756
rect 8866 56588 8876 56644
rect 8932 56588 9660 56644
rect 9716 56588 10220 56644
rect 10276 56588 10286 56644
rect 14466 56588 14476 56644
rect 14532 56588 15596 56644
rect 15652 56588 15662 56644
rect 24434 56588 24444 56644
rect 24500 56588 25340 56644
rect 25396 56588 25406 56644
rect 31602 56588 31612 56644
rect 31668 56588 32508 56644
rect 32564 56588 33180 56644
rect 33236 56588 33246 56644
rect 34402 56588 34412 56644
rect 34468 56588 34860 56644
rect 34916 56588 34926 56644
rect 37090 56588 37100 56644
rect 37156 56588 37660 56644
rect 37716 56588 37726 56644
rect 38322 56588 38332 56644
rect 38388 56588 40236 56644
rect 40292 56588 40302 56644
rect 41010 56588 41020 56644
rect 41076 56588 46732 56644
rect 46788 56588 46798 56644
rect 23986 56476 23996 56532
rect 24052 56476 32284 56532
rect 32340 56476 33068 56532
rect 33124 56476 37996 56532
rect 38052 56476 38062 56532
rect 44258 56476 44268 56532
rect 44324 56476 44334 56532
rect 19826 56420 19836 56476
rect 19892 56420 19940 56476
rect 19996 56420 20044 56476
rect 20100 56420 20110 56476
rect 9314 56364 9324 56420
rect 9380 56364 10332 56420
rect 10388 56364 10780 56420
rect 10836 56364 10846 56420
rect 18946 56364 18956 56420
rect 19012 56364 19022 56420
rect 6402 56252 6412 56308
rect 6468 56252 7084 56308
rect 7140 56252 7150 56308
rect 15922 56252 15932 56308
rect 15988 56252 17388 56308
rect 17444 56252 17454 56308
rect 15138 56140 15148 56196
rect 15204 56140 16716 56196
rect 16772 56140 16782 56196
rect 6962 56028 6972 56084
rect 7028 56028 8092 56084
rect 8148 56028 8158 56084
rect 9538 56028 9548 56084
rect 9604 56028 10108 56084
rect 10164 56028 10892 56084
rect 10948 56028 10958 56084
rect 18956 55860 19012 56364
rect 44268 56308 44324 56476
rect 50546 56420 50556 56476
rect 50612 56420 50660 56476
rect 50716 56420 50764 56476
rect 50820 56420 50830 56476
rect 45462 56364 45500 56420
rect 45556 56364 46396 56420
rect 46452 56364 46462 56420
rect 24434 56252 24444 56308
rect 24500 56252 25228 56308
rect 25284 56252 25294 56308
rect 43810 56252 43820 56308
rect 43876 56252 45388 56308
rect 45444 56252 45454 56308
rect 47282 56252 47292 56308
rect 47348 56252 48636 56308
rect 48692 56252 49980 56308
rect 50036 56252 50046 56308
rect 31490 56140 31500 56196
rect 31556 56140 31836 56196
rect 31892 56140 31902 56196
rect 34290 56140 34300 56196
rect 34356 56140 39116 56196
rect 39172 56140 39182 56196
rect 42662 56140 42700 56196
rect 42756 56140 42766 56196
rect 44034 56140 44044 56196
rect 44100 56140 47852 56196
rect 47908 56140 48972 56196
rect 49028 56140 49038 56196
rect 20738 56028 20748 56084
rect 20804 56028 22540 56084
rect 22596 56028 23548 56084
rect 23604 56028 23614 56084
rect 32386 56028 32396 56084
rect 32452 56028 33516 56084
rect 33572 56028 33964 56084
rect 34020 56028 34412 56084
rect 34468 56028 34478 56084
rect 42914 56028 42924 56084
rect 42980 56028 43932 56084
rect 43988 56028 44716 56084
rect 44772 56028 44782 56084
rect 46946 56028 46956 56084
rect 47012 56028 47628 56084
rect 47684 56028 47694 56084
rect 48066 56028 48076 56084
rect 48132 56028 48860 56084
rect 48916 56028 48926 56084
rect 27346 55916 27356 55972
rect 27412 55916 28028 55972
rect 28084 55916 28094 55972
rect 40338 55916 40348 55972
rect 40404 55916 42476 55972
rect 42532 55916 42542 55972
rect 6626 55804 6636 55860
rect 6692 55804 7868 55860
rect 7924 55804 7934 55860
rect 18946 55804 18956 55860
rect 19012 55804 19022 55860
rect 4466 55636 4476 55692
rect 4532 55636 4580 55692
rect 4636 55636 4684 55692
rect 4740 55636 4750 55692
rect 35186 55636 35196 55692
rect 35252 55636 35300 55692
rect 35356 55636 35404 55692
rect 35460 55636 35470 55692
rect 18386 55468 18396 55524
rect 18452 55468 21980 55524
rect 22036 55468 22046 55524
rect 27766 55468 27804 55524
rect 27860 55468 27870 55524
rect 30034 55468 30044 55524
rect 30100 55468 32060 55524
rect 32116 55468 32126 55524
rect 36306 55468 36316 55524
rect 36372 55468 36988 55524
rect 37044 55468 37054 55524
rect 43810 55468 43820 55524
rect 43876 55468 45836 55524
rect 45892 55468 45902 55524
rect 13458 55356 13468 55412
rect 13524 55356 15260 55412
rect 15316 55356 15326 55412
rect 20514 55356 20524 55412
rect 20580 55356 21308 55412
rect 21364 55356 21374 55412
rect 25554 55356 25564 55412
rect 25620 55356 26236 55412
rect 26292 55356 27244 55412
rect 27300 55356 27310 55412
rect 28578 55356 28588 55412
rect 28644 55356 29932 55412
rect 29988 55356 29998 55412
rect 30370 55356 30380 55412
rect 30436 55356 33292 55412
rect 33348 55356 33964 55412
rect 34020 55356 38668 55412
rect 38724 55356 38734 55412
rect 39788 55356 42364 55412
rect 42420 55356 43372 55412
rect 43428 55356 43438 55412
rect 39788 55300 39844 55356
rect 18610 55244 18620 55300
rect 18676 55244 20300 55300
rect 20356 55244 20366 55300
rect 20626 55244 20636 55300
rect 20692 55244 22316 55300
rect 22372 55244 22988 55300
rect 23044 55244 23054 55300
rect 26338 55244 26348 55300
rect 26404 55244 30492 55300
rect 30548 55244 34972 55300
rect 35028 55244 35038 55300
rect 38612 55244 39844 55300
rect 40796 55244 41580 55300
rect 41636 55244 42588 55300
rect 42644 55244 42654 55300
rect 38612 55188 38668 55244
rect 10658 55132 10668 55188
rect 10724 55132 11452 55188
rect 11508 55132 11518 55188
rect 19842 55132 19852 55188
rect 19908 55132 20524 55188
rect 20580 55132 20590 55188
rect 25890 55132 25900 55188
rect 25956 55132 25966 55188
rect 28354 55132 28364 55188
rect 28420 55132 30772 55188
rect 34402 55132 34412 55188
rect 34468 55132 38668 55188
rect 25900 55076 25956 55132
rect 30716 55076 30772 55132
rect 17350 55020 17388 55076
rect 17444 55020 18396 55076
rect 18452 55020 18462 55076
rect 19394 55020 19404 55076
rect 19460 55020 20300 55076
rect 20356 55020 20366 55076
rect 25900 55020 27916 55076
rect 27972 55020 29148 55076
rect 29204 55020 29214 55076
rect 30706 55020 30716 55076
rect 30772 55020 31276 55076
rect 31332 55020 33852 55076
rect 33908 55020 33918 55076
rect 35634 55020 35644 55076
rect 35700 55020 35710 55076
rect 35858 55020 35868 55076
rect 35924 55020 37100 55076
rect 37156 55020 37166 55076
rect 35644 54964 35700 55020
rect 40796 54964 40852 55244
rect 41010 55132 41020 55188
rect 41076 55132 42252 55188
rect 42308 55132 42318 55188
rect 41766 55020 41804 55076
rect 41860 55020 41870 55076
rect 42354 55020 42364 55076
rect 42420 55020 43036 55076
rect 43092 55020 43932 55076
rect 43988 55020 43998 55076
rect 49970 55020 49980 55076
rect 50036 55020 50876 55076
rect 50932 55020 50942 55076
rect 25330 54908 25340 54964
rect 25396 54908 26460 54964
rect 26516 54908 26526 54964
rect 29810 54908 29820 54964
rect 29876 54908 40852 54964
rect 41804 54964 41860 55020
rect 41804 54908 42924 54964
rect 42980 54908 42990 54964
rect 19826 54852 19836 54908
rect 19892 54852 19940 54908
rect 19996 54852 20044 54908
rect 20100 54852 20110 54908
rect 50546 54852 50556 54908
rect 50612 54852 50660 54908
rect 50716 54852 50764 54908
rect 50820 54852 50830 54908
rect 23986 54796 23996 54852
rect 24052 54796 27020 54852
rect 27076 54796 27086 54852
rect 29922 54796 29932 54852
rect 29988 54796 31164 54852
rect 31220 54796 31230 54852
rect 34066 54796 34076 54852
rect 34132 54796 34412 54852
rect 34468 54796 34478 54852
rect 7634 54684 7644 54740
rect 7700 54684 8652 54740
rect 8708 54684 8718 54740
rect 24210 54684 24220 54740
rect 24276 54684 26460 54740
rect 26516 54684 26526 54740
rect 30818 54684 30828 54740
rect 30884 54684 31836 54740
rect 31892 54684 34860 54740
rect 34916 54684 34926 54740
rect 47954 54684 47964 54740
rect 48020 54684 49532 54740
rect 49588 54684 49598 54740
rect 15138 54572 15148 54628
rect 15204 54572 16492 54628
rect 16548 54572 16558 54628
rect 24882 54572 24892 54628
rect 24948 54572 29148 54628
rect 29204 54572 30156 54628
rect 30212 54572 30222 54628
rect 24546 54460 24556 54516
rect 24612 54460 26124 54516
rect 26180 54460 26190 54516
rect 26898 54460 26908 54516
rect 26964 54460 27916 54516
rect 27972 54460 27982 54516
rect 30482 54460 30492 54516
rect 30548 54460 30940 54516
rect 30996 54460 32172 54516
rect 32228 54460 32238 54516
rect 34626 54460 34636 54516
rect 34692 54460 36428 54516
rect 36484 54460 39676 54516
rect 39732 54460 39900 54516
rect 39956 54460 39966 54516
rect 41010 54460 41020 54516
rect 41076 54460 44156 54516
rect 44212 54460 45164 54516
rect 45220 54460 45500 54516
rect 45556 54460 45566 54516
rect 48514 54460 48524 54516
rect 48580 54460 49868 54516
rect 49924 54460 49934 54516
rect 1698 54348 1708 54404
rect 1764 54348 2492 54404
rect 2548 54348 2558 54404
rect 27010 54348 27020 54404
rect 27076 54348 28364 54404
rect 28420 54348 31612 54404
rect 31668 54348 31678 54404
rect 33282 54348 33292 54404
rect 33348 54348 34972 54404
rect 35028 54348 35038 54404
rect 42130 54348 42140 54404
rect 42196 54348 43820 54404
rect 43876 54348 43886 54404
rect 48738 54348 48748 54404
rect 48804 54348 49308 54404
rect 49364 54348 49374 54404
rect 11218 54236 11228 54292
rect 11284 54236 12460 54292
rect 12516 54236 12526 54292
rect 24658 54236 24668 54292
rect 24724 54236 25452 54292
rect 25508 54236 25518 54292
rect 34738 54236 34748 54292
rect 34804 54236 35084 54292
rect 35140 54236 35150 54292
rect 35410 54236 35420 54292
rect 35476 54236 35756 54292
rect 35812 54236 35822 54292
rect 16258 54124 16268 54180
rect 16324 54124 16604 54180
rect 16660 54124 17500 54180
rect 17556 54124 27244 54180
rect 27300 54124 27310 54180
rect 4466 54068 4476 54124
rect 4532 54068 4580 54124
rect 4636 54068 4684 54124
rect 4740 54068 4750 54124
rect 35186 54068 35196 54124
rect 35252 54068 35300 54124
rect 35356 54068 35404 54124
rect 35460 54068 35470 54124
rect 24770 53900 24780 53956
rect 24836 53900 26124 53956
rect 26180 53900 26190 53956
rect 28550 53900 28588 53956
rect 28644 53900 28654 53956
rect 35746 53900 35756 53956
rect 35812 53900 36428 53956
rect 36484 53900 37884 53956
rect 37940 53900 37950 53956
rect 47618 53900 47628 53956
rect 47684 53900 48524 53956
rect 48580 53900 49756 53956
rect 49812 53900 49822 53956
rect 0 53844 800 53872
rect 0 53788 1708 53844
rect 1764 53788 1774 53844
rect 5282 53788 5292 53844
rect 5348 53788 6636 53844
rect 6692 53788 6702 53844
rect 16370 53788 16380 53844
rect 16436 53788 16446 53844
rect 22082 53788 22092 53844
rect 22148 53788 26684 53844
rect 26740 53788 26750 53844
rect 27122 53788 27132 53844
rect 27188 53788 27916 53844
rect 27972 53788 27982 53844
rect 35074 53788 35084 53844
rect 35140 53788 35980 53844
rect 36036 53788 36204 53844
rect 36260 53788 36270 53844
rect 46722 53788 46732 53844
rect 46788 53788 47852 53844
rect 47908 53788 47918 53844
rect 48626 53788 48636 53844
rect 48692 53788 49420 53844
rect 49476 53788 49486 53844
rect 0 53760 800 53788
rect 16380 53732 16436 53788
rect 9426 53676 9436 53732
rect 9492 53676 10556 53732
rect 10612 53676 10622 53732
rect 16380 53676 17948 53732
rect 18004 53676 21308 53732
rect 21364 53676 21374 53732
rect 23314 53676 23324 53732
rect 23380 53676 24444 53732
rect 24500 53676 24510 53732
rect 28018 53676 28028 53732
rect 28084 53676 29484 53732
rect 29540 53676 30268 53732
rect 30324 53676 31052 53732
rect 31108 53676 31118 53732
rect 36530 53676 36540 53732
rect 36596 53676 38220 53732
rect 38276 53676 38286 53732
rect 38612 53676 40124 53732
rect 40180 53676 40796 53732
rect 40852 53676 40862 53732
rect 29698 53564 29708 53620
rect 29764 53564 30044 53620
rect 30100 53564 30110 53620
rect 33170 53564 33180 53620
rect 33236 53564 34412 53620
rect 34468 53564 36764 53620
rect 36820 53564 36830 53620
rect 6626 53452 6636 53508
rect 6692 53452 8092 53508
rect 8148 53452 8158 53508
rect 16146 53452 16156 53508
rect 16212 53452 16604 53508
rect 16660 53452 16670 53508
rect 20066 53452 20076 53508
rect 20132 53452 21868 53508
rect 21924 53452 21934 53508
rect 25778 53452 25788 53508
rect 25844 53452 26572 53508
rect 26628 53452 26638 53508
rect 28242 53452 28252 53508
rect 28308 53452 29932 53508
rect 29988 53452 29998 53508
rect 31602 53452 31612 53508
rect 31668 53452 34076 53508
rect 34132 53452 34860 53508
rect 34916 53452 34926 53508
rect 36194 53452 36204 53508
rect 36260 53452 37324 53508
rect 37380 53452 37390 53508
rect 38612 53396 38668 53676
rect 42476 53564 42700 53620
rect 42756 53564 42766 53620
rect 43810 53564 43820 53620
rect 43876 53564 44828 53620
rect 44884 53564 44894 53620
rect 49634 53564 49644 53620
rect 49700 53564 50316 53620
rect 50372 53564 50876 53620
rect 50932 53564 50942 53620
rect 42476 53508 42532 53564
rect 41346 53452 41356 53508
rect 41412 53452 42252 53508
rect 42308 53452 42318 53508
rect 42466 53452 42476 53508
rect 42532 53452 42542 53508
rect 46610 53452 46620 53508
rect 46676 53452 47516 53508
rect 47572 53452 47582 53508
rect 26852 53340 38668 53396
rect 19826 53284 19836 53340
rect 19892 53284 19940 53340
rect 19996 53284 20044 53340
rect 20100 53284 20110 53340
rect 26852 53284 26908 53340
rect 50546 53284 50556 53340
rect 50612 53284 50660 53340
rect 50716 53284 50764 53340
rect 50820 53284 50830 53340
rect 26674 53228 26684 53284
rect 26740 53228 26908 53284
rect 28364 53228 30940 53284
rect 30996 53228 31006 53284
rect 34738 53228 34748 53284
rect 34804 53228 35420 53284
rect 35476 53228 35486 53284
rect 43362 53228 43372 53284
rect 43428 53228 43708 53284
rect 43764 53228 45052 53284
rect 45108 53228 45948 53284
rect 46004 53228 47180 53284
rect 47236 53228 47246 53284
rect 49074 53228 49084 53284
rect 49140 53228 50204 53284
rect 50260 53228 50270 53284
rect 0 53172 800 53200
rect 28364 53172 28420 53228
rect 0 53116 1708 53172
rect 1764 53116 2492 53172
rect 2548 53116 2558 53172
rect 6962 53116 6972 53172
rect 7028 53116 8428 53172
rect 8484 53116 8494 53172
rect 8642 53116 8652 53172
rect 8708 53116 11676 53172
rect 11732 53116 11742 53172
rect 18050 53116 18060 53172
rect 18116 53116 21028 53172
rect 22978 53116 22988 53172
rect 23044 53116 24220 53172
rect 24276 53116 24286 53172
rect 26852 53116 28364 53172
rect 28420 53116 28430 53172
rect 30034 53116 30044 53172
rect 30100 53116 30828 53172
rect 30884 53116 30894 53172
rect 32274 53116 32284 53172
rect 32340 53116 33068 53172
rect 33124 53116 33134 53172
rect 35186 53116 35196 53172
rect 35252 53116 36764 53172
rect 36820 53116 36830 53172
rect 37426 53116 37436 53172
rect 37492 53116 37996 53172
rect 38052 53116 40460 53172
rect 40516 53116 41244 53172
rect 41300 53116 41804 53172
rect 41860 53116 41870 53172
rect 42354 53116 42364 53172
rect 42420 53116 43148 53172
rect 43204 53116 43214 53172
rect 46498 53116 46508 53172
rect 46564 53116 46956 53172
rect 47012 53116 47022 53172
rect 0 53088 800 53116
rect 20972 53060 21028 53116
rect 26852 53060 26908 53116
rect 1586 53004 1596 53060
rect 1652 53004 2044 53060
rect 2100 53004 2110 53060
rect 6738 53004 6748 53060
rect 6804 53004 7756 53060
rect 7812 53004 7822 53060
rect 12674 53004 12684 53060
rect 12740 53004 13580 53060
rect 13636 53004 13646 53060
rect 16716 53004 20748 53060
rect 20804 53004 20814 53060
rect 20962 53004 20972 53060
rect 21028 53004 21038 53060
rect 26002 53004 26012 53060
rect 26068 53004 26908 53060
rect 27468 53004 29036 53060
rect 29092 53004 30156 53060
rect 30212 53004 30222 53060
rect 33394 53004 33404 53060
rect 33460 53004 36092 53060
rect 36148 53004 36158 53060
rect 37090 53004 37100 53060
rect 37156 53004 41020 53060
rect 41076 53004 41086 53060
rect 41794 53004 41804 53060
rect 41860 53004 42588 53060
rect 42644 53004 42654 53060
rect 45378 53004 45388 53060
rect 45444 53004 48076 53060
rect 48132 53004 48142 53060
rect 16716 52948 16772 53004
rect 27468 52948 27524 53004
rect 8306 52892 8316 52948
rect 8372 52892 9660 52948
rect 9716 52892 11116 52948
rect 11172 52892 11182 52948
rect 12002 52892 12012 52948
rect 12068 52892 16716 52948
rect 16772 52892 16782 52948
rect 19170 52892 19180 52948
rect 19236 52892 21196 52948
rect 21252 52892 21262 52948
rect 22194 52892 22204 52948
rect 22260 52892 22764 52948
rect 22820 52892 22830 52948
rect 23202 52892 23212 52948
rect 23268 52892 23996 52948
rect 24052 52892 24444 52948
rect 24500 52892 24510 52948
rect 26898 52892 26908 52948
rect 26964 52892 27468 52948
rect 27524 52892 27534 52948
rect 27906 52892 27916 52948
rect 27972 52892 29260 52948
rect 29316 52892 29326 52948
rect 31378 52892 31388 52948
rect 31444 52892 32396 52948
rect 32452 52892 32462 52948
rect 35634 52892 35644 52948
rect 35700 52892 37212 52948
rect 37268 52892 37278 52948
rect 37538 52892 37548 52948
rect 37604 52892 39564 52948
rect 39620 52892 39630 52948
rect 42690 52892 42700 52948
rect 42756 52892 42812 52948
rect 42868 52892 42878 52948
rect 46498 52892 46508 52948
rect 46564 52892 47180 52948
rect 47236 52892 47246 52948
rect 42700 52836 42756 52892
rect 13906 52780 13916 52836
rect 13972 52780 14700 52836
rect 14756 52780 15596 52836
rect 15652 52780 15662 52836
rect 18162 52780 18172 52836
rect 18228 52780 20524 52836
rect 20580 52780 20590 52836
rect 25218 52780 25228 52836
rect 25284 52780 27356 52836
rect 27412 52780 27422 52836
rect 34962 52780 34972 52836
rect 35028 52780 35868 52836
rect 35924 52780 35934 52836
rect 36194 52780 36204 52836
rect 36260 52780 36540 52836
rect 36596 52780 42756 52836
rect 45042 52780 45052 52836
rect 45108 52780 47292 52836
rect 47348 52780 47358 52836
rect 13794 52668 13804 52724
rect 13860 52668 14588 52724
rect 14644 52668 14654 52724
rect 15092 52668 15484 52724
rect 15540 52668 15550 52724
rect 20962 52668 20972 52724
rect 21028 52668 21868 52724
rect 21924 52668 21934 52724
rect 24210 52668 24220 52724
rect 24276 52668 25340 52724
rect 25396 52668 26236 52724
rect 26292 52668 26796 52724
rect 26852 52668 26862 52724
rect 28354 52668 28364 52724
rect 28420 52668 29036 52724
rect 29092 52668 29102 52724
rect 30370 52668 30380 52724
rect 30436 52668 30716 52724
rect 30772 52668 30782 52724
rect 31378 52668 31388 52724
rect 31444 52668 31724 52724
rect 31780 52668 31790 52724
rect 49074 52668 49084 52724
rect 49140 52668 50092 52724
rect 50148 52668 50158 52724
rect 15092 52612 15148 52668
rect 14130 52556 14140 52612
rect 14196 52556 15148 52612
rect 15362 52556 15372 52612
rect 15428 52556 16604 52612
rect 16660 52556 16670 52612
rect 20738 52556 20748 52612
rect 20804 52556 25676 52612
rect 25732 52556 25742 52612
rect 28242 52556 28252 52612
rect 28308 52556 29596 52612
rect 29652 52556 29662 52612
rect 0 52500 800 52528
rect 4466 52500 4476 52556
rect 4532 52500 4580 52556
rect 4636 52500 4684 52556
rect 4740 52500 4750 52556
rect 23996 52500 24052 52556
rect 35186 52500 35196 52556
rect 35252 52500 35300 52556
rect 35356 52500 35404 52556
rect 35460 52500 35470 52556
rect 0 52444 1708 52500
rect 1764 52444 2492 52500
rect 2548 52444 2558 52500
rect 23986 52444 23996 52500
rect 24052 52444 24062 52500
rect 27234 52444 27244 52500
rect 27300 52444 27916 52500
rect 27972 52444 27982 52500
rect 29138 52444 29148 52500
rect 29204 52444 29484 52500
rect 29540 52444 29550 52500
rect 0 52416 800 52444
rect 6514 52332 6524 52388
rect 6580 52332 8092 52388
rect 8148 52332 8158 52388
rect 20290 52332 20300 52388
rect 20356 52332 31892 52388
rect 5282 52220 5292 52276
rect 5348 52220 6636 52276
rect 6692 52220 6702 52276
rect 21410 52220 21420 52276
rect 21476 52220 21532 52276
rect 21588 52220 21598 52276
rect 22754 52220 22764 52276
rect 22820 52220 23548 52276
rect 23604 52220 27244 52276
rect 27300 52220 27310 52276
rect 28578 52220 28588 52276
rect 28644 52220 28812 52276
rect 28868 52220 29148 52276
rect 29204 52220 29214 52276
rect 31836 52164 31892 52332
rect 33282 52220 33292 52276
rect 33348 52220 33516 52276
rect 33572 52220 33582 52276
rect 38658 52220 38668 52276
rect 38724 52220 38892 52276
rect 38948 52220 38958 52276
rect 46946 52220 46956 52276
rect 47012 52220 48636 52276
rect 48692 52220 48702 52276
rect 11442 52108 11452 52164
rect 11508 52108 12572 52164
rect 12628 52108 13020 52164
rect 13076 52108 13692 52164
rect 13748 52108 13758 52164
rect 14578 52108 14588 52164
rect 14644 52108 16604 52164
rect 16660 52108 17500 52164
rect 17556 52108 17566 52164
rect 18722 52108 18732 52164
rect 18788 52108 19964 52164
rect 20020 52108 21644 52164
rect 21700 52108 21710 52164
rect 24210 52108 24220 52164
rect 24276 52108 24892 52164
rect 24948 52108 26348 52164
rect 26404 52108 26414 52164
rect 31826 52108 31836 52164
rect 31892 52108 38108 52164
rect 38164 52108 38174 52164
rect 38434 52108 38444 52164
rect 38500 52108 38668 52164
rect 38724 52108 40908 52164
rect 40964 52108 40974 52164
rect 42578 52108 42588 52164
rect 42644 52108 44268 52164
rect 44324 52108 49420 52164
rect 49476 52108 49486 52164
rect 17042 51996 17052 52052
rect 17108 51996 18172 52052
rect 18228 51996 18238 52052
rect 23090 51996 23100 52052
rect 23156 51996 23436 52052
rect 23492 51996 25116 52052
rect 25172 51996 25182 52052
rect 26450 51996 26460 52052
rect 26516 51996 28476 52052
rect 28532 51996 28542 52052
rect 30930 51996 30940 52052
rect 30996 51996 31332 52052
rect 39218 51996 39228 52052
rect 39284 51996 39452 52052
rect 39508 51996 39518 52052
rect 44146 51996 44156 52052
rect 44212 51996 45500 52052
rect 45556 51996 45566 52052
rect 31276 51940 31332 51996
rect 18610 51884 18620 51940
rect 18676 51884 19404 51940
rect 19460 51884 19470 51940
rect 29922 51884 29932 51940
rect 29988 51884 31052 51940
rect 31108 51884 31118 51940
rect 31276 51884 32620 51940
rect 32676 51884 34412 51940
rect 34468 51884 34478 51940
rect 0 51828 800 51856
rect 0 51772 1708 51828
rect 1764 51772 2492 51828
rect 2548 51772 2558 51828
rect 17938 51772 17948 51828
rect 18004 51772 18844 51828
rect 18900 51772 18910 51828
rect 33954 51772 33964 51828
rect 34020 51772 34748 51828
rect 34804 51772 34814 51828
rect 0 51744 800 51772
rect 19826 51716 19836 51772
rect 19892 51716 19940 51772
rect 19996 51716 20044 51772
rect 20100 51716 20110 51772
rect 50546 51716 50556 51772
rect 50612 51716 50660 51772
rect 50716 51716 50764 51772
rect 50820 51716 50830 51772
rect 32722 51660 32732 51716
rect 32788 51660 34076 51716
rect 34132 51660 34142 51716
rect 38770 51660 38780 51716
rect 38836 51660 39564 51716
rect 39620 51660 39630 51716
rect 19058 51548 19068 51604
rect 19124 51548 19740 51604
rect 19796 51548 19806 51604
rect 20514 51548 20524 51604
rect 20580 51548 22092 51604
rect 22148 51548 22158 51604
rect 22642 51548 22652 51604
rect 22708 51548 23772 51604
rect 23828 51548 23838 51604
rect 33954 51548 33964 51604
rect 34020 51548 34030 51604
rect 38994 51548 39004 51604
rect 39060 51548 39228 51604
rect 39284 51548 39294 51604
rect 47058 51548 47068 51604
rect 47124 51548 48860 51604
rect 48916 51548 48926 51604
rect 49298 51548 49308 51604
rect 49364 51548 49756 51604
rect 49812 51548 49822 51604
rect 33964 51492 34020 51548
rect 11778 51436 11788 51492
rect 11844 51436 14028 51492
rect 14084 51436 14094 51492
rect 16482 51436 16492 51492
rect 16548 51436 16828 51492
rect 16884 51436 17388 51492
rect 17444 51436 17454 51492
rect 18834 51436 18844 51492
rect 18900 51436 19964 51492
rect 20020 51436 20030 51492
rect 21186 51436 21196 51492
rect 21252 51436 22876 51492
rect 22932 51436 23212 51492
rect 23268 51436 23278 51492
rect 23548 51436 35644 51492
rect 35700 51436 35710 51492
rect 37986 51436 37996 51492
rect 38052 51436 41804 51492
rect 41860 51436 41870 51492
rect 45378 51436 45388 51492
rect 45444 51436 45724 51492
rect 45780 51436 45790 51492
rect 46722 51436 46732 51492
rect 46788 51436 48972 51492
rect 49028 51436 49038 51492
rect 21858 51324 21868 51380
rect 21924 51324 23324 51380
rect 23380 51324 23390 51380
rect 23548 51268 23604 51436
rect 45724 51380 45780 51436
rect 23734 51324 23772 51380
rect 23828 51324 24220 51380
rect 24276 51324 24286 51380
rect 37874 51324 37884 51380
rect 37940 51324 38892 51380
rect 38948 51324 38958 51380
rect 39414 51324 39452 51380
rect 39508 51324 39518 51380
rect 39890 51324 39900 51380
rect 39956 51324 40012 51380
rect 40068 51324 40078 51380
rect 45724 51324 47068 51380
rect 47124 51324 47404 51380
rect 47460 51324 47470 51380
rect 19282 51212 19292 51268
rect 19348 51212 20300 51268
rect 20356 51212 23604 51268
rect 31378 51212 31388 51268
rect 31444 51212 31836 51268
rect 31892 51212 31902 51268
rect 36082 51212 36092 51268
rect 36148 51212 36764 51268
rect 36820 51212 36830 51268
rect 40002 51212 40012 51268
rect 40068 51212 41356 51268
rect 41412 51212 41422 51268
rect 43810 51212 43820 51268
rect 43876 51212 46396 51268
rect 46452 51212 46462 51268
rect 0 51156 800 51184
rect 0 51100 1708 51156
rect 1764 51100 2940 51156
rect 2996 51100 3006 51156
rect 20626 51100 20636 51156
rect 20692 51100 22204 51156
rect 22260 51100 22270 51156
rect 37986 51100 37996 51156
rect 38052 51100 38668 51156
rect 39638 51100 39676 51156
rect 39732 51100 39742 51156
rect 48066 51100 48076 51156
rect 48132 51100 49196 51156
rect 49252 51100 49262 51156
rect 0 51072 800 51100
rect 38612 51044 38668 51100
rect 21410 50988 21420 51044
rect 21476 50988 23436 51044
rect 23492 50988 23502 51044
rect 38612 50988 39228 51044
rect 39284 50988 39294 51044
rect 4466 50932 4476 50988
rect 4532 50932 4580 50988
rect 4636 50932 4684 50988
rect 4740 50932 4750 50988
rect 35186 50932 35196 50988
rect 35252 50932 35300 50988
rect 35356 50932 35404 50988
rect 35460 50932 35470 50988
rect 20626 50876 20636 50932
rect 20692 50876 21532 50932
rect 21588 50876 21598 50932
rect 38882 50876 38892 50932
rect 38948 50876 39564 50932
rect 39620 50876 41916 50932
rect 41972 50876 41982 50932
rect 10098 50764 10108 50820
rect 10164 50764 12236 50820
rect 12292 50764 17500 50820
rect 17556 50764 17566 50820
rect 18386 50764 18396 50820
rect 18452 50764 19516 50820
rect 19572 50764 21420 50820
rect 21476 50764 21486 50820
rect 22306 50764 22316 50820
rect 22372 50764 23324 50820
rect 23380 50764 29484 50820
rect 29540 50764 33852 50820
rect 33908 50764 36988 50820
rect 37044 50764 37212 50820
rect 37268 50764 37278 50820
rect 2034 50652 2044 50708
rect 2100 50652 5404 50708
rect 5460 50652 5470 50708
rect 14578 50652 14588 50708
rect 14644 50652 15708 50708
rect 15764 50652 15774 50708
rect 20178 50652 20188 50708
rect 20244 50652 26908 50708
rect 26964 50652 26974 50708
rect 41346 50652 41356 50708
rect 41412 50652 41692 50708
rect 41748 50652 41758 50708
rect 42354 50652 42364 50708
rect 42420 50652 46732 50708
rect 46788 50652 47516 50708
rect 47572 50652 47582 50708
rect 1474 50540 1484 50596
rect 1540 50540 2716 50596
rect 2772 50540 2782 50596
rect 9762 50540 9772 50596
rect 9828 50540 11228 50596
rect 11284 50540 11294 50596
rect 12338 50540 12348 50596
rect 12404 50540 12908 50596
rect 12964 50540 12974 50596
rect 13122 50540 13132 50596
rect 13188 50540 17164 50596
rect 17220 50540 18060 50596
rect 18116 50540 18126 50596
rect 20738 50540 20748 50596
rect 20804 50540 22092 50596
rect 22148 50540 22158 50596
rect 0 50484 800 50512
rect 0 50428 2380 50484
rect 2436 50428 3164 50484
rect 3220 50428 3230 50484
rect 7074 50428 7084 50484
rect 7140 50428 7308 50484
rect 7364 50428 7374 50484
rect 7858 50428 7868 50484
rect 7924 50428 8764 50484
rect 8820 50428 9436 50484
rect 9492 50428 9884 50484
rect 9940 50428 9950 50484
rect 10882 50428 10892 50484
rect 10948 50428 12796 50484
rect 12852 50428 12862 50484
rect 13458 50428 13468 50484
rect 13524 50428 13916 50484
rect 13972 50428 13982 50484
rect 15810 50428 15820 50484
rect 15876 50428 16940 50484
rect 16996 50428 20076 50484
rect 20132 50428 23660 50484
rect 23716 50428 23726 50484
rect 0 50400 800 50428
rect 26572 50372 26628 50652
rect 28242 50540 28252 50596
rect 28308 50540 33404 50596
rect 33460 50540 33470 50596
rect 43474 50540 43484 50596
rect 43540 50540 44716 50596
rect 44772 50540 44782 50596
rect 38098 50428 38108 50484
rect 38164 50428 41132 50484
rect 41188 50428 41198 50484
rect 1810 50316 1820 50372
rect 1876 50316 2492 50372
rect 2548 50316 2558 50372
rect 7746 50316 7756 50372
rect 7812 50316 8316 50372
rect 8372 50316 9996 50372
rect 10052 50316 10062 50372
rect 12002 50316 12012 50372
rect 12068 50316 13132 50372
rect 13188 50316 13198 50372
rect 14690 50316 14700 50372
rect 14756 50316 16604 50372
rect 16660 50316 16670 50372
rect 25330 50316 25340 50372
rect 25396 50316 26236 50372
rect 26292 50316 26302 50372
rect 26562 50316 26572 50372
rect 26628 50316 26638 50372
rect 31154 50316 31164 50372
rect 31220 50316 31892 50372
rect 47170 50316 47180 50372
rect 47236 50316 49308 50372
rect 49364 50316 49980 50372
rect 50036 50316 51660 50372
rect 51716 50316 51726 50372
rect 31836 50260 31892 50316
rect 31826 50204 31836 50260
rect 31892 50204 31902 50260
rect 39330 50204 39340 50260
rect 39396 50204 40236 50260
rect 40292 50204 42700 50260
rect 42756 50204 42766 50260
rect 19826 50148 19836 50204
rect 19892 50148 19940 50204
rect 19996 50148 20044 50204
rect 20100 50148 20110 50204
rect 50546 50148 50556 50204
rect 50612 50148 50660 50204
rect 50716 50148 50764 50204
rect 50820 50148 50830 50204
rect 16940 50092 17276 50148
rect 17332 50092 17342 50148
rect 7186 49980 7196 50036
rect 7252 49980 8316 50036
rect 8372 49980 8382 50036
rect 14242 49980 14252 50036
rect 14308 49980 15596 50036
rect 15652 49980 16268 50036
rect 16324 49980 16334 50036
rect 0 49812 800 49840
rect 0 49756 1820 49812
rect 1876 49756 1886 49812
rect 9650 49756 9660 49812
rect 9716 49756 11788 49812
rect 11844 49756 12796 49812
rect 12852 49756 12862 49812
rect 15474 49756 15484 49812
rect 15540 49756 16492 49812
rect 16548 49756 16558 49812
rect 0 49728 800 49756
rect 1698 49644 1708 49700
rect 1764 49644 2492 49700
rect 2548 49644 2558 49700
rect 10322 49644 10332 49700
rect 10388 49644 13580 49700
rect 13636 49644 13646 49700
rect 16940 49476 16996 50092
rect 27458 49980 27468 50036
rect 27524 49980 28140 50036
rect 28196 49980 28206 50036
rect 36530 49980 36540 50036
rect 36596 49980 37548 50036
rect 37604 49980 37996 50036
rect 38052 49980 38062 50036
rect 40226 49980 40236 50036
rect 40292 49980 43148 50036
rect 43204 49980 43214 50036
rect 43810 49980 43820 50036
rect 43876 49980 43886 50036
rect 45910 49980 45948 50036
rect 46004 49980 46014 50036
rect 30370 49868 30380 49924
rect 30436 49868 31164 49924
rect 31220 49868 31230 49924
rect 38210 49868 38220 49924
rect 38276 49868 38668 49924
rect 38724 49868 39228 49924
rect 39284 49868 39294 49924
rect 43820 49812 43876 49980
rect 26338 49756 26348 49812
rect 26404 49756 26908 49812
rect 26964 49756 26974 49812
rect 27234 49756 27244 49812
rect 27300 49756 28700 49812
rect 28756 49756 28766 49812
rect 30146 49756 30156 49812
rect 30212 49756 30716 49812
rect 30772 49756 31388 49812
rect 31444 49756 31454 49812
rect 35298 49756 35308 49812
rect 35364 49756 37100 49812
rect 37156 49756 37166 49812
rect 39974 49756 40012 49812
rect 40068 49756 40078 49812
rect 43474 49756 43484 49812
rect 43540 49756 44268 49812
rect 44324 49756 44334 49812
rect 20066 49644 20076 49700
rect 20132 49644 20412 49700
rect 20468 49644 20478 49700
rect 38658 49644 38668 49700
rect 38724 49644 39340 49700
rect 39396 49644 39406 49700
rect 17798 49532 17836 49588
rect 17892 49532 17902 49588
rect 24322 49532 24332 49588
rect 24388 49532 25228 49588
rect 25284 49532 25294 49588
rect 42130 49532 42140 49588
rect 42196 49532 42924 49588
rect 42980 49532 42990 49588
rect 16930 49420 16940 49476
rect 16996 49420 17006 49476
rect 4466 49364 4476 49420
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4740 49364 4750 49420
rect 35186 49364 35196 49420
rect 35252 49364 35300 49420
rect 35356 49364 35404 49420
rect 35460 49364 35470 49420
rect 20738 49308 20748 49364
rect 20804 49308 21196 49364
rect 21252 49308 21262 49364
rect 30594 49308 30604 49364
rect 30660 49308 31388 49364
rect 31444 49308 31454 49364
rect 2034 49196 2044 49252
rect 2100 49196 10892 49252
rect 10948 49196 10958 49252
rect 11442 49196 11452 49252
rect 11508 49196 12572 49252
rect 12628 49196 12638 49252
rect 0 49140 800 49168
rect 0 49084 1708 49140
rect 1764 49084 1774 49140
rect 4834 49084 4844 49140
rect 4900 49084 5628 49140
rect 5684 49084 5694 49140
rect 8530 49084 8540 49140
rect 8596 49084 8988 49140
rect 9044 49084 9054 49140
rect 26450 49084 26460 49140
rect 26516 49084 26684 49140
rect 26740 49084 26908 49140
rect 39554 49084 39564 49140
rect 39620 49084 40236 49140
rect 40292 49084 40302 49140
rect 0 49056 800 49084
rect 11218 48972 11228 49028
rect 11284 48972 13916 49028
rect 13972 48972 13982 49028
rect 14690 48972 14700 49028
rect 14756 48972 15260 49028
rect 15316 48972 15326 49028
rect 16482 48972 16492 49028
rect 16548 48972 18284 49028
rect 18340 48972 18350 49028
rect 4274 48860 4284 48916
rect 4340 48860 4732 48916
rect 4788 48860 8428 48916
rect 8484 48860 8494 48916
rect 10546 48860 10556 48916
rect 10612 48860 13692 48916
rect 13748 48860 13758 48916
rect 17714 48860 17724 48916
rect 17780 48860 18060 48916
rect 18116 48860 18126 48916
rect 7410 48748 7420 48804
rect 7476 48748 8876 48804
rect 8932 48748 8942 48804
rect 11666 48748 11676 48804
rect 11732 48748 12012 48804
rect 12068 48748 12796 48804
rect 12852 48748 12862 48804
rect 15026 48748 15036 48804
rect 15092 48748 18844 48804
rect 18900 48748 18910 48804
rect 26852 48748 26908 49084
rect 29026 48972 29036 49028
rect 29092 48972 29820 49028
rect 29876 48972 29886 49028
rect 31602 48972 31612 49028
rect 31668 48972 33404 49028
rect 33460 48972 34636 49028
rect 34692 48972 34702 49028
rect 35746 48972 35756 49028
rect 35812 48972 36204 49028
rect 36260 48972 38108 49028
rect 38164 48972 39900 49028
rect 39956 48972 39966 49028
rect 41122 48972 41132 49028
rect 41188 48972 42028 49028
rect 42084 48972 42094 49028
rect 30482 48860 30492 48916
rect 30548 48860 32620 48916
rect 32676 48860 32686 48916
rect 33730 48860 33740 48916
rect 33796 48860 34300 48916
rect 34356 48860 39788 48916
rect 39844 48860 41468 48916
rect 41524 48860 41534 48916
rect 42242 48860 42252 48916
rect 42308 48860 43596 48916
rect 43652 48860 43662 48916
rect 46498 48860 46508 48916
rect 46564 48860 47852 48916
rect 47908 48860 47918 48916
rect 26964 48748 26974 48804
rect 29250 48748 29260 48804
rect 29316 48748 31948 48804
rect 32004 48748 34748 48804
rect 34804 48748 34814 48804
rect 36418 48748 36428 48804
rect 36484 48748 37212 48804
rect 37268 48748 37278 48804
rect 37874 48748 37884 48804
rect 37940 48748 38668 48804
rect 38724 48748 38734 48804
rect 39106 48748 39116 48804
rect 39172 48748 41020 48804
rect 41076 48748 41086 48804
rect 41570 48748 41580 48804
rect 41636 48748 42924 48804
rect 42980 48748 42990 48804
rect 43138 48748 43148 48804
rect 43204 48748 43932 48804
rect 43988 48748 43998 48804
rect 44146 48748 44156 48804
rect 44212 48748 45276 48804
rect 45332 48748 45342 48804
rect 46610 48748 46620 48804
rect 46676 48748 48748 48804
rect 48804 48748 50316 48804
rect 50372 48748 50382 48804
rect 18162 48636 18172 48692
rect 18228 48636 18620 48692
rect 18676 48636 18686 48692
rect 37090 48636 37100 48692
rect 37156 48636 37436 48692
rect 37492 48636 37502 48692
rect 38210 48636 38220 48692
rect 38276 48636 39676 48692
rect 39732 48636 39742 48692
rect 19826 48580 19836 48636
rect 19892 48580 19940 48636
rect 19996 48580 20044 48636
rect 20100 48580 20110 48636
rect 50546 48580 50556 48636
rect 50612 48580 50660 48636
rect 50716 48580 50764 48636
rect 50820 48580 50830 48636
rect 34402 48524 34412 48580
rect 34468 48524 36204 48580
rect 36260 48524 36270 48580
rect 41794 48524 41804 48580
rect 41860 48524 45388 48580
rect 45444 48524 46396 48580
rect 46452 48524 46462 48580
rect 0 48468 800 48496
rect 0 48412 1932 48468
rect 1988 48412 1998 48468
rect 6402 48412 6412 48468
rect 6468 48412 7084 48468
rect 7140 48412 7150 48468
rect 23762 48412 23772 48468
rect 23828 48412 24220 48468
rect 24276 48412 24780 48468
rect 24836 48412 24846 48468
rect 37538 48412 37548 48468
rect 37604 48412 38332 48468
rect 38388 48412 38398 48468
rect 39106 48412 39116 48468
rect 39172 48412 40012 48468
rect 40068 48412 40078 48468
rect 42354 48412 42364 48468
rect 42420 48412 43820 48468
rect 43876 48412 43886 48468
rect 44818 48412 44828 48468
rect 44884 48412 45500 48468
rect 45556 48412 45566 48468
rect 0 48384 800 48412
rect 7186 48300 7196 48356
rect 7252 48300 7756 48356
rect 7812 48300 7822 48356
rect 8642 48300 8652 48356
rect 8708 48300 8988 48356
rect 9044 48300 10108 48356
rect 10164 48300 10174 48356
rect 16818 48300 16828 48356
rect 16884 48300 17388 48356
rect 17444 48300 17454 48356
rect 31378 48300 31388 48356
rect 31444 48300 33068 48356
rect 33124 48300 33134 48356
rect 38434 48300 38444 48356
rect 38500 48300 40460 48356
rect 40516 48300 40526 48356
rect 42466 48300 42476 48356
rect 42532 48300 43260 48356
rect 43316 48300 43326 48356
rect 46386 48300 46396 48356
rect 46452 48300 52332 48356
rect 52388 48300 52398 48356
rect 12898 48188 12908 48244
rect 12964 48188 12974 48244
rect 21522 48188 21532 48244
rect 21588 48188 22428 48244
rect 22484 48188 22494 48244
rect 29922 48188 29932 48244
rect 29988 48188 30716 48244
rect 30772 48188 30782 48244
rect 32050 48188 32060 48244
rect 32116 48188 32732 48244
rect 32788 48188 33292 48244
rect 33348 48188 33358 48244
rect 39330 48188 39340 48244
rect 39396 48188 40236 48244
rect 40292 48188 40796 48244
rect 40852 48188 40862 48244
rect 41458 48188 41468 48244
rect 41524 48188 41916 48244
rect 41972 48188 46172 48244
rect 46228 48188 46238 48244
rect 12908 48132 12964 48188
rect 10098 48076 10108 48132
rect 10164 48076 11116 48132
rect 11172 48076 11182 48132
rect 12450 48076 12460 48132
rect 12516 48076 15708 48132
rect 15764 48076 15774 48132
rect 20962 48076 20972 48132
rect 21028 48076 21756 48132
rect 21812 48076 21822 48132
rect 23650 48076 23660 48132
rect 23716 48076 24780 48132
rect 24836 48076 25116 48132
rect 25172 48076 27244 48132
rect 27300 48076 27310 48132
rect 35746 48076 35756 48132
rect 35812 48076 36876 48132
rect 36932 48076 39228 48132
rect 39284 48076 39294 48132
rect 40450 48076 40460 48132
rect 40516 48076 40908 48132
rect 40964 48076 40974 48132
rect 43922 48076 43932 48132
rect 43988 48076 48188 48132
rect 48244 48076 48254 48132
rect 1922 47964 1932 48020
rect 1988 47964 1998 48020
rect 6290 47964 6300 48020
rect 6356 47964 6860 48020
rect 6916 47964 7420 48020
rect 7476 47964 7486 48020
rect 34738 47964 34748 48020
rect 34804 47964 37772 48020
rect 37828 47964 37838 48020
rect 42924 47964 43596 48020
rect 43652 47964 44380 48020
rect 44436 47964 44446 48020
rect 0 47796 800 47824
rect 1932 47796 1988 47964
rect 42924 47908 42980 47964
rect 18498 47852 18508 47908
rect 18564 47852 19068 47908
rect 19124 47852 24668 47908
rect 24724 47852 33516 47908
rect 33572 47852 33582 47908
rect 33814 47852 33852 47908
rect 33908 47852 33918 47908
rect 37314 47852 37324 47908
rect 37380 47852 42924 47908
rect 42980 47852 42990 47908
rect 4466 47796 4476 47852
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4740 47796 4750 47852
rect 35186 47796 35196 47852
rect 35252 47796 35300 47852
rect 35356 47796 35404 47852
rect 35460 47796 35470 47852
rect 0 47740 1988 47796
rect 17826 47740 17836 47796
rect 17892 47740 18060 47796
rect 18116 47740 18126 47796
rect 27234 47740 27244 47796
rect 27300 47740 27804 47796
rect 27860 47740 27870 47796
rect 0 47712 800 47740
rect 14466 47628 14476 47684
rect 14532 47628 15820 47684
rect 15876 47628 15886 47684
rect 21074 47628 21084 47684
rect 21140 47628 21756 47684
rect 21812 47628 21822 47684
rect 30716 47628 32508 47684
rect 32564 47628 34300 47684
rect 34356 47628 35980 47684
rect 36036 47628 36046 47684
rect 37202 47628 37212 47684
rect 37268 47628 38108 47684
rect 38164 47628 38174 47684
rect 30716 47572 30772 47628
rect 16258 47516 16268 47572
rect 16324 47516 17948 47572
rect 18004 47516 18014 47572
rect 21410 47516 21420 47572
rect 21476 47516 21980 47572
rect 22036 47516 22046 47572
rect 22418 47516 22428 47572
rect 22484 47516 23716 47572
rect 28914 47516 28924 47572
rect 28980 47516 30716 47572
rect 30772 47516 30782 47572
rect 36988 47516 38892 47572
rect 38948 47516 38958 47572
rect 39554 47516 39564 47572
rect 39620 47516 40572 47572
rect 40628 47516 40638 47572
rect 44034 47516 44044 47572
rect 44100 47516 45164 47572
rect 45220 47516 48300 47572
rect 48356 47516 48366 47572
rect 48738 47516 48748 47572
rect 48804 47516 49756 47572
rect 49812 47516 49822 47572
rect 4834 47404 4844 47460
rect 4900 47404 18508 47460
rect 18564 47404 22652 47460
rect 22708 47404 22718 47460
rect 23660 47348 23716 47516
rect 36988 47460 37044 47516
rect 48748 47460 48804 47516
rect 26786 47404 26796 47460
rect 26852 47404 28028 47460
rect 28084 47404 28094 47460
rect 29810 47404 29820 47460
rect 29876 47404 30492 47460
rect 30548 47404 31836 47460
rect 31892 47404 31902 47460
rect 32498 47404 32508 47460
rect 32564 47404 32732 47460
rect 32788 47404 32798 47460
rect 34412 47404 34972 47460
rect 35028 47404 36988 47460
rect 37044 47404 37054 47460
rect 38434 47404 38444 47460
rect 38500 47404 38668 47460
rect 38724 47404 41020 47460
rect 41076 47404 41086 47460
rect 45714 47404 45724 47460
rect 45780 47404 46620 47460
rect 46676 47404 47180 47460
rect 47236 47404 47246 47460
rect 47730 47404 47740 47460
rect 47796 47404 48804 47460
rect 16034 47292 16044 47348
rect 16100 47292 20076 47348
rect 20132 47292 20142 47348
rect 20962 47292 20972 47348
rect 21028 47292 23100 47348
rect 23156 47292 23166 47348
rect 23650 47292 23660 47348
rect 23716 47292 24220 47348
rect 24276 47292 24286 47348
rect 27570 47292 27580 47348
rect 27636 47292 28140 47348
rect 28196 47292 28206 47348
rect 29586 47292 29596 47348
rect 29652 47292 31612 47348
rect 31668 47292 31678 47348
rect 34412 47236 34468 47404
rect 47740 47348 47796 47404
rect 39778 47292 39788 47348
rect 39844 47292 41132 47348
rect 41188 47292 41198 47348
rect 42914 47292 42924 47348
rect 42980 47292 44492 47348
rect 44548 47292 44558 47348
rect 45938 47292 45948 47348
rect 46004 47292 47796 47348
rect 10546 47180 10556 47236
rect 10612 47180 11676 47236
rect 11732 47180 11742 47236
rect 12226 47180 12236 47236
rect 12292 47180 16268 47236
rect 16324 47180 16334 47236
rect 17378 47180 17388 47236
rect 17444 47180 19628 47236
rect 19684 47180 19694 47236
rect 23874 47180 23884 47236
rect 23940 47180 24444 47236
rect 24500 47180 25228 47236
rect 25284 47180 25294 47236
rect 28242 47180 28252 47236
rect 28308 47180 28318 47236
rect 29026 47180 29036 47236
rect 29092 47180 32508 47236
rect 32564 47180 32574 47236
rect 34402 47180 34412 47236
rect 34468 47180 34478 47236
rect 34962 47180 34972 47236
rect 35028 47180 37996 47236
rect 38052 47180 38062 47236
rect 38322 47180 38332 47236
rect 38388 47180 41580 47236
rect 41636 47180 43260 47236
rect 43316 47180 43326 47236
rect 43922 47180 43932 47236
rect 43988 47180 46956 47236
rect 47012 47180 47022 47236
rect 0 47124 800 47152
rect 0 47068 1932 47124
rect 1988 47068 1998 47124
rect 0 47040 800 47068
rect 19826 47012 19836 47068
rect 19892 47012 19940 47068
rect 19996 47012 20044 47068
rect 20100 47012 20110 47068
rect 28252 47012 28308 47180
rect 29362 47068 29372 47124
rect 29428 47068 29708 47124
rect 29764 47068 29774 47124
rect 30146 47068 30156 47124
rect 30212 47068 31276 47124
rect 31332 47068 32060 47124
rect 32116 47068 32126 47124
rect 32844 47068 33516 47124
rect 33572 47068 33582 47124
rect 36866 47068 36876 47124
rect 36932 47068 41916 47124
rect 41972 47068 41982 47124
rect 45938 47068 45948 47124
rect 46004 47068 46396 47124
rect 46452 47068 46462 47124
rect 32844 47012 32900 47068
rect 50546 47012 50556 47068
rect 50612 47012 50660 47068
rect 50716 47012 50764 47068
rect 50820 47012 50830 47068
rect 4610 46956 4620 47012
rect 4676 46956 5292 47012
rect 5348 46956 5852 47012
rect 5908 46956 5918 47012
rect 10322 46956 10332 47012
rect 10388 46956 11228 47012
rect 11284 46956 11294 47012
rect 26562 46956 26572 47012
rect 26628 46956 28476 47012
rect 28532 46956 28542 47012
rect 32834 46956 32844 47012
rect 32900 46956 32910 47012
rect 33058 46956 33068 47012
rect 33124 46956 33964 47012
rect 34020 46956 34030 47012
rect 34178 46956 34188 47012
rect 34244 46956 34636 47012
rect 34692 46956 34702 47012
rect 39442 46956 39452 47012
rect 39508 46956 41132 47012
rect 41188 46956 41198 47012
rect 42354 46956 42364 47012
rect 42420 46956 43260 47012
rect 43316 46956 43708 47012
rect 43764 46956 43774 47012
rect 44258 46956 44268 47012
rect 44324 46956 45052 47012
rect 45108 46956 45118 47012
rect 6402 46844 6412 46900
rect 6468 46844 7756 46900
rect 7812 46844 7822 46900
rect 8418 46844 8428 46900
rect 8484 46844 21812 46900
rect 22082 46844 22092 46900
rect 22148 46844 22428 46900
rect 22484 46844 22494 46900
rect 27122 46844 27132 46900
rect 27188 46844 27692 46900
rect 27748 46844 27758 46900
rect 28690 46844 28700 46900
rect 28756 46844 29260 46900
rect 29316 46844 32284 46900
rect 32340 46844 36204 46900
rect 36260 46844 36270 46900
rect 41346 46844 41356 46900
rect 41412 46844 43820 46900
rect 43876 46844 44604 46900
rect 44660 46844 44670 46900
rect 46274 46844 46284 46900
rect 46340 46844 46732 46900
rect 46788 46844 46798 46900
rect 2034 46732 2044 46788
rect 2100 46732 12124 46788
rect 12180 46732 12190 46788
rect 21756 46676 21812 46844
rect 34066 46732 34076 46788
rect 34132 46732 34972 46788
rect 35028 46732 35038 46788
rect 42578 46732 42588 46788
rect 42644 46732 42654 46788
rect 47058 46732 47068 46788
rect 47124 46732 47628 46788
rect 47684 46732 47694 46788
rect 21746 46620 21756 46676
rect 21812 46620 25340 46676
rect 25396 46620 25788 46676
rect 25844 46620 25854 46676
rect 34178 46620 34188 46676
rect 34244 46620 35196 46676
rect 35252 46620 37212 46676
rect 37268 46620 37278 46676
rect 42588 46564 42644 46732
rect 42914 46620 42924 46676
rect 42980 46620 43484 46676
rect 43540 46620 43550 46676
rect 46050 46620 46060 46676
rect 46116 46620 47404 46676
rect 47460 46620 47470 46676
rect 5282 46508 5292 46564
rect 5348 46508 8092 46564
rect 8148 46508 8158 46564
rect 20626 46508 20636 46564
rect 20692 46508 22428 46564
rect 22484 46508 22494 46564
rect 25554 46508 25564 46564
rect 25620 46508 27580 46564
rect 27636 46508 27646 46564
rect 33730 46508 33740 46564
rect 33796 46508 34636 46564
rect 34692 46508 36764 46564
rect 36820 46508 36830 46564
rect 42588 46508 42812 46564
rect 42868 46508 42878 46564
rect 47506 46508 47516 46564
rect 47572 46508 48300 46564
rect 48356 46508 48366 46564
rect 0 46452 800 46480
rect 59200 46452 60000 46480
rect 0 46396 1708 46452
rect 1764 46396 2940 46452
rect 2996 46396 3006 46452
rect 9538 46396 9548 46452
rect 9604 46396 10220 46452
rect 10276 46396 11564 46452
rect 11620 46396 11630 46452
rect 23538 46396 23548 46452
rect 23604 46396 25228 46452
rect 25284 46396 25294 46452
rect 32050 46396 32060 46452
rect 32116 46396 33180 46452
rect 33236 46396 36988 46452
rect 37044 46396 37054 46452
rect 43698 46396 43708 46452
rect 43764 46396 44828 46452
rect 44884 46396 44894 46452
rect 55346 46396 55356 46452
rect 55412 46396 60000 46452
rect 0 46368 800 46396
rect 59200 46368 60000 46396
rect 5394 46284 5404 46340
rect 5460 46284 10444 46340
rect 10500 46284 10510 46340
rect 27906 46284 27916 46340
rect 27972 46284 28700 46340
rect 28756 46284 28766 46340
rect 36194 46284 36204 46340
rect 36260 46284 45388 46340
rect 45444 46284 45454 46340
rect 47618 46284 47628 46340
rect 47684 46284 47694 46340
rect 4466 46228 4476 46284
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4740 46228 4750 46284
rect 28700 46228 28756 46284
rect 35186 46228 35196 46284
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35460 46228 35470 46284
rect 7970 46172 7980 46228
rect 8036 46172 8046 46228
rect 14914 46172 14924 46228
rect 14980 46172 25788 46228
rect 25844 46172 25854 46228
rect 28700 46172 29260 46228
rect 29316 46172 29326 46228
rect 0 45780 800 45808
rect 7980 45780 8036 46172
rect 10658 45948 10668 46004
rect 10724 45948 11340 46004
rect 11396 45948 11406 46004
rect 17154 45948 17164 46004
rect 17220 45948 20748 46004
rect 20804 45948 20814 46004
rect 33730 45948 33740 46004
rect 33796 45948 33964 46004
rect 34020 45948 34030 46004
rect 35410 45948 35420 46004
rect 35476 45948 36428 46004
rect 36484 45948 36494 46004
rect 37762 45948 37772 46004
rect 37828 45948 38556 46004
rect 38612 45948 40908 46004
rect 40964 45948 40974 46004
rect 47628 45892 47684 46284
rect 10770 45836 10780 45892
rect 10836 45836 11116 45892
rect 11172 45836 11182 45892
rect 22530 45836 22540 45892
rect 22596 45836 23772 45892
rect 23828 45836 24892 45892
rect 24948 45836 24958 45892
rect 33618 45836 33628 45892
rect 33684 45836 34076 45892
rect 34132 45836 34142 45892
rect 34626 45836 34636 45892
rect 34692 45836 35868 45892
rect 35924 45836 35934 45892
rect 43474 45836 43484 45892
rect 43540 45836 45052 45892
rect 45108 45836 45118 45892
rect 45266 45836 45276 45892
rect 45332 45836 46396 45892
rect 46452 45836 47964 45892
rect 48020 45836 48030 45892
rect 51090 45836 51100 45892
rect 51156 45836 55580 45892
rect 55636 45836 55646 45892
rect 59200 45780 60000 45808
rect 0 45724 2380 45780
rect 2436 45724 3164 45780
rect 3220 45724 3230 45780
rect 6514 45724 6524 45780
rect 6580 45724 7532 45780
rect 7588 45724 8036 45780
rect 8418 45724 8428 45780
rect 8484 45724 8764 45780
rect 8820 45724 8988 45780
rect 9044 45724 9054 45780
rect 9538 45724 9548 45780
rect 9604 45724 11228 45780
rect 11284 45724 11294 45780
rect 12786 45724 12796 45780
rect 12852 45724 14476 45780
rect 14532 45724 14542 45780
rect 27010 45724 27020 45780
rect 27076 45724 27356 45780
rect 27412 45724 28476 45780
rect 28532 45724 30380 45780
rect 30436 45724 30446 45780
rect 33394 45724 33404 45780
rect 33460 45724 34972 45780
rect 35028 45724 35038 45780
rect 55010 45724 55020 45780
rect 55076 45724 60000 45780
rect 0 45696 800 45724
rect 59200 45696 60000 45724
rect 2034 45612 2044 45668
rect 2100 45612 2110 45668
rect 6626 45612 6636 45668
rect 6692 45612 7644 45668
rect 7700 45612 7710 45668
rect 19170 45612 19180 45668
rect 19236 45612 20076 45668
rect 20132 45612 21308 45668
rect 21364 45612 21756 45668
rect 21812 45612 21822 45668
rect 22054 45612 22092 45668
rect 22148 45612 22158 45668
rect 23090 45612 23100 45668
rect 23156 45612 23324 45668
rect 23380 45612 23390 45668
rect 31938 45612 31948 45668
rect 32004 45612 35308 45668
rect 35364 45612 35374 45668
rect 2044 45444 2100 45612
rect 6850 45500 6860 45556
rect 6916 45500 7756 45556
rect 7812 45500 7822 45556
rect 8082 45500 8092 45556
rect 8148 45500 8876 45556
rect 8932 45500 8942 45556
rect 33506 45500 33516 45556
rect 33572 45500 35532 45556
rect 35588 45500 36204 45556
rect 36260 45500 36270 45556
rect 19826 45444 19836 45500
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 20100 45444 20110 45500
rect 50546 45444 50556 45500
rect 50612 45444 50660 45500
rect 50716 45444 50764 45500
rect 50820 45444 50830 45500
rect 2044 45388 17724 45444
rect 17780 45388 17790 45444
rect 20962 45388 20972 45444
rect 21028 45388 21868 45444
rect 21924 45388 21934 45444
rect 33954 45388 33964 45444
rect 34020 45388 34636 45444
rect 34692 45388 34702 45444
rect 37202 45388 37212 45444
rect 37268 45388 37772 45444
rect 37828 45388 37838 45444
rect 38612 45388 41804 45444
rect 41860 45388 41870 45444
rect 7970 45276 7980 45332
rect 8036 45276 8652 45332
rect 8708 45276 8718 45332
rect 16594 45276 16604 45332
rect 16660 45276 18284 45332
rect 18340 45276 18956 45332
rect 19012 45276 19022 45332
rect 19282 45276 19292 45332
rect 19348 45276 21420 45332
rect 21476 45276 21486 45332
rect 24658 45276 24668 45332
rect 24724 45276 25564 45332
rect 25620 45276 25630 45332
rect 28690 45276 28700 45332
rect 28756 45276 32396 45332
rect 32452 45276 32462 45332
rect 33730 45276 33740 45332
rect 33796 45276 34748 45332
rect 34804 45276 34814 45332
rect 37090 45276 37100 45332
rect 37156 45276 38108 45332
rect 38164 45276 38174 45332
rect 2034 45164 2044 45220
rect 2100 45164 9772 45220
rect 9828 45164 9838 45220
rect 18162 45164 18172 45220
rect 18228 45164 18844 45220
rect 18900 45164 18910 45220
rect 28578 45164 28588 45220
rect 28644 45164 29372 45220
rect 29428 45164 29438 45220
rect 31266 45164 31276 45220
rect 31332 45164 33964 45220
rect 34020 45164 34030 45220
rect 34962 45164 34972 45220
rect 35028 45164 37436 45220
rect 37492 45164 37502 45220
rect 0 45108 800 45136
rect 0 45052 1820 45108
rect 1876 45052 2268 45108
rect 2324 45052 2334 45108
rect 12674 45052 12684 45108
rect 12740 45052 14364 45108
rect 14420 45052 14430 45108
rect 20626 45052 20636 45108
rect 20692 45052 21308 45108
rect 21364 45052 21374 45108
rect 23202 45052 23212 45108
rect 23268 45052 24444 45108
rect 24500 45052 25340 45108
rect 25396 45052 25406 45108
rect 28690 45052 28700 45108
rect 28756 45052 29148 45108
rect 29204 45052 29214 45108
rect 31042 45052 31052 45108
rect 31108 45052 32284 45108
rect 32340 45052 32350 45108
rect 0 45024 800 45052
rect 1698 44940 1708 44996
rect 1764 44940 2492 44996
rect 2548 44940 2558 44996
rect 12562 44940 12572 44996
rect 12628 44940 13020 44996
rect 13076 44940 13086 44996
rect 13570 44940 13580 44996
rect 13636 44940 14476 44996
rect 14532 44940 14542 44996
rect 28354 44940 28364 44996
rect 28420 44940 29596 44996
rect 29652 44940 29662 44996
rect 30930 44940 30940 44996
rect 30996 44940 31612 44996
rect 31668 44940 31678 44996
rect 38612 44884 38668 45388
rect 44146 45276 44156 45332
rect 44212 45276 44940 45332
rect 44996 45276 45006 45332
rect 45154 45276 45164 45332
rect 45220 45276 45948 45332
rect 46004 45276 46014 45332
rect 45164 45220 45220 45276
rect 42914 45164 42924 45220
rect 42980 45164 43708 45220
rect 43764 45164 43774 45220
rect 44034 45164 44044 45220
rect 44100 45164 45220 45220
rect 59200 45108 60000 45136
rect 44818 45052 44828 45108
rect 44884 45052 45612 45108
rect 45668 45052 45678 45108
rect 57922 45052 57932 45108
rect 57988 45052 60000 45108
rect 59200 45024 60000 45052
rect 43362 44940 43372 44996
rect 43428 44940 43820 44996
rect 43876 44940 43886 44996
rect 1922 44828 1932 44884
rect 1988 44828 9660 44884
rect 9716 44828 9726 44884
rect 12450 44828 12460 44884
rect 12516 44828 12684 44884
rect 12740 44828 13244 44884
rect 13300 44828 13310 44884
rect 31490 44828 31500 44884
rect 31556 44828 38668 44884
rect 34178 44716 34188 44772
rect 34244 44716 35028 44772
rect 4466 44660 4476 44716
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4740 44660 4750 44716
rect 34972 44660 35028 44716
rect 35186 44660 35196 44716
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35460 44660 35470 44716
rect 5170 44604 5180 44660
rect 5236 44604 15148 44660
rect 34962 44604 34972 44660
rect 35028 44604 35038 44660
rect 15092 44548 15148 44604
rect 3378 44492 3388 44548
rect 3444 44492 11116 44548
rect 11172 44492 11182 44548
rect 15092 44492 19292 44548
rect 19348 44492 21532 44548
rect 21588 44492 22092 44548
rect 22148 44492 22158 44548
rect 25106 44492 25116 44548
rect 25172 44492 25182 44548
rect 27132 44492 27468 44548
rect 27524 44492 27534 44548
rect 34402 44492 34412 44548
rect 34468 44492 34748 44548
rect 34804 44492 34814 44548
rect 41346 44492 41356 44548
rect 41412 44492 52220 44548
rect 52276 44492 52286 44548
rect 0 44436 800 44464
rect 25116 44436 25172 44492
rect 0 44380 1708 44436
rect 1764 44380 1774 44436
rect 2706 44380 2716 44436
rect 2772 44380 11900 44436
rect 11956 44380 11966 44436
rect 24098 44380 24108 44436
rect 24164 44380 25172 44436
rect 0 44352 800 44380
rect 10210 44268 10220 44324
rect 10276 44268 17612 44324
rect 17668 44268 22652 44324
rect 22708 44268 23212 44324
rect 23268 44268 23278 44324
rect 27132 44212 27188 44492
rect 59200 44436 60000 44464
rect 33394 44380 33404 44436
rect 33460 44380 34076 44436
rect 34132 44380 34142 44436
rect 34486 44380 34524 44436
rect 34580 44380 34590 44436
rect 35858 44380 35868 44436
rect 35924 44380 42812 44436
rect 42868 44380 42878 44436
rect 57810 44380 57820 44436
rect 57876 44380 60000 44436
rect 59200 44352 60000 44380
rect 35298 44268 35308 44324
rect 35364 44268 44940 44324
rect 44996 44268 45006 44324
rect 46834 44268 46844 44324
rect 46900 44268 48412 44324
rect 48468 44268 49644 44324
rect 49700 44268 49710 44324
rect 51650 44268 51660 44324
rect 51716 44268 55580 44324
rect 55636 44268 55646 44324
rect 7410 44156 7420 44212
rect 7476 44156 8988 44212
rect 9044 44156 9054 44212
rect 11890 44156 11900 44212
rect 11956 44156 12796 44212
rect 12852 44156 13244 44212
rect 13300 44156 13310 44212
rect 20178 44156 20188 44212
rect 20244 44156 20748 44212
rect 20804 44156 20814 44212
rect 24210 44156 24220 44212
rect 24276 44156 24286 44212
rect 27122 44156 27132 44212
rect 27188 44156 27198 44212
rect 32386 44156 32396 44212
rect 32452 44156 35084 44212
rect 35140 44156 37100 44212
rect 37156 44156 37166 44212
rect 38630 44156 38668 44212
rect 38724 44156 38734 44212
rect 40674 44156 40684 44212
rect 40740 44156 41580 44212
rect 41636 44156 42140 44212
rect 42196 44156 42206 44212
rect 47506 44156 47516 44212
rect 47572 44156 48860 44212
rect 48916 44156 48926 44212
rect 2034 44044 2044 44100
rect 2100 44044 6636 44100
rect 6692 44044 6702 44100
rect 12114 44044 12124 44100
rect 12180 44044 12460 44100
rect 12516 44044 12526 44100
rect 17826 44044 17836 44100
rect 17892 44044 18732 44100
rect 18788 44044 18798 44100
rect 20066 44044 20076 44100
rect 20132 44044 21532 44100
rect 21588 44044 21598 44100
rect 12338 43932 12348 43988
rect 12404 43932 12796 43988
rect 12852 43932 12862 43988
rect 16930 43932 16940 43988
rect 16996 43932 17500 43988
rect 17556 43932 18620 43988
rect 18676 43932 19404 43988
rect 19460 43932 19470 43988
rect 19826 43876 19836 43932
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 20100 43876 20110 43932
rect 9538 43820 9548 43876
rect 9604 43820 19684 43876
rect 0 43764 800 43792
rect 19628 43764 19684 43820
rect 24220 43764 24276 44156
rect 26422 44044 26460 44100
rect 26516 44044 26526 44100
rect 28466 44044 28476 44100
rect 28532 44044 29260 44100
rect 29316 44044 29326 44100
rect 50546 43876 50556 43932
rect 50612 43876 50660 43932
rect 50716 43876 50764 43932
rect 50820 43876 50830 43932
rect 33954 43820 33964 43876
rect 34020 43820 35308 43876
rect 35364 43820 35374 43876
rect 0 43708 1708 43764
rect 1764 43708 2492 43764
rect 2548 43708 2558 43764
rect 6402 43708 6412 43764
rect 6468 43708 7644 43764
rect 7700 43708 7710 43764
rect 11330 43708 11340 43764
rect 11396 43708 12236 43764
rect 12292 43708 12302 43764
rect 12786 43708 12796 43764
rect 12852 43708 13692 43764
rect 13748 43708 15932 43764
rect 15988 43708 15998 43764
rect 19628 43708 20188 43764
rect 20244 43708 20254 43764
rect 24220 43708 24332 43764
rect 24388 43708 24398 43764
rect 31490 43708 31500 43764
rect 31556 43708 32284 43764
rect 32340 43708 32350 43764
rect 0 43680 800 43708
rect 33964 43652 34020 43820
rect 59200 43764 60000 43792
rect 46050 43708 46060 43764
rect 46116 43708 46844 43764
rect 46900 43708 46910 43764
rect 50642 43708 50652 43764
rect 50708 43708 51660 43764
rect 51716 43708 51726 43764
rect 57922 43708 57932 43764
rect 57988 43708 60000 43764
rect 59200 43680 60000 43708
rect 1474 43596 1484 43652
rect 1540 43596 9884 43652
rect 9940 43596 9950 43652
rect 11442 43596 11452 43652
rect 11508 43596 12348 43652
rect 12404 43596 12414 43652
rect 17714 43596 17724 43652
rect 17780 43596 18396 43652
rect 18452 43596 18462 43652
rect 20486 43596 20524 43652
rect 20580 43596 20590 43652
rect 25106 43596 25116 43652
rect 25172 43596 28924 43652
rect 28980 43596 29596 43652
rect 29652 43596 29662 43652
rect 32610 43596 32620 43652
rect 32676 43596 34020 43652
rect 35970 43596 35980 43652
rect 36036 43596 38668 43652
rect 38882 43596 38892 43652
rect 38948 43596 39564 43652
rect 39620 43596 39630 43652
rect 38612 43540 38668 43596
rect 11666 43484 11676 43540
rect 11732 43484 12236 43540
rect 12292 43484 12302 43540
rect 16818 43484 16828 43540
rect 16884 43484 18172 43540
rect 18228 43484 18238 43540
rect 19142 43484 19180 43540
rect 19236 43484 19246 43540
rect 23314 43484 23324 43540
rect 23380 43484 23884 43540
rect 23940 43484 23950 43540
rect 27570 43484 27580 43540
rect 27636 43484 29932 43540
rect 29988 43484 33740 43540
rect 33796 43484 38332 43540
rect 38388 43484 38398 43540
rect 38612 43484 42924 43540
rect 42980 43484 42990 43540
rect 2146 43372 2156 43428
rect 2212 43372 10444 43428
rect 10500 43372 10510 43428
rect 11890 43372 11900 43428
rect 11956 43372 12908 43428
rect 12964 43372 12974 43428
rect 26338 43372 26348 43428
rect 26404 43372 26796 43428
rect 26852 43372 26862 43428
rect 30370 43372 30380 43428
rect 30436 43372 30940 43428
rect 30996 43372 31006 43428
rect 35186 43372 35196 43428
rect 35252 43372 36876 43428
rect 36932 43372 36942 43428
rect 38770 43372 38780 43428
rect 38836 43372 40908 43428
rect 40964 43372 40974 43428
rect 1922 43260 1932 43316
rect 1988 43260 1998 43316
rect 12114 43260 12124 43316
rect 12180 43260 13020 43316
rect 13076 43260 14028 43316
rect 14084 43260 14094 43316
rect 16594 43260 16604 43316
rect 16660 43260 18172 43316
rect 18228 43260 18238 43316
rect 21298 43260 21308 43316
rect 21364 43260 21644 43316
rect 21700 43260 22204 43316
rect 22260 43260 22270 43316
rect 33170 43260 33180 43316
rect 33236 43260 52108 43316
rect 52164 43260 52174 43316
rect 0 43092 800 43120
rect 1932 43092 1988 43260
rect 9762 43148 9772 43204
rect 9828 43148 19180 43204
rect 19236 43148 19740 43204
rect 19796 43148 19806 43204
rect 24994 43148 25004 43204
rect 25060 43148 26012 43204
rect 26068 43148 26348 43204
rect 26404 43148 26414 43204
rect 34066 43148 34076 43204
rect 34132 43148 34524 43204
rect 34580 43148 34590 43204
rect 37986 43148 37996 43204
rect 38052 43148 38668 43204
rect 38724 43148 41580 43204
rect 41636 43148 41646 43204
rect 42578 43148 42588 43204
rect 42644 43148 45612 43204
rect 45668 43148 46284 43204
rect 46340 43148 47292 43204
rect 47348 43148 48748 43204
rect 48804 43148 48814 43204
rect 4466 43092 4476 43148
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4740 43092 4750 43148
rect 35186 43092 35196 43148
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35460 43092 35470 43148
rect 41580 43092 41636 43148
rect 59200 43092 60000 43120
rect 0 43036 1988 43092
rect 41580 43036 42700 43092
rect 42756 43036 42766 43092
rect 57922 43036 57932 43092
rect 57988 43036 60000 43092
rect 0 43008 800 43036
rect 59200 43008 60000 43036
rect 4834 42924 4844 42980
rect 4900 42924 20188 42980
rect 20244 42924 20748 42980
rect 20804 42924 22036 42980
rect 23090 42924 23100 42980
rect 23156 42924 23324 42980
rect 23380 42924 23390 42980
rect 45042 42924 45052 42980
rect 45108 42924 53228 42980
rect 53284 42924 53294 42980
rect 21980 42868 22036 42924
rect 2818 42812 2828 42868
rect 2884 42812 9324 42868
rect 9380 42812 10220 42868
rect 10276 42812 10286 42868
rect 21970 42812 21980 42868
rect 22036 42812 22046 42868
rect 23762 42812 23772 42868
rect 23828 42812 27916 42868
rect 27972 42812 27982 42868
rect 32498 42812 32508 42868
rect 32564 42812 33180 42868
rect 33236 42812 33246 42868
rect 37874 42812 37884 42868
rect 37940 42812 39116 42868
rect 39172 42812 43708 42868
rect 47618 42812 47628 42868
rect 47684 42812 49868 42868
rect 49924 42812 50204 42868
rect 50260 42812 50270 42868
rect 43652 42756 43708 42812
rect 18834 42700 18844 42756
rect 18900 42700 19964 42756
rect 20020 42700 21084 42756
rect 21140 42700 21150 42756
rect 24322 42700 24332 42756
rect 24388 42700 25284 42756
rect 29586 42700 29596 42756
rect 29652 42700 30716 42756
rect 30772 42700 31612 42756
rect 31668 42700 31678 42756
rect 32732 42700 33628 42756
rect 33684 42700 34636 42756
rect 34692 42700 34702 42756
rect 37314 42700 37324 42756
rect 37380 42700 37660 42756
rect 37716 42700 37726 42756
rect 38322 42700 38332 42756
rect 38388 42700 39676 42756
rect 39732 42700 40572 42756
rect 40628 42700 41356 42756
rect 41412 42700 41422 42756
rect 43652 42700 45668 42756
rect 46946 42700 46956 42756
rect 47012 42700 47852 42756
rect 47908 42700 48188 42756
rect 48244 42700 48254 42756
rect 53778 42700 53788 42756
rect 53844 42700 55580 42756
rect 55636 42700 55646 42756
rect 25228 42644 25284 42700
rect 32732 42644 32788 42700
rect 12002 42588 12012 42644
rect 12068 42588 13916 42644
rect 13972 42588 13982 42644
rect 23762 42588 23772 42644
rect 23828 42588 24556 42644
rect 24612 42588 24622 42644
rect 25218 42588 25228 42644
rect 25284 42588 26012 42644
rect 26068 42588 26078 42644
rect 26674 42588 26684 42644
rect 26740 42588 32732 42644
rect 32788 42588 32798 42644
rect 33394 42588 33404 42644
rect 33460 42588 34188 42644
rect 34244 42588 35084 42644
rect 35140 42588 35150 42644
rect 36418 42588 36428 42644
rect 36484 42588 38780 42644
rect 38836 42588 39228 42644
rect 39284 42588 39294 42644
rect 40226 42588 40236 42644
rect 40292 42588 41020 42644
rect 41076 42588 41916 42644
rect 41972 42588 44828 42644
rect 44884 42588 45388 42644
rect 45444 42588 45454 42644
rect 45612 42532 45668 42700
rect 10210 42476 10220 42532
rect 10276 42476 11004 42532
rect 11060 42476 11070 42532
rect 18610 42476 18620 42532
rect 18676 42476 21700 42532
rect 23874 42476 23884 42532
rect 23940 42476 24668 42532
rect 24724 42476 24734 42532
rect 25890 42476 25900 42532
rect 25956 42476 26348 42532
rect 26404 42476 26414 42532
rect 26898 42476 26908 42532
rect 26964 42476 28252 42532
rect 28308 42476 28318 42532
rect 29586 42476 29596 42532
rect 29652 42476 30156 42532
rect 30212 42476 31388 42532
rect 31444 42476 37324 42532
rect 37380 42476 37390 42532
rect 40786 42476 40796 42532
rect 40852 42476 42252 42532
rect 42308 42476 42318 42532
rect 45154 42476 45164 42532
rect 45220 42476 46172 42532
rect 46228 42476 46238 42532
rect 0 42420 800 42448
rect 21644 42420 21700 42476
rect 47628 42420 47684 42700
rect 49522 42476 49532 42532
rect 49588 42476 50540 42532
rect 50596 42476 50606 42532
rect 59200 42420 60000 42448
rect 0 42364 1708 42420
rect 1764 42364 2492 42420
rect 2548 42364 2558 42420
rect 21634 42364 21644 42420
rect 21700 42364 22540 42420
rect 22596 42364 36764 42420
rect 36820 42364 36830 42420
rect 47618 42364 47628 42420
rect 47684 42364 47694 42420
rect 57922 42364 57932 42420
rect 57988 42364 60000 42420
rect 0 42336 800 42364
rect 19826 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20110 42364
rect 50546 42308 50556 42364
rect 50612 42308 50660 42364
rect 50716 42308 50764 42364
rect 50820 42308 50830 42364
rect 59200 42336 60000 42364
rect 2034 42252 2044 42308
rect 2100 42252 2110 42308
rect 25778 42252 25788 42308
rect 25844 42252 27580 42308
rect 27636 42252 27646 42308
rect 47058 42252 47068 42308
rect 47124 42252 47460 42308
rect 2044 42084 2100 42252
rect 9986 42140 9996 42196
rect 10052 42140 24780 42196
rect 24836 42140 24846 42196
rect 46508 42140 47180 42196
rect 47236 42140 47246 42196
rect 2044 42028 10444 42084
rect 10500 42028 10510 42084
rect 17826 42028 17836 42084
rect 17892 42028 21308 42084
rect 21364 42028 21374 42084
rect 24546 42028 24556 42084
rect 24612 42028 25228 42084
rect 25284 42028 25294 42084
rect 27234 42028 27244 42084
rect 27300 42028 28476 42084
rect 28532 42028 29708 42084
rect 29764 42028 29774 42084
rect 46508 41972 46564 42140
rect 47404 41972 47460 42252
rect 49298 42028 49308 42084
rect 49364 42028 50316 42084
rect 50372 42028 50382 42084
rect 51650 42028 51660 42084
rect 51716 42028 52668 42084
rect 52724 42028 52734 42084
rect 2034 41916 2044 41972
rect 2100 41916 9884 41972
rect 9940 41916 9950 41972
rect 21970 41916 21980 41972
rect 22036 41916 23660 41972
rect 23716 41916 23726 41972
rect 27122 41916 27132 41972
rect 27188 41916 27692 41972
rect 27748 41916 27758 41972
rect 29810 41916 29820 41972
rect 29876 41916 30492 41972
rect 30548 41916 30558 41972
rect 33282 41916 33292 41972
rect 33348 41916 33628 41972
rect 33684 41916 34860 41972
rect 34916 41916 34926 41972
rect 36754 41916 36764 41972
rect 36820 41916 37324 41972
rect 37380 41916 37548 41972
rect 37604 41916 37614 41972
rect 39666 41916 39676 41972
rect 39732 41916 39742 41972
rect 41458 41916 41468 41972
rect 41524 41916 42924 41972
rect 42980 41916 42990 41972
rect 46498 41916 46508 41972
rect 46564 41916 46574 41972
rect 47404 41916 49084 41972
rect 49140 41916 49150 41972
rect 52098 41916 52108 41972
rect 52164 41916 55468 41972
rect 55524 41916 55534 41972
rect 39676 41860 39732 41916
rect 6626 41804 6636 41860
rect 6692 41804 10556 41860
rect 10612 41804 10622 41860
rect 22642 41804 22652 41860
rect 22708 41804 22988 41860
rect 23044 41804 23054 41860
rect 24434 41804 24444 41860
rect 24500 41804 25340 41860
rect 25396 41804 25406 41860
rect 29334 41804 29372 41860
rect 29428 41804 29438 41860
rect 30818 41804 30828 41860
rect 30884 41804 31948 41860
rect 32004 41804 39732 41860
rect 41010 41804 41020 41860
rect 41076 41804 41580 41860
rect 41636 41804 41646 41860
rect 0 41748 800 41776
rect 59200 41748 60000 41776
rect 0 41692 1708 41748
rect 1764 41692 2492 41748
rect 2548 41692 2558 41748
rect 9874 41692 9884 41748
rect 9940 41692 10892 41748
rect 10948 41692 10958 41748
rect 24780 41692 25004 41748
rect 25060 41692 25452 41748
rect 25508 41692 35644 41748
rect 35700 41692 37660 41748
rect 37716 41692 37726 41748
rect 55346 41692 55356 41748
rect 55412 41692 60000 41748
rect 0 41664 800 41692
rect 4466 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4750 41580
rect 24780 41524 24836 41692
rect 59200 41664 60000 41692
rect 29446 41580 29484 41636
rect 29540 41580 29550 41636
rect 35186 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35470 41580
rect 24770 41468 24780 41524
rect 24836 41468 24846 41524
rect 28476 41468 33404 41524
rect 33460 41468 33470 41524
rect 33842 41468 33852 41524
rect 33908 41468 33964 41524
rect 34020 41468 34030 41524
rect 38612 41468 53228 41524
rect 53284 41468 53294 41524
rect 28476 41412 28532 41468
rect 38612 41412 38668 41468
rect 1586 41356 1596 41412
rect 1652 41356 10108 41412
rect 10164 41356 10174 41412
rect 10434 41356 10444 41412
rect 10500 41356 10780 41412
rect 10836 41356 10846 41412
rect 21522 41356 21532 41412
rect 21588 41356 28532 41412
rect 28690 41356 28700 41412
rect 28756 41356 29148 41412
rect 29204 41356 38668 41412
rect 41122 41356 41132 41412
rect 41188 41356 43036 41412
rect 43092 41356 43102 41412
rect 43652 41356 46732 41412
rect 46788 41356 46798 41412
rect 49522 41356 49532 41412
rect 49588 41356 50988 41412
rect 51044 41356 51054 41412
rect 43652 41300 43708 41356
rect 21970 41244 21980 41300
rect 22036 41244 24444 41300
rect 24500 41244 25116 41300
rect 25172 41244 25182 41300
rect 25442 41244 25452 41300
rect 25508 41244 27468 41300
rect 27524 41244 27534 41300
rect 28018 41244 28028 41300
rect 28084 41244 38108 41300
rect 38164 41244 38556 41300
rect 38612 41244 38622 41300
rect 39666 41244 39676 41300
rect 39732 41244 43708 41300
rect 19954 41132 19964 41188
rect 20020 41132 23100 41188
rect 23156 41132 23166 41188
rect 24444 41132 26460 41188
rect 26516 41132 27580 41188
rect 27636 41132 27646 41188
rect 0 41076 800 41104
rect 24444 41076 24500 41132
rect 28028 41076 28084 41244
rect 29250 41132 29260 41188
rect 29316 41132 29484 41188
rect 29540 41132 29550 41188
rect 33394 41132 33404 41188
rect 33460 41132 34188 41188
rect 34244 41132 35196 41188
rect 35252 41132 35262 41188
rect 43362 41132 43372 41188
rect 43428 41132 45164 41188
rect 45220 41132 49196 41188
rect 49252 41132 49262 41188
rect 59200 41076 60000 41104
rect 0 41020 1708 41076
rect 1764 41020 2492 41076
rect 2548 41020 2558 41076
rect 2706 41020 2716 41076
rect 2772 41020 9772 41076
rect 9828 41020 9838 41076
rect 11554 41020 11564 41076
rect 11620 41020 11630 41076
rect 12226 41020 12236 41076
rect 12292 41020 12684 41076
rect 12740 41020 12750 41076
rect 15698 41020 15708 41076
rect 15764 41020 22652 41076
rect 22708 41020 22718 41076
rect 22978 41020 22988 41076
rect 23044 41020 24500 41076
rect 24658 41020 24668 41076
rect 24724 41020 25564 41076
rect 25620 41020 26012 41076
rect 26068 41020 26078 41076
rect 26852 41020 27020 41076
rect 27076 41020 28084 41076
rect 30370 41020 30380 41076
rect 30436 41020 31276 41076
rect 31332 41020 31342 41076
rect 57922 41020 57932 41076
rect 57988 41020 60000 41076
rect 0 40992 800 41020
rect 11564 40964 11620 41020
rect 26852 40964 26908 41020
rect 59200 40992 60000 41020
rect 2034 40908 2044 40964
rect 2100 40908 11620 40964
rect 19842 40908 19852 40964
rect 19908 40908 20748 40964
rect 20804 40908 21420 40964
rect 21476 40908 21868 40964
rect 21924 40908 21934 40964
rect 23650 40908 23660 40964
rect 23716 40908 25452 40964
rect 25508 40908 25518 40964
rect 26114 40908 26124 40964
rect 26180 40908 26908 40964
rect 34290 40908 34300 40964
rect 34356 40908 34748 40964
rect 34804 40908 34972 40964
rect 35028 40908 35868 40964
rect 35924 40908 35934 40964
rect 49186 40908 49196 40964
rect 49252 40908 51436 40964
rect 51492 40908 51502 40964
rect 29922 40796 29932 40852
rect 29988 40796 30380 40852
rect 30436 40796 30446 40852
rect 35522 40796 35532 40852
rect 35588 40796 39788 40852
rect 39844 40796 39854 40852
rect 19826 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20110 40796
rect 50546 40740 50556 40796
rect 50612 40740 50660 40796
rect 50716 40740 50764 40796
rect 50820 40740 50830 40796
rect 16818 40684 16828 40740
rect 16884 40684 17836 40740
rect 17892 40684 17902 40740
rect 25106 40684 25116 40740
rect 25172 40684 26012 40740
rect 26068 40684 29820 40740
rect 29876 40684 29886 40740
rect 43652 40684 45052 40740
rect 45108 40684 45118 40740
rect 43652 40628 43708 40684
rect 4162 40572 4172 40628
rect 4228 40572 9436 40628
rect 9492 40572 9502 40628
rect 12674 40572 12684 40628
rect 12740 40572 18508 40628
rect 18564 40572 19068 40628
rect 19124 40572 19134 40628
rect 20402 40572 20412 40628
rect 20468 40572 21084 40628
rect 21140 40572 21150 40628
rect 23090 40572 23100 40628
rect 23156 40572 23884 40628
rect 23940 40572 24332 40628
rect 24388 40572 24398 40628
rect 34738 40572 34748 40628
rect 34804 40572 35308 40628
rect 35364 40572 35374 40628
rect 36306 40572 36316 40628
rect 36372 40572 37212 40628
rect 37268 40572 43708 40628
rect 45266 40572 45276 40628
rect 45332 40572 53508 40628
rect 8764 40460 22764 40516
rect 22820 40460 23436 40516
rect 23492 40460 25452 40516
rect 25508 40460 25788 40516
rect 25844 40460 25854 40516
rect 30566 40460 30604 40516
rect 30660 40460 30670 40516
rect 34178 40460 34188 40516
rect 34244 40460 35756 40516
rect 35812 40460 35822 40516
rect 48514 40460 48524 40516
rect 48580 40460 48860 40516
rect 48916 40460 48926 40516
rect 0 40404 800 40432
rect 0 40348 2380 40404
rect 2436 40348 3164 40404
rect 3220 40348 3230 40404
rect 0 40320 800 40348
rect 8764 40292 8820 40460
rect 53452 40404 53508 40572
rect 59200 40404 60000 40432
rect 9426 40348 9436 40404
rect 9492 40348 26460 40404
rect 26516 40348 27244 40404
rect 27300 40348 27310 40404
rect 32050 40348 32060 40404
rect 32116 40348 33964 40404
rect 34020 40348 34030 40404
rect 34402 40348 34412 40404
rect 34468 40348 34748 40404
rect 34804 40348 34814 40404
rect 35186 40348 35196 40404
rect 35252 40348 36204 40404
rect 36260 40348 36270 40404
rect 38994 40348 39004 40404
rect 39060 40348 39564 40404
rect 39620 40348 40908 40404
rect 40964 40348 40974 40404
rect 41570 40348 41580 40404
rect 41636 40348 42028 40404
rect 42084 40348 42094 40404
rect 43026 40348 43036 40404
rect 43092 40348 44940 40404
rect 44996 40348 48636 40404
rect 48692 40348 48702 40404
rect 53442 40348 53452 40404
rect 53508 40348 53518 40404
rect 55010 40348 55020 40404
rect 55076 40348 60000 40404
rect 59200 40320 60000 40348
rect 2034 40236 2044 40292
rect 2100 40236 8820 40292
rect 17042 40236 17052 40292
rect 17108 40236 18284 40292
rect 18340 40236 18350 40292
rect 23874 40236 23884 40292
rect 23940 40236 25116 40292
rect 25172 40236 25182 40292
rect 37874 40236 37884 40292
rect 37940 40236 38780 40292
rect 38836 40236 38846 40292
rect 47730 40236 47740 40292
rect 47796 40236 52108 40292
rect 52164 40236 52174 40292
rect 30482 40124 30492 40180
rect 30548 40124 30558 40180
rect 46162 40124 46172 40180
rect 46228 40124 46956 40180
rect 47012 40124 47022 40180
rect 53778 40124 53788 40180
rect 53844 40124 53854 40180
rect 16258 40012 16268 40068
rect 16324 40012 19628 40068
rect 19684 40012 19694 40068
rect 4466 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4750 40012
rect 5842 39900 5852 39956
rect 5908 39900 11228 39956
rect 11284 39900 11294 39956
rect 15026 39900 15036 39956
rect 15092 39900 17948 39956
rect 18004 39900 18014 39956
rect 30492 39844 30548 40124
rect 53788 40068 53844 40124
rect 43474 40012 43484 40068
rect 43540 40012 44156 40068
rect 44212 40012 53844 40068
rect 35186 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35470 40012
rect 4274 39788 4284 39844
rect 4340 39788 13916 39844
rect 13972 39788 15148 39844
rect 20178 39788 20188 39844
rect 20244 39788 20748 39844
rect 20804 39788 21532 39844
rect 21588 39788 30548 39844
rect 32386 39788 32396 39844
rect 32452 39788 55468 39844
rect 55524 39788 55534 39844
rect 0 39732 800 39760
rect 15092 39732 15148 39788
rect 59200 39732 60000 39760
rect 0 39676 1708 39732
rect 1764 39676 2940 39732
rect 2996 39676 3006 39732
rect 12898 39676 12908 39732
rect 12964 39676 13580 39732
rect 13636 39676 13646 39732
rect 15092 39676 16828 39732
rect 16884 39676 17388 39732
rect 17444 39676 17454 39732
rect 18722 39676 18732 39732
rect 18788 39676 19964 39732
rect 20020 39676 20030 39732
rect 23202 39676 23212 39732
rect 23268 39676 24332 39732
rect 24388 39676 24398 39732
rect 41458 39676 41468 39732
rect 41524 39676 43372 39732
rect 43428 39676 43438 39732
rect 55346 39676 55356 39732
rect 55412 39676 60000 39732
rect 0 39648 800 39676
rect 59200 39648 60000 39676
rect 6738 39564 6748 39620
rect 6804 39564 10444 39620
rect 10500 39564 10510 39620
rect 10994 39564 11004 39620
rect 11060 39564 15260 39620
rect 15316 39564 15326 39620
rect 17490 39564 17500 39620
rect 17556 39564 19516 39620
rect 19572 39564 19582 39620
rect 26786 39564 26796 39620
rect 2034 39452 2044 39508
rect 2100 39452 10556 39508
rect 10612 39452 10622 39508
rect 26852 39396 26908 39620
rect 29586 39564 29596 39620
rect 29652 39564 31388 39620
rect 31444 39564 32172 39620
rect 32228 39564 32238 39620
rect 43026 39564 43036 39620
rect 43092 39564 43932 39620
rect 43988 39564 55580 39620
rect 55636 39564 55646 39620
rect 30044 39508 30100 39564
rect 29782 39452 29820 39508
rect 29876 39452 29886 39508
rect 30034 39452 30044 39508
rect 30100 39452 30110 39508
rect 31826 39452 31836 39508
rect 31892 39452 32396 39508
rect 32452 39452 32462 39508
rect 36082 39452 36092 39508
rect 36148 39452 36876 39508
rect 36932 39452 45164 39508
rect 45220 39452 45230 39508
rect 11890 39340 11900 39396
rect 11956 39340 13468 39396
rect 13524 39340 13534 39396
rect 14018 39340 14028 39396
rect 14084 39340 17052 39396
rect 17108 39340 17118 39396
rect 25554 39340 25564 39396
rect 25620 39340 27468 39396
rect 27524 39340 27534 39396
rect 29362 39340 29372 39396
rect 29428 39340 30380 39396
rect 30436 39340 30446 39396
rect 40898 39340 40908 39396
rect 40964 39340 41356 39396
rect 41412 39340 41422 39396
rect 46386 39340 46396 39396
rect 46452 39340 47628 39396
rect 47684 39340 47694 39396
rect 30146 39228 30156 39284
rect 30212 39228 30716 39284
rect 30772 39228 32508 39284
rect 32564 39228 40684 39284
rect 40740 39228 45388 39284
rect 45444 39228 45454 39284
rect 19826 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20110 39228
rect 50546 39172 50556 39228
rect 50612 39172 50660 39228
rect 50716 39172 50764 39228
rect 50820 39172 50830 39228
rect 14588 39116 15036 39172
rect 15092 39116 15932 39172
rect 15988 39116 15998 39172
rect 17042 39116 17052 39172
rect 17108 39116 19292 39172
rect 19348 39116 19358 39172
rect 20738 39116 20748 39172
rect 20804 39116 21868 39172
rect 21924 39116 21934 39172
rect 0 39060 800 39088
rect 14588 39060 14644 39116
rect 59200 39060 60000 39088
rect 0 39004 1708 39060
rect 1764 39004 2492 39060
rect 2548 39004 2558 39060
rect 14578 39004 14588 39060
rect 14644 39004 14654 39060
rect 15250 39004 15260 39060
rect 15316 39004 16044 39060
rect 16100 39004 16110 39060
rect 24658 39004 24668 39060
rect 24724 39004 25452 39060
rect 25508 39004 25518 39060
rect 31714 39004 31724 39060
rect 31780 39004 32172 39060
rect 32228 39004 32238 39060
rect 38210 39004 38220 39060
rect 38276 39004 39788 39060
rect 39844 39004 39854 39060
rect 40898 39004 40908 39060
rect 40964 39004 45276 39060
rect 45332 39004 45342 39060
rect 45602 39004 45612 39060
rect 45668 39004 46620 39060
rect 46676 39004 49084 39060
rect 49140 39004 49756 39060
rect 49812 39004 49822 39060
rect 57922 39004 57932 39060
rect 57988 39004 60000 39060
rect 0 38976 800 39004
rect 59200 38976 60000 39004
rect 20132 38892 20860 38948
rect 20916 38892 21084 38948
rect 21140 38892 23660 38948
rect 23716 38892 23726 38948
rect 29362 38892 29372 38948
rect 29428 38892 29596 38948
rect 29652 38892 29662 38948
rect 39442 38892 39452 38948
rect 39508 38892 40012 38948
rect 40068 38892 52668 38948
rect 52724 38892 52734 38948
rect 9762 38668 9772 38724
rect 9828 38668 10668 38724
rect 10724 38668 10734 38724
rect 12674 38668 12684 38724
rect 12740 38668 14028 38724
rect 14084 38668 14364 38724
rect 14420 38668 14430 38724
rect 20132 38612 20188 38892
rect 1922 38556 1932 38612
rect 1988 38556 1998 38612
rect 14242 38556 14252 38612
rect 14308 38556 15596 38612
rect 15652 38556 15662 38612
rect 19842 38556 19852 38612
rect 19908 38556 20188 38612
rect 22204 38780 24332 38836
rect 24388 38780 24398 38836
rect 39666 38780 39676 38836
rect 39732 38780 41132 38836
rect 41188 38780 41198 38836
rect 0 38388 800 38416
rect 1932 38388 1988 38556
rect 22204 38500 22260 38780
rect 23650 38668 23660 38724
rect 23716 38668 24556 38724
rect 24612 38668 24622 38724
rect 27458 38668 27468 38724
rect 27524 38668 28700 38724
rect 28756 38668 28766 38724
rect 38322 38668 38332 38724
rect 38388 38668 38892 38724
rect 38948 38668 42028 38724
rect 42084 38668 43260 38724
rect 43316 38668 43326 38724
rect 29698 38556 29708 38612
rect 29764 38556 30604 38612
rect 30660 38556 32172 38612
rect 32228 38556 33292 38612
rect 33348 38556 33358 38612
rect 33516 38556 35532 38612
rect 35588 38556 35598 38612
rect 55346 38556 55356 38612
rect 20514 38444 20524 38500
rect 20580 38444 22260 38500
rect 4466 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4750 38444
rect 33516 38388 33572 38556
rect 35186 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35470 38444
rect 55412 38388 55468 38612
rect 59200 38388 60000 38416
rect 0 38332 1988 38388
rect 14466 38332 14476 38388
rect 14532 38332 19516 38388
rect 19572 38332 19582 38388
rect 21746 38332 21756 38388
rect 21812 38332 22988 38388
rect 23044 38332 23884 38388
rect 23940 38332 33572 38388
rect 55412 38332 60000 38388
rect 0 38304 800 38332
rect 59200 38304 60000 38332
rect 10770 38220 10780 38276
rect 10836 38220 13468 38276
rect 13524 38220 13534 38276
rect 15698 38220 15708 38276
rect 15764 38220 18284 38276
rect 18340 38220 18350 38276
rect 20962 38220 20972 38276
rect 21028 38220 22092 38276
rect 22148 38220 22158 38276
rect 31602 38220 31612 38276
rect 31668 38220 33852 38276
rect 33908 38220 33918 38276
rect 34598 38220 34636 38276
rect 34692 38220 34702 38276
rect 11666 38108 11676 38164
rect 11732 38108 14588 38164
rect 14644 38108 14654 38164
rect 21858 38108 21868 38164
rect 21924 38108 22092 38164
rect 22148 38108 22158 38164
rect 27906 38108 27916 38164
rect 27972 38108 29372 38164
rect 29428 38108 29438 38164
rect 30146 38108 30156 38164
rect 30212 38108 30828 38164
rect 30884 38108 30894 38164
rect 33506 38108 33516 38164
rect 33572 38108 33964 38164
rect 34020 38108 53228 38164
rect 53284 38108 53294 38164
rect 8418 37996 8428 38052
rect 8484 37996 9100 38052
rect 9156 37996 11228 38052
rect 11284 37996 11788 38052
rect 11844 37996 11854 38052
rect 15092 37996 15708 38052
rect 15764 37996 15774 38052
rect 17490 37996 17500 38052
rect 17556 37996 17836 38052
rect 17892 37996 18844 38052
rect 18900 37996 18910 38052
rect 20402 37996 20412 38052
rect 20468 37996 21644 38052
rect 21700 37996 21710 38052
rect 23062 37996 23100 38052
rect 23156 37996 23166 38052
rect 23314 37996 23324 38052
rect 23380 37996 24220 38052
rect 24276 37996 24286 38052
rect 33814 37996 33852 38052
rect 33908 37996 33918 38052
rect 45154 37996 45164 38052
rect 45220 37996 55356 38052
rect 55412 37996 55422 38052
rect 15092 37828 15148 37996
rect 15474 37884 15484 37940
rect 15540 37884 17388 37940
rect 17444 37884 18060 37940
rect 18116 37884 18126 37940
rect 24994 37884 25004 37940
rect 25060 37884 26236 37940
rect 26292 37884 26302 37940
rect 33926 37884 33964 37940
rect 34020 37884 34030 37940
rect 2034 37772 2044 37828
rect 2100 37772 15148 37828
rect 20850 37772 20860 37828
rect 20916 37772 23324 37828
rect 23380 37772 23390 37828
rect 26898 37772 26908 37828
rect 26964 37772 34524 37828
rect 34580 37772 35420 37828
rect 35476 37772 41468 37828
rect 41524 37772 41534 37828
rect 42578 37772 42588 37828
rect 42644 37772 43708 37828
rect 43764 37772 43774 37828
rect 47618 37772 47628 37828
rect 47684 37772 48412 37828
rect 48468 37772 48478 37828
rect 0 37716 800 37744
rect 59200 37716 60000 37744
rect 0 37660 1708 37716
rect 1764 37660 2492 37716
rect 2548 37660 2558 37716
rect 2706 37660 2716 37716
rect 2772 37660 6748 37716
rect 6804 37660 6814 37716
rect 19282 37660 19292 37716
rect 19348 37660 19358 37716
rect 27234 37660 27244 37716
rect 27300 37660 28252 37716
rect 28308 37660 28318 37716
rect 57922 37660 57932 37716
rect 57988 37660 60000 37716
rect 0 37632 800 37660
rect 19292 37492 19348 37660
rect 19826 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20110 37660
rect 50546 37604 50556 37660
rect 50612 37604 50660 37660
rect 50716 37604 50764 37660
rect 50820 37604 50830 37660
rect 59200 37632 60000 37660
rect 22054 37548 22092 37604
rect 22148 37548 22158 37604
rect 24098 37548 24108 37604
rect 24164 37548 31164 37604
rect 31220 37548 31230 37604
rect 14354 37436 14364 37492
rect 14420 37436 15372 37492
rect 15428 37436 15438 37492
rect 15810 37436 15820 37492
rect 15876 37436 16828 37492
rect 16884 37436 16894 37492
rect 17938 37436 17948 37492
rect 18004 37436 18956 37492
rect 19012 37436 19022 37492
rect 19292 37436 20076 37492
rect 20132 37436 20142 37492
rect 20514 37436 20524 37492
rect 20580 37436 21308 37492
rect 21364 37436 24444 37492
rect 24500 37436 26124 37492
rect 26180 37436 26190 37492
rect 27122 37436 27132 37492
rect 27188 37436 27468 37492
rect 27524 37436 29372 37492
rect 29428 37436 29438 37492
rect 30146 37436 30156 37492
rect 30212 37436 30222 37492
rect 41458 37436 41468 37492
rect 41524 37436 42812 37492
rect 42868 37436 42878 37492
rect 47730 37436 47740 37492
rect 47796 37436 48076 37492
rect 48132 37436 49308 37492
rect 49364 37436 49374 37492
rect 30156 37380 30212 37436
rect 11778 37324 11788 37380
rect 11844 37324 13468 37380
rect 13524 37324 13534 37380
rect 15092 37324 27020 37380
rect 27076 37324 30212 37380
rect 30482 37324 30492 37380
rect 30548 37324 31388 37380
rect 31444 37324 31454 37380
rect 11890 37212 11900 37268
rect 11956 37212 12236 37268
rect 12292 37212 13692 37268
rect 13748 37212 13758 37268
rect 15092 37156 15148 37324
rect 20066 37212 20076 37268
rect 20132 37212 21196 37268
rect 21252 37212 21262 37268
rect 22194 37212 22204 37268
rect 22260 37212 22652 37268
rect 22708 37212 24668 37268
rect 24724 37212 24734 37268
rect 25442 37212 25452 37268
rect 25508 37212 25788 37268
rect 25844 37212 26068 37268
rect 41346 37212 41356 37268
rect 41412 37212 41916 37268
rect 41972 37212 45164 37268
rect 45220 37212 45230 37268
rect 48514 37212 48524 37268
rect 48580 37212 49308 37268
rect 49364 37212 53452 37268
rect 53508 37212 53518 37268
rect 7868 37100 15148 37156
rect 18050 37100 18060 37156
rect 18116 37100 18396 37156
rect 18452 37100 18462 37156
rect 18610 37100 18620 37156
rect 18676 37100 20860 37156
rect 20916 37100 20926 37156
rect 21634 37100 21644 37156
rect 21700 37100 22540 37156
rect 22596 37100 23100 37156
rect 23156 37100 23166 37156
rect 25330 37100 25340 37156
rect 25396 37100 25676 37156
rect 25732 37100 25742 37156
rect 0 37044 800 37072
rect 0 36988 1708 37044
rect 1764 36988 2492 37044
rect 2548 36988 2558 37044
rect 0 36960 800 36988
rect 7868 36932 7924 37100
rect 26012 37044 26068 37212
rect 45826 37100 45836 37156
rect 45892 37100 46508 37156
rect 46564 37100 46574 37156
rect 46834 37100 46844 37156
rect 46900 37100 47964 37156
rect 48020 37100 52668 37156
rect 52724 37100 52734 37156
rect 59200 37044 60000 37072
rect 9202 36988 9212 37044
rect 9268 36988 10220 37044
rect 10276 36988 10286 37044
rect 18844 36988 20188 37044
rect 20244 36988 20972 37044
rect 21028 36988 21038 37044
rect 26012 36988 27468 37044
rect 27524 36988 27534 37044
rect 31154 36988 31164 37044
rect 31220 36988 32620 37044
rect 32676 36988 32686 37044
rect 41682 36988 41692 37044
rect 41748 36988 43260 37044
rect 43316 36988 43326 37044
rect 43810 36988 43820 37044
rect 43876 36988 44716 37044
rect 44772 36988 53844 37044
rect 55346 36988 55356 37044
rect 55412 36988 60000 37044
rect 18844 36932 18900 36988
rect 53788 36932 53844 36988
rect 59200 36960 60000 36988
rect 4834 36876 4844 36932
rect 4900 36876 7924 36932
rect 17490 36876 17500 36932
rect 17556 36876 18844 36932
rect 18900 36876 18910 36932
rect 20486 36876 20524 36932
rect 20580 36876 20590 36932
rect 40338 36876 40348 36932
rect 40404 36876 41132 36932
rect 41188 36876 41198 36932
rect 42354 36876 42364 36932
rect 42420 36876 44940 36932
rect 44996 36876 45006 36932
rect 53788 36876 55580 36932
rect 55636 36876 55646 36932
rect 4466 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4750 36876
rect 35186 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35470 36876
rect 16370 36652 16380 36708
rect 16436 36652 18284 36708
rect 18340 36652 18350 36708
rect 20626 36652 20636 36708
rect 20692 36652 26460 36708
rect 26516 36652 26526 36708
rect 49186 36652 49196 36708
rect 49252 36652 50428 36708
rect 50484 36652 50494 36708
rect 1922 36540 1932 36596
rect 1988 36540 1998 36596
rect 16482 36540 16492 36596
rect 16548 36540 16558 36596
rect 16706 36540 16716 36596
rect 16772 36540 17724 36596
rect 17780 36540 17790 36596
rect 22642 36540 22652 36596
rect 22708 36540 23548 36596
rect 23604 36540 23614 36596
rect 26338 36540 26348 36596
rect 26404 36540 27468 36596
rect 27524 36540 27534 36596
rect 43474 36540 43484 36596
rect 43540 36540 44380 36596
rect 44436 36540 44446 36596
rect 0 36372 800 36400
rect 1932 36372 1988 36540
rect 4162 36428 4172 36484
rect 4228 36428 4844 36484
rect 4900 36428 4910 36484
rect 0 36316 1988 36372
rect 0 36288 800 36316
rect 16492 36260 16548 36540
rect 21298 36428 21308 36484
rect 21364 36428 23996 36484
rect 24052 36428 24062 36484
rect 27234 36428 27244 36484
rect 27300 36428 28140 36484
rect 28196 36428 28206 36484
rect 29810 36428 29820 36484
rect 29876 36428 30380 36484
rect 30436 36428 30828 36484
rect 30884 36428 30894 36484
rect 42802 36428 42812 36484
rect 42868 36428 45164 36484
rect 45220 36428 45230 36484
rect 52098 36428 52108 36484
rect 52164 36428 52780 36484
rect 52836 36428 52846 36484
rect 59200 36372 60000 36400
rect 32946 36316 32956 36372
rect 33012 36316 33516 36372
rect 33572 36316 33582 36372
rect 38434 36316 38444 36372
rect 38500 36316 38780 36372
rect 38836 36316 38846 36372
rect 55234 36316 55244 36372
rect 55300 36316 60000 36372
rect 59200 36288 60000 36316
rect 15372 36204 16548 36260
rect 20626 36204 20636 36260
rect 20692 36204 22428 36260
rect 22484 36204 22494 36260
rect 24882 36204 24892 36260
rect 24948 36204 25228 36260
rect 25284 36204 25294 36260
rect 29138 36204 29148 36260
rect 29204 36204 30380 36260
rect 30436 36204 30716 36260
rect 30772 36204 30782 36260
rect 41570 36204 41580 36260
rect 41636 36204 43372 36260
rect 43428 36204 43438 36260
rect 47954 36204 47964 36260
rect 48020 36204 50876 36260
rect 50932 36204 50942 36260
rect 15372 36148 15428 36204
rect 15362 36092 15372 36148
rect 15428 36092 15438 36148
rect 28578 36092 28588 36148
rect 28644 36092 30156 36148
rect 30212 36092 38444 36148
rect 38500 36092 38510 36148
rect 19826 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20110 36092
rect 26450 35980 26460 36036
rect 26516 35980 27020 36036
rect 27076 35980 27356 36036
rect 27412 35980 27916 36036
rect 27972 35980 27982 36036
rect 22978 35868 22988 35924
rect 23044 35868 23548 35924
rect 23604 35868 23772 35924
rect 23828 35868 23838 35924
rect 23986 35868 23996 35924
rect 24052 35868 24090 35924
rect 26002 35868 26012 35924
rect 26068 35868 26908 35924
rect 26964 35868 26974 35924
rect 28588 35812 28644 36092
rect 50546 36036 50556 36092
rect 50612 36036 50660 36092
rect 50716 36036 50764 36092
rect 50820 36036 50830 36092
rect 33618 35980 33628 36036
rect 33684 35980 34412 36036
rect 34468 35980 34478 36036
rect 41010 35980 41020 36036
rect 41076 35980 48188 36036
rect 48244 35980 48254 36036
rect 33730 35868 33740 35924
rect 33796 35868 34748 35924
rect 34804 35868 35644 35924
rect 35700 35868 35710 35924
rect 38210 35868 38220 35924
rect 38276 35868 39788 35924
rect 39844 35868 39854 35924
rect 40114 35868 40124 35924
rect 40180 35868 42700 35924
rect 42756 35868 42766 35924
rect 45154 35868 45164 35924
rect 45220 35868 45500 35924
rect 45556 35868 45566 35924
rect 45826 35868 45836 35924
rect 45892 35868 46284 35924
rect 46340 35868 48076 35924
rect 48132 35868 48142 35924
rect 49074 35868 49084 35924
rect 49140 35868 49420 35924
rect 49476 35868 49486 35924
rect 2034 35756 2044 35812
rect 2100 35756 11004 35812
rect 11060 35756 11070 35812
rect 19170 35756 19180 35812
rect 19236 35756 19404 35812
rect 19460 35756 28644 35812
rect 34514 35756 34524 35812
rect 34580 35756 35084 35812
rect 35140 35756 36540 35812
rect 36596 35756 52108 35812
rect 52164 35756 52174 35812
rect 0 35700 800 35728
rect 59200 35700 60000 35728
rect 0 35644 1708 35700
rect 1764 35644 2492 35700
rect 2548 35644 2558 35700
rect 3332 35644 10780 35700
rect 10836 35644 10846 35700
rect 16482 35644 16492 35700
rect 16548 35644 16940 35700
rect 16996 35644 17388 35700
rect 17444 35644 17454 35700
rect 21410 35644 21420 35700
rect 21476 35644 21980 35700
rect 22036 35644 22764 35700
rect 22820 35644 22830 35700
rect 28130 35644 28140 35700
rect 28196 35644 29260 35700
rect 29316 35644 29326 35700
rect 34290 35644 34300 35700
rect 34356 35644 35532 35700
rect 35588 35644 37212 35700
rect 37268 35644 37278 35700
rect 39890 35644 39900 35700
rect 39956 35644 40908 35700
rect 40964 35644 40974 35700
rect 44258 35644 44268 35700
rect 44324 35644 49868 35700
rect 49924 35644 49934 35700
rect 55010 35644 55020 35700
rect 55076 35644 60000 35700
rect 0 35616 800 35644
rect 3332 35588 3388 35644
rect 59200 35616 60000 35644
rect 2146 35532 2156 35588
rect 2212 35532 3388 35588
rect 18722 35532 18732 35588
rect 18788 35532 19740 35588
rect 19796 35532 21868 35588
rect 21924 35532 21934 35588
rect 34710 35532 34748 35588
rect 34804 35532 34814 35588
rect 42242 35532 42252 35588
rect 42308 35532 44716 35588
rect 44772 35532 46172 35588
rect 46228 35532 46238 35588
rect 50530 35532 50540 35588
rect 50596 35532 51660 35588
rect 51716 35532 55468 35588
rect 55524 35532 55534 35588
rect 9090 35420 9100 35476
rect 9156 35420 10108 35476
rect 10164 35420 10174 35476
rect 10322 35420 10332 35476
rect 10388 35420 11116 35476
rect 11172 35420 11182 35476
rect 11330 35420 11340 35476
rect 11396 35420 12348 35476
rect 12404 35420 12414 35476
rect 17602 35420 17612 35476
rect 17668 35420 19404 35476
rect 19460 35420 19470 35476
rect 15250 35308 15260 35364
rect 15316 35308 16716 35364
rect 16772 35308 16782 35364
rect 4466 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4750 35308
rect 21868 35252 21924 35532
rect 32498 35420 32508 35476
rect 32564 35420 33180 35476
rect 33236 35420 38668 35476
rect 42578 35420 42588 35476
rect 42644 35420 44156 35476
rect 44212 35420 44222 35476
rect 45378 35420 45388 35476
rect 45444 35420 46396 35476
rect 46452 35420 48748 35476
rect 48804 35420 48814 35476
rect 48972 35420 53228 35476
rect 53284 35420 53294 35476
rect 38612 35364 38668 35420
rect 48972 35364 49028 35420
rect 24882 35308 24892 35364
rect 24948 35308 31164 35364
rect 31220 35308 31230 35364
rect 38612 35308 49028 35364
rect 49858 35308 49868 35364
rect 49924 35308 53956 35364
rect 35186 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35470 35308
rect 21868 35196 26572 35252
rect 26628 35196 31276 35252
rect 31332 35196 31342 35252
rect 16818 35084 16828 35140
rect 16884 35084 18956 35140
rect 19012 35084 19022 35140
rect 24518 35084 24556 35140
rect 24612 35084 24622 35140
rect 27346 35084 27356 35140
rect 27412 35084 28476 35140
rect 28532 35084 28542 35140
rect 35858 35084 35868 35140
rect 35924 35084 37100 35140
rect 37156 35084 37166 35140
rect 0 35028 800 35056
rect 0 34972 2380 35028
rect 2436 34972 3164 35028
rect 3220 34972 3230 35028
rect 11218 34972 11228 35028
rect 11284 34972 13020 35028
rect 13076 34972 13086 35028
rect 23202 34972 23212 35028
rect 23268 34972 30268 35028
rect 30324 34972 30604 35028
rect 30660 34972 30670 35028
rect 38770 34972 38780 35028
rect 38836 34972 38846 35028
rect 0 34944 800 34972
rect 3332 34860 12012 34916
rect 12068 34860 12078 34916
rect 16370 34860 16380 34916
rect 16436 34860 17164 34916
rect 17220 34860 17230 34916
rect 26898 34860 26908 34916
rect 26964 34860 27580 34916
rect 27636 34860 27646 34916
rect 3332 34692 3388 34860
rect 38780 34804 38836 34972
rect 53900 34916 53956 35308
rect 55234 35084 55244 35140
rect 55300 35084 56588 35140
rect 56644 35084 56654 35140
rect 59200 35028 60000 35056
rect 55346 34972 55356 35028
rect 55412 34972 60000 35028
rect 59200 34944 60000 34972
rect 40450 34860 40460 34916
rect 40516 34860 40796 34916
rect 40852 34860 43988 34916
rect 47730 34860 47740 34916
rect 47796 34860 48860 34916
rect 48916 34860 48926 34916
rect 53900 34860 55580 34916
rect 55636 34860 55646 34916
rect 43932 34804 43988 34860
rect 20738 34748 20748 34804
rect 20804 34748 21756 34804
rect 21812 34748 21822 34804
rect 28018 34748 28028 34804
rect 28084 34748 29260 34804
rect 29316 34748 29326 34804
rect 31602 34748 31612 34804
rect 31668 34748 31948 34804
rect 32004 34748 33180 34804
rect 33236 34748 35420 34804
rect 35476 34748 35756 34804
rect 35812 34748 35822 34804
rect 38780 34748 39676 34804
rect 39732 34748 40124 34804
rect 40180 34748 40190 34804
rect 40898 34748 40908 34804
rect 40964 34748 43148 34804
rect 43204 34748 43214 34804
rect 43922 34748 43932 34804
rect 43988 34748 44828 34804
rect 44884 34748 44894 34804
rect 2034 34636 2044 34692
rect 2100 34636 3388 34692
rect 12114 34636 12124 34692
rect 12180 34636 12908 34692
rect 12964 34636 17388 34692
rect 17444 34636 17454 34692
rect 27234 34636 27244 34692
rect 27300 34636 29596 34692
rect 29652 34636 29662 34692
rect 33282 34636 33292 34692
rect 33348 34636 33852 34692
rect 33908 34636 33918 34692
rect 35298 34636 35308 34692
rect 35364 34636 36428 34692
rect 36484 34636 38220 34692
rect 38276 34636 38286 34692
rect 38770 34636 38780 34692
rect 38836 34636 39340 34692
rect 39396 34636 39406 34692
rect 42354 34636 42364 34692
rect 42420 34636 43596 34692
rect 43652 34636 43662 34692
rect 45938 34636 45948 34692
rect 46004 34636 46844 34692
rect 46900 34636 47516 34692
rect 47572 34636 47582 34692
rect 48178 34636 48188 34692
rect 48244 34636 55244 34692
rect 55300 34636 55310 34692
rect 41122 34524 41132 34580
rect 41188 34524 41468 34580
rect 41524 34524 41534 34580
rect 41794 34524 41804 34580
rect 41860 34524 42700 34580
rect 42756 34524 42766 34580
rect 19826 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20110 34524
rect 50546 34468 50556 34524
rect 50612 34468 50660 34524
rect 50716 34468 50764 34524
rect 50820 34468 50830 34524
rect 25190 34412 25228 34468
rect 25284 34412 25294 34468
rect 27692 34412 33852 34468
rect 33908 34412 34188 34468
rect 34244 34412 34254 34468
rect 40114 34412 40124 34468
rect 40180 34412 45724 34468
rect 45780 34412 45790 34468
rect 0 34356 800 34384
rect 27692 34356 27748 34412
rect 59200 34356 60000 34384
rect 0 34300 1708 34356
rect 1764 34300 2940 34356
rect 2996 34300 3006 34356
rect 15698 34300 15708 34356
rect 15764 34300 16156 34356
rect 16212 34300 16222 34356
rect 27458 34300 27468 34356
rect 27524 34300 27692 34356
rect 27748 34300 27758 34356
rect 28466 34300 28476 34356
rect 28532 34300 28924 34356
rect 28980 34300 29820 34356
rect 29876 34300 29886 34356
rect 34402 34300 34412 34356
rect 34468 34300 35756 34356
rect 35812 34300 35822 34356
rect 47618 34300 47628 34356
rect 47684 34300 48188 34356
rect 48244 34300 48254 34356
rect 57922 34300 57932 34356
rect 57988 34300 60000 34356
rect 0 34272 800 34300
rect 59200 34272 60000 34300
rect 28354 34188 28364 34244
rect 28420 34188 29484 34244
rect 29540 34188 29550 34244
rect 32610 34188 32620 34244
rect 32676 34188 36988 34244
rect 37044 34188 37054 34244
rect 39330 34188 39340 34244
rect 39396 34188 40908 34244
rect 40964 34188 40974 34244
rect 45602 34188 45612 34244
rect 45668 34188 46732 34244
rect 46788 34188 46798 34244
rect 47954 34188 47964 34244
rect 48020 34188 49532 34244
rect 49588 34188 49598 34244
rect 11778 34076 11788 34132
rect 11844 34076 13580 34132
rect 13636 34076 13646 34132
rect 23650 34076 23660 34132
rect 23716 34076 24444 34132
rect 24500 34076 24510 34132
rect 24770 34076 24780 34132
rect 24836 34076 25452 34132
rect 25508 34076 25518 34132
rect 25666 34076 25676 34132
rect 25732 34076 26908 34132
rect 26964 34076 26974 34132
rect 40674 34076 40684 34132
rect 40740 34076 41020 34132
rect 41076 34076 41086 34132
rect 4274 33964 4284 34020
rect 4340 33964 4732 34020
rect 4788 33964 22652 34020
rect 22708 33964 23212 34020
rect 23268 33964 23278 34020
rect 24658 33964 24668 34020
rect 24724 33964 25788 34020
rect 25844 33964 25854 34020
rect 28550 33964 28588 34020
rect 28644 33964 28654 34020
rect 29698 33964 29708 34020
rect 29764 33964 32060 34020
rect 32116 33964 32396 34020
rect 32452 33964 32462 34020
rect 35074 33964 35084 34020
rect 35140 33964 37212 34020
rect 37268 33964 38332 34020
rect 38388 33964 38398 34020
rect 48178 33964 48188 34020
rect 48244 33964 48412 34020
rect 48468 33964 48478 34020
rect 50978 33964 50988 34020
rect 51044 33964 51660 34020
rect 51716 33964 53452 34020
rect 53508 33964 53518 34020
rect 1922 33852 1932 33908
rect 1988 33852 1998 33908
rect 10210 33852 10220 33908
rect 10276 33852 11116 33908
rect 11172 33852 11182 33908
rect 14914 33852 14924 33908
rect 14980 33852 16156 33908
rect 16212 33852 16222 33908
rect 44370 33852 44380 33908
rect 44436 33852 50428 33908
rect 55346 33852 55356 33908
rect 0 33684 800 33712
rect 1932 33684 1988 33852
rect 25218 33740 25228 33796
rect 25284 33740 26460 33796
rect 26516 33740 26526 33796
rect 48178 33740 48188 33796
rect 48244 33740 48636 33796
rect 48692 33740 48702 33796
rect 4466 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4750 33740
rect 35186 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35470 33740
rect 50372 33684 50428 33852
rect 55412 33684 55468 33908
rect 59200 33684 60000 33712
rect 0 33628 1988 33684
rect 19842 33628 19852 33684
rect 19908 33628 20412 33684
rect 20468 33628 20478 33684
rect 29250 33628 29260 33684
rect 29316 33628 33628 33684
rect 33684 33628 33694 33684
rect 47058 33628 47068 33684
rect 47124 33628 48748 33684
rect 48804 33628 48814 33684
rect 50372 33628 53452 33684
rect 53508 33628 53518 33684
rect 55412 33628 60000 33684
rect 0 33600 800 33628
rect 14690 33516 14700 33572
rect 14756 33516 15260 33572
rect 15316 33516 15326 33572
rect 15474 33516 15484 33572
rect 15540 33516 16268 33572
rect 16324 33516 16334 33572
rect 18498 33516 18508 33572
rect 18564 33516 20636 33572
rect 20692 33516 21196 33572
rect 21252 33516 21262 33572
rect 27458 33516 27468 33572
rect 27524 33516 28476 33572
rect 28532 33516 28542 33572
rect 30930 33516 30940 33572
rect 30996 33516 31836 33572
rect 31892 33516 31902 33572
rect 15484 33460 15540 33516
rect 33628 33460 33684 33628
rect 59200 33600 60000 33628
rect 35522 33516 35532 33572
rect 35588 33516 37436 33572
rect 37492 33516 37502 33572
rect 15026 33404 15036 33460
rect 15092 33404 15540 33460
rect 17602 33404 17612 33460
rect 17668 33404 18060 33460
rect 18116 33404 19292 33460
rect 19348 33404 21980 33460
rect 22036 33404 22046 33460
rect 31266 33404 31276 33460
rect 31332 33404 31500 33460
rect 31556 33404 32620 33460
rect 32676 33404 32686 33460
rect 33628 33404 35140 33460
rect 35858 33404 35868 33460
rect 35924 33404 36652 33460
rect 36708 33404 37548 33460
rect 37604 33404 37614 33460
rect 46274 33404 46284 33460
rect 46340 33404 49532 33460
rect 49588 33404 50092 33460
rect 50148 33404 50652 33460
rect 50708 33404 50718 33460
rect 35084 33348 35140 33404
rect 18834 33292 18844 33348
rect 18900 33292 19628 33348
rect 19684 33292 19694 33348
rect 22418 33292 22428 33348
rect 22484 33292 22876 33348
rect 22932 33292 22942 33348
rect 26908 33292 27580 33348
rect 27636 33292 30044 33348
rect 30100 33292 30110 33348
rect 31154 33292 31164 33348
rect 31220 33292 32284 33348
rect 32340 33292 32350 33348
rect 33618 33292 33628 33348
rect 33684 33292 34076 33348
rect 34132 33292 34142 33348
rect 35074 33292 35084 33348
rect 35140 33292 37660 33348
rect 37716 33292 37726 33348
rect 47954 33292 47964 33348
rect 48020 33292 48748 33348
rect 48804 33292 48814 33348
rect 55412 33292 55580 33348
rect 55636 33292 55646 33348
rect 16930 33180 16940 33236
rect 16996 33180 20412 33236
rect 20468 33180 24892 33236
rect 24948 33180 24958 33236
rect 26908 33124 26964 33292
rect 27122 33180 27132 33236
rect 27188 33180 29372 33236
rect 29428 33180 29438 33236
rect 32834 33180 32844 33236
rect 32900 33180 55356 33236
rect 55412 33180 55468 33292
rect 2034 33068 2044 33124
rect 2100 33068 11788 33124
rect 11844 33068 11854 33124
rect 15092 33068 23100 33124
rect 23156 33068 26572 33124
rect 26628 33068 26638 33124
rect 26898 33068 26908 33124
rect 26964 33068 26974 33124
rect 28466 33068 28476 33124
rect 28532 33068 29148 33124
rect 29204 33068 29214 33124
rect 29586 33068 29596 33124
rect 29652 33068 30380 33124
rect 30436 33068 30446 33124
rect 34178 33068 34188 33124
rect 34244 33068 35532 33124
rect 35588 33068 35980 33124
rect 36036 33068 36046 33124
rect 38434 33068 38444 33124
rect 38500 33068 40684 33124
rect 40740 33068 41020 33124
rect 41076 33068 41086 33124
rect 44146 33068 44156 33124
rect 44212 33068 44940 33124
rect 44996 33068 46284 33124
rect 46340 33068 46350 33124
rect 0 33012 800 33040
rect 15092 33012 15148 33068
rect 59200 33012 60000 33040
rect 0 32956 1708 33012
rect 1764 32956 2492 33012
rect 2548 32956 2558 33012
rect 5058 32956 5068 33012
rect 5124 32956 15148 33012
rect 57922 32956 57932 33012
rect 57988 32956 60000 33012
rect 0 32928 800 32956
rect 19826 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20110 32956
rect 50546 32900 50556 32956
rect 50612 32900 50660 32956
rect 50716 32900 50764 32956
rect 50820 32900 50830 32956
rect 59200 32928 60000 32956
rect 27906 32844 27916 32900
rect 27972 32844 31164 32900
rect 31220 32844 31724 32900
rect 31780 32844 35196 32900
rect 35252 32844 35262 32900
rect 24210 32732 24220 32788
rect 24276 32732 25116 32788
rect 25172 32732 25182 32788
rect 25750 32732 25788 32788
rect 25844 32732 25854 32788
rect 30146 32732 30156 32788
rect 30212 32732 31276 32788
rect 31332 32732 31342 32788
rect 32162 32732 32172 32788
rect 32228 32732 34188 32788
rect 34244 32732 34412 32788
rect 34468 32732 34478 32788
rect 34636 32732 43036 32788
rect 43092 32732 43708 32788
rect 43764 32732 43774 32788
rect 50372 32732 53228 32788
rect 53284 32732 53294 32788
rect 34636 32676 34692 32732
rect 50372 32676 50428 32732
rect 20514 32620 20524 32676
rect 20580 32620 21532 32676
rect 21588 32620 21598 32676
rect 21970 32620 21980 32676
rect 22036 32620 22540 32676
rect 22596 32620 22606 32676
rect 24882 32620 24892 32676
rect 24948 32620 26236 32676
rect 26292 32620 30828 32676
rect 30884 32620 31836 32676
rect 31892 32620 31902 32676
rect 32396 32620 34692 32676
rect 38098 32620 38108 32676
rect 38164 32620 50428 32676
rect 11106 32508 11116 32564
rect 11172 32508 13580 32564
rect 13636 32508 13646 32564
rect 17714 32508 17724 32564
rect 17780 32508 18508 32564
rect 18564 32508 18574 32564
rect 24434 32508 24444 32564
rect 24500 32508 25452 32564
rect 25508 32508 26348 32564
rect 26404 32508 26414 32564
rect 30370 32508 30380 32564
rect 30436 32508 32172 32564
rect 32228 32508 32238 32564
rect 32396 32452 32452 32620
rect 34290 32508 34300 32564
rect 34356 32508 35644 32564
rect 35700 32508 35710 32564
rect 12450 32396 12460 32452
rect 12516 32396 13468 32452
rect 13524 32396 13534 32452
rect 15092 32396 15596 32452
rect 15652 32396 18844 32452
rect 18900 32396 18910 32452
rect 26002 32396 26012 32452
rect 26068 32396 27020 32452
rect 27076 32396 27086 32452
rect 30706 32396 30716 32452
rect 30772 32396 31388 32452
rect 31444 32396 31612 32452
rect 31668 32396 32452 32452
rect 35644 32452 35700 32508
rect 35644 32396 36540 32452
rect 36596 32396 37324 32452
rect 37380 32396 37390 32452
rect 48514 32396 48524 32452
rect 48580 32396 48860 32452
rect 48916 32396 49196 32452
rect 49252 32396 49262 32452
rect 0 32340 800 32368
rect 15092 32340 15148 32396
rect 59200 32340 60000 32368
rect 0 32284 1708 32340
rect 1764 32284 2492 32340
rect 2548 32284 2558 32340
rect 9986 32284 9996 32340
rect 10052 32284 12012 32340
rect 12068 32284 12078 32340
rect 14690 32284 14700 32340
rect 14756 32284 15148 32340
rect 34738 32284 34748 32340
rect 34804 32284 37100 32340
rect 37156 32284 39900 32340
rect 39956 32284 39966 32340
rect 55346 32284 55356 32340
rect 55412 32284 60000 32340
rect 0 32256 800 32284
rect 59200 32256 60000 32284
rect 11330 32172 11340 32228
rect 11396 32172 14028 32228
rect 14084 32172 14094 32228
rect 21270 32172 21308 32228
rect 21364 32172 21374 32228
rect 22754 32172 22764 32228
rect 22820 32172 23436 32228
rect 23492 32172 31948 32228
rect 32004 32172 32014 32228
rect 36082 32172 36092 32228
rect 36148 32172 36988 32228
rect 37044 32172 37054 32228
rect 4466 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4750 32172
rect 35186 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35470 32172
rect 11666 31948 11676 32004
rect 11732 31948 12684 32004
rect 12740 31948 12750 32004
rect 24210 31948 24220 32004
rect 24276 31948 25340 32004
rect 25396 31948 25406 32004
rect 26002 31948 26012 32004
rect 26068 31948 26684 32004
rect 26740 31948 29372 32004
rect 29428 31948 29932 32004
rect 29988 31948 29998 32004
rect 32050 31948 32060 32004
rect 32116 31948 33292 32004
rect 33348 31948 33358 32004
rect 35410 31948 35420 32004
rect 35476 31948 36428 32004
rect 36484 31948 36494 32004
rect 39414 31948 39452 32004
rect 39508 31948 39518 32004
rect 1922 31836 1932 31892
rect 1988 31836 1998 31892
rect 15372 31836 16716 31892
rect 16772 31836 17500 31892
rect 17556 31836 17566 31892
rect 17826 31836 17836 31892
rect 17892 31836 23100 31892
rect 23156 31836 23996 31892
rect 24052 31836 24062 31892
rect 27682 31836 27692 31892
rect 27748 31836 28364 31892
rect 28420 31836 29484 31892
rect 29540 31836 29550 31892
rect 38210 31836 38220 31892
rect 38276 31836 39004 31892
rect 39060 31836 39070 31892
rect 43138 31836 43148 31892
rect 43204 31836 44044 31892
rect 44100 31836 44110 31892
rect 49410 31836 49420 31892
rect 49476 31836 50540 31892
rect 50596 31836 50606 31892
rect 0 31668 800 31696
rect 1932 31668 1988 31836
rect 15372 31780 15428 31836
rect 4162 31724 4172 31780
rect 4228 31724 4844 31780
rect 4900 31724 4910 31780
rect 14466 31724 14476 31780
rect 14532 31724 15372 31780
rect 15428 31724 15438 31780
rect 15810 31724 15820 31780
rect 15876 31724 16604 31780
rect 16660 31724 16670 31780
rect 19170 31724 19180 31780
rect 19236 31724 19628 31780
rect 19684 31724 19694 31780
rect 25666 31724 25676 31780
rect 25732 31724 25900 31780
rect 25956 31724 25966 31780
rect 28102 31724 28140 31780
rect 28196 31724 28206 31780
rect 29362 31724 29372 31780
rect 29428 31724 30268 31780
rect 30324 31724 31500 31780
rect 31556 31724 31566 31780
rect 35634 31724 35644 31780
rect 35700 31724 36316 31780
rect 36372 31724 37548 31780
rect 37604 31724 37614 31780
rect 42802 31724 42812 31780
rect 42868 31724 43260 31780
rect 43316 31724 43326 31780
rect 59200 31668 60000 31696
rect 0 31612 1988 31668
rect 14130 31612 14140 31668
rect 14196 31612 16044 31668
rect 16100 31612 16110 31668
rect 26898 31612 26908 31668
rect 26964 31612 28588 31668
rect 28644 31612 28654 31668
rect 45154 31612 45164 31668
rect 45220 31612 46508 31668
rect 46564 31612 46574 31668
rect 57922 31612 57932 31668
rect 57988 31612 60000 31668
rect 0 31584 800 31612
rect 59200 31584 60000 31612
rect 2034 31500 2044 31556
rect 2100 31500 10108 31556
rect 10164 31500 10174 31556
rect 12338 31500 12348 31556
rect 12404 31500 12684 31556
rect 12740 31500 13692 31556
rect 13748 31500 13758 31556
rect 15026 31500 15036 31556
rect 15092 31500 16380 31556
rect 16436 31500 17612 31556
rect 17668 31500 17678 31556
rect 22530 31500 22540 31556
rect 22596 31500 25452 31556
rect 25508 31500 25518 31556
rect 25666 31500 25676 31556
rect 25732 31500 26236 31556
rect 26292 31500 26302 31556
rect 27794 31500 27804 31556
rect 27860 31500 29148 31556
rect 29204 31500 29214 31556
rect 29362 31500 29372 31556
rect 29428 31500 29932 31556
rect 29988 31500 33068 31556
rect 33124 31500 33134 31556
rect 33730 31500 33740 31556
rect 33796 31500 35532 31556
rect 35588 31500 36316 31556
rect 36372 31500 36382 31556
rect 38854 31500 38892 31556
rect 38948 31500 38958 31556
rect 14018 31388 14028 31444
rect 14084 31388 15596 31444
rect 15652 31388 15662 31444
rect 24546 31388 24556 31444
rect 24612 31388 26348 31444
rect 26404 31388 26414 31444
rect 26852 31388 27356 31444
rect 27412 31388 28140 31444
rect 28196 31388 28206 31444
rect 19826 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20110 31388
rect 22866 31276 22876 31332
rect 22932 31276 23548 31332
rect 23604 31276 23614 31332
rect 23986 31276 23996 31332
rect 24052 31276 25228 31332
rect 25284 31276 25294 31332
rect 25750 31276 25788 31332
rect 25844 31276 25854 31332
rect 26852 31220 26908 31388
rect 50546 31332 50556 31388
rect 50612 31332 50660 31388
rect 50716 31332 50764 31388
rect 50820 31332 50830 31388
rect 27682 31276 27692 31332
rect 27748 31276 30492 31332
rect 30548 31276 30558 31332
rect 2034 31164 2044 31220
rect 2100 31164 5852 31220
rect 5908 31164 5918 31220
rect 9538 31164 9548 31220
rect 9604 31164 26908 31220
rect 31490 31164 31500 31220
rect 31556 31164 33404 31220
rect 33460 31164 33470 31220
rect 39890 31164 39900 31220
rect 39956 31164 41244 31220
rect 41300 31164 41310 31220
rect 42802 31164 42812 31220
rect 42868 31164 42878 31220
rect 46274 31164 46284 31220
rect 46340 31164 46350 31220
rect 48066 31164 48076 31220
rect 48132 31164 48636 31220
rect 48692 31164 48702 31220
rect 42812 31108 42868 31164
rect 16594 31052 16604 31108
rect 16660 31052 17500 31108
rect 17556 31052 17566 31108
rect 22978 31052 22988 31108
rect 23044 31052 23054 31108
rect 30930 31052 30940 31108
rect 30996 31052 31276 31108
rect 31332 31052 31342 31108
rect 33842 31052 33852 31108
rect 33908 31052 35420 31108
rect 35476 31052 35486 31108
rect 36418 31052 36428 31108
rect 36484 31052 36988 31108
rect 37044 31052 37054 31108
rect 41132 31052 42868 31108
rect 0 30996 800 31024
rect 0 30940 1708 30996
rect 1764 30940 2492 30996
rect 2548 30940 2558 30996
rect 10546 30940 10556 30996
rect 10612 30940 12124 30996
rect 12180 30940 12190 30996
rect 0 30912 800 30940
rect 22988 30884 23044 31052
rect 23762 30940 23772 30996
rect 23828 30940 24444 30996
rect 24500 30940 27132 30996
rect 27188 30940 27198 30996
rect 28690 30940 28700 30996
rect 28756 30940 31164 30996
rect 31220 30940 31230 30996
rect 38098 30940 38108 30996
rect 38164 30940 38780 30996
rect 38836 30940 39340 30996
rect 39396 30940 39406 30996
rect 2370 30828 2380 30884
rect 2436 30828 3164 30884
rect 3220 30828 3230 30884
rect 12786 30828 12796 30884
rect 12852 30828 14028 30884
rect 14084 30828 14094 30884
rect 21522 30828 21532 30884
rect 21588 30828 23212 30884
rect 23268 30828 23278 30884
rect 26338 30828 26348 30884
rect 26404 30828 26572 30884
rect 26628 30828 27244 30884
rect 27300 30828 27310 30884
rect 38322 30828 38332 30884
rect 38388 30828 39452 30884
rect 39508 30828 39518 30884
rect 41132 30772 41188 31052
rect 42476 30996 42532 31052
rect 46284 30996 46340 31164
rect 47618 31052 47628 31108
rect 47684 31052 50764 31108
rect 50820 31052 51324 31108
rect 51380 31052 51390 31108
rect 59200 30996 60000 31024
rect 41346 30940 41356 30996
rect 41412 30940 41422 30996
rect 42466 30940 42476 30996
rect 42532 30940 42542 30996
rect 43138 30940 43148 30996
rect 43204 30940 45164 30996
rect 45220 30940 47404 30996
rect 47460 30940 47470 30996
rect 55010 30940 55020 30996
rect 55076 30940 60000 30996
rect 8978 30716 8988 30772
rect 9044 30716 10332 30772
rect 10388 30716 10398 30772
rect 10770 30716 10780 30772
rect 10836 30716 11676 30772
rect 11732 30716 11742 30772
rect 16258 30716 16268 30772
rect 16324 30716 17500 30772
rect 17556 30716 17566 30772
rect 35746 30716 35756 30772
rect 35812 30716 36204 30772
rect 36260 30716 36270 30772
rect 36978 30716 36988 30772
rect 37044 30716 41188 30772
rect 41356 30772 41412 30940
rect 59200 30912 60000 30940
rect 45826 30828 45836 30884
rect 45892 30828 46508 30884
rect 46564 30828 46574 30884
rect 41356 30716 42252 30772
rect 42308 30716 42924 30772
rect 42980 30716 43260 30772
rect 43316 30716 43326 30772
rect 45154 30716 45164 30772
rect 45220 30716 47628 30772
rect 47684 30716 47694 30772
rect 9986 30604 9996 30660
rect 10052 30604 25340 30660
rect 25396 30604 25406 30660
rect 39554 30604 39564 30660
rect 39620 30604 43148 30660
rect 43204 30604 43214 30660
rect 4466 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4750 30604
rect 35186 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35470 30604
rect 2034 30492 2044 30548
rect 2100 30492 3388 30548
rect 24658 30492 24668 30548
rect 24724 30492 28812 30548
rect 28868 30492 28878 30548
rect 35718 30492 35756 30548
rect 35812 30492 35822 30548
rect 45602 30492 45612 30548
rect 45668 30492 45948 30548
rect 46004 30492 46620 30548
rect 46676 30492 46686 30548
rect 3332 30436 3388 30492
rect 2706 30380 2716 30436
rect 2772 30380 2782 30436
rect 3332 30380 8484 30436
rect 25778 30380 25788 30436
rect 25844 30380 26796 30436
rect 26852 30380 26862 30436
rect 32610 30380 32620 30436
rect 32676 30380 47180 30436
rect 47236 30380 47246 30436
rect 0 30324 800 30352
rect 2716 30324 2772 30380
rect 0 30268 2380 30324
rect 2436 30268 2446 30324
rect 2716 30268 5124 30324
rect 0 30240 800 30268
rect 5068 30100 5124 30268
rect 8428 30212 8484 30380
rect 59200 30324 60000 30352
rect 19366 30268 19404 30324
rect 19460 30268 19470 30324
rect 31826 30268 31836 30324
rect 31892 30268 32508 30324
rect 32564 30268 33068 30324
rect 33124 30268 33134 30324
rect 33618 30268 33628 30324
rect 33684 30268 34748 30324
rect 34804 30268 45052 30324
rect 45108 30268 46060 30324
rect 46116 30268 46126 30324
rect 48402 30268 48412 30324
rect 48468 30268 49868 30324
rect 49924 30268 49934 30324
rect 55346 30268 55356 30324
rect 55412 30268 60000 30324
rect 59200 30240 60000 30268
rect 8428 30156 13020 30212
rect 13076 30156 13086 30212
rect 21746 30156 21756 30212
rect 21812 30156 22316 30212
rect 22372 30156 22382 30212
rect 22530 30156 22540 30212
rect 22596 30156 24108 30212
rect 24164 30156 24174 30212
rect 27458 30156 27468 30212
rect 27524 30156 28588 30212
rect 28644 30156 30268 30212
rect 30324 30156 31164 30212
rect 31220 30156 31230 30212
rect 33394 30156 33404 30212
rect 33460 30156 34076 30212
rect 34132 30156 34142 30212
rect 38882 30156 38892 30212
rect 38948 30156 39228 30212
rect 39284 30156 39294 30212
rect 40562 30156 40572 30212
rect 40628 30156 43260 30212
rect 43316 30156 43326 30212
rect 44930 30156 44940 30212
rect 44996 30156 46844 30212
rect 46900 30156 46910 30212
rect 47954 30156 47964 30212
rect 48020 30156 48748 30212
rect 48804 30156 48814 30212
rect 49410 30156 49420 30212
rect 49476 30156 50428 30212
rect 50484 30156 50494 30212
rect 22540 30100 22596 30156
rect 5068 30044 10108 30100
rect 10164 30044 10174 30100
rect 18946 30044 18956 30100
rect 19012 30044 22596 30100
rect 27234 30044 27244 30100
rect 27300 30044 31724 30100
rect 31780 30044 31790 30100
rect 38322 30044 38332 30100
rect 38388 30044 40012 30100
rect 40068 30044 40078 30100
rect 40786 30044 40796 30100
rect 40852 30044 42140 30100
rect 42196 30044 42206 30100
rect 46134 30044 46172 30100
rect 46228 30044 46238 30100
rect 46722 30044 46732 30100
rect 46788 30044 47292 30100
rect 47348 30044 47628 30100
rect 47684 30044 47694 30100
rect 47842 30044 47852 30100
rect 47908 30044 50764 30100
rect 50820 30044 50830 30100
rect 19058 29932 19068 29988
rect 19124 29932 20076 29988
rect 20132 29932 20142 29988
rect 22194 29932 22204 29988
rect 22260 29932 23212 29988
rect 23268 29932 23278 29988
rect 23762 29932 23772 29988
rect 23828 29932 24556 29988
rect 24612 29932 25116 29988
rect 25172 29932 25182 29988
rect 27682 29932 27692 29988
rect 27748 29932 28364 29988
rect 28420 29932 29820 29988
rect 29876 29932 29886 29988
rect 37090 29932 37100 29988
rect 37156 29932 38556 29988
rect 38612 29932 38622 29988
rect 38780 29876 38836 30044
rect 39330 29932 39340 29988
rect 39396 29932 40460 29988
rect 40516 29932 40526 29988
rect 41458 29932 41468 29988
rect 41524 29932 42700 29988
rect 42756 29932 42766 29988
rect 45266 29932 45276 29988
rect 45332 29932 45948 29988
rect 46004 29932 46014 29988
rect 48962 29932 48972 29988
rect 49028 29932 50204 29988
rect 50260 29932 50270 29988
rect 50372 29932 50652 29988
rect 50708 29932 50718 29988
rect 21858 29820 21868 29876
rect 21924 29820 22540 29876
rect 22596 29820 22606 29876
rect 29026 29820 29036 29876
rect 29092 29820 33068 29876
rect 33124 29820 33628 29876
rect 33684 29820 34076 29876
rect 34132 29820 34142 29876
rect 38770 29820 38780 29876
rect 38836 29820 38846 29876
rect 38994 29820 39004 29876
rect 39060 29820 39788 29876
rect 39844 29820 39854 29876
rect 41346 29820 41356 29876
rect 41412 29820 42812 29876
rect 42868 29820 42878 29876
rect 46834 29820 46844 29876
rect 46900 29820 47740 29876
rect 47796 29820 49644 29876
rect 49700 29820 49710 29876
rect 50306 29820 50316 29876
rect 50372 29820 50428 29932
rect 19826 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20110 29820
rect 50316 29764 50372 29820
rect 50546 29764 50556 29820
rect 50612 29764 50660 29820
rect 50716 29764 50764 29820
rect 50820 29764 50830 29820
rect 31602 29708 31612 29764
rect 31668 29708 32732 29764
rect 32788 29708 32798 29764
rect 47618 29708 47628 29764
rect 47684 29708 50372 29764
rect 0 29652 800 29680
rect 0 29596 1708 29652
rect 1764 29596 2940 29652
rect 2996 29596 3006 29652
rect 11218 29596 11228 29652
rect 11284 29596 14028 29652
rect 14084 29596 14094 29652
rect 21298 29596 21308 29652
rect 21364 29596 21756 29652
rect 21812 29596 21822 29652
rect 30930 29596 30940 29652
rect 30996 29596 32284 29652
rect 32340 29596 32844 29652
rect 32900 29596 32910 29652
rect 36642 29596 36652 29652
rect 36708 29596 44380 29652
rect 44436 29596 45388 29652
rect 45444 29596 45454 29652
rect 46498 29596 46508 29652
rect 46564 29596 48076 29652
rect 48132 29596 48412 29652
rect 48468 29596 48478 29652
rect 0 29568 800 29596
rect 2034 29484 2044 29540
rect 2100 29484 16716 29540
rect 16772 29484 16782 29540
rect 25862 29484 25900 29540
rect 25956 29484 25966 29540
rect 29474 29484 29484 29540
rect 29540 29484 30492 29540
rect 30548 29484 30558 29540
rect 31490 29484 31500 29540
rect 31556 29484 34412 29540
rect 34468 29484 34478 29540
rect 37426 29484 37436 29540
rect 37492 29484 41132 29540
rect 41188 29484 41198 29540
rect 47394 29484 47404 29540
rect 47460 29484 47964 29540
rect 48020 29484 48030 29540
rect 10546 29372 10556 29428
rect 10612 29372 11340 29428
rect 11396 29372 12796 29428
rect 12852 29372 12862 29428
rect 14242 29372 14252 29428
rect 14308 29372 15148 29428
rect 24770 29372 24780 29428
rect 24836 29372 25788 29428
rect 25844 29372 25854 29428
rect 29250 29372 29260 29428
rect 29316 29372 30044 29428
rect 30100 29372 30110 29428
rect 31042 29372 31052 29428
rect 31108 29372 31948 29428
rect 32004 29372 32172 29428
rect 32228 29372 32238 29428
rect 34962 29372 34972 29428
rect 35028 29372 35644 29428
rect 35700 29372 35710 29428
rect 36082 29372 36092 29428
rect 36148 29372 37212 29428
rect 37268 29372 37278 29428
rect 37538 29372 37548 29428
rect 37604 29372 38332 29428
rect 38388 29372 38398 29428
rect 40450 29372 40460 29428
rect 40516 29372 46172 29428
rect 46228 29372 48860 29428
rect 48916 29372 48926 29428
rect 15092 29316 15148 29372
rect 37212 29316 37268 29372
rect 10770 29260 10780 29316
rect 10836 29260 12236 29316
rect 12292 29260 13692 29316
rect 13748 29260 13758 29316
rect 15092 29260 15932 29316
rect 15988 29260 15998 29316
rect 24658 29260 24668 29316
rect 24724 29260 25676 29316
rect 25732 29260 25742 29316
rect 29922 29260 29932 29316
rect 29988 29260 31388 29316
rect 31444 29260 31454 29316
rect 37212 29260 38108 29316
rect 38164 29260 38174 29316
rect 8978 29148 8988 29204
rect 9044 29148 10332 29204
rect 10388 29148 10398 29204
rect 13570 29148 13580 29204
rect 13636 29148 14252 29204
rect 14308 29148 14318 29204
rect 16034 29148 16044 29204
rect 16100 29148 16604 29204
rect 16660 29148 16670 29204
rect 22642 29148 22652 29204
rect 22708 29148 24444 29204
rect 24500 29148 24510 29204
rect 25330 29148 25340 29204
rect 25396 29148 26684 29204
rect 26740 29148 26750 29204
rect 39414 29148 39452 29204
rect 39508 29148 40012 29204
rect 40068 29148 40078 29204
rect 44258 29148 44268 29204
rect 44324 29148 45836 29204
rect 45892 29148 45902 29204
rect 46050 29148 46060 29204
rect 46116 29148 46508 29204
rect 46564 29148 46574 29204
rect 22082 29036 22092 29092
rect 22148 29036 23436 29092
rect 23492 29036 23502 29092
rect 0 28980 800 29008
rect 4466 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4750 29036
rect 35186 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35470 29036
rect 0 28924 1708 28980
rect 1764 28924 2492 28980
rect 2548 28924 2558 28980
rect 0 28896 800 28924
rect 9986 28812 9996 28868
rect 10052 28812 13468 28868
rect 13524 28812 13534 28868
rect 34524 28812 36316 28868
rect 36372 28812 37548 28868
rect 37604 28812 37614 28868
rect 16146 28700 16156 28756
rect 16212 28700 16604 28756
rect 16660 28700 16670 28756
rect 17154 28700 17164 28756
rect 17220 28700 18956 28756
rect 19012 28700 19022 28756
rect 20402 28700 20412 28756
rect 20468 28700 23212 28756
rect 23268 28700 23278 28756
rect 23772 28700 24108 28756
rect 24164 28700 24174 28756
rect 29810 28700 29820 28756
rect 29876 28700 31164 28756
rect 31220 28700 31230 28756
rect 23772 28644 23828 28700
rect 34524 28644 34580 28812
rect 35532 28700 36428 28756
rect 36484 28700 36494 28756
rect 38322 28700 38332 28756
rect 38388 28700 38668 28756
rect 38724 28700 41132 28756
rect 41188 28700 47852 28756
rect 47908 28700 47918 28756
rect 35532 28644 35588 28700
rect 2034 28588 2044 28644
rect 2100 28588 8316 28644
rect 8372 28588 8382 28644
rect 11778 28588 11788 28644
rect 11844 28588 13468 28644
rect 13524 28588 13534 28644
rect 14242 28588 14252 28644
rect 14308 28588 15372 28644
rect 15428 28588 17500 28644
rect 17556 28588 19068 28644
rect 19124 28588 19134 28644
rect 19618 28588 19628 28644
rect 19684 28588 21868 28644
rect 21924 28588 23828 28644
rect 23986 28588 23996 28644
rect 24052 28588 26572 28644
rect 26628 28588 26638 28644
rect 30594 28588 30604 28644
rect 30660 28588 32284 28644
rect 32340 28588 32350 28644
rect 32722 28588 32732 28644
rect 32788 28588 34524 28644
rect 34580 28588 34590 28644
rect 34962 28588 34972 28644
rect 35028 28588 35532 28644
rect 35588 28588 35598 28644
rect 35858 28588 35868 28644
rect 35924 28588 36988 28644
rect 37044 28588 37054 28644
rect 40226 28588 40236 28644
rect 40292 28588 41020 28644
rect 41076 28588 42700 28644
rect 42756 28588 42766 28644
rect 15026 28476 15036 28532
rect 15092 28476 15820 28532
rect 15876 28476 15886 28532
rect 21980 28476 22092 28532
rect 22148 28476 22158 28532
rect 23090 28476 23100 28532
rect 23156 28476 23436 28532
rect 23492 28476 25452 28532
rect 25508 28476 25518 28532
rect 29138 28476 29148 28532
rect 29204 28476 30940 28532
rect 30996 28476 37100 28532
rect 37156 28476 37166 28532
rect 38612 28476 39116 28532
rect 39172 28476 39182 28532
rect 21980 28420 22036 28476
rect 38612 28420 38668 28476
rect 21970 28364 21980 28420
rect 22036 28364 22046 28420
rect 22194 28364 22204 28420
rect 22260 28364 26236 28420
rect 26292 28364 26302 28420
rect 28578 28364 28588 28420
rect 28644 28364 29260 28420
rect 29316 28364 29326 28420
rect 30146 28364 30156 28420
rect 30212 28364 31164 28420
rect 31220 28364 31230 28420
rect 33730 28364 33740 28420
rect 33796 28364 34188 28420
rect 34244 28364 38108 28420
rect 38164 28364 38668 28420
rect 43474 28364 43484 28420
rect 43540 28364 44044 28420
rect 44100 28364 44110 28420
rect 0 28308 800 28336
rect 0 28252 1708 28308
rect 1764 28252 2492 28308
rect 2548 28252 2558 28308
rect 32610 28252 32620 28308
rect 32676 28252 32686 28308
rect 0 28224 800 28252
rect 19826 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20110 28252
rect 32620 28196 32676 28252
rect 50546 28196 50556 28252
rect 50612 28196 50660 28252
rect 50716 28196 50764 28252
rect 50820 28196 50830 28252
rect 21074 28140 21084 28196
rect 21140 28140 24724 28196
rect 32162 28140 32172 28196
rect 32228 28140 32676 28196
rect 34962 28140 34972 28196
rect 35028 28140 35196 28196
rect 35252 28140 35262 28196
rect 36642 28140 36652 28196
rect 36708 28140 36988 28196
rect 37044 28140 37054 28196
rect 42466 28140 42476 28196
rect 42532 28140 43484 28196
rect 43540 28140 43550 28196
rect 21084 28084 21140 28140
rect 24668 28084 24724 28140
rect 12786 28028 12796 28084
rect 12852 28028 14364 28084
rect 14420 28028 14924 28084
rect 14980 28028 14990 28084
rect 16706 28028 16716 28084
rect 16772 28028 17500 28084
rect 17556 28028 21140 28084
rect 22530 28028 22540 28084
rect 22596 28028 23324 28084
rect 23380 28028 23390 28084
rect 24658 28028 24668 28084
rect 24724 28028 25228 28084
rect 25284 28028 25294 28084
rect 25890 28028 25900 28084
rect 25956 28028 26796 28084
rect 26852 28028 27132 28084
rect 27188 28028 27198 28084
rect 27906 28028 27916 28084
rect 27972 28028 29484 28084
rect 29540 28028 29708 28084
rect 29764 28028 30604 28084
rect 30660 28028 38668 28084
rect 40002 28028 40012 28084
rect 40068 28028 40908 28084
rect 40964 28028 40974 28084
rect 45154 28028 45164 28084
rect 45220 28028 45724 28084
rect 45780 28028 45790 28084
rect 38612 27972 38668 28028
rect 2034 27916 2044 27972
rect 2100 27916 8988 27972
rect 9044 27916 9054 27972
rect 21522 27916 21532 27972
rect 21588 27916 23548 27972
rect 23604 27916 23614 27972
rect 29810 27916 29820 27972
rect 29876 27916 30156 27972
rect 30212 27916 32284 27972
rect 32340 27916 32350 27972
rect 36614 27916 36652 27972
rect 36708 27916 36718 27972
rect 38612 27916 39788 27972
rect 39844 27916 45388 27972
rect 45444 27916 45454 27972
rect 12338 27804 12348 27860
rect 12404 27804 15596 27860
rect 15652 27804 15662 27860
rect 22978 27804 22988 27860
rect 23044 27804 25564 27860
rect 25620 27804 25630 27860
rect 29026 27804 29036 27860
rect 29092 27804 30268 27860
rect 30324 27804 30334 27860
rect 32610 27804 32620 27860
rect 32676 27804 33516 27860
rect 33572 27804 33582 27860
rect 40338 27804 40348 27860
rect 40404 27804 41244 27860
rect 41300 27804 41692 27860
rect 41748 27804 41758 27860
rect 48066 27804 48076 27860
rect 48132 27804 48748 27860
rect 48804 27804 48814 27860
rect 12562 27692 12572 27748
rect 12628 27692 15148 27748
rect 15204 27692 15214 27748
rect 19842 27692 19852 27748
rect 19908 27692 22428 27748
rect 22484 27692 22494 27748
rect 27570 27692 27580 27748
rect 27636 27692 28476 27748
rect 28532 27692 28542 27748
rect 46834 27692 46844 27748
rect 46900 27692 47964 27748
rect 48020 27692 48030 27748
rect 0 27636 800 27664
rect 0 27580 1708 27636
rect 1764 27580 2492 27636
rect 2548 27580 2558 27636
rect 2706 27580 2716 27636
rect 2772 27580 13692 27636
rect 13748 27580 13758 27636
rect 21634 27580 21644 27636
rect 21700 27580 22540 27636
rect 22596 27580 23212 27636
rect 23268 27580 23278 27636
rect 41234 27580 41244 27636
rect 41300 27580 45052 27636
rect 45108 27580 45118 27636
rect 0 27552 800 27580
rect 21970 27468 21980 27524
rect 22036 27468 22428 27524
rect 22484 27468 25228 27524
rect 25284 27468 25294 27524
rect 4466 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4750 27468
rect 35186 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35470 27468
rect 8306 27356 8316 27412
rect 8372 27356 17612 27412
rect 17668 27356 17678 27412
rect 20738 27356 20748 27412
rect 20804 27356 23324 27412
rect 23380 27356 23390 27412
rect 33282 27356 33292 27412
rect 33348 27356 34412 27412
rect 34468 27356 34478 27412
rect 34710 27356 34748 27412
rect 34804 27356 34814 27412
rect 12114 27244 12124 27300
rect 12180 27244 12796 27300
rect 12852 27244 14140 27300
rect 14196 27244 14206 27300
rect 23398 27244 23436 27300
rect 23492 27244 23502 27300
rect 23958 27244 23996 27300
rect 24052 27244 24062 27300
rect 24210 27244 24220 27300
rect 24276 27244 25116 27300
rect 25172 27244 25900 27300
rect 25956 27244 26348 27300
rect 26404 27244 26414 27300
rect 33730 27244 33740 27300
rect 33796 27244 35196 27300
rect 35252 27244 35262 27300
rect 43474 27244 43484 27300
rect 43540 27244 43932 27300
rect 43988 27244 44492 27300
rect 44548 27244 44558 27300
rect 11218 27132 11228 27188
rect 11284 27132 12572 27188
rect 12628 27132 12638 27188
rect 20850 27132 20860 27188
rect 20916 27132 22204 27188
rect 22260 27132 22270 27188
rect 22642 27132 22652 27188
rect 22708 27132 24108 27188
rect 24164 27132 24174 27188
rect 25442 27132 25452 27188
rect 25508 27132 32508 27188
rect 32564 27132 41580 27188
rect 41636 27132 42476 27188
rect 42532 27132 46172 27188
rect 46228 27132 46238 27188
rect 46722 27132 46732 27188
rect 46788 27132 47740 27188
rect 47796 27132 48524 27188
rect 48580 27132 50428 27188
rect 50484 27132 50494 27188
rect 14018 27020 14028 27076
rect 14084 27020 14094 27076
rect 14466 27020 14476 27076
rect 14532 27020 15484 27076
rect 15540 27020 15550 27076
rect 23538 27020 23548 27076
rect 23604 27020 24220 27076
rect 24276 27020 24286 27076
rect 27682 27020 27692 27076
rect 27748 27020 33292 27076
rect 33348 27020 33358 27076
rect 34178 27020 34188 27076
rect 34244 27020 34524 27076
rect 34580 27020 34590 27076
rect 34850 27020 34860 27076
rect 34916 27020 35756 27076
rect 35812 27020 35822 27076
rect 37324 27020 37772 27076
rect 37828 27020 37838 27076
rect 38546 27020 38556 27076
rect 38612 27020 39396 27076
rect 40338 27020 40348 27076
rect 40404 27020 42140 27076
rect 42196 27020 43260 27076
rect 43316 27020 43326 27076
rect 46050 27020 46060 27076
rect 46116 27020 47404 27076
rect 47460 27020 47470 27076
rect 0 26964 800 26992
rect 14028 26964 14084 27020
rect 37324 26964 37380 27020
rect 0 26908 1708 26964
rect 1764 26908 2492 26964
rect 2548 26908 2558 26964
rect 6514 26908 6524 26964
rect 6580 26908 8428 26964
rect 8484 26908 8494 26964
rect 13570 26908 13580 26964
rect 13636 26908 14084 26964
rect 16258 26908 16268 26964
rect 16324 26908 16940 26964
rect 16996 26908 17006 26964
rect 18274 26908 18284 26964
rect 18340 26908 18732 26964
rect 18788 26908 20076 26964
rect 20132 26908 20142 26964
rect 21298 26908 21308 26964
rect 21364 26908 24108 26964
rect 24164 26908 24556 26964
rect 24612 26908 24622 26964
rect 26338 26908 26348 26964
rect 26404 26908 28140 26964
rect 28196 26908 28206 26964
rect 34738 26908 34748 26964
rect 34804 26908 35308 26964
rect 35364 26908 35374 26964
rect 35522 26908 35532 26964
rect 35588 26908 36316 26964
rect 36372 26908 37324 26964
rect 37380 26908 37390 26964
rect 37538 26908 37548 26964
rect 37604 26908 39116 26964
rect 39172 26908 39182 26964
rect 39340 26908 39396 27020
rect 48178 26908 48188 26964
rect 48244 26908 48972 26964
rect 49028 26908 49038 26964
rect 49746 26908 49756 26964
rect 49812 26908 50652 26964
rect 50708 26908 50718 26964
rect 0 26880 800 26908
rect 39330 26852 39340 26908
rect 39396 26852 39406 26908
rect 1932 26796 2044 26852
rect 2100 26796 2110 26852
rect 2370 26796 2380 26852
rect 2436 26796 3164 26852
rect 3220 26796 3230 26852
rect 18498 26796 18508 26852
rect 18564 26796 19068 26852
rect 19124 26796 19134 26852
rect 22418 26796 22428 26852
rect 22484 26796 23884 26852
rect 23940 26796 23950 26852
rect 37986 26796 37996 26852
rect 38052 26796 39004 26852
rect 39060 26796 39070 26852
rect 40002 26796 40012 26852
rect 40068 26796 42028 26852
rect 42084 26796 42094 26852
rect 44930 26796 44940 26852
rect 44996 26796 45612 26852
rect 45668 26796 45678 26852
rect 45826 26796 45836 26852
rect 45892 26796 46508 26852
rect 46564 26796 46574 26852
rect 1932 26628 1988 26796
rect 2146 26684 2156 26740
rect 2212 26684 19180 26740
rect 19236 26684 19246 26740
rect 19826 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20110 26684
rect 50546 26628 50556 26684
rect 50612 26628 50660 26684
rect 50716 26628 50764 26684
rect 50820 26628 50830 26684
rect 1932 26572 17612 26628
rect 17668 26572 17678 26628
rect 18834 26572 18844 26628
rect 18900 26572 19628 26628
rect 19684 26572 19694 26628
rect 28018 26572 28028 26628
rect 28084 26572 37212 26628
rect 37268 26572 38332 26628
rect 38388 26572 38398 26628
rect 11106 26460 11116 26516
rect 11172 26460 12012 26516
rect 12068 26460 12078 26516
rect 15362 26460 15372 26516
rect 15428 26460 16604 26516
rect 16660 26460 16670 26516
rect 23398 26460 23436 26516
rect 23492 26460 23502 26516
rect 23650 26460 23660 26516
rect 23716 26460 24780 26516
rect 24836 26460 25116 26516
rect 25172 26460 25182 26516
rect 25974 26460 26012 26516
rect 26068 26460 26078 26516
rect 26786 26460 26796 26516
rect 26852 26460 27132 26516
rect 27188 26460 27198 26516
rect 48066 26460 48076 26516
rect 48132 26460 49644 26516
rect 49700 26460 49710 26516
rect 11666 26348 11676 26404
rect 11732 26348 13020 26404
rect 13076 26348 14700 26404
rect 14756 26348 14766 26404
rect 19058 26348 19068 26404
rect 19124 26348 21532 26404
rect 21588 26348 21598 26404
rect 21756 26348 23324 26404
rect 23380 26348 25452 26404
rect 25508 26348 25518 26404
rect 25778 26348 25788 26404
rect 25844 26348 27580 26404
rect 27636 26348 29260 26404
rect 29316 26348 29326 26404
rect 35186 26348 35196 26404
rect 35252 26348 39340 26404
rect 39396 26348 39406 26404
rect 48374 26348 48412 26404
rect 48468 26348 48478 26404
rect 0 26292 800 26320
rect 21756 26292 21812 26348
rect 0 26236 2380 26292
rect 2436 26236 2446 26292
rect 17378 26236 17388 26292
rect 17444 26236 18060 26292
rect 18116 26236 20412 26292
rect 20468 26236 20478 26292
rect 21634 26236 21644 26292
rect 21700 26236 21812 26292
rect 22306 26236 22316 26292
rect 22372 26236 24220 26292
rect 24276 26236 24286 26292
rect 33282 26236 33292 26292
rect 33348 26236 34300 26292
rect 34356 26236 34366 26292
rect 36082 26236 36092 26292
rect 36148 26236 36316 26292
rect 36372 26236 37884 26292
rect 37940 26236 37950 26292
rect 42354 26236 42364 26292
rect 42420 26236 43148 26292
rect 43204 26236 47068 26292
rect 47124 26236 47740 26292
rect 47796 26236 47806 26292
rect 48066 26236 48076 26292
rect 48132 26236 48748 26292
rect 48804 26236 49532 26292
rect 49588 26236 49598 26292
rect 0 26208 800 26236
rect 1698 26124 1708 26180
rect 1764 26124 2940 26180
rect 2996 26124 3006 26180
rect 16146 26124 16156 26180
rect 16212 26124 16492 26180
rect 16548 26124 18508 26180
rect 18564 26124 18574 26180
rect 19170 26124 19180 26180
rect 19236 26124 20636 26180
rect 20692 26124 20702 26180
rect 26852 26124 27244 26180
rect 27300 26124 30716 26180
rect 30772 26124 30782 26180
rect 33394 26124 33404 26180
rect 33460 26124 34748 26180
rect 34804 26124 34972 26180
rect 35028 26124 35038 26180
rect 35858 26124 35868 26180
rect 35924 26124 36876 26180
rect 36932 26124 36942 26180
rect 42690 26124 42700 26180
rect 42756 26124 43932 26180
rect 43988 26124 43998 26180
rect 48486 26124 48524 26180
rect 48580 26124 48590 26180
rect 26852 26068 26908 26124
rect 11330 26012 11340 26068
rect 11396 26012 14924 26068
rect 14980 26012 15820 26068
rect 15876 26012 15886 26068
rect 17042 26012 17052 26068
rect 17108 26012 17948 26068
rect 18004 26012 18014 26068
rect 18162 26012 18172 26068
rect 18228 26012 20972 26068
rect 21028 26012 21038 26068
rect 26562 26012 26572 26068
rect 26628 26012 26908 26068
rect 45266 26012 45276 26068
rect 45332 26012 57036 26068
rect 57092 26012 57102 26068
rect 15148 25900 26348 25956
rect 26404 25900 26414 25956
rect 42914 25900 42924 25956
rect 42980 25900 46620 25956
rect 46676 25900 46686 25956
rect 48066 25900 48076 25956
rect 48132 25900 50316 25956
rect 50372 25900 50382 25956
rect 4466 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4750 25900
rect 15148 25732 15204 25900
rect 35186 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35470 25900
rect 19730 25788 19740 25844
rect 19796 25788 23100 25844
rect 23156 25788 23166 25844
rect 24434 25788 24444 25844
rect 24500 25788 28140 25844
rect 28196 25788 28206 25844
rect 12786 25676 12796 25732
rect 12852 25676 13468 25732
rect 13524 25676 13534 25732
rect 14914 25676 14924 25732
rect 14980 25676 15148 25732
rect 15204 25676 15214 25732
rect 18172 25676 26460 25732
rect 26516 25676 26526 25732
rect 0 25620 800 25648
rect 18172 25620 18228 25676
rect 0 25564 1708 25620
rect 1764 25564 1774 25620
rect 14690 25564 14700 25620
rect 14756 25564 18228 25620
rect 18386 25564 18396 25620
rect 18452 25564 19516 25620
rect 19572 25564 21644 25620
rect 21700 25564 21710 25620
rect 23986 25564 23996 25620
rect 24052 25564 24332 25620
rect 24388 25564 24398 25620
rect 0 25536 800 25564
rect 2034 25452 2044 25508
rect 2100 25452 10444 25508
rect 10500 25452 10510 25508
rect 14242 25452 14252 25508
rect 14308 25452 15372 25508
rect 15428 25452 15438 25508
rect 16818 25452 16828 25508
rect 16884 25452 18732 25508
rect 18788 25452 19404 25508
rect 19460 25452 19470 25508
rect 27682 25452 27692 25508
rect 27748 25452 28140 25508
rect 28196 25452 28206 25508
rect 30706 25452 30716 25508
rect 30772 25452 36204 25508
rect 36260 25452 36270 25508
rect 28130 25340 28140 25396
rect 28196 25340 28364 25396
rect 28420 25340 28430 25396
rect 30482 25340 30492 25396
rect 30548 25340 31724 25396
rect 31780 25340 31790 25396
rect 32162 25340 32172 25396
rect 32228 25340 34188 25396
rect 34244 25340 34254 25396
rect 57586 25340 57596 25396
rect 57652 25340 58156 25396
rect 58212 25340 58222 25396
rect 20178 25228 20188 25284
rect 20244 25228 21532 25284
rect 21588 25228 21598 25284
rect 33842 25228 33852 25284
rect 33908 25228 35868 25284
rect 35924 25228 40236 25284
rect 40292 25228 41020 25284
rect 41076 25228 41086 25284
rect 43586 25228 43596 25284
rect 43652 25228 44940 25284
rect 44996 25228 45006 25284
rect 55412 25228 57820 25284
rect 57876 25228 57886 25284
rect 21858 25116 21868 25172
rect 21924 25116 22764 25172
rect 22820 25116 22830 25172
rect 44370 25116 44380 25172
rect 44436 25116 45836 25172
rect 45892 25116 46844 25172
rect 46900 25116 46910 25172
rect 19826 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20110 25116
rect 50546 25060 50556 25116
rect 50612 25060 50660 25116
rect 50716 25060 50764 25116
rect 50820 25060 50830 25116
rect 12898 25004 12908 25060
rect 12964 25004 14252 25060
rect 14308 25004 14318 25060
rect 25442 25004 25452 25060
rect 25508 25004 26572 25060
rect 26628 25004 31052 25060
rect 31108 25004 31118 25060
rect 31714 25004 31724 25060
rect 31780 25004 33964 25060
rect 34020 25004 34748 25060
rect 34804 25004 35196 25060
rect 35252 25004 35262 25060
rect 36754 25004 36764 25060
rect 36820 25004 46956 25060
rect 47012 25004 47022 25060
rect 0 24948 800 24976
rect 55412 24948 55468 25228
rect 59200 24948 60000 24976
rect 0 24892 1708 24948
rect 1764 24892 2492 24948
rect 2548 24892 2558 24948
rect 10210 24892 10220 24948
rect 10276 24892 11228 24948
rect 11284 24892 14588 24948
rect 14644 24892 14654 24948
rect 22082 24892 22092 24948
rect 22148 24892 24556 24948
rect 24612 24892 24622 24948
rect 34066 24892 34076 24948
rect 34132 24892 34748 24948
rect 34804 24892 34814 24948
rect 43362 24892 43372 24948
rect 43428 24892 55468 24948
rect 57026 24892 57036 24948
rect 57092 24892 57820 24948
rect 57876 24892 57886 24948
rect 58146 24892 58156 24948
rect 58212 24892 60000 24948
rect 0 24864 800 24892
rect 59200 24864 60000 24892
rect 8306 24780 8316 24836
rect 8372 24780 10108 24836
rect 10164 24780 10174 24836
rect 23874 24780 23884 24836
rect 23940 24780 24556 24836
rect 24612 24780 24622 24836
rect 26852 24780 31500 24836
rect 31556 24780 31566 24836
rect 33282 24780 33292 24836
rect 33348 24780 33460 24836
rect 33954 24780 33964 24836
rect 34020 24780 34860 24836
rect 34916 24780 34926 24836
rect 44146 24780 44156 24836
rect 44212 24780 44828 24836
rect 44884 24780 44894 24836
rect 48178 24780 48188 24836
rect 48244 24780 49868 24836
rect 49924 24780 49934 24836
rect 26852 24724 26908 24780
rect 8978 24668 8988 24724
rect 9044 24668 11788 24724
rect 11844 24668 11854 24724
rect 21410 24668 21420 24724
rect 21476 24668 26908 24724
rect 30258 24668 30268 24724
rect 30324 24668 31948 24724
rect 32004 24668 33068 24724
rect 33124 24668 33134 24724
rect 33404 24612 33460 24780
rect 49410 24668 49420 24724
rect 49476 24668 50540 24724
rect 50596 24668 50606 24724
rect 6290 24556 6300 24612
rect 6356 24556 8764 24612
rect 8820 24556 8830 24612
rect 11106 24556 11116 24612
rect 11172 24556 11676 24612
rect 11732 24556 11742 24612
rect 17714 24556 17724 24612
rect 17780 24556 21868 24612
rect 21924 24556 21934 24612
rect 29026 24556 29036 24612
rect 29092 24556 31948 24612
rect 32004 24556 32396 24612
rect 32452 24556 32462 24612
rect 33394 24556 33404 24612
rect 33460 24556 33470 24612
rect 34178 24556 34188 24612
rect 34244 24556 34636 24612
rect 34692 24556 34702 24612
rect 43698 24556 43708 24612
rect 43764 24556 44716 24612
rect 44772 24556 44782 24612
rect 20290 24444 20300 24500
rect 20356 24444 20748 24500
rect 20804 24444 22652 24500
rect 22708 24444 23884 24500
rect 23940 24444 23950 24500
rect 43026 24444 43036 24500
rect 43092 24444 43596 24500
rect 43652 24444 43662 24500
rect 0 24276 800 24304
rect 4466 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4750 24332
rect 35186 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35470 24332
rect 59200 24276 60000 24304
rect 0 24220 1708 24276
rect 1764 24220 2492 24276
rect 2548 24220 2558 24276
rect 58146 24220 58156 24276
rect 58212 24220 60000 24276
rect 0 24192 800 24220
rect 59200 24192 60000 24220
rect 34626 24108 34636 24164
rect 34692 24108 35084 24164
rect 35140 24108 37100 24164
rect 37156 24108 38780 24164
rect 38836 24108 40460 24164
rect 40516 24108 40526 24164
rect 11218 23996 11228 24052
rect 11284 23996 12124 24052
rect 12180 23996 12190 24052
rect 22978 23996 22988 24052
rect 23044 23996 23660 24052
rect 23716 23996 25116 24052
rect 25172 23996 25182 24052
rect 26114 23996 26124 24052
rect 26180 23996 28252 24052
rect 28308 23996 28318 24052
rect 32722 23996 32732 24052
rect 32788 23996 33292 24052
rect 33348 23996 33358 24052
rect 39106 23996 39116 24052
rect 39172 23996 40348 24052
rect 40404 23996 41692 24052
rect 41748 23996 41758 24052
rect 7634 23884 7644 23940
rect 7700 23884 9324 23940
rect 9380 23884 11788 23940
rect 11844 23884 11854 23940
rect 15026 23884 15036 23940
rect 15092 23884 17276 23940
rect 17332 23884 17724 23940
rect 17780 23884 17790 23940
rect 19058 23884 19068 23940
rect 19124 23884 37436 23940
rect 37492 23884 37996 23940
rect 38052 23884 39228 23940
rect 39284 23884 40236 23940
rect 40292 23884 40302 23940
rect 47282 23884 47292 23940
rect 47348 23884 48860 23940
rect 48916 23884 50092 23940
rect 50148 23884 50988 23940
rect 51044 23884 51054 23940
rect 2034 23772 2044 23828
rect 2100 23772 6972 23828
rect 7028 23772 7038 23828
rect 8082 23772 8092 23828
rect 8148 23772 8764 23828
rect 8820 23772 8830 23828
rect 12114 23772 12124 23828
rect 12180 23772 12908 23828
rect 12964 23772 13692 23828
rect 13748 23772 13758 23828
rect 24434 23772 24444 23828
rect 24500 23772 25564 23828
rect 25620 23772 25630 23828
rect 28578 23772 28588 23828
rect 28644 23772 29596 23828
rect 29652 23772 29662 23828
rect 32274 23772 32284 23828
rect 32340 23772 33740 23828
rect 33796 23772 36988 23828
rect 37044 23772 37054 23828
rect 37314 23772 37324 23828
rect 37380 23772 38668 23828
rect 38724 23772 38734 23828
rect 41234 23772 41244 23828
rect 41300 23772 43932 23828
rect 43988 23772 43998 23828
rect 46834 23772 46844 23828
rect 46900 23772 47852 23828
rect 47908 23772 47918 23828
rect 49410 23772 49420 23828
rect 49476 23772 49868 23828
rect 49924 23772 50428 23828
rect 50484 23772 50494 23828
rect 9986 23660 9996 23716
rect 10052 23660 11228 23716
rect 11284 23660 12348 23716
rect 12404 23660 12414 23716
rect 15586 23660 15596 23716
rect 15652 23660 20356 23716
rect 29922 23660 29932 23716
rect 29988 23660 31164 23716
rect 31220 23660 34524 23716
rect 34580 23660 35196 23716
rect 35252 23660 35262 23716
rect 42802 23660 42812 23716
rect 42868 23660 44044 23716
rect 44100 23660 44110 23716
rect 50194 23660 50204 23716
rect 50260 23660 50652 23716
rect 50708 23660 50718 23716
rect 55412 23660 57820 23716
rect 57876 23660 57886 23716
rect 0 23604 800 23632
rect 20300 23604 20356 23660
rect 0 23548 1708 23604
rect 1764 23548 2492 23604
rect 2548 23548 2558 23604
rect 7746 23548 7756 23604
rect 7812 23548 9212 23604
rect 9268 23548 9660 23604
rect 9716 23548 9726 23604
rect 20290 23548 20300 23604
rect 20356 23548 20636 23604
rect 20692 23548 20702 23604
rect 35746 23548 35756 23604
rect 35812 23548 36764 23604
rect 36820 23548 36830 23604
rect 42018 23548 42028 23604
rect 42084 23548 43372 23604
rect 43428 23548 44156 23604
rect 44212 23548 47068 23604
rect 47124 23548 47134 23604
rect 49634 23548 49644 23604
rect 49700 23548 50316 23604
rect 50372 23548 50382 23604
rect 0 23520 800 23548
rect 19826 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20110 23548
rect 50546 23492 50556 23548
rect 50612 23492 50660 23548
rect 50716 23492 50764 23548
rect 50820 23492 50830 23548
rect 7186 23436 7196 23492
rect 7252 23436 10332 23492
rect 10388 23436 10398 23492
rect 21634 23436 21644 23492
rect 21700 23436 22260 23492
rect 26450 23436 26460 23492
rect 26516 23436 27188 23492
rect 27458 23436 27468 23492
rect 27524 23436 28252 23492
rect 28308 23436 28318 23492
rect 43250 23436 43260 23492
rect 43316 23436 44940 23492
rect 44996 23436 45836 23492
rect 45892 23436 45902 23492
rect 49858 23436 49868 23492
rect 49924 23436 50204 23492
rect 50260 23436 50270 23492
rect 22204 23380 22260 23436
rect 27132 23380 27188 23436
rect 55412 23380 55468 23660
rect 59200 23604 60000 23632
rect 57586 23548 57596 23604
rect 57652 23548 58156 23604
rect 58212 23548 60000 23604
rect 59200 23520 60000 23548
rect 13794 23324 13804 23380
rect 13860 23324 14364 23380
rect 14420 23324 16156 23380
rect 16212 23324 16222 23380
rect 21830 23324 21868 23380
rect 21924 23324 21934 23380
rect 22194 23324 22204 23380
rect 22260 23324 22988 23380
rect 23044 23324 23054 23380
rect 26338 23324 26348 23380
rect 26404 23324 26908 23380
rect 27132 23324 27356 23380
rect 27412 23324 27422 23380
rect 43026 23324 43036 23380
rect 43092 23324 44604 23380
rect 44660 23324 44670 23380
rect 46386 23324 46396 23380
rect 46452 23324 55468 23380
rect 26852 23268 26908 23324
rect 18498 23212 18508 23268
rect 18564 23212 20972 23268
rect 21028 23212 22652 23268
rect 22708 23212 24556 23268
rect 24612 23212 24622 23268
rect 26852 23212 27692 23268
rect 27748 23212 28364 23268
rect 28420 23212 28430 23268
rect 31826 23212 31836 23268
rect 31892 23212 35644 23268
rect 35700 23212 36316 23268
rect 36372 23212 36382 23268
rect 39778 23212 39788 23268
rect 39844 23212 41580 23268
rect 41636 23212 42924 23268
rect 42980 23212 42990 23268
rect 45266 23212 45276 23268
rect 45332 23212 47852 23268
rect 47908 23212 47918 23268
rect 2146 23100 2156 23156
rect 2212 23100 9772 23156
rect 9828 23100 9838 23156
rect 12226 23100 12236 23156
rect 12292 23100 13020 23156
rect 13076 23100 13468 23156
rect 13524 23100 13534 23156
rect 20290 23100 20300 23156
rect 20356 23100 22540 23156
rect 22596 23100 23548 23156
rect 23604 23100 25340 23156
rect 25396 23100 25406 23156
rect 27122 23100 27132 23156
rect 27188 23100 27804 23156
rect 27860 23100 27870 23156
rect 41458 23100 41468 23156
rect 41524 23100 42140 23156
rect 42196 23100 42206 23156
rect 42578 23100 42588 23156
rect 42644 23100 43148 23156
rect 43204 23100 44940 23156
rect 44996 23100 45006 23156
rect 45826 23100 45836 23156
rect 45892 23100 47292 23156
rect 47348 23100 47358 23156
rect 6066 22988 6076 23044
rect 6132 22988 6972 23044
rect 7028 22988 7038 23044
rect 22866 22988 22876 23044
rect 22932 22988 23772 23044
rect 23828 22988 23838 23044
rect 26114 22988 26124 23044
rect 26180 22988 26908 23044
rect 26964 22988 26974 23044
rect 27234 22988 27244 23044
rect 27300 22988 27804 23044
rect 27860 22988 27870 23044
rect 28914 22988 28924 23044
rect 28980 22988 30156 23044
rect 30212 22988 30828 23044
rect 30884 22988 30894 23044
rect 46162 22988 46172 23044
rect 46228 22988 48748 23044
rect 48804 22988 48814 23044
rect 0 22932 800 22960
rect 0 22876 1708 22932
rect 1764 22876 2492 22932
rect 2548 22876 2558 22932
rect 14914 22876 14924 22932
rect 14980 22876 14990 22932
rect 37100 22876 40908 22932
rect 40964 22876 41244 22932
rect 41300 22876 41310 22932
rect 43474 22876 43484 22932
rect 43540 22876 43932 22932
rect 43988 22876 43998 22932
rect 0 22848 800 22876
rect 4466 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4750 22764
rect 14924 22484 14980 22876
rect 37100 22820 37156 22876
rect 19618 22764 19628 22820
rect 19684 22764 20524 22820
rect 20580 22764 20590 22820
rect 27122 22764 27132 22820
rect 27188 22764 27356 22820
rect 27412 22764 27422 22820
rect 36418 22764 36428 22820
rect 36484 22764 37100 22820
rect 37156 22764 37166 22820
rect 35186 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35470 22764
rect 23202 22652 23212 22708
rect 23268 22652 26572 22708
rect 26628 22652 31164 22708
rect 31220 22652 31230 22708
rect 24546 22540 24556 22596
rect 24612 22540 40796 22596
rect 40852 22540 40862 22596
rect 7074 22428 7084 22484
rect 7140 22428 7756 22484
rect 7812 22428 7822 22484
rect 8418 22428 8428 22484
rect 8484 22428 8988 22484
rect 9044 22428 11788 22484
rect 11844 22428 11854 22484
rect 14914 22428 14924 22484
rect 14980 22428 14990 22484
rect 23426 22428 23436 22484
rect 23492 22428 24332 22484
rect 24388 22428 24398 22484
rect 26338 22428 26348 22484
rect 26404 22428 26796 22484
rect 26852 22428 28140 22484
rect 28196 22428 28206 22484
rect 30706 22428 30716 22484
rect 30772 22428 33180 22484
rect 33236 22428 33246 22484
rect 35634 22428 35644 22484
rect 35700 22428 36764 22484
rect 36820 22428 36830 22484
rect 38994 22428 39004 22484
rect 39060 22428 42140 22484
rect 42196 22428 42812 22484
rect 42868 22428 42878 22484
rect 2034 22316 2044 22372
rect 2100 22316 10108 22372
rect 10164 22316 10174 22372
rect 18386 22316 18396 22372
rect 18452 22316 19628 22372
rect 19684 22316 21420 22372
rect 21476 22316 21486 22372
rect 22754 22316 22764 22372
rect 22820 22316 25228 22372
rect 25284 22316 25676 22372
rect 25732 22316 27692 22372
rect 27748 22316 27758 22372
rect 30818 22316 30828 22372
rect 30884 22316 32396 22372
rect 32452 22316 32462 22372
rect 36306 22316 36316 22372
rect 36372 22316 37548 22372
rect 37604 22316 37614 22372
rect 44818 22316 44828 22372
rect 44884 22316 46172 22372
rect 46228 22316 46238 22372
rect 47506 22316 47516 22372
rect 47572 22316 48972 22372
rect 49028 22316 49038 22372
rect 0 22260 800 22288
rect 0 22204 1708 22260
rect 1764 22204 2492 22260
rect 2548 22204 2558 22260
rect 57586 22204 57596 22260
rect 57652 22204 58156 22260
rect 58212 22204 58222 22260
rect 0 22176 800 22204
rect 10994 22092 11004 22148
rect 11060 22092 13468 22148
rect 13524 22092 13534 22148
rect 31826 22092 31836 22148
rect 31892 22092 32396 22148
rect 32452 22092 32462 22148
rect 45266 22092 45276 22148
rect 45332 22092 45948 22148
rect 46004 22092 46508 22148
rect 46564 22092 46574 22148
rect 55412 22092 57820 22148
rect 57876 22092 57886 22148
rect 9986 21980 9996 22036
rect 10052 21980 11228 22036
rect 11284 21980 13916 22036
rect 13972 21980 15148 22036
rect 15204 21980 15214 22036
rect 29138 21980 29148 22036
rect 29204 21980 30268 22036
rect 30324 21980 30334 22036
rect 45042 21980 45052 22036
rect 45108 21980 46620 22036
rect 46676 21980 46686 22036
rect 19826 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20110 21980
rect 50546 21924 50556 21980
rect 50612 21924 50660 21980
rect 50716 21924 50764 21980
rect 50820 21924 50830 21980
rect 55412 21924 55468 22092
rect 24882 21868 24892 21924
rect 24948 21868 27244 21924
rect 27300 21868 27310 21924
rect 27794 21868 27804 21924
rect 27860 21868 29876 21924
rect 34402 21868 34412 21924
rect 34468 21868 36876 21924
rect 36932 21868 40796 21924
rect 40852 21868 40862 21924
rect 41010 21868 41020 21924
rect 41076 21868 41916 21924
rect 41972 21868 42588 21924
rect 42644 21868 42654 21924
rect 43586 21868 43596 21924
rect 43652 21868 44604 21924
rect 44660 21868 44670 21924
rect 53778 21868 53788 21924
rect 53844 21868 55468 21924
rect 1820 21756 2380 21812
rect 2436 21756 3164 21812
rect 3220 21756 3230 21812
rect 18162 21756 18172 21812
rect 18228 21756 19068 21812
rect 19124 21756 19134 21812
rect 23090 21756 23100 21812
rect 23156 21756 28588 21812
rect 28644 21756 28654 21812
rect 0 21588 800 21616
rect 1820 21588 1876 21756
rect 29820 21700 29876 21868
rect 31154 21756 31164 21812
rect 31220 21756 33068 21812
rect 33124 21756 33134 21812
rect 34962 21756 34972 21812
rect 35028 21756 35868 21812
rect 35924 21756 37996 21812
rect 38052 21756 38062 21812
rect 38322 21756 38332 21812
rect 38388 21756 40124 21812
rect 40180 21756 40190 21812
rect 41458 21756 41468 21812
rect 41524 21756 42140 21812
rect 42196 21756 42206 21812
rect 2034 21644 2044 21700
rect 2100 21644 14308 21700
rect 17714 21644 17724 21700
rect 17780 21644 19516 21700
rect 19572 21644 21868 21700
rect 21924 21644 23324 21700
rect 23380 21644 23390 21700
rect 24434 21644 24444 21700
rect 24500 21644 25004 21700
rect 25060 21644 25452 21700
rect 25508 21644 26012 21700
rect 26068 21644 26078 21700
rect 27010 21644 27020 21700
rect 27076 21644 27086 21700
rect 29820 21644 36428 21700
rect 36484 21644 42252 21700
rect 42308 21644 42318 21700
rect 0 21532 1876 21588
rect 2146 21532 2156 21588
rect 2212 21532 6524 21588
rect 6580 21532 6590 21588
rect 7858 21532 7868 21588
rect 7924 21532 9212 21588
rect 9268 21532 9278 21588
rect 0 21504 800 21532
rect 14252 21476 14308 21644
rect 23538 21532 23548 21588
rect 23604 21532 24332 21588
rect 24388 21532 24398 21588
rect 24556 21532 26460 21588
rect 26516 21532 26526 21588
rect 24556 21476 24612 21532
rect 27020 21476 27076 21644
rect 59200 21588 60000 21616
rect 30482 21532 30492 21588
rect 30548 21532 31500 21588
rect 31556 21532 31566 21588
rect 34962 21532 34972 21588
rect 35028 21532 35196 21588
rect 35252 21532 35262 21588
rect 38546 21532 38556 21588
rect 38612 21532 40012 21588
rect 40068 21532 40460 21588
rect 40516 21532 40526 21588
rect 46162 21532 46172 21588
rect 46228 21532 46844 21588
rect 46900 21532 47292 21588
rect 47348 21532 47358 21588
rect 58146 21532 58156 21588
rect 58212 21532 60000 21588
rect 59200 21504 60000 21532
rect 1698 21420 1708 21476
rect 1764 21420 2940 21476
rect 2996 21420 3006 21476
rect 8978 21420 8988 21476
rect 9044 21420 9660 21476
rect 9716 21420 9726 21476
rect 14242 21420 14252 21476
rect 14308 21420 14318 21476
rect 20402 21420 20412 21476
rect 20468 21420 22316 21476
rect 22372 21420 22382 21476
rect 24098 21420 24108 21476
rect 24164 21420 24612 21476
rect 25554 21420 25564 21476
rect 25620 21420 26684 21476
rect 26740 21420 26750 21476
rect 27010 21420 27020 21476
rect 27076 21420 27086 21476
rect 30034 21420 30044 21476
rect 30100 21420 30604 21476
rect 30660 21420 30670 21476
rect 38098 21420 38108 21476
rect 38164 21420 38892 21476
rect 38948 21420 38958 21476
rect 6850 21308 6860 21364
rect 6916 21308 9548 21364
rect 9604 21308 9614 21364
rect 28690 21308 28700 21364
rect 28756 21308 30492 21364
rect 30548 21308 30558 21364
rect 23986 21196 23996 21252
rect 24052 21196 30380 21252
rect 30436 21196 30446 21252
rect 48402 21196 48412 21252
rect 48468 21196 49644 21252
rect 49700 21196 49710 21252
rect 4466 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4750 21196
rect 35186 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35470 21196
rect 6738 20972 6748 21028
rect 6804 20972 10108 21028
rect 10164 20972 10174 21028
rect 45938 20972 45948 21028
rect 46004 20972 46284 21028
rect 46340 20972 46350 21028
rect 0 20916 800 20944
rect 0 20860 1708 20916
rect 1764 20860 1774 20916
rect 8978 20860 8988 20916
rect 9044 20860 10332 20916
rect 10388 20860 10398 20916
rect 16818 20860 16828 20916
rect 16884 20860 17724 20916
rect 17780 20860 17790 20916
rect 22530 20860 22540 20916
rect 22596 20860 23324 20916
rect 23380 20860 23390 20916
rect 41346 20860 41356 20916
rect 41412 20860 44044 20916
rect 44100 20860 44110 20916
rect 0 20832 800 20860
rect 9202 20748 9212 20804
rect 9268 20748 10556 20804
rect 10612 20748 10622 20804
rect 14802 20748 14812 20804
rect 14868 20748 16156 20804
rect 16212 20748 16222 20804
rect 28242 20748 28252 20804
rect 28308 20748 28588 20804
rect 28644 20748 28654 20804
rect 40338 20748 40348 20804
rect 40404 20748 41580 20804
rect 41636 20748 42924 20804
rect 42980 20748 42990 20804
rect 47842 20748 47852 20804
rect 47908 20748 50092 20804
rect 50148 20748 50158 20804
rect 6290 20636 6300 20692
rect 6356 20636 9324 20692
rect 9380 20636 9390 20692
rect 16034 20636 16044 20692
rect 16100 20636 17612 20692
rect 17668 20636 17678 20692
rect 28914 20636 28924 20692
rect 28980 20636 34300 20692
rect 34356 20636 34972 20692
rect 35028 20636 35038 20692
rect 41234 20636 41244 20692
rect 41300 20636 41468 20692
rect 41524 20636 42364 20692
rect 42420 20636 42430 20692
rect 27766 20524 27804 20580
rect 27860 20524 31500 20580
rect 31556 20524 31566 20580
rect 33506 20524 33516 20580
rect 33572 20524 35756 20580
rect 35812 20524 37100 20580
rect 37156 20524 37166 20580
rect 37650 20524 37660 20580
rect 37716 20524 40684 20580
rect 40740 20524 40750 20580
rect 41122 20524 41132 20580
rect 41188 20524 45388 20580
rect 45444 20524 46844 20580
rect 46900 20524 47180 20580
rect 47236 20524 47246 20580
rect 26786 20412 26796 20468
rect 26852 20412 28252 20468
rect 28308 20412 28318 20468
rect 19826 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20110 20412
rect 50546 20356 50556 20412
rect 50612 20356 50660 20412
rect 50716 20356 50764 20412
rect 50820 20356 50830 20412
rect 33590 20300 33628 20356
rect 33684 20300 33694 20356
rect 35634 20300 35644 20356
rect 35700 20300 36092 20356
rect 36148 20300 36158 20356
rect 43586 20300 43596 20356
rect 43652 20300 45500 20356
rect 45556 20300 45566 20356
rect 0 20244 800 20272
rect 0 20188 1708 20244
rect 1764 20188 2492 20244
rect 2548 20188 2558 20244
rect 16706 20188 16716 20244
rect 16772 20188 19292 20244
rect 19348 20188 19358 20244
rect 24546 20188 24556 20244
rect 24612 20188 25340 20244
rect 25396 20188 26908 20244
rect 29698 20188 29708 20244
rect 29764 20188 31276 20244
rect 31332 20188 31342 20244
rect 34290 20188 34300 20244
rect 34356 20188 34860 20244
rect 34916 20188 35084 20244
rect 35140 20188 35150 20244
rect 38098 20188 38108 20244
rect 38164 20188 42476 20244
rect 42532 20188 46508 20244
rect 46564 20188 46574 20244
rect 0 20160 800 20188
rect 26852 20132 26908 20188
rect 2034 20076 2044 20132
rect 2100 20076 9548 20132
rect 9604 20076 9614 20132
rect 12226 20076 12236 20132
rect 12292 20076 13468 20132
rect 13524 20076 13534 20132
rect 13682 20076 13692 20132
rect 13748 20076 15036 20132
rect 15092 20076 16044 20132
rect 16100 20076 17612 20132
rect 17668 20076 17678 20132
rect 19618 20076 19628 20132
rect 19684 20076 20860 20132
rect 20916 20076 20926 20132
rect 26852 20076 31724 20132
rect 31780 20076 31790 20132
rect 34066 20076 34076 20132
rect 34132 20076 39452 20132
rect 39508 20076 39518 20132
rect 41692 20020 41748 20188
rect 43362 20076 43372 20132
rect 43428 20076 53788 20132
rect 53844 20076 53854 20132
rect 15362 19964 15372 20020
rect 15428 19964 16604 20020
rect 16660 19964 16670 20020
rect 19506 19964 19516 20020
rect 19572 19964 19964 20020
rect 20020 19964 20412 20020
rect 20468 19964 20478 20020
rect 21410 19964 21420 20020
rect 21476 19964 21868 20020
rect 21924 19964 21934 20020
rect 24770 19964 24780 20020
rect 24836 19964 25676 20020
rect 25732 19964 25742 20020
rect 30370 19964 30380 20020
rect 30436 19964 31164 20020
rect 31220 19964 31230 20020
rect 34850 19964 34860 20020
rect 34916 19964 38668 20020
rect 41682 19964 41692 20020
rect 41748 19964 41758 20020
rect 44482 19964 44492 20020
rect 44548 19964 46284 20020
rect 46340 19964 46350 20020
rect 7970 19852 7980 19908
rect 8036 19852 8988 19908
rect 9044 19852 11452 19908
rect 11508 19852 11518 19908
rect 15698 19852 15708 19908
rect 15764 19852 18620 19908
rect 18676 19852 18686 19908
rect 27234 19852 27244 19908
rect 27300 19852 27692 19908
rect 27748 19852 27758 19908
rect 31378 19852 31388 19908
rect 31444 19852 31948 19908
rect 32004 19852 33516 19908
rect 33572 19852 33582 19908
rect 38612 19796 38668 19964
rect 44370 19852 44380 19908
rect 44436 19852 46060 19908
rect 46116 19852 47292 19908
rect 47348 19852 47358 19908
rect 2706 19740 2716 19796
rect 2772 19740 13916 19796
rect 13972 19740 13982 19796
rect 14578 19740 14588 19796
rect 14644 19740 17388 19796
rect 17444 19740 17454 19796
rect 34738 19740 34748 19796
rect 34804 19740 34814 19796
rect 38612 19740 39900 19796
rect 39956 19740 39966 19796
rect 40226 19740 40236 19796
rect 40292 19740 42588 19796
rect 42644 19740 42654 19796
rect 7186 19628 7196 19684
rect 7252 19628 11004 19684
rect 11060 19628 14252 19684
rect 14308 19628 15708 19684
rect 15764 19628 15774 19684
rect 16594 19628 16604 19684
rect 16660 19628 17836 19684
rect 17892 19628 17902 19684
rect 0 19572 800 19600
rect 4466 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4750 19628
rect 0 19516 1708 19572
rect 1764 19516 2492 19572
rect 2548 19516 2558 19572
rect 12338 19516 12348 19572
rect 12404 19516 17724 19572
rect 17780 19516 17790 19572
rect 0 19488 800 19516
rect 34748 19460 34804 19740
rect 37202 19628 37212 19684
rect 37268 19628 43708 19684
rect 43764 19628 47628 19684
rect 47684 19628 48860 19684
rect 48916 19628 48926 19684
rect 35186 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35470 19628
rect 13570 19404 13580 19460
rect 13636 19404 16828 19460
rect 16884 19404 16894 19460
rect 26002 19404 26012 19460
rect 26068 19404 27244 19460
rect 27300 19404 27692 19460
rect 27748 19404 27758 19460
rect 34748 19404 35308 19460
rect 35364 19404 35644 19460
rect 35700 19404 35710 19460
rect 36194 19404 36204 19460
rect 36260 19404 37100 19460
rect 37156 19404 37166 19460
rect 13122 19292 13132 19348
rect 13188 19292 14588 19348
rect 14644 19292 15484 19348
rect 15540 19292 15550 19348
rect 17938 19292 17948 19348
rect 18004 19292 19852 19348
rect 19908 19292 21756 19348
rect 21812 19292 21822 19348
rect 25666 19292 25676 19348
rect 25732 19292 26460 19348
rect 26516 19292 26526 19348
rect 34962 19292 34972 19348
rect 35028 19292 35420 19348
rect 35476 19292 36092 19348
rect 36148 19292 36652 19348
rect 36708 19292 37660 19348
rect 37716 19292 37726 19348
rect 41570 19292 41580 19348
rect 41636 19292 42700 19348
rect 42756 19292 42766 19348
rect 47730 19292 47740 19348
rect 47796 19292 48076 19348
rect 48132 19292 48142 19348
rect 9650 19180 9660 19236
rect 9716 19180 11900 19236
rect 11956 19180 12684 19236
rect 12740 19180 12750 19236
rect 15026 19180 15036 19236
rect 15092 19180 16940 19236
rect 16996 19180 17006 19236
rect 21858 19180 21868 19236
rect 21924 19180 24780 19236
rect 24836 19180 24846 19236
rect 27458 19180 27468 19236
rect 27524 19180 28140 19236
rect 28196 19180 28206 19236
rect 35746 19180 35756 19236
rect 35812 19180 38108 19236
rect 38164 19180 38174 19236
rect 40786 19180 40796 19236
rect 40852 19180 42588 19236
rect 42644 19180 45500 19236
rect 45556 19180 45566 19236
rect 7858 19068 7868 19124
rect 7924 19068 8764 19124
rect 8820 19068 11452 19124
rect 11508 19068 11518 19124
rect 12898 19068 12908 19124
rect 12964 19068 16156 19124
rect 16212 19068 16222 19124
rect 20738 19068 20748 19124
rect 20804 19068 21868 19124
rect 21924 19068 22204 19124
rect 22260 19068 22270 19124
rect 22418 19068 22428 19124
rect 22484 19068 23548 19124
rect 23604 19068 23614 19124
rect 25442 19068 25452 19124
rect 25508 19068 26908 19124
rect 26964 19068 26974 19124
rect 31826 19068 31836 19124
rect 31892 19068 37100 19124
rect 37156 19068 38556 19124
rect 38612 19068 38622 19124
rect 41794 19068 41804 19124
rect 41860 19068 42924 19124
rect 42980 19068 42990 19124
rect 44034 19068 44044 19124
rect 44100 19068 44940 19124
rect 44996 19068 45006 19124
rect 16818 18956 16828 19012
rect 16884 18956 17500 19012
rect 17556 18956 17566 19012
rect 22082 18956 22092 19012
rect 22148 18956 22876 19012
rect 22932 18956 22942 19012
rect 25666 18956 25676 19012
rect 25732 18956 26124 19012
rect 26180 18956 26190 19012
rect 26450 18956 26460 19012
rect 26516 18956 27804 19012
rect 27860 18956 27870 19012
rect 29586 18956 29596 19012
rect 29652 18956 30492 19012
rect 30548 18956 30558 19012
rect 36502 18956 36540 19012
rect 36596 18956 36606 19012
rect 42242 18956 42252 19012
rect 42308 18956 43148 19012
rect 43204 18956 43214 19012
rect 43922 18956 43932 19012
rect 43988 18956 44716 19012
rect 44772 18956 44782 19012
rect 46358 18956 46396 19012
rect 46452 18956 46462 19012
rect 34402 18844 34412 18900
rect 34468 18844 35084 18900
rect 35140 18844 35150 18900
rect 42802 18844 42812 18900
rect 42868 18844 43372 18900
rect 43428 18844 43438 18900
rect 19826 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20110 18844
rect 50546 18788 50556 18844
rect 50612 18788 50660 18844
rect 50716 18788 50764 18844
rect 50820 18788 50830 18844
rect 23650 18732 23660 18788
rect 23716 18732 24668 18788
rect 24724 18732 28812 18788
rect 28868 18732 28878 18788
rect 34486 18732 34524 18788
rect 34580 18732 34590 18788
rect 35644 18732 36316 18788
rect 36372 18732 36382 18788
rect 40226 18732 40236 18788
rect 40292 18732 40684 18788
rect 40740 18732 40750 18788
rect 35644 18676 35700 18732
rect 8866 18620 8876 18676
rect 8932 18620 9884 18676
rect 9940 18620 10276 18676
rect 24546 18620 24556 18676
rect 24612 18620 25228 18676
rect 25284 18620 25294 18676
rect 25890 18620 25900 18676
rect 25956 18620 27356 18676
rect 27412 18620 27422 18676
rect 27794 18620 27804 18676
rect 27860 18620 33068 18676
rect 33124 18620 33134 18676
rect 35634 18620 35644 18676
rect 35700 18620 35710 18676
rect 40338 18620 40348 18676
rect 40404 18620 40796 18676
rect 40852 18620 40862 18676
rect 42578 18620 42588 18676
rect 42644 18620 43820 18676
rect 43876 18620 43886 18676
rect 47058 18620 47068 18676
rect 47124 18620 48076 18676
rect 48132 18620 48142 18676
rect 10220 18452 10276 18620
rect 28140 18564 28196 18620
rect 11554 18508 11564 18564
rect 11620 18508 12348 18564
rect 12404 18508 12414 18564
rect 22530 18508 22540 18564
rect 22596 18508 23100 18564
rect 23156 18508 23772 18564
rect 23828 18508 23838 18564
rect 26226 18508 26236 18564
rect 26292 18508 26908 18564
rect 26964 18508 27468 18564
rect 27524 18508 27534 18564
rect 28130 18508 28140 18564
rect 28196 18508 28206 18564
rect 29698 18508 29708 18564
rect 29764 18508 30380 18564
rect 30436 18508 30446 18564
rect 33964 18508 35420 18564
rect 35476 18508 35486 18564
rect 36082 18508 36092 18564
rect 36148 18508 37324 18564
rect 37380 18508 37390 18564
rect 40226 18508 40236 18564
rect 40292 18508 40908 18564
rect 40964 18508 40974 18564
rect 42914 18508 42924 18564
rect 42980 18508 43596 18564
rect 43652 18508 43662 18564
rect 45490 18508 45500 18564
rect 45556 18508 46844 18564
rect 46900 18508 46910 18564
rect 33964 18452 34020 18508
rect 6066 18396 6076 18452
rect 6132 18396 7084 18452
rect 7140 18396 8316 18452
rect 8372 18396 9884 18452
rect 9940 18396 9950 18452
rect 10220 18396 11340 18452
rect 11396 18396 11676 18452
rect 11732 18396 11742 18452
rect 16482 18396 16492 18452
rect 16548 18396 17388 18452
rect 17444 18396 17454 18452
rect 19730 18396 19740 18452
rect 19796 18396 20748 18452
rect 20804 18396 21084 18452
rect 21140 18396 21150 18452
rect 23314 18396 23324 18452
rect 23380 18396 24332 18452
rect 24388 18396 24398 18452
rect 30258 18396 30268 18452
rect 30324 18396 31500 18452
rect 31556 18396 32284 18452
rect 32340 18396 32350 18452
rect 32834 18396 32844 18452
rect 32900 18396 33740 18452
rect 33796 18396 33806 18452
rect 33954 18396 33964 18452
rect 34020 18396 34030 18452
rect 36642 18396 36652 18452
rect 36708 18396 39116 18452
rect 39172 18396 39182 18452
rect 39330 18396 39340 18452
rect 39396 18396 42140 18452
rect 42196 18396 42206 18452
rect 43362 18396 43372 18452
rect 43428 18396 45276 18452
rect 45332 18396 45342 18452
rect 2034 18284 2044 18340
rect 2100 18284 6524 18340
rect 6580 18284 6590 18340
rect 8194 18284 8204 18340
rect 8260 18284 10556 18340
rect 10612 18284 10622 18340
rect 16258 18284 16268 18340
rect 16324 18284 18060 18340
rect 18116 18284 18126 18340
rect 18274 18284 18284 18340
rect 18340 18284 19292 18340
rect 19348 18284 19358 18340
rect 22754 18284 22764 18340
rect 22820 18284 24108 18340
rect 24164 18284 24174 18340
rect 33618 18284 33628 18340
rect 33684 18284 34188 18340
rect 34244 18284 34254 18340
rect 35074 18284 35084 18340
rect 35140 18284 35756 18340
rect 35812 18284 35822 18340
rect 37202 18284 37212 18340
rect 37268 18284 37660 18340
rect 37716 18284 37726 18340
rect 0 18228 800 18256
rect 39116 18228 39172 18396
rect 40002 18284 40012 18340
rect 40068 18284 41020 18340
rect 41076 18284 41086 18340
rect 46274 18284 46284 18340
rect 46340 18284 47516 18340
rect 47572 18284 48300 18340
rect 48356 18284 48748 18340
rect 48804 18284 49756 18340
rect 49812 18284 49822 18340
rect 0 18172 1708 18228
rect 1764 18172 2492 18228
rect 2548 18172 2558 18228
rect 7858 18172 7868 18228
rect 7924 18172 10444 18228
rect 10500 18172 10510 18228
rect 14354 18172 14364 18228
rect 14420 18172 15596 18228
rect 15652 18172 16492 18228
rect 16548 18172 16558 18228
rect 24210 18172 24220 18228
rect 24276 18172 25004 18228
rect 25060 18172 25340 18228
rect 25396 18172 25406 18228
rect 25778 18172 25788 18228
rect 25844 18172 28588 18228
rect 28644 18172 29260 18228
rect 29316 18172 29326 18228
rect 33394 18172 33404 18228
rect 33460 18172 34524 18228
rect 34580 18172 34590 18228
rect 34962 18172 34972 18228
rect 35028 18172 35644 18228
rect 35700 18172 35980 18228
rect 36036 18172 36046 18228
rect 39116 18172 45724 18228
rect 45780 18172 45790 18228
rect 0 18144 800 18172
rect 25788 18116 25844 18172
rect 6962 18060 6972 18116
rect 7028 18060 9548 18116
rect 9604 18060 9614 18116
rect 12114 18060 12124 18116
rect 12180 18060 12908 18116
rect 12964 18060 13692 18116
rect 13748 18060 13758 18116
rect 15922 18060 15932 18116
rect 15988 18060 16380 18116
rect 16436 18060 16446 18116
rect 21522 18060 21532 18116
rect 21588 18060 22204 18116
rect 22260 18060 25844 18116
rect 33842 18060 33852 18116
rect 33908 18060 34412 18116
rect 34468 18060 34478 18116
rect 35858 18060 35868 18116
rect 35924 18060 36988 18116
rect 37044 18060 37054 18116
rect 38322 18060 38332 18116
rect 38388 18060 39228 18116
rect 39284 18060 39294 18116
rect 4466 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4750 18060
rect 23212 18004 23268 18060
rect 35186 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35470 18060
rect 23202 17948 23212 18004
rect 23268 17948 23278 18004
rect 37874 17948 37884 18004
rect 37940 17948 38892 18004
rect 38948 17948 38958 18004
rect 41570 17948 41580 18004
rect 41636 17948 43036 18004
rect 43092 17948 44604 18004
rect 44660 17948 46956 18004
rect 47012 17948 47022 18004
rect 17938 17836 17948 17892
rect 18004 17836 18956 17892
rect 19012 17836 19022 17892
rect 46610 17836 46620 17892
rect 46676 17836 47628 17892
rect 47684 17836 47694 17892
rect 48402 17836 48412 17892
rect 48468 17836 48972 17892
rect 49028 17836 49038 17892
rect 9762 17724 9772 17780
rect 9828 17724 11116 17780
rect 11172 17724 11182 17780
rect 17714 17724 17724 17780
rect 17780 17724 20076 17780
rect 20132 17724 20142 17780
rect 23874 17724 23884 17780
rect 23940 17724 25340 17780
rect 25396 17724 28364 17780
rect 28420 17724 28430 17780
rect 29922 17724 29932 17780
rect 29988 17724 30828 17780
rect 30884 17724 30894 17780
rect 33170 17724 33180 17780
rect 33236 17724 33628 17780
rect 33684 17724 36652 17780
rect 36708 17724 36718 17780
rect 38658 17724 38668 17780
rect 38724 17724 39564 17780
rect 39620 17724 39630 17780
rect 41794 17724 41804 17780
rect 41860 17724 43036 17780
rect 43092 17724 43932 17780
rect 43988 17724 43998 17780
rect 46358 17724 46396 17780
rect 46452 17724 46462 17780
rect 18050 17612 18060 17668
rect 18116 17612 19292 17668
rect 19348 17612 20188 17668
rect 20244 17612 20254 17668
rect 0 17556 800 17584
rect 0 17500 1708 17556
rect 1764 17500 2492 17556
rect 2548 17500 2558 17556
rect 2706 17500 2716 17556
rect 2772 17500 7420 17556
rect 7476 17500 7486 17556
rect 11106 17500 11116 17556
rect 11172 17500 11452 17556
rect 11508 17500 12348 17556
rect 12404 17500 12414 17556
rect 0 17472 800 17500
rect 2034 17388 2044 17444
rect 2100 17388 5180 17444
rect 5236 17388 5246 17444
rect 16482 17388 16492 17444
rect 16548 17388 18620 17444
rect 18676 17388 20188 17444
rect 20244 17388 20254 17444
rect 2146 17276 2156 17332
rect 2212 17276 13692 17332
rect 13748 17276 13758 17332
rect 19826 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20110 17276
rect 28364 17220 28420 17724
rect 31378 17612 31388 17668
rect 31444 17612 32284 17668
rect 32340 17612 32844 17668
rect 32900 17612 34076 17668
rect 34132 17612 35196 17668
rect 35252 17612 35262 17668
rect 35420 17612 36092 17668
rect 36148 17612 36540 17668
rect 36596 17612 36606 17668
rect 47730 17612 47740 17668
rect 47796 17612 48188 17668
rect 48244 17612 48748 17668
rect 48804 17612 48814 17668
rect 29810 17500 29820 17556
rect 29876 17500 31612 17556
rect 31668 17500 31678 17556
rect 34514 17500 34524 17556
rect 34580 17500 34748 17556
rect 34804 17500 34814 17556
rect 35420 17444 35476 17612
rect 36978 17500 36988 17556
rect 37044 17500 37324 17556
rect 37380 17500 43372 17556
rect 43428 17500 43438 17556
rect 45714 17500 45724 17556
rect 45780 17500 47404 17556
rect 47460 17500 48076 17556
rect 48132 17500 48142 17556
rect 31378 17388 31388 17444
rect 31444 17388 35476 17444
rect 36166 17388 36204 17444
rect 36260 17388 36270 17444
rect 40786 17388 40796 17444
rect 40852 17388 42812 17444
rect 42868 17388 42878 17444
rect 45378 17388 45388 17444
rect 45444 17388 46284 17444
rect 46340 17388 46350 17444
rect 47618 17388 47628 17444
rect 47684 17388 48860 17444
rect 48916 17388 48926 17444
rect 35634 17276 35644 17332
rect 35700 17276 45052 17332
rect 45108 17276 46732 17332
rect 46788 17276 46798 17332
rect 50546 17220 50556 17276
rect 50612 17220 50660 17276
rect 50716 17220 50764 17276
rect 50820 17220 50830 17276
rect 11330 17164 11340 17220
rect 11396 17164 12124 17220
rect 12180 17164 12190 17220
rect 23538 17164 23548 17220
rect 23604 17164 24108 17220
rect 24164 17164 24444 17220
rect 24500 17164 24510 17220
rect 28364 17164 30268 17220
rect 30324 17164 31388 17220
rect 31444 17164 31454 17220
rect 32050 17164 32060 17220
rect 32116 17164 33180 17220
rect 33236 17164 33246 17220
rect 33506 17164 33516 17220
rect 33572 17164 36540 17220
rect 36596 17164 39676 17220
rect 39732 17164 46396 17220
rect 46452 17164 46462 17220
rect 30818 17052 30828 17108
rect 30884 17052 31948 17108
rect 32004 17052 32014 17108
rect 34178 17052 34188 17108
rect 34244 17052 35756 17108
rect 35812 17052 36204 17108
rect 36260 17052 36270 17108
rect 36642 17052 36652 17108
rect 36708 17052 36988 17108
rect 37044 17052 37054 17108
rect 37650 17052 37660 17108
rect 37716 17052 39228 17108
rect 39284 17052 40124 17108
rect 40180 17052 40190 17108
rect 41346 17052 41356 17108
rect 41412 17052 41580 17108
rect 41636 17052 41646 17108
rect 44930 17052 44940 17108
rect 44996 17052 46060 17108
rect 46116 17052 46126 17108
rect 48290 17052 48300 17108
rect 48356 17052 49308 17108
rect 49364 17052 49374 17108
rect 36540 16940 37212 16996
rect 37268 16940 37278 16996
rect 39106 16940 39116 16996
rect 39172 16940 39452 16996
rect 39508 16940 41692 16996
rect 41748 16940 41758 16996
rect 43698 16940 43708 16996
rect 43764 16940 45276 16996
rect 45332 16940 45342 16996
rect 49186 16940 49196 16996
rect 49252 16940 50876 16996
rect 50932 16940 50942 16996
rect 0 16884 800 16912
rect 36540 16884 36596 16940
rect 0 16828 2380 16884
rect 2436 16828 3164 16884
rect 3220 16828 3230 16884
rect 8978 16828 8988 16884
rect 9044 16828 11228 16884
rect 11284 16828 11294 16884
rect 17490 16828 17500 16884
rect 17556 16828 18284 16884
rect 18340 16828 18350 16884
rect 30594 16828 30604 16884
rect 30660 16828 31948 16884
rect 32004 16828 32014 16884
rect 34738 16828 34748 16884
rect 34804 16828 35644 16884
rect 35700 16828 35710 16884
rect 36530 16828 36540 16884
rect 36596 16828 36606 16884
rect 37090 16828 37100 16884
rect 37156 16828 38556 16884
rect 38612 16828 39340 16884
rect 39396 16828 39406 16884
rect 40338 16828 40348 16884
rect 40404 16828 42028 16884
rect 42084 16828 42094 16884
rect 44818 16828 44828 16884
rect 44884 16828 46620 16884
rect 46676 16828 46686 16884
rect 0 16800 800 16828
rect 2034 16716 2044 16772
rect 2100 16716 6916 16772
rect 8866 16716 8876 16772
rect 8932 16716 10108 16772
rect 10164 16716 10174 16772
rect 22194 16716 22204 16772
rect 22260 16716 23660 16772
rect 23716 16716 23726 16772
rect 26450 16716 26460 16772
rect 26516 16716 27020 16772
rect 27076 16716 27916 16772
rect 27972 16716 27982 16772
rect 28690 16716 28700 16772
rect 28756 16716 34188 16772
rect 34244 16716 34254 16772
rect 45154 16716 45164 16772
rect 45220 16716 45612 16772
rect 45668 16716 45678 16772
rect 6860 16548 6916 16716
rect 8754 16604 8764 16660
rect 8820 16604 10220 16660
rect 10276 16604 10286 16660
rect 24770 16604 24780 16660
rect 24836 16604 25340 16660
rect 25396 16604 25406 16660
rect 26226 16604 26236 16660
rect 26292 16604 26796 16660
rect 26852 16604 27692 16660
rect 27748 16604 27758 16660
rect 30034 16604 30044 16660
rect 30100 16604 31724 16660
rect 31780 16604 31790 16660
rect 35410 16604 35420 16660
rect 35476 16604 36540 16660
rect 36596 16604 36606 16660
rect 40898 16604 40908 16660
rect 40964 16604 42028 16660
rect 42084 16604 42094 16660
rect 42802 16604 42812 16660
rect 42868 16604 48412 16660
rect 48468 16604 48478 16660
rect 6860 16492 10332 16548
rect 10388 16492 10398 16548
rect 4466 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4750 16492
rect 35186 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35470 16492
rect 17266 16268 17276 16324
rect 17332 16268 18956 16324
rect 19012 16268 19022 16324
rect 0 16212 800 16240
rect 0 16156 1820 16212
rect 1876 16156 1886 16212
rect 18610 16156 18620 16212
rect 18676 16156 19516 16212
rect 19572 16156 19582 16212
rect 21858 16156 21868 16212
rect 21924 16156 22652 16212
rect 22708 16156 22718 16212
rect 29026 16156 29036 16212
rect 29092 16156 30604 16212
rect 30660 16156 32620 16212
rect 32676 16156 32686 16212
rect 46722 16156 46732 16212
rect 46788 16156 47292 16212
rect 47348 16156 47740 16212
rect 47796 16156 49980 16212
rect 50036 16156 50046 16212
rect 0 16128 800 16156
rect 28914 16044 28924 16100
rect 28980 16044 29260 16100
rect 29316 16044 29326 16100
rect 34738 16044 34748 16100
rect 34804 16044 35644 16100
rect 35700 16044 35710 16100
rect 40226 16044 40236 16100
rect 40292 16044 41804 16100
rect 41860 16044 41870 16100
rect 43474 16044 43484 16100
rect 43540 16044 45052 16100
rect 45108 16044 45118 16100
rect 45602 16044 45612 16100
rect 45668 16044 46620 16100
rect 46676 16044 46686 16100
rect 48402 16044 48412 16100
rect 48468 16044 49756 16100
rect 49812 16044 49822 16100
rect 15138 15932 15148 15988
rect 15204 15932 16604 15988
rect 16660 15932 16670 15988
rect 25442 15932 25452 15988
rect 25508 15932 26236 15988
rect 26292 15932 26302 15988
rect 26562 15932 26572 15988
rect 26628 15932 27804 15988
rect 27860 15932 27870 15988
rect 31714 15932 31724 15988
rect 31780 15932 36372 15988
rect 38546 15932 38556 15988
rect 38612 15932 39228 15988
rect 39284 15932 39294 15988
rect 40898 15932 40908 15988
rect 40964 15932 41916 15988
rect 41972 15932 41982 15988
rect 48066 15932 48076 15988
rect 48132 15932 49420 15988
rect 49476 15932 49486 15988
rect 36316 15876 36372 15932
rect 50372 15876 50428 16100
rect 50484 16044 50494 16100
rect 12786 15820 12796 15876
rect 12852 15820 13692 15876
rect 13748 15820 13758 15876
rect 27682 15820 27692 15876
rect 27748 15820 29036 15876
rect 29092 15820 29102 15876
rect 31938 15820 31948 15876
rect 32004 15820 33068 15876
rect 33124 15820 33134 15876
rect 35970 15820 35980 15876
rect 36036 15820 36092 15876
rect 36148 15820 36158 15876
rect 36306 15820 36316 15876
rect 36372 15820 36382 15876
rect 37314 15820 37324 15876
rect 37380 15820 38444 15876
rect 38500 15820 38510 15876
rect 40674 15820 40684 15876
rect 40740 15820 41020 15876
rect 41076 15820 41086 15876
rect 46050 15820 46060 15876
rect 46116 15820 48748 15876
rect 48804 15820 48814 15876
rect 48962 15820 48972 15876
rect 49028 15820 49532 15876
rect 49588 15820 50428 15876
rect 29586 15708 29596 15764
rect 29652 15708 32172 15764
rect 32228 15708 32844 15764
rect 32900 15708 32910 15764
rect 47618 15708 47628 15764
rect 47684 15708 47694 15764
rect 19826 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20110 15708
rect 47628 15652 47684 15708
rect 50546 15652 50556 15708
rect 50612 15652 50660 15708
rect 50716 15652 50764 15708
rect 50820 15652 50830 15708
rect 18946 15596 18956 15652
rect 19012 15596 19628 15652
rect 19684 15596 19694 15652
rect 22642 15596 22652 15652
rect 22708 15596 30044 15652
rect 30100 15596 30110 15652
rect 32050 15596 32060 15652
rect 32116 15596 33404 15652
rect 33460 15596 35196 15652
rect 35252 15596 35980 15652
rect 36036 15596 36046 15652
rect 47628 15596 49028 15652
rect 16370 15484 16380 15540
rect 16436 15484 19068 15540
rect 19124 15484 19134 15540
rect 22978 15484 22988 15540
rect 23044 15484 23660 15540
rect 23716 15484 23726 15540
rect 23874 15484 23884 15540
rect 23940 15484 24668 15540
rect 24724 15484 29148 15540
rect 29204 15484 29214 15540
rect 29362 15484 29372 15540
rect 29428 15484 33292 15540
rect 33348 15484 33358 15540
rect 47842 15484 47852 15540
rect 47908 15484 48748 15540
rect 48804 15484 48814 15540
rect 30818 15372 30828 15428
rect 30884 15372 33068 15428
rect 33124 15372 33134 15428
rect 39778 15372 39788 15428
rect 39844 15372 41580 15428
rect 41636 15372 41646 15428
rect 43922 15372 43932 15428
rect 43988 15372 44940 15428
rect 44996 15372 45006 15428
rect 47394 15372 47404 15428
rect 47460 15372 48076 15428
rect 48132 15372 48142 15428
rect 14466 15260 14476 15316
rect 14532 15260 17836 15316
rect 17892 15260 18508 15316
rect 18564 15260 18574 15316
rect 23314 15260 23324 15316
rect 23380 15260 25228 15316
rect 25284 15260 27244 15316
rect 27300 15260 27310 15316
rect 28354 15260 28364 15316
rect 28420 15260 29260 15316
rect 29316 15260 29326 15316
rect 32498 15260 32508 15316
rect 32564 15260 33516 15316
rect 33572 15260 33582 15316
rect 33954 15260 33964 15316
rect 34020 15260 35308 15316
rect 35364 15260 35374 15316
rect 36306 15260 36316 15316
rect 36372 15260 37884 15316
rect 37940 15260 37950 15316
rect 40002 15260 40012 15316
rect 40068 15260 40460 15316
rect 40516 15260 41916 15316
rect 41972 15260 41982 15316
rect 28364 15204 28420 15260
rect 48972 15204 49028 15596
rect 25676 15148 28420 15204
rect 31490 15148 31500 15204
rect 31556 15148 33180 15204
rect 33236 15148 33246 15204
rect 35634 15148 35644 15204
rect 35700 15148 42700 15204
rect 42756 15148 42766 15204
rect 45154 15148 45164 15204
rect 45220 15148 46508 15204
rect 46564 15148 46574 15204
rect 48962 15148 48972 15204
rect 49028 15148 49038 15204
rect 25676 15092 25732 15148
rect 23202 15036 23212 15092
rect 23268 15036 24332 15092
rect 24388 15036 24398 15092
rect 25666 15036 25676 15092
rect 25732 15036 25742 15092
rect 28130 15036 28140 15092
rect 28196 15036 28588 15092
rect 28644 15036 28654 15092
rect 33628 15036 35420 15092
rect 35476 15036 35980 15092
rect 36036 15036 36046 15092
rect 41682 15036 41692 15092
rect 41748 15036 42364 15092
rect 42420 15036 42430 15092
rect 47954 15036 47964 15092
rect 48020 15036 49420 15092
rect 49476 15036 51660 15092
rect 51716 15036 52780 15092
rect 52836 15036 52846 15092
rect 33628 14980 33684 15036
rect 23762 14924 23772 14980
rect 23828 14924 24444 14980
rect 24500 14924 24510 14980
rect 33618 14924 33628 14980
rect 33684 14924 33694 14980
rect 37874 14924 37884 14980
rect 37940 14924 39564 14980
rect 39620 14924 39900 14980
rect 39956 14924 39966 14980
rect 4466 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4750 14924
rect 35186 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35470 14924
rect 30258 14812 30268 14868
rect 30324 14812 31948 14868
rect 32004 14812 34748 14868
rect 34804 14812 34814 14868
rect 40226 14812 40236 14868
rect 40292 14812 41580 14868
rect 41636 14812 43036 14868
rect 43092 14812 43102 14868
rect 23538 14700 23548 14756
rect 23604 14700 24108 14756
rect 24164 14700 25228 14756
rect 25284 14700 25294 14756
rect 35074 14700 35084 14756
rect 35140 14700 35308 14756
rect 28130 14588 28140 14644
rect 28196 14588 28700 14644
rect 28756 14588 28766 14644
rect 35252 14532 35308 14700
rect 42998 14588 43036 14644
rect 43092 14588 43102 14644
rect 44818 14588 44828 14644
rect 44884 14588 45500 14644
rect 45556 14588 45566 14644
rect 5170 14476 5180 14532
rect 5236 14476 9772 14532
rect 9828 14476 9838 14532
rect 11218 14476 11228 14532
rect 11284 14476 11900 14532
rect 11956 14476 11966 14532
rect 29922 14476 29932 14532
rect 29988 14476 30604 14532
rect 30660 14476 31276 14532
rect 31332 14476 31342 14532
rect 35252 14476 35756 14532
rect 35812 14476 37044 14532
rect 38322 14476 38332 14532
rect 38388 14476 38668 14532
rect 38724 14476 38734 14532
rect 47058 14476 47068 14532
rect 47124 14476 49868 14532
rect 49924 14476 49934 14532
rect 36988 14420 37044 14476
rect 24434 14364 24444 14420
rect 24500 14364 25116 14420
rect 25172 14364 25182 14420
rect 25778 14364 25788 14420
rect 25844 14364 26572 14420
rect 26628 14364 26638 14420
rect 29698 14364 29708 14420
rect 29764 14364 30828 14420
rect 30884 14364 31164 14420
rect 31220 14364 31230 14420
rect 35522 14364 35532 14420
rect 35588 14364 35644 14420
rect 35700 14364 35710 14420
rect 36978 14364 36988 14420
rect 37044 14364 37324 14420
rect 37380 14364 37390 14420
rect 37986 14364 37996 14420
rect 38052 14364 38780 14420
rect 38836 14364 38846 14420
rect 19282 14252 19292 14308
rect 19348 14252 21308 14308
rect 21364 14252 21374 14308
rect 22530 14252 22540 14308
rect 22596 14252 24220 14308
rect 24276 14252 24286 14308
rect 35074 14252 35084 14308
rect 35140 14252 37212 14308
rect 37268 14252 37278 14308
rect 38994 14252 39004 14308
rect 39060 14252 39900 14308
rect 39956 14252 43484 14308
rect 43540 14252 43550 14308
rect 19826 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20110 14140
rect 50546 14084 50556 14140
rect 50612 14084 50660 14140
rect 50716 14084 50764 14140
rect 50820 14084 50830 14140
rect 38210 13916 38220 13972
rect 38276 13916 38780 13972
rect 38836 13916 38846 13972
rect 41458 13916 41468 13972
rect 41524 13916 42476 13972
rect 42532 13916 43036 13972
rect 43092 13916 43484 13972
rect 43540 13916 43550 13972
rect 47842 13916 47852 13972
rect 47908 13916 49196 13972
rect 49252 13916 49262 13972
rect 33394 13804 33404 13860
rect 33460 13804 34300 13860
rect 34356 13804 34972 13860
rect 35028 13804 35038 13860
rect 35186 13804 35196 13860
rect 35252 13804 36764 13860
rect 36820 13804 40796 13860
rect 40852 13804 41132 13860
rect 41188 13804 43708 13860
rect 46722 13804 46732 13860
rect 46788 13804 47628 13860
rect 47684 13804 47694 13860
rect 43652 13748 43708 13804
rect 24658 13692 24668 13748
rect 24724 13692 25340 13748
rect 25396 13692 25900 13748
rect 25956 13692 26348 13748
rect 26404 13692 26414 13748
rect 34524 13692 35084 13748
rect 35140 13692 35150 13748
rect 37426 13692 37436 13748
rect 37492 13692 37502 13748
rect 38434 13692 38444 13748
rect 38500 13692 39004 13748
rect 39060 13692 39070 13748
rect 43652 13692 45612 13748
rect 45668 13692 45678 13748
rect 46732 13692 48972 13748
rect 49028 13692 49038 13748
rect 34524 13636 34580 13692
rect 21410 13580 21420 13636
rect 21476 13580 22652 13636
rect 22708 13580 22718 13636
rect 27318 13580 27356 13636
rect 27412 13580 27422 13636
rect 29026 13580 29036 13636
rect 29092 13580 29596 13636
rect 29652 13580 29662 13636
rect 34066 13580 34076 13636
rect 34132 13580 34580 13636
rect 37436 13636 37492 13692
rect 46732 13636 46788 13692
rect 37436 13580 37604 13636
rect 37986 13580 37996 13636
rect 38052 13580 38892 13636
rect 38948 13580 38958 13636
rect 46722 13580 46732 13636
rect 46788 13580 46798 13636
rect 47058 13580 47068 13636
rect 47124 13580 47404 13636
rect 47460 13580 47470 13636
rect 48402 13580 48412 13636
rect 48468 13580 48860 13636
rect 48916 13580 48926 13636
rect 28578 13468 28588 13524
rect 28644 13468 30268 13524
rect 30324 13468 31388 13524
rect 31444 13468 37324 13524
rect 37380 13468 37390 13524
rect 28588 13412 28644 13468
rect 26898 13356 26908 13412
rect 26964 13356 27132 13412
rect 27188 13356 28644 13412
rect 37548 13412 37604 13580
rect 38098 13468 38108 13524
rect 38164 13468 38668 13524
rect 38724 13468 38734 13524
rect 46274 13468 46284 13524
rect 46340 13468 46844 13524
rect 46900 13468 46910 13524
rect 37548 13356 37660 13412
rect 37716 13356 37726 13412
rect 4466 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4750 13356
rect 35186 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35470 13356
rect 26674 13244 26684 13300
rect 26740 13244 28700 13300
rect 28756 13244 28766 13300
rect 48514 13244 48524 13300
rect 48580 13244 48860 13300
rect 48916 13244 49420 13300
rect 49476 13244 49486 13300
rect 21522 13132 21532 13188
rect 21588 13132 22092 13188
rect 22148 13132 22158 13188
rect 20738 13020 20748 13076
rect 20804 13020 22540 13076
rect 22596 13020 22606 13076
rect 28242 13020 28252 13076
rect 28308 13020 29372 13076
rect 29428 13020 29438 13076
rect 35858 13020 35868 13076
rect 35924 13020 36204 13076
rect 36260 13020 36764 13076
rect 36820 13020 36830 13076
rect 44594 13020 44604 13076
rect 44660 13020 45500 13076
rect 45556 13020 45566 13076
rect 21746 12908 21756 12964
rect 21812 12908 22988 12964
rect 23044 12908 23996 12964
rect 24052 12908 25340 12964
rect 25396 12908 25406 12964
rect 31490 12908 31500 12964
rect 31556 12908 32508 12964
rect 32564 12908 32574 12964
rect 22306 12796 22316 12852
rect 22372 12796 23436 12852
rect 23492 12796 33964 12852
rect 34020 12796 34188 12852
rect 34244 12796 36316 12852
rect 36372 12796 36382 12852
rect 37314 12796 37324 12852
rect 37380 12796 37772 12852
rect 37828 12796 43932 12852
rect 43988 12796 43998 12852
rect 47170 12796 47180 12852
rect 47236 12796 47740 12852
rect 47796 12796 47806 12852
rect 19826 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20110 12572
rect 50546 12516 50556 12572
rect 50612 12516 50660 12572
rect 50716 12516 50764 12572
rect 50820 12516 50830 12572
rect 19954 12348 19964 12404
rect 20020 12348 20860 12404
rect 20916 12348 20926 12404
rect 32498 12348 32508 12404
rect 32564 12348 33292 12404
rect 33348 12348 33358 12404
rect 37314 12348 37324 12404
rect 37380 12348 40236 12404
rect 40292 12348 40302 12404
rect 42578 12348 42588 12404
rect 42644 12348 45724 12404
rect 45780 12348 45790 12404
rect 45938 12348 45948 12404
rect 46004 12348 46508 12404
rect 46564 12348 47852 12404
rect 47908 12348 48860 12404
rect 48916 12348 48926 12404
rect 19506 12236 19516 12292
rect 19572 12236 23100 12292
rect 23156 12236 23772 12292
rect 23828 12236 23838 12292
rect 24994 12236 25004 12292
rect 25060 12236 28196 12292
rect 31266 12236 31276 12292
rect 31332 12236 32284 12292
rect 32340 12236 32350 12292
rect 19394 12124 19404 12180
rect 19460 12124 20300 12180
rect 20356 12124 21644 12180
rect 21700 12124 21710 12180
rect 24658 12124 24668 12180
rect 24724 12124 25452 12180
rect 25508 12124 26460 12180
rect 26516 12124 26526 12180
rect 28140 12068 28196 12236
rect 29698 12124 29708 12180
rect 29764 12124 30828 12180
rect 30884 12124 31612 12180
rect 31668 12124 31678 12180
rect 37426 12124 37436 12180
rect 37492 12124 38892 12180
rect 38948 12124 38958 12180
rect 39554 12124 39564 12180
rect 39620 12124 40572 12180
rect 40628 12124 41244 12180
rect 41300 12124 41310 12180
rect 26114 12012 26124 12068
rect 26180 12012 26908 12068
rect 26964 12012 26974 12068
rect 28130 12012 28140 12068
rect 28196 12012 28206 12068
rect 35298 12012 35308 12068
rect 35364 12012 35756 12068
rect 35812 12012 35822 12068
rect 36194 12012 36204 12068
rect 36260 12012 37660 12068
rect 37716 12012 38108 12068
rect 38164 12012 38174 12068
rect 38612 12012 42812 12068
rect 42868 12012 42878 12068
rect 43250 12012 43260 12068
rect 43316 12012 44380 12068
rect 44436 12012 47404 12068
rect 47460 12012 47470 12068
rect 26852 11844 26908 12012
rect 38612 11956 38668 12012
rect 32610 11900 32620 11956
rect 32676 11900 33180 11956
rect 33236 11900 34748 11956
rect 34804 11900 38668 11956
rect 20962 11788 20972 11844
rect 21028 11788 21980 11844
rect 22036 11788 24108 11844
rect 24164 11788 25228 11844
rect 25284 11788 25294 11844
rect 26852 11788 32004 11844
rect 4466 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4750 11788
rect 31948 11732 32004 11788
rect 35186 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35470 11788
rect 31938 11676 31948 11732
rect 32004 11676 32116 11732
rect 37202 11676 37212 11732
rect 37268 11676 38556 11732
rect 38612 11676 39340 11732
rect 39396 11676 39406 11732
rect 32060 11620 32116 11676
rect 32060 11564 38668 11620
rect 40338 11564 40348 11620
rect 40404 11564 41468 11620
rect 41524 11564 41534 11620
rect 44146 11564 44156 11620
rect 44212 11564 45276 11620
rect 45332 11564 45342 11620
rect 38612 11508 38668 11564
rect 18386 11452 18396 11508
rect 18452 11452 24668 11508
rect 24724 11452 24734 11508
rect 37314 11452 37324 11508
rect 37380 11452 37996 11508
rect 38052 11452 38062 11508
rect 38612 11452 39900 11508
rect 39956 11452 43708 11508
rect 37996 11396 38052 11452
rect 43652 11396 43708 11452
rect 18722 11340 18732 11396
rect 18788 11340 20300 11396
rect 20356 11340 20366 11396
rect 28018 11340 28028 11396
rect 28084 11340 29372 11396
rect 29428 11340 30716 11396
rect 30772 11340 30782 11396
rect 31042 11340 31052 11396
rect 31108 11340 33740 11396
rect 33796 11340 33806 11396
rect 37996 11340 42588 11396
rect 42644 11340 42654 11396
rect 43652 11340 44380 11396
rect 44436 11340 44828 11396
rect 44884 11340 44894 11396
rect 21858 11228 21868 11284
rect 21924 11228 25340 11284
rect 25396 11228 25406 11284
rect 29250 11228 29260 11284
rect 29316 11228 31948 11284
rect 32004 11228 32014 11284
rect 38322 11228 38332 11284
rect 38388 11228 38780 11284
rect 38836 11228 39676 11284
rect 39732 11228 40908 11284
rect 40964 11228 40974 11284
rect 45490 11228 45500 11284
rect 45556 11228 46060 11284
rect 46116 11228 46126 11284
rect 19842 11116 19852 11172
rect 19908 11116 25004 11172
rect 25060 11116 25070 11172
rect 37090 11116 37100 11172
rect 37156 11116 40796 11172
rect 40852 11116 42140 11172
rect 42196 11116 42206 11172
rect 45378 11116 45388 11172
rect 45444 11116 45836 11172
rect 45892 11116 45902 11172
rect 38098 11004 38108 11060
rect 38164 11004 40012 11060
rect 40068 11004 40078 11060
rect 19826 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20110 11004
rect 50546 10948 50556 11004
rect 50612 10948 50660 11004
rect 50716 10948 50764 11004
rect 50820 10948 50830 11004
rect 30706 10668 30716 10724
rect 30772 10668 33068 10724
rect 33124 10668 33134 10724
rect 35746 10668 35756 10724
rect 35812 10668 36764 10724
rect 36820 10668 36830 10724
rect 25442 10556 25452 10612
rect 25508 10556 27020 10612
rect 27076 10556 27086 10612
rect 35634 10556 35644 10612
rect 35700 10556 37212 10612
rect 37268 10556 37278 10612
rect 41906 10556 41916 10612
rect 41972 10556 46508 10612
rect 46564 10556 46574 10612
rect 33730 10444 33740 10500
rect 33796 10444 34748 10500
rect 34804 10444 37660 10500
rect 37716 10444 37726 10500
rect 41570 10444 41580 10500
rect 41636 10444 44828 10500
rect 44884 10444 44894 10500
rect 34962 10332 34972 10388
rect 35028 10332 36204 10388
rect 36260 10332 36270 10388
rect 42354 10220 42364 10276
rect 42420 10220 42812 10276
rect 42868 10220 43036 10276
rect 43092 10220 43102 10276
rect 4466 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4750 10220
rect 35186 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35470 10220
rect 30818 10108 30828 10164
rect 30884 10108 32396 10164
rect 32452 10108 32462 10164
rect 38546 10108 38556 10164
rect 38612 10108 38780 10164
rect 38836 10108 38846 10164
rect 43586 10108 43596 10164
rect 43652 10108 44156 10164
rect 44212 10108 44222 10164
rect 25106 9996 25116 10052
rect 25172 9996 25564 10052
rect 25620 9996 26572 10052
rect 26628 9996 26638 10052
rect 28130 9996 28140 10052
rect 28196 9996 28812 10052
rect 28868 9996 28878 10052
rect 27906 9884 27916 9940
rect 27972 9884 29260 9940
rect 29316 9884 29326 9940
rect 33170 9884 33180 9940
rect 33236 9884 33516 9940
rect 33572 9884 33582 9940
rect 36418 9884 36428 9940
rect 36484 9884 36988 9940
rect 37044 9884 37054 9940
rect 28690 9772 28700 9828
rect 28756 9772 31276 9828
rect 31332 9772 31342 9828
rect 32498 9772 32508 9828
rect 32564 9772 33628 9828
rect 33684 9772 34188 9828
rect 34244 9772 34254 9828
rect 22978 9660 22988 9716
rect 23044 9660 24444 9716
rect 24500 9660 24510 9716
rect 21634 9548 21644 9604
rect 21700 9548 29708 9604
rect 29764 9548 30380 9604
rect 30436 9548 38892 9604
rect 38948 9548 40908 9604
rect 40964 9548 40974 9604
rect 37762 9436 37772 9492
rect 37828 9436 38108 9492
rect 38164 9436 38174 9492
rect 19826 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20110 9436
rect 50546 9380 50556 9436
rect 50612 9380 50660 9436
rect 50716 9380 50764 9436
rect 50820 9380 50830 9436
rect 36194 9212 36204 9268
rect 36260 9212 38332 9268
rect 38388 9212 39228 9268
rect 39284 9212 41916 9268
rect 41972 9212 41982 9268
rect 19618 9100 19628 9156
rect 19684 9100 22988 9156
rect 23044 9100 23054 9156
rect 38434 9100 38444 9156
rect 38500 9100 39676 9156
rect 39732 9100 39742 9156
rect 23874 8988 23884 9044
rect 23940 8988 25004 9044
rect 25060 8988 26236 9044
rect 26292 8988 26302 9044
rect 27794 8988 27804 9044
rect 27860 8988 28364 9044
rect 28420 8988 28430 9044
rect 40226 8988 40236 9044
rect 40292 8988 41356 9044
rect 41412 8988 41422 9044
rect 42252 8988 42364 9044
rect 42420 8988 44828 9044
rect 44884 8988 44894 9044
rect 20514 8876 20524 8932
rect 20580 8876 22988 8932
rect 23044 8876 23054 8932
rect 23426 8876 23436 8932
rect 23492 8876 24220 8932
rect 24276 8876 24286 8932
rect 30818 8876 30828 8932
rect 30884 8876 31612 8932
rect 31668 8876 33180 8932
rect 33236 8876 36316 8932
rect 36372 8876 36988 8932
rect 37044 8876 37054 8932
rect 4466 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4750 8652
rect 35186 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35470 8652
rect 42252 8372 42308 8988
rect 40338 8316 40348 8372
rect 40404 8316 42308 8372
rect 46162 8316 46172 8372
rect 46228 8316 47852 8372
rect 47908 8316 47918 8372
rect 41458 8204 41468 8260
rect 41524 8204 42364 8260
rect 42420 8204 43596 8260
rect 43652 8204 43662 8260
rect 36418 8092 36428 8148
rect 36484 8092 37772 8148
rect 37828 8092 37838 8148
rect 43362 8092 43372 8148
rect 43428 8092 44268 8148
rect 44324 8092 44334 8148
rect 19826 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20110 7868
rect 50546 7812 50556 7868
rect 50612 7812 50660 7868
rect 50716 7812 50764 7868
rect 50820 7812 50830 7868
rect 43698 7644 43708 7700
rect 43764 7644 45612 7700
rect 45668 7644 45678 7700
rect 45266 7532 45276 7588
rect 45332 7532 46172 7588
rect 46228 7532 46238 7588
rect 44258 7308 44268 7364
rect 44324 7308 45164 7364
rect 45220 7308 45612 7364
rect 45668 7308 45678 7364
rect 42130 7196 42140 7252
rect 42196 7196 43148 7252
rect 43204 7196 43214 7252
rect 4466 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4750 7084
rect 35186 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35470 7084
rect 45154 6972 45164 7028
rect 45220 6972 46060 7028
rect 46116 6972 46126 7028
rect 19826 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20110 6300
rect 50546 6244 50556 6300
rect 50612 6244 50660 6300
rect 50716 6244 50764 6300
rect 50820 6244 50830 6300
rect 42578 6076 42588 6132
rect 42644 6076 43708 6132
rect 43764 6076 43774 6132
rect 4466 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4750 5516
rect 35186 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35470 5516
rect 34850 4956 34860 5012
rect 34916 4956 38220 5012
rect 38276 4956 38286 5012
rect 19826 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20110 4732
rect 50546 4676 50556 4732
rect 50612 4676 50660 4732
rect 50716 4676 50764 4732
rect 50820 4676 50830 4732
rect 25106 4284 25116 4340
rect 25172 4284 27244 4340
rect 27300 4284 27310 4340
rect 27122 4060 27132 4116
rect 27188 4060 28140 4116
rect 28196 4060 28206 4116
rect 4466 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4750 3948
rect 35186 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35470 3948
rect 26226 3612 26236 3668
rect 26292 3612 29372 3668
rect 29428 3612 29438 3668
rect 27234 3500 27244 3556
rect 27300 3500 28364 3556
rect 28420 3500 28430 3556
rect 13458 3388 13468 3444
rect 13524 3388 16380 3444
rect 16436 3388 16446 3444
rect 17714 3388 17724 3444
rect 17780 3388 19180 3444
rect 19236 3388 19246 3444
rect 19618 3388 19628 3444
rect 19684 3388 19852 3444
rect 19908 3388 19918 3444
rect 20178 3388 20188 3444
rect 20244 3388 21868 3444
rect 21924 3388 21934 3444
rect 26786 3388 26796 3444
rect 26852 3388 27580 3444
rect 27636 3388 27646 3444
rect 34150 3388 34188 3444
rect 34244 3388 34254 3444
rect 36278 3388 36316 3444
rect 36372 3388 36382 3444
rect 37202 3388 37212 3444
rect 37268 3388 37884 3444
rect 37940 3388 37950 3444
rect 43026 3388 43036 3444
rect 43092 3388 43372 3444
rect 43428 3388 43932 3444
rect 43988 3388 43998 3444
rect 19826 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20110 3164
rect 50546 3108 50556 3164
rect 50612 3108 50660 3164
rect 50716 3108 50764 3164
rect 50820 3108 50830 3164
<< via3 >>
rect 19836 76804 19892 76860
rect 19940 76804 19996 76860
rect 20044 76804 20100 76860
rect 50556 76804 50612 76860
rect 50660 76804 50716 76860
rect 50764 76804 50820 76860
rect 4476 76020 4532 76076
rect 4580 76020 4636 76076
rect 4684 76020 4740 76076
rect 35196 76020 35252 76076
rect 35300 76020 35356 76076
rect 35404 76020 35460 76076
rect 19836 75236 19892 75292
rect 19940 75236 19996 75292
rect 20044 75236 20100 75292
rect 50556 75236 50612 75292
rect 50660 75236 50716 75292
rect 50764 75236 50820 75292
rect 4476 74452 4532 74508
rect 4580 74452 4636 74508
rect 4684 74452 4740 74508
rect 35196 74452 35252 74508
rect 35300 74452 35356 74508
rect 35404 74452 35460 74508
rect 19836 73668 19892 73724
rect 19940 73668 19996 73724
rect 20044 73668 20100 73724
rect 50556 73668 50612 73724
rect 50660 73668 50716 73724
rect 50764 73668 50820 73724
rect 4476 72884 4532 72940
rect 4580 72884 4636 72940
rect 4684 72884 4740 72940
rect 35196 72884 35252 72940
rect 35300 72884 35356 72940
rect 35404 72884 35460 72940
rect 19836 72100 19892 72156
rect 19940 72100 19996 72156
rect 20044 72100 20100 72156
rect 50556 72100 50612 72156
rect 50660 72100 50716 72156
rect 50764 72100 50820 72156
rect 4476 71316 4532 71372
rect 4580 71316 4636 71372
rect 4684 71316 4740 71372
rect 35196 71316 35252 71372
rect 35300 71316 35356 71372
rect 35404 71316 35460 71372
rect 19836 70532 19892 70588
rect 19940 70532 19996 70588
rect 20044 70532 20100 70588
rect 50556 70532 50612 70588
rect 50660 70532 50716 70588
rect 50764 70532 50820 70588
rect 4476 69748 4532 69804
rect 4580 69748 4636 69804
rect 4684 69748 4740 69804
rect 35196 69748 35252 69804
rect 35300 69748 35356 69804
rect 35404 69748 35460 69804
rect 29260 69132 29316 69188
rect 42140 69132 42196 69188
rect 19836 68964 19892 69020
rect 19940 68964 19996 69020
rect 20044 68964 20100 69020
rect 50556 68964 50612 69020
rect 50660 68964 50716 69020
rect 50764 68964 50820 69020
rect 4476 68180 4532 68236
rect 4580 68180 4636 68236
rect 4684 68180 4740 68236
rect 35196 68180 35252 68236
rect 35300 68180 35356 68236
rect 35404 68180 35460 68236
rect 25452 67788 25508 67844
rect 42140 67452 42196 67508
rect 19836 67396 19892 67452
rect 19940 67396 19996 67452
rect 20044 67396 20100 67452
rect 50556 67396 50612 67452
rect 50660 67396 50716 67452
rect 50764 67396 50820 67452
rect 29260 67228 29316 67284
rect 39452 66780 39508 66836
rect 4476 66612 4532 66668
rect 4580 66612 4636 66668
rect 4684 66612 4740 66668
rect 35196 66612 35252 66668
rect 35300 66612 35356 66668
rect 35404 66612 35460 66668
rect 34188 66444 34244 66500
rect 41244 66220 41300 66276
rect 25452 66108 25508 66164
rect 19836 65828 19892 65884
rect 19940 65828 19996 65884
rect 20044 65828 20100 65884
rect 50556 65828 50612 65884
rect 50660 65828 50716 65884
rect 50764 65828 50820 65884
rect 4476 65044 4532 65100
rect 4580 65044 4636 65100
rect 4684 65044 4740 65100
rect 35196 65044 35252 65100
rect 35300 65044 35356 65100
rect 35404 65044 35460 65100
rect 19836 64260 19892 64316
rect 19940 64260 19996 64316
rect 20044 64260 20100 64316
rect 50556 64260 50612 64316
rect 50660 64260 50716 64316
rect 50764 64260 50820 64316
rect 41244 64092 41300 64148
rect 34188 63980 34244 64036
rect 4476 63476 4532 63532
rect 4580 63476 4636 63532
rect 4684 63476 4740 63532
rect 35196 63476 35252 63532
rect 35300 63476 35356 63532
rect 35404 63476 35460 63532
rect 40012 63420 40068 63476
rect 44268 62860 44324 62916
rect 19836 62692 19892 62748
rect 19940 62692 19996 62748
rect 20044 62692 20100 62748
rect 50556 62692 50612 62748
rect 50660 62692 50716 62748
rect 50764 62692 50820 62748
rect 43260 62524 43316 62580
rect 40012 62076 40068 62132
rect 4476 61908 4532 61964
rect 4580 61908 4636 61964
rect 4684 61908 4740 61964
rect 34188 61964 34244 62020
rect 35196 61908 35252 61964
rect 35300 61908 35356 61964
rect 35404 61908 35460 61964
rect 28476 61292 28532 61348
rect 42588 61180 42644 61236
rect 19836 61124 19892 61180
rect 19940 61124 19996 61180
rect 20044 61124 20100 61180
rect 50556 61124 50612 61180
rect 50660 61124 50716 61180
rect 50764 61124 50820 61180
rect 33964 61068 34020 61124
rect 42140 61068 42196 61124
rect 4476 60340 4532 60396
rect 4580 60340 4636 60396
rect 4684 60340 4740 60396
rect 35196 60340 35252 60396
rect 35300 60340 35356 60396
rect 35404 60340 35460 60396
rect 39340 60396 39396 60452
rect 19836 59556 19892 59612
rect 19940 59556 19996 59612
rect 20044 59556 20100 59612
rect 39452 59612 39508 59668
rect 50556 59556 50612 59612
rect 50660 59556 50716 59612
rect 50764 59556 50820 59612
rect 21532 59500 21588 59556
rect 39340 59388 39396 59444
rect 28476 59276 28532 59332
rect 4476 58772 4532 58828
rect 4580 58772 4636 58828
rect 4684 58772 4740 58828
rect 35196 58772 35252 58828
rect 35300 58772 35356 58828
rect 35404 58772 35460 58828
rect 43260 58940 43316 58996
rect 44268 58940 44324 58996
rect 42588 58828 42644 58884
rect 45948 58604 46004 58660
rect 44940 58044 44996 58100
rect 19836 57988 19892 58044
rect 19940 57988 19996 58044
rect 20044 57988 20100 58044
rect 50556 57988 50612 58044
rect 50660 57988 50716 58044
rect 50764 57988 50820 58044
rect 44940 57820 44996 57876
rect 23996 57708 24052 57764
rect 4476 57204 4532 57260
rect 4580 57204 4636 57260
rect 4684 57204 4740 57260
rect 35196 57204 35252 57260
rect 35300 57204 35356 57260
rect 35404 57204 35460 57260
rect 33964 56924 34020 56980
rect 19836 56420 19892 56476
rect 19940 56420 19996 56476
rect 20044 56420 20100 56476
rect 50556 56420 50612 56476
rect 50660 56420 50716 56476
rect 50764 56420 50820 56476
rect 45500 56364 45556 56420
rect 42700 56140 42756 56196
rect 4476 55636 4532 55692
rect 4580 55636 4636 55692
rect 4684 55636 4740 55692
rect 35196 55636 35252 55692
rect 35300 55636 35356 55692
rect 35404 55636 35460 55692
rect 27804 55468 27860 55524
rect 17388 55020 17444 55076
rect 33852 55020 33908 55076
rect 41804 55020 41860 55076
rect 19836 54852 19892 54908
rect 19940 54852 19996 54908
rect 20044 54852 20100 54908
rect 50556 54852 50612 54908
rect 50660 54852 50716 54908
rect 50764 54852 50820 54908
rect 23996 54796 24052 54852
rect 39676 54460 39732 54516
rect 4476 54068 4532 54124
rect 4580 54068 4636 54124
rect 4684 54068 4740 54124
rect 35196 54068 35252 54124
rect 35300 54068 35356 54124
rect 35404 54068 35460 54124
rect 28588 53900 28644 53956
rect 19836 53284 19892 53340
rect 19940 53284 19996 53340
rect 20044 53284 20100 53340
rect 50556 53284 50612 53340
rect 50660 53284 50716 53340
rect 50764 53284 50820 53340
rect 41804 53004 41860 53060
rect 42700 52892 42756 52948
rect 26796 52668 26852 52724
rect 4476 52500 4532 52556
rect 4580 52500 4636 52556
rect 4684 52500 4740 52556
rect 35196 52500 35252 52556
rect 35300 52500 35356 52556
rect 35404 52500 35460 52556
rect 21532 52220 21588 52276
rect 38668 52108 38724 52164
rect 39452 51996 39508 52052
rect 19836 51716 19892 51772
rect 19940 51716 19996 51772
rect 20044 51716 20100 51772
rect 50556 51716 50612 51772
rect 50660 51716 50716 51772
rect 50764 51716 50820 51772
rect 33964 51548 34020 51604
rect 23772 51324 23828 51380
rect 39452 51324 39508 51380
rect 40012 51324 40068 51380
rect 39676 51100 39732 51156
rect 4476 50932 4532 50988
rect 4580 50932 4636 50988
rect 4684 50932 4740 50988
rect 35196 50932 35252 50988
rect 35300 50932 35356 50988
rect 35404 50932 35460 50988
rect 21532 50876 21588 50932
rect 19836 50148 19892 50204
rect 19940 50148 19996 50204
rect 20044 50148 20100 50204
rect 50556 50148 50612 50204
rect 50660 50148 50716 50204
rect 50764 50148 50820 50204
rect 45948 49980 46004 50036
rect 40012 49756 40068 49812
rect 17836 49532 17892 49588
rect 4476 49364 4532 49420
rect 4580 49364 4636 49420
rect 4684 49364 4740 49420
rect 35196 49364 35252 49420
rect 35300 49364 35356 49420
rect 35404 49364 35460 49420
rect 31948 48748 32004 48804
rect 19836 48580 19892 48636
rect 19940 48580 19996 48636
rect 20044 48580 20100 48636
rect 50556 48580 50612 48636
rect 50660 48580 50716 48636
rect 50764 48580 50820 48636
rect 45500 48412 45556 48468
rect 33852 47852 33908 47908
rect 4476 47796 4532 47852
rect 4580 47796 4636 47852
rect 4684 47796 4740 47852
rect 35196 47796 35252 47852
rect 35300 47796 35356 47852
rect 35404 47796 35460 47852
rect 17836 47740 17892 47796
rect 27804 47740 27860 47796
rect 19836 47012 19892 47068
rect 19940 47012 19996 47068
rect 20044 47012 20100 47068
rect 36876 47068 36932 47124
rect 50556 47012 50612 47068
rect 50660 47012 50716 47068
rect 50764 47012 50820 47068
rect 34636 46956 34692 47012
rect 4476 46228 4532 46284
rect 4580 46228 4636 46284
rect 4684 46228 4740 46284
rect 35196 46228 35252 46284
rect 35300 46228 35356 46284
rect 35404 46228 35460 46284
rect 33964 45948 34020 46004
rect 22092 45612 22148 45668
rect 23100 45612 23156 45668
rect 19836 45444 19892 45500
rect 19940 45444 19996 45500
rect 20044 45444 20100 45500
rect 50556 45444 50612 45500
rect 50660 45444 50716 45500
rect 50764 45444 50820 45500
rect 4476 44660 4532 44716
rect 4580 44660 4636 44716
rect 4684 44660 4740 44716
rect 35196 44660 35252 44716
rect 35300 44660 35356 44716
rect 35404 44660 35460 44716
rect 34748 44492 34804 44548
rect 34524 44380 34580 44436
rect 38668 44156 38724 44212
rect 19836 43876 19892 43932
rect 19940 43876 19996 43932
rect 20044 43876 20100 43932
rect 26460 44044 26516 44100
rect 29260 44044 29316 44100
rect 50556 43876 50612 43932
rect 50660 43876 50716 43932
rect 50764 43876 50820 43932
rect 20524 43596 20580 43652
rect 19180 43484 19236 43540
rect 36876 43372 36932 43428
rect 34524 43148 34580 43204
rect 4476 43092 4532 43148
rect 4580 43092 4636 43148
rect 4684 43092 4740 43148
rect 35196 43092 35252 43148
rect 35300 43092 35356 43148
rect 35404 43092 35460 43148
rect 23772 42812 23828 42868
rect 25900 42476 25956 42532
rect 19836 42308 19892 42364
rect 19940 42308 19996 42364
rect 20044 42308 20100 42364
rect 50556 42308 50612 42364
rect 50660 42308 50716 42364
rect 50764 42308 50820 42364
rect 29820 41916 29876 41972
rect 33628 41916 33684 41972
rect 29372 41804 29428 41860
rect 4476 41524 4532 41580
rect 4580 41524 4636 41580
rect 4684 41524 4740 41580
rect 29484 41580 29540 41636
rect 35196 41524 35252 41580
rect 35300 41524 35356 41580
rect 35404 41524 35460 41580
rect 33852 41468 33908 41524
rect 29484 41132 29540 41188
rect 26012 41020 26068 41076
rect 34972 40908 35028 40964
rect 19836 40740 19892 40796
rect 19940 40740 19996 40796
rect 20044 40740 20100 40796
rect 50556 40740 50612 40796
rect 50660 40740 50716 40796
rect 50764 40740 50820 40796
rect 29820 40684 29876 40740
rect 30604 40460 30660 40516
rect 4476 39956 4532 40012
rect 4580 39956 4636 40012
rect 4684 39956 4740 40012
rect 35196 39956 35252 40012
rect 35300 39956 35356 40012
rect 35404 39956 35460 40012
rect 29820 39452 29876 39508
rect 19836 39172 19892 39228
rect 19940 39172 19996 39228
rect 20044 39172 20100 39228
rect 50556 39172 50612 39228
rect 50660 39172 50716 39228
rect 50764 39172 50820 39228
rect 29372 38892 29428 38948
rect 4476 38388 4532 38444
rect 4580 38388 4636 38444
rect 4684 38388 4740 38444
rect 35196 38388 35252 38444
rect 35300 38388 35356 38444
rect 35404 38388 35460 38444
rect 34636 38220 34692 38276
rect 22092 38108 22148 38164
rect 23100 37996 23156 38052
rect 33852 37996 33908 38052
rect 33964 37884 34020 37940
rect 19836 37604 19892 37660
rect 19940 37604 19996 37660
rect 20044 37604 20100 37660
rect 50556 37604 50612 37660
rect 50660 37604 50716 37660
rect 50764 37604 50820 37660
rect 22092 37548 22148 37604
rect 20524 36876 20580 36932
rect 4476 36820 4532 36876
rect 4580 36820 4636 36876
rect 4684 36820 4740 36876
rect 35196 36820 35252 36876
rect 35300 36820 35356 36876
rect 35404 36820 35460 36876
rect 23996 36428 24052 36484
rect 19836 36036 19892 36092
rect 19940 36036 19996 36092
rect 20044 36036 20100 36092
rect 23772 35868 23828 35924
rect 23996 35868 24052 35924
rect 50556 36036 50612 36092
rect 50660 36036 50716 36092
rect 50764 36036 50820 36092
rect 19180 35756 19236 35812
rect 29260 35644 29316 35700
rect 34748 35532 34804 35588
rect 46172 35532 46228 35588
rect 4476 35252 4532 35308
rect 4580 35252 4636 35308
rect 4684 35252 4740 35308
rect 35196 35252 35252 35308
rect 35300 35252 35356 35308
rect 35404 35252 35460 35308
rect 24556 35084 24612 35140
rect 17388 34636 17444 34692
rect 19836 34468 19892 34524
rect 19940 34468 19996 34524
rect 20044 34468 20100 34524
rect 50556 34468 50612 34524
rect 50660 34468 50716 34524
rect 50764 34468 50820 34524
rect 25228 34412 25284 34468
rect 35756 34300 35812 34356
rect 28588 33964 28644 34020
rect 48412 33964 48468 34020
rect 4476 33684 4532 33740
rect 4580 33684 4636 33740
rect 4684 33684 4740 33740
rect 35196 33684 35252 33740
rect 35300 33684 35356 33740
rect 35404 33684 35460 33740
rect 33628 33628 33684 33684
rect 36652 33404 36708 33460
rect 19836 32900 19892 32956
rect 19940 32900 19996 32956
rect 20044 32900 20100 32956
rect 50556 32900 50612 32956
rect 50660 32900 50716 32956
rect 50764 32900 50820 32956
rect 25788 32732 25844 32788
rect 48524 32396 48580 32452
rect 21308 32172 21364 32228
rect 31948 32172 32004 32228
rect 4476 32116 4532 32172
rect 4580 32116 4636 32172
rect 4684 32116 4740 32172
rect 35196 32116 35252 32172
rect 35300 32116 35356 32172
rect 35404 32116 35460 32172
rect 25340 31948 25396 32004
rect 39452 31948 39508 32004
rect 28140 31724 28196 31780
rect 38892 31500 38948 31556
rect 19836 31332 19892 31388
rect 19940 31332 19996 31388
rect 20044 31332 20100 31388
rect 25228 31276 25284 31332
rect 25788 31276 25844 31332
rect 50556 31332 50612 31388
rect 50660 31332 50716 31388
rect 50764 31332 50820 31388
rect 4476 30548 4532 30604
rect 4580 30548 4636 30604
rect 4684 30548 4740 30604
rect 35196 30548 35252 30604
rect 35300 30548 35356 30604
rect 35404 30548 35460 30604
rect 35756 30492 35812 30548
rect 19404 30268 19460 30324
rect 38892 30156 38948 30212
rect 46172 30044 46228 30100
rect 47628 30044 47684 30100
rect 25116 29932 25172 29988
rect 19836 29764 19892 29820
rect 19940 29764 19996 29820
rect 20044 29764 20100 29820
rect 50556 29764 50612 29820
rect 50660 29764 50716 29820
rect 50764 29764 50820 29820
rect 47628 29708 47684 29764
rect 21308 29596 21364 29652
rect 25900 29484 25956 29540
rect 25340 29148 25396 29204
rect 39452 29148 39508 29204
rect 4476 28980 4532 29036
rect 4580 28980 4636 29036
rect 4684 28980 4740 29036
rect 35196 28980 35252 29036
rect 35300 28980 35356 29036
rect 35404 28980 35460 29036
rect 22092 28476 22148 28532
rect 19836 28196 19892 28252
rect 19940 28196 19996 28252
rect 20044 28196 20100 28252
rect 50556 28196 50612 28252
rect 50660 28196 50716 28252
rect 50764 28196 50820 28252
rect 26796 28028 26852 28084
rect 36652 27916 36708 27972
rect 4476 27412 4532 27468
rect 4580 27412 4636 27468
rect 4684 27412 4740 27468
rect 35196 27412 35252 27468
rect 35300 27412 35356 27468
rect 35404 27412 35460 27468
rect 34748 27356 34804 27412
rect 23436 27244 23492 27300
rect 23996 27244 24052 27300
rect 19836 26628 19892 26684
rect 19940 26628 19996 26684
rect 20044 26628 20100 26684
rect 50556 26628 50612 26684
rect 50660 26628 50716 26684
rect 50764 26628 50820 26684
rect 23436 26460 23492 26516
rect 26012 26460 26068 26516
rect 48412 26348 48468 26404
rect 36316 26236 36372 26292
rect 30716 26124 30772 26180
rect 48524 26124 48580 26180
rect 4476 25844 4532 25900
rect 4580 25844 4636 25900
rect 4684 25844 4740 25900
rect 35196 25844 35252 25900
rect 35300 25844 35356 25900
rect 35404 25844 35460 25900
rect 26460 25676 26516 25732
rect 23996 25564 24052 25620
rect 19404 25452 19460 25508
rect 30716 25452 30772 25508
rect 28140 25340 28196 25396
rect 34188 25340 34244 25396
rect 19836 25060 19892 25116
rect 19940 25060 19996 25116
rect 20044 25060 20100 25116
rect 50556 25060 50612 25116
rect 50660 25060 50716 25116
rect 50764 25060 50820 25116
rect 36764 25004 36820 25060
rect 34748 24892 34804 24948
rect 24556 24780 24612 24836
rect 31948 24556 32004 24612
rect 34188 24556 34244 24612
rect 4476 24276 4532 24332
rect 4580 24276 4636 24332
rect 4684 24276 4740 24332
rect 35196 24276 35252 24332
rect 35300 24276 35356 24332
rect 35404 24276 35460 24332
rect 36764 23548 36820 23604
rect 19836 23492 19892 23548
rect 19940 23492 19996 23548
rect 20044 23492 20100 23548
rect 50556 23492 50612 23548
rect 50660 23492 50716 23548
rect 50764 23492 50820 23548
rect 21868 23324 21924 23380
rect 27804 22988 27860 23044
rect 4476 22708 4532 22764
rect 4580 22708 4636 22764
rect 4684 22708 4740 22764
rect 27356 22764 27412 22820
rect 35196 22708 35252 22764
rect 35300 22708 35356 22764
rect 35404 22708 35460 22764
rect 19628 22316 19684 22372
rect 19836 21924 19892 21980
rect 19940 21924 19996 21980
rect 20044 21924 20100 21980
rect 50556 21924 50612 21980
rect 50660 21924 50716 21980
rect 50764 21924 50820 21980
rect 34972 21532 35028 21588
rect 4476 21140 4532 21196
rect 4580 21140 4636 21196
rect 4684 21140 4740 21196
rect 35196 21140 35252 21196
rect 35300 21140 35356 21196
rect 35404 21140 35460 21196
rect 34972 20636 35028 20692
rect 27804 20524 27860 20580
rect 19836 20356 19892 20412
rect 19940 20356 19996 20412
rect 20044 20356 20100 20412
rect 50556 20356 50612 20412
rect 50660 20356 50716 20412
rect 50764 20356 50820 20412
rect 33628 20300 33684 20356
rect 4476 19572 4532 19628
rect 4580 19572 4636 19628
rect 4684 19572 4740 19628
rect 35196 19572 35252 19628
rect 35300 19572 35356 19628
rect 35404 19572 35460 19628
rect 21868 19068 21924 19124
rect 36540 18956 36596 19012
rect 46396 18956 46452 19012
rect 19836 18788 19892 18844
rect 19940 18788 19996 18844
rect 20044 18788 20100 18844
rect 50556 18788 50612 18844
rect 50660 18788 50716 18844
rect 50764 18788 50820 18844
rect 34524 18732 34580 18788
rect 33628 18284 33684 18340
rect 34524 18172 34580 18228
rect 35644 18172 35700 18228
rect 4476 18004 4532 18060
rect 4580 18004 4636 18060
rect 4684 18004 4740 18060
rect 35196 18004 35252 18060
rect 35300 18004 35356 18060
rect 35404 18004 35460 18060
rect 43036 17948 43092 18004
rect 46396 17724 46452 17780
rect 19836 17220 19892 17276
rect 19940 17220 19996 17276
rect 20044 17220 20100 17276
rect 36092 17612 36148 17668
rect 36204 17388 36260 17444
rect 50556 17220 50612 17276
rect 50660 17220 50716 17276
rect 50764 17220 50820 17276
rect 36540 16604 36596 16660
rect 4476 16436 4532 16492
rect 4580 16436 4636 16492
rect 4684 16436 4740 16492
rect 35196 16436 35252 16492
rect 35300 16436 35356 16492
rect 35404 16436 35460 16492
rect 31948 15820 32004 15876
rect 36092 15820 36148 15876
rect 19836 15652 19892 15708
rect 19940 15652 19996 15708
rect 20044 15652 20100 15708
rect 50556 15652 50612 15708
rect 50660 15652 50716 15708
rect 50764 15652 50820 15708
rect 4476 14868 4532 14924
rect 4580 14868 4636 14924
rect 4684 14868 4740 14924
rect 35196 14868 35252 14924
rect 35300 14868 35356 14924
rect 35404 14868 35460 14924
rect 31948 14812 32004 14868
rect 43036 14588 43092 14644
rect 35644 14364 35700 14420
rect 19836 14084 19892 14140
rect 19940 14084 19996 14140
rect 20044 14084 20100 14140
rect 50556 14084 50612 14140
rect 50660 14084 50716 14140
rect 50764 14084 50820 14140
rect 36764 13804 36820 13860
rect 27356 13580 27412 13636
rect 4476 13300 4532 13356
rect 4580 13300 4636 13356
rect 4684 13300 4740 13356
rect 35196 13300 35252 13356
rect 35300 13300 35356 13356
rect 35404 13300 35460 13356
rect 36204 13020 36260 13076
rect 19836 12516 19892 12572
rect 19940 12516 19996 12572
rect 20044 12516 20100 12572
rect 50556 12516 50612 12572
rect 50660 12516 50716 12572
rect 50764 12516 50820 12572
rect 4476 11732 4532 11788
rect 4580 11732 4636 11788
rect 4684 11732 4740 11788
rect 35196 11732 35252 11788
rect 35300 11732 35356 11788
rect 35404 11732 35460 11788
rect 19836 10948 19892 11004
rect 19940 10948 19996 11004
rect 20044 10948 20100 11004
rect 50556 10948 50612 11004
rect 50660 10948 50716 11004
rect 50764 10948 50820 11004
rect 4476 10164 4532 10220
rect 4580 10164 4636 10220
rect 4684 10164 4740 10220
rect 35196 10164 35252 10220
rect 35300 10164 35356 10220
rect 35404 10164 35460 10220
rect 19836 9380 19892 9436
rect 19940 9380 19996 9436
rect 20044 9380 20100 9436
rect 50556 9380 50612 9436
rect 50660 9380 50716 9436
rect 50764 9380 50820 9436
rect 4476 8596 4532 8652
rect 4580 8596 4636 8652
rect 4684 8596 4740 8652
rect 35196 8596 35252 8652
rect 35300 8596 35356 8652
rect 35404 8596 35460 8652
rect 19836 7812 19892 7868
rect 19940 7812 19996 7868
rect 20044 7812 20100 7868
rect 50556 7812 50612 7868
rect 50660 7812 50716 7868
rect 50764 7812 50820 7868
rect 4476 7028 4532 7084
rect 4580 7028 4636 7084
rect 4684 7028 4740 7084
rect 35196 7028 35252 7084
rect 35300 7028 35356 7084
rect 35404 7028 35460 7084
rect 19836 6244 19892 6300
rect 19940 6244 19996 6300
rect 20044 6244 20100 6300
rect 50556 6244 50612 6300
rect 50660 6244 50716 6300
rect 50764 6244 50820 6300
rect 4476 5460 4532 5516
rect 4580 5460 4636 5516
rect 4684 5460 4740 5516
rect 35196 5460 35252 5516
rect 35300 5460 35356 5516
rect 35404 5460 35460 5516
rect 19836 4676 19892 4732
rect 19940 4676 19996 4732
rect 20044 4676 20100 4732
rect 50556 4676 50612 4732
rect 50660 4676 50716 4732
rect 50764 4676 50820 4732
rect 25116 4284 25172 4340
rect 4476 3892 4532 3948
rect 4580 3892 4636 3948
rect 4684 3892 4740 3948
rect 35196 3892 35252 3948
rect 35300 3892 35356 3948
rect 35404 3892 35460 3948
rect 19628 3388 19684 3444
rect 34188 3388 34244 3444
rect 36316 3388 36372 3444
rect 19836 3108 19892 3164
rect 19940 3108 19996 3164
rect 20044 3108 20100 3164
rect 50556 3108 50612 3164
rect 50660 3108 50716 3164
rect 50764 3108 50820 3164
<< metal4 >>
rect 4448 76076 4768 76892
rect 4448 76020 4476 76076
rect 4532 76020 4580 76076
rect 4636 76020 4684 76076
rect 4740 76020 4768 76076
rect 4448 74508 4768 76020
rect 4448 74452 4476 74508
rect 4532 74452 4580 74508
rect 4636 74452 4684 74508
rect 4740 74452 4768 74508
rect 4448 72940 4768 74452
rect 4448 72884 4476 72940
rect 4532 72884 4580 72940
rect 4636 72884 4684 72940
rect 4740 72884 4768 72940
rect 4448 71372 4768 72884
rect 4448 71316 4476 71372
rect 4532 71316 4580 71372
rect 4636 71316 4684 71372
rect 4740 71316 4768 71372
rect 4448 69804 4768 71316
rect 4448 69748 4476 69804
rect 4532 69748 4580 69804
rect 4636 69748 4684 69804
rect 4740 69748 4768 69804
rect 4448 68236 4768 69748
rect 4448 68180 4476 68236
rect 4532 68180 4580 68236
rect 4636 68180 4684 68236
rect 4740 68180 4768 68236
rect 4448 66668 4768 68180
rect 4448 66612 4476 66668
rect 4532 66612 4580 66668
rect 4636 66612 4684 66668
rect 4740 66612 4768 66668
rect 4448 65100 4768 66612
rect 4448 65044 4476 65100
rect 4532 65044 4580 65100
rect 4636 65044 4684 65100
rect 4740 65044 4768 65100
rect 4448 63532 4768 65044
rect 4448 63476 4476 63532
rect 4532 63476 4580 63532
rect 4636 63476 4684 63532
rect 4740 63476 4768 63532
rect 4448 61964 4768 63476
rect 4448 61908 4476 61964
rect 4532 61908 4580 61964
rect 4636 61908 4684 61964
rect 4740 61908 4768 61964
rect 4448 60396 4768 61908
rect 4448 60340 4476 60396
rect 4532 60340 4580 60396
rect 4636 60340 4684 60396
rect 4740 60340 4768 60396
rect 4448 58828 4768 60340
rect 4448 58772 4476 58828
rect 4532 58772 4580 58828
rect 4636 58772 4684 58828
rect 4740 58772 4768 58828
rect 4448 57260 4768 58772
rect 4448 57204 4476 57260
rect 4532 57204 4580 57260
rect 4636 57204 4684 57260
rect 4740 57204 4768 57260
rect 4448 55692 4768 57204
rect 4448 55636 4476 55692
rect 4532 55636 4580 55692
rect 4636 55636 4684 55692
rect 4740 55636 4768 55692
rect 4448 54124 4768 55636
rect 19808 76860 20128 76892
rect 19808 76804 19836 76860
rect 19892 76804 19940 76860
rect 19996 76804 20044 76860
rect 20100 76804 20128 76860
rect 19808 75292 20128 76804
rect 19808 75236 19836 75292
rect 19892 75236 19940 75292
rect 19996 75236 20044 75292
rect 20100 75236 20128 75292
rect 19808 73724 20128 75236
rect 19808 73668 19836 73724
rect 19892 73668 19940 73724
rect 19996 73668 20044 73724
rect 20100 73668 20128 73724
rect 19808 72156 20128 73668
rect 19808 72100 19836 72156
rect 19892 72100 19940 72156
rect 19996 72100 20044 72156
rect 20100 72100 20128 72156
rect 19808 70588 20128 72100
rect 19808 70532 19836 70588
rect 19892 70532 19940 70588
rect 19996 70532 20044 70588
rect 20100 70532 20128 70588
rect 19808 69020 20128 70532
rect 35168 76076 35488 76892
rect 35168 76020 35196 76076
rect 35252 76020 35300 76076
rect 35356 76020 35404 76076
rect 35460 76020 35488 76076
rect 35168 74508 35488 76020
rect 35168 74452 35196 74508
rect 35252 74452 35300 74508
rect 35356 74452 35404 74508
rect 35460 74452 35488 74508
rect 35168 72940 35488 74452
rect 35168 72884 35196 72940
rect 35252 72884 35300 72940
rect 35356 72884 35404 72940
rect 35460 72884 35488 72940
rect 35168 71372 35488 72884
rect 35168 71316 35196 71372
rect 35252 71316 35300 71372
rect 35356 71316 35404 71372
rect 35460 71316 35488 71372
rect 35168 69804 35488 71316
rect 35168 69748 35196 69804
rect 35252 69748 35300 69804
rect 35356 69748 35404 69804
rect 35460 69748 35488 69804
rect 19808 68964 19836 69020
rect 19892 68964 19940 69020
rect 19996 68964 20044 69020
rect 20100 68964 20128 69020
rect 19808 67452 20128 68964
rect 29260 69188 29316 69198
rect 19808 67396 19836 67452
rect 19892 67396 19940 67452
rect 19996 67396 20044 67452
rect 20100 67396 20128 67452
rect 19808 65884 20128 67396
rect 25452 67844 25508 67854
rect 25452 66164 25508 67788
rect 29260 67284 29316 69132
rect 29260 67218 29316 67228
rect 35168 68236 35488 69748
rect 50528 76860 50848 76892
rect 50528 76804 50556 76860
rect 50612 76804 50660 76860
rect 50716 76804 50764 76860
rect 50820 76804 50848 76860
rect 50528 75292 50848 76804
rect 50528 75236 50556 75292
rect 50612 75236 50660 75292
rect 50716 75236 50764 75292
rect 50820 75236 50848 75292
rect 50528 73724 50848 75236
rect 50528 73668 50556 73724
rect 50612 73668 50660 73724
rect 50716 73668 50764 73724
rect 50820 73668 50848 73724
rect 50528 72156 50848 73668
rect 50528 72100 50556 72156
rect 50612 72100 50660 72156
rect 50716 72100 50764 72156
rect 50820 72100 50848 72156
rect 50528 70588 50848 72100
rect 50528 70532 50556 70588
rect 50612 70532 50660 70588
rect 50716 70532 50764 70588
rect 50820 70532 50848 70588
rect 35168 68180 35196 68236
rect 35252 68180 35300 68236
rect 35356 68180 35404 68236
rect 35460 68180 35488 68236
rect 35168 66668 35488 68180
rect 42140 69188 42196 69198
rect 42140 67508 42196 69132
rect 35168 66612 35196 66668
rect 35252 66612 35300 66668
rect 35356 66612 35404 66668
rect 35460 66612 35488 66668
rect 25452 66098 25508 66108
rect 34188 66500 34244 66510
rect 19808 65828 19836 65884
rect 19892 65828 19940 65884
rect 19996 65828 20044 65884
rect 20100 65828 20128 65884
rect 19808 64316 20128 65828
rect 19808 64260 19836 64316
rect 19892 64260 19940 64316
rect 19996 64260 20044 64316
rect 20100 64260 20128 64316
rect 19808 62748 20128 64260
rect 19808 62692 19836 62748
rect 19892 62692 19940 62748
rect 19996 62692 20044 62748
rect 20100 62692 20128 62748
rect 19808 61180 20128 62692
rect 34188 64036 34244 66444
rect 34188 62020 34244 63980
rect 34188 61954 34244 61964
rect 35168 65100 35488 66612
rect 35168 65044 35196 65100
rect 35252 65044 35300 65100
rect 35356 65044 35404 65100
rect 35460 65044 35488 65100
rect 35168 63532 35488 65044
rect 35168 63476 35196 63532
rect 35252 63476 35300 63532
rect 35356 63476 35404 63532
rect 35460 63476 35488 63532
rect 35168 61964 35488 63476
rect 35168 61908 35196 61964
rect 35252 61908 35300 61964
rect 35356 61908 35404 61964
rect 35460 61908 35488 61964
rect 19808 61124 19836 61180
rect 19892 61124 19940 61180
rect 19996 61124 20044 61180
rect 20100 61124 20128 61180
rect 19808 59612 20128 61124
rect 19808 59556 19836 59612
rect 19892 59556 19940 59612
rect 19996 59556 20044 59612
rect 20100 59556 20128 59612
rect 28476 61348 28532 61358
rect 19808 58044 20128 59556
rect 19808 57988 19836 58044
rect 19892 57988 19940 58044
rect 19996 57988 20044 58044
rect 20100 57988 20128 58044
rect 19808 56476 20128 57988
rect 19808 56420 19836 56476
rect 19892 56420 19940 56476
rect 19996 56420 20044 56476
rect 20100 56420 20128 56476
rect 4448 54068 4476 54124
rect 4532 54068 4580 54124
rect 4636 54068 4684 54124
rect 4740 54068 4768 54124
rect 4448 52556 4768 54068
rect 4448 52500 4476 52556
rect 4532 52500 4580 52556
rect 4636 52500 4684 52556
rect 4740 52500 4768 52556
rect 4448 50988 4768 52500
rect 4448 50932 4476 50988
rect 4532 50932 4580 50988
rect 4636 50932 4684 50988
rect 4740 50932 4768 50988
rect 4448 49420 4768 50932
rect 4448 49364 4476 49420
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4740 49364 4768 49420
rect 4448 47852 4768 49364
rect 4448 47796 4476 47852
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4740 47796 4768 47852
rect 4448 46284 4768 47796
rect 4448 46228 4476 46284
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4740 46228 4768 46284
rect 4448 44716 4768 46228
rect 4448 44660 4476 44716
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4740 44660 4768 44716
rect 4448 43148 4768 44660
rect 4448 43092 4476 43148
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4740 43092 4768 43148
rect 4448 41580 4768 43092
rect 4448 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4768 41580
rect 4448 40012 4768 41524
rect 4448 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4768 40012
rect 4448 38444 4768 39956
rect 4448 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4768 38444
rect 4448 36876 4768 38388
rect 4448 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4768 36876
rect 4448 35308 4768 36820
rect 4448 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4768 35308
rect 4448 33740 4768 35252
rect 17388 55076 17444 55086
rect 17388 34692 17444 55020
rect 19808 54908 20128 56420
rect 19808 54852 19836 54908
rect 19892 54852 19940 54908
rect 19996 54852 20044 54908
rect 20100 54852 20128 54908
rect 19808 53340 20128 54852
rect 19808 53284 19836 53340
rect 19892 53284 19940 53340
rect 19996 53284 20044 53340
rect 20100 53284 20128 53340
rect 19808 51772 20128 53284
rect 19808 51716 19836 51772
rect 19892 51716 19940 51772
rect 19996 51716 20044 51772
rect 20100 51716 20128 51772
rect 19808 50204 20128 51716
rect 21532 59556 21588 59566
rect 21532 52276 21588 59500
rect 28476 59332 28532 61292
rect 28476 59266 28532 59276
rect 33964 61124 34020 61134
rect 21532 50932 21588 52220
rect 23996 57764 24052 57774
rect 23996 54852 24052 57708
rect 33964 56980 34020 61068
rect 21532 50866 21588 50876
rect 23772 51380 23828 51390
rect 19808 50148 19836 50204
rect 19892 50148 19940 50204
rect 19996 50148 20044 50204
rect 20100 50148 20128 50204
rect 17836 49588 17892 49598
rect 17836 47796 17892 49532
rect 17836 47730 17892 47740
rect 19808 48636 20128 50148
rect 19808 48580 19836 48636
rect 19892 48580 19940 48636
rect 19996 48580 20044 48636
rect 20100 48580 20128 48636
rect 19808 47068 20128 48580
rect 19808 47012 19836 47068
rect 19892 47012 19940 47068
rect 19996 47012 20044 47068
rect 20100 47012 20128 47068
rect 19808 45500 20128 47012
rect 19808 45444 19836 45500
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 20100 45444 20128 45500
rect 19808 43932 20128 45444
rect 19808 43876 19836 43932
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 20100 43876 20128 43932
rect 19180 43540 19236 43550
rect 19180 35812 19236 43484
rect 19180 35746 19236 35756
rect 19808 42364 20128 43876
rect 22092 45668 22148 45678
rect 19808 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20128 42364
rect 19808 40796 20128 42308
rect 19808 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20128 40796
rect 19808 39228 20128 40740
rect 19808 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20128 39228
rect 19808 37660 20128 39172
rect 19808 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20128 37660
rect 19808 36092 20128 37604
rect 20524 43652 20580 43662
rect 20524 36932 20580 43596
rect 22092 38164 22148 45612
rect 22092 38098 22148 38108
rect 23100 45668 23156 45678
rect 23100 38052 23156 45612
rect 23100 37986 23156 37996
rect 23772 42868 23828 51324
rect 20524 36866 20580 36876
rect 22092 37604 22148 37614
rect 19808 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20128 36092
rect 17388 34626 17444 34636
rect 4448 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4768 33740
rect 4448 32172 4768 33684
rect 4448 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4768 32172
rect 4448 30604 4768 32116
rect 4448 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4768 30604
rect 4448 29036 4768 30548
rect 19808 34524 20128 36036
rect 19808 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20128 34524
rect 19808 32956 20128 34468
rect 19808 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20128 32956
rect 19808 31388 20128 32900
rect 19808 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20128 31388
rect 4448 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4768 29036
rect 4448 27468 4768 28980
rect 4448 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4768 27468
rect 4448 25900 4768 27412
rect 4448 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4768 25900
rect 4448 24332 4768 25844
rect 19404 30324 19460 30334
rect 19404 25508 19460 30268
rect 19404 25442 19460 25452
rect 19808 29820 20128 31332
rect 19808 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20128 29820
rect 19808 28252 20128 29764
rect 21308 32228 21364 32238
rect 21308 29652 21364 32172
rect 21308 29586 21364 29596
rect 22092 28532 22148 37548
rect 23772 35924 23828 42812
rect 23772 35858 23828 35868
rect 23996 36484 24052 54796
rect 27804 55524 27860 55534
rect 26796 52724 26852 52734
rect 26460 44100 26516 44110
rect 23996 35924 24052 36428
rect 23996 35858 24052 35868
rect 25900 42532 25956 42542
rect 22092 28466 22148 28476
rect 24556 35140 24612 35150
rect 19808 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20128 28252
rect 19808 26684 20128 28196
rect 19808 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20128 26684
rect 4448 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4768 24332
rect 4448 22764 4768 24276
rect 4448 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4768 22764
rect 4448 21196 4768 22708
rect 19808 25116 20128 26628
rect 23436 27300 23492 27310
rect 23436 26516 23492 27244
rect 23436 26450 23492 26460
rect 23996 27300 24052 27310
rect 23996 25620 24052 27244
rect 23996 25554 24052 25564
rect 19808 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20128 25116
rect 19808 23548 20128 25060
rect 24556 24836 24612 35084
rect 25228 34468 25284 34478
rect 25228 31332 25284 34412
rect 25788 32788 25844 32798
rect 25228 31266 25284 31276
rect 25340 32004 25396 32014
rect 24556 24770 24612 24780
rect 25116 29988 25172 29998
rect 19808 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20128 23548
rect 4448 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4768 21196
rect 4448 19628 4768 21140
rect 4448 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4768 19628
rect 4448 18060 4768 19572
rect 4448 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4768 18060
rect 4448 16492 4768 18004
rect 4448 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4768 16492
rect 4448 14924 4768 16436
rect 4448 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4768 14924
rect 4448 13356 4768 14868
rect 4448 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4768 13356
rect 4448 11788 4768 13300
rect 4448 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4768 11788
rect 4448 10220 4768 11732
rect 4448 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4768 10220
rect 4448 8652 4768 10164
rect 4448 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4768 8652
rect 4448 7084 4768 8596
rect 4448 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4768 7084
rect 4448 5516 4768 7028
rect 4448 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4768 5516
rect 4448 3948 4768 5460
rect 4448 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4768 3948
rect 4448 3076 4768 3892
rect 19628 22372 19684 22382
rect 19628 3444 19684 22316
rect 19628 3378 19684 3388
rect 19808 21980 20128 23492
rect 19808 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20128 21980
rect 19808 20412 20128 21924
rect 19808 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20128 20412
rect 19808 18844 20128 20356
rect 21868 23380 21924 23390
rect 21868 19124 21924 23324
rect 21868 19058 21924 19068
rect 19808 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20128 18844
rect 19808 17276 20128 18788
rect 19808 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20128 17276
rect 19808 15708 20128 17220
rect 19808 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20128 15708
rect 19808 14140 20128 15652
rect 19808 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20128 14140
rect 19808 12572 20128 14084
rect 19808 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20128 12572
rect 19808 11004 20128 12516
rect 19808 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20128 11004
rect 19808 9436 20128 10948
rect 19808 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20128 9436
rect 19808 7868 20128 9380
rect 19808 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20128 7868
rect 19808 6300 20128 7812
rect 19808 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20128 6300
rect 19808 4732 20128 6244
rect 19808 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20128 4732
rect 19808 3164 20128 4676
rect 25116 4340 25172 29932
rect 25340 29204 25396 31948
rect 25788 31332 25844 32732
rect 25788 31266 25844 31276
rect 25900 29540 25956 42476
rect 25900 29474 25956 29484
rect 26012 41076 26068 41086
rect 25340 29138 25396 29148
rect 26012 26516 26068 41020
rect 26012 26450 26068 26460
rect 26460 25732 26516 44044
rect 26796 28084 26852 52668
rect 27804 47796 27860 55468
rect 33852 55076 33908 55086
rect 27804 47730 27860 47740
rect 28588 53956 28644 53966
rect 28588 34020 28644 53900
rect 31948 48804 32004 48814
rect 29260 44100 29316 44110
rect 29260 35700 29316 44044
rect 29820 41972 29876 41982
rect 29372 41860 29428 41870
rect 29372 38948 29428 41804
rect 29484 41636 29540 41646
rect 29484 41188 29540 41580
rect 29484 41122 29540 41132
rect 29820 40740 29876 41916
rect 29820 39508 29876 40684
rect 29820 39442 29876 39452
rect 30604 40516 30660 40526
rect 29372 38882 29428 38892
rect 30604 38668 30660 40460
rect 30604 38612 30772 38668
rect 29260 35634 29316 35644
rect 28588 33954 28644 33964
rect 26796 28018 26852 28028
rect 28140 31780 28196 31790
rect 26460 25666 26516 25676
rect 28140 25396 28196 31724
rect 30716 26180 30772 38612
rect 30716 25508 30772 26124
rect 30716 25442 30772 25452
rect 31948 32228 32004 48748
rect 33852 47908 33908 55020
rect 33964 51604 34020 56924
rect 33964 51538 34020 51548
rect 35168 60396 35488 61908
rect 39452 66836 39508 66846
rect 35168 60340 35196 60396
rect 35252 60340 35300 60396
rect 35356 60340 35404 60396
rect 35460 60340 35488 60396
rect 35168 58828 35488 60340
rect 39340 60452 39396 60462
rect 39340 59444 39396 60396
rect 39452 59668 39508 66780
rect 41244 66276 41300 66286
rect 41244 64148 41300 66220
rect 41244 64082 41300 64092
rect 40012 63476 40068 63486
rect 40012 62132 40068 63420
rect 40012 62066 40068 62076
rect 42140 61124 42196 67452
rect 50528 69020 50848 70532
rect 50528 68964 50556 69020
rect 50612 68964 50660 69020
rect 50716 68964 50764 69020
rect 50820 68964 50848 69020
rect 50528 67452 50848 68964
rect 50528 67396 50556 67452
rect 50612 67396 50660 67452
rect 50716 67396 50764 67452
rect 50820 67396 50848 67452
rect 50528 65884 50848 67396
rect 50528 65828 50556 65884
rect 50612 65828 50660 65884
rect 50716 65828 50764 65884
rect 50820 65828 50848 65884
rect 50528 64316 50848 65828
rect 50528 64260 50556 64316
rect 50612 64260 50660 64316
rect 50716 64260 50764 64316
rect 50820 64260 50848 64316
rect 44268 62916 44324 62926
rect 43260 62580 43316 62590
rect 42140 61058 42196 61068
rect 42588 61236 42644 61246
rect 39452 59602 39508 59612
rect 39340 59378 39396 59388
rect 35168 58772 35196 58828
rect 35252 58772 35300 58828
rect 35356 58772 35404 58828
rect 35460 58772 35488 58828
rect 42588 58884 42644 61180
rect 43260 58996 43316 62524
rect 43260 58930 43316 58940
rect 44268 58996 44324 62860
rect 44268 58930 44324 58940
rect 50528 62748 50848 64260
rect 50528 62692 50556 62748
rect 50612 62692 50660 62748
rect 50716 62692 50764 62748
rect 50820 62692 50848 62748
rect 50528 61180 50848 62692
rect 50528 61124 50556 61180
rect 50612 61124 50660 61180
rect 50716 61124 50764 61180
rect 50820 61124 50848 61180
rect 50528 59612 50848 61124
rect 50528 59556 50556 59612
rect 50612 59556 50660 59612
rect 50716 59556 50764 59612
rect 50820 59556 50848 59612
rect 42588 58818 42644 58828
rect 35168 57260 35488 58772
rect 45948 58660 46004 58670
rect 44940 58100 44996 58110
rect 44940 57876 44996 58044
rect 44940 57810 44996 57820
rect 35168 57204 35196 57260
rect 35252 57204 35300 57260
rect 35356 57204 35404 57260
rect 35460 57204 35488 57260
rect 35168 55692 35488 57204
rect 45500 56420 45556 56430
rect 35168 55636 35196 55692
rect 35252 55636 35300 55692
rect 35356 55636 35404 55692
rect 35460 55636 35488 55692
rect 35168 54124 35488 55636
rect 42700 56196 42756 56206
rect 41804 55076 41860 55086
rect 35168 54068 35196 54124
rect 35252 54068 35300 54124
rect 35356 54068 35404 54124
rect 35460 54068 35488 54124
rect 35168 52556 35488 54068
rect 35168 52500 35196 52556
rect 35252 52500 35300 52556
rect 35356 52500 35404 52556
rect 35460 52500 35488 52556
rect 33852 47842 33908 47852
rect 35168 50988 35488 52500
rect 39676 54516 39732 54526
rect 35168 50932 35196 50988
rect 35252 50932 35300 50988
rect 35356 50932 35404 50988
rect 35460 50932 35488 50988
rect 35168 49420 35488 50932
rect 35168 49364 35196 49420
rect 35252 49364 35300 49420
rect 35356 49364 35404 49420
rect 35460 49364 35488 49420
rect 35168 47852 35488 49364
rect 35168 47796 35196 47852
rect 35252 47796 35300 47852
rect 35356 47796 35404 47852
rect 35460 47796 35488 47852
rect 34636 47012 34692 47022
rect 33964 46004 34020 46014
rect 33628 41972 33684 41982
rect 33628 33684 33684 41916
rect 33852 41524 33908 41534
rect 33852 38052 33908 41468
rect 33852 37986 33908 37996
rect 33964 37940 34020 45948
rect 34524 44436 34580 44446
rect 34524 43204 34580 44380
rect 34524 43138 34580 43148
rect 34636 38276 34692 46956
rect 35168 46284 35488 47796
rect 38668 52164 38724 52174
rect 35168 46228 35196 46284
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35460 46228 35488 46284
rect 35168 44716 35488 46228
rect 35168 44660 35196 44716
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35460 44660 35488 44716
rect 34636 38210 34692 38220
rect 34748 44548 34804 44558
rect 33964 37874 34020 37884
rect 34748 35588 34804 44492
rect 35168 43148 35488 44660
rect 36876 47124 36932 47134
rect 36876 43428 36932 47068
rect 38668 44212 38724 52108
rect 39452 52052 39508 52062
rect 39452 51380 39508 51996
rect 39452 51314 39508 51324
rect 39676 51156 39732 54460
rect 41804 53060 41860 55020
rect 41804 52994 41860 53004
rect 42700 52948 42756 56140
rect 42700 52882 42756 52892
rect 39676 51090 39732 51100
rect 40012 51380 40068 51390
rect 40012 49812 40068 51324
rect 40012 49746 40068 49756
rect 45500 48468 45556 56364
rect 45948 50036 46004 58604
rect 45948 49970 46004 49980
rect 50528 58044 50848 59556
rect 50528 57988 50556 58044
rect 50612 57988 50660 58044
rect 50716 57988 50764 58044
rect 50820 57988 50848 58044
rect 50528 56476 50848 57988
rect 50528 56420 50556 56476
rect 50612 56420 50660 56476
rect 50716 56420 50764 56476
rect 50820 56420 50848 56476
rect 50528 54908 50848 56420
rect 50528 54852 50556 54908
rect 50612 54852 50660 54908
rect 50716 54852 50764 54908
rect 50820 54852 50848 54908
rect 50528 53340 50848 54852
rect 50528 53284 50556 53340
rect 50612 53284 50660 53340
rect 50716 53284 50764 53340
rect 50820 53284 50848 53340
rect 50528 51772 50848 53284
rect 50528 51716 50556 51772
rect 50612 51716 50660 51772
rect 50716 51716 50764 51772
rect 50820 51716 50848 51772
rect 50528 50204 50848 51716
rect 50528 50148 50556 50204
rect 50612 50148 50660 50204
rect 50716 50148 50764 50204
rect 50820 50148 50848 50204
rect 45500 48402 45556 48412
rect 50528 48636 50848 50148
rect 50528 48580 50556 48636
rect 50612 48580 50660 48636
rect 50716 48580 50764 48636
rect 50820 48580 50848 48636
rect 38668 44146 38724 44156
rect 50528 47068 50848 48580
rect 50528 47012 50556 47068
rect 50612 47012 50660 47068
rect 50716 47012 50764 47068
rect 50820 47012 50848 47068
rect 50528 45500 50848 47012
rect 50528 45444 50556 45500
rect 50612 45444 50660 45500
rect 50716 45444 50764 45500
rect 50820 45444 50848 45500
rect 36876 43362 36932 43372
rect 50528 43932 50848 45444
rect 50528 43876 50556 43932
rect 50612 43876 50660 43932
rect 50716 43876 50764 43932
rect 50820 43876 50848 43932
rect 35168 43092 35196 43148
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35460 43092 35488 43148
rect 35168 41580 35488 43092
rect 35168 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35488 41580
rect 34748 35522 34804 35532
rect 34972 40964 35028 40974
rect 33628 33618 33684 33628
rect 28140 25330 28196 25340
rect 31948 24612 32004 32172
rect 34748 27412 34804 27422
rect 31948 24546 32004 24556
rect 34188 25396 34244 25406
rect 34188 24612 34244 25340
rect 34748 24948 34804 27356
rect 34748 24882 34804 24892
rect 27804 23044 27860 23054
rect 27356 22820 27412 22830
rect 27356 13636 27412 22764
rect 27804 20580 27860 22988
rect 27804 20514 27860 20524
rect 33628 20356 33684 20366
rect 33628 18340 33684 20300
rect 33628 18274 33684 18284
rect 31948 15876 32004 15886
rect 31948 14868 32004 15820
rect 31948 14802 32004 14812
rect 27356 13570 27412 13580
rect 25116 4274 25172 4284
rect 34188 3444 34244 24556
rect 34972 21588 35028 40908
rect 34972 20692 35028 21532
rect 34972 20626 35028 20636
rect 35168 40012 35488 41524
rect 35168 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35488 40012
rect 35168 38444 35488 39956
rect 35168 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35488 38444
rect 35168 36876 35488 38388
rect 35168 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35488 36876
rect 35168 35308 35488 36820
rect 50528 42364 50848 43876
rect 50528 42308 50556 42364
rect 50612 42308 50660 42364
rect 50716 42308 50764 42364
rect 50820 42308 50848 42364
rect 50528 40796 50848 42308
rect 50528 40740 50556 40796
rect 50612 40740 50660 40796
rect 50716 40740 50764 40796
rect 50820 40740 50848 40796
rect 50528 39228 50848 40740
rect 50528 39172 50556 39228
rect 50612 39172 50660 39228
rect 50716 39172 50764 39228
rect 50820 39172 50848 39228
rect 50528 37660 50848 39172
rect 50528 37604 50556 37660
rect 50612 37604 50660 37660
rect 50716 37604 50764 37660
rect 50820 37604 50848 37660
rect 50528 36092 50848 37604
rect 50528 36036 50556 36092
rect 50612 36036 50660 36092
rect 50716 36036 50764 36092
rect 50820 36036 50848 36092
rect 35168 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35488 35308
rect 35168 33740 35488 35252
rect 46172 35588 46228 35598
rect 35168 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35488 33740
rect 35168 32172 35488 33684
rect 35168 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35488 32172
rect 35168 30604 35488 32116
rect 35168 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35488 30604
rect 35168 29036 35488 30548
rect 35756 34356 35812 34366
rect 35756 30548 35812 34300
rect 35756 30482 35812 30492
rect 36652 33460 36708 33470
rect 35168 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35488 29036
rect 35168 27468 35488 28980
rect 36652 27972 36708 33404
rect 39452 32004 39508 32014
rect 38892 31556 38948 31566
rect 38892 30212 38948 31500
rect 38892 30146 38948 30156
rect 39452 29204 39508 31948
rect 46172 30100 46228 35532
rect 50528 34524 50848 36036
rect 50528 34468 50556 34524
rect 50612 34468 50660 34524
rect 50716 34468 50764 34524
rect 50820 34468 50848 34524
rect 48412 34020 48468 34030
rect 46172 30034 46228 30044
rect 47628 30100 47684 30110
rect 47628 29764 47684 30044
rect 47628 29698 47684 29708
rect 39452 29138 39508 29148
rect 36652 27906 36708 27916
rect 35168 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35488 27468
rect 35168 25900 35488 27412
rect 48412 26404 48468 33964
rect 50528 32956 50848 34468
rect 50528 32900 50556 32956
rect 50612 32900 50660 32956
rect 50716 32900 50764 32956
rect 50820 32900 50848 32956
rect 48412 26338 48468 26348
rect 48524 32452 48580 32462
rect 35168 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35488 25900
rect 35168 24332 35488 25844
rect 35168 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35488 24332
rect 35168 22764 35488 24276
rect 35168 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35488 22764
rect 35168 21196 35488 22708
rect 35168 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35488 21196
rect 35168 19628 35488 21140
rect 35168 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35488 19628
rect 34524 18788 34580 18798
rect 34524 18228 34580 18732
rect 34524 18162 34580 18172
rect 34188 3378 34244 3388
rect 35168 18060 35488 19572
rect 36316 26292 36372 26302
rect 35168 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35488 18060
rect 35168 16492 35488 18004
rect 35168 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35488 16492
rect 35168 14924 35488 16436
rect 35168 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35488 14924
rect 35168 13356 35488 14868
rect 35644 18228 35700 18238
rect 35644 14420 35700 18172
rect 36092 17668 36148 17678
rect 36092 15876 36148 17612
rect 36092 15810 36148 15820
rect 36204 17444 36260 17454
rect 35644 14354 35700 14364
rect 35168 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35488 13356
rect 35168 11788 35488 13300
rect 36204 13076 36260 17388
rect 36204 13010 36260 13020
rect 35168 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35488 11788
rect 35168 10220 35488 11732
rect 35168 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35488 10220
rect 35168 8652 35488 10164
rect 35168 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35488 8652
rect 35168 7084 35488 8596
rect 35168 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35488 7084
rect 35168 5516 35488 7028
rect 35168 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35488 5516
rect 35168 3948 35488 5460
rect 35168 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35488 3948
rect 19808 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20128 3164
rect 19808 3076 20128 3108
rect 35168 3076 35488 3892
rect 36316 3444 36372 26236
rect 48524 26180 48580 32396
rect 48524 26114 48580 26124
rect 50528 31388 50848 32900
rect 50528 31332 50556 31388
rect 50612 31332 50660 31388
rect 50716 31332 50764 31388
rect 50820 31332 50848 31388
rect 50528 29820 50848 31332
rect 50528 29764 50556 29820
rect 50612 29764 50660 29820
rect 50716 29764 50764 29820
rect 50820 29764 50848 29820
rect 50528 28252 50848 29764
rect 50528 28196 50556 28252
rect 50612 28196 50660 28252
rect 50716 28196 50764 28252
rect 50820 28196 50848 28252
rect 50528 26684 50848 28196
rect 50528 26628 50556 26684
rect 50612 26628 50660 26684
rect 50716 26628 50764 26684
rect 50820 26628 50848 26684
rect 50528 25116 50848 26628
rect 36764 25060 36820 25070
rect 36764 23604 36820 25004
rect 36540 19012 36596 19022
rect 36540 16660 36596 18956
rect 36540 16594 36596 16604
rect 36764 13860 36820 23548
rect 50528 25060 50556 25116
rect 50612 25060 50660 25116
rect 50716 25060 50764 25116
rect 50820 25060 50848 25116
rect 50528 23548 50848 25060
rect 50528 23492 50556 23548
rect 50612 23492 50660 23548
rect 50716 23492 50764 23548
rect 50820 23492 50848 23548
rect 50528 21980 50848 23492
rect 50528 21924 50556 21980
rect 50612 21924 50660 21980
rect 50716 21924 50764 21980
rect 50820 21924 50848 21980
rect 50528 20412 50848 21924
rect 50528 20356 50556 20412
rect 50612 20356 50660 20412
rect 50716 20356 50764 20412
rect 50820 20356 50848 20412
rect 46396 19012 46452 19022
rect 43036 18004 43092 18014
rect 43036 14644 43092 17948
rect 46396 17780 46452 18956
rect 46396 17714 46452 17724
rect 50528 18844 50848 20356
rect 50528 18788 50556 18844
rect 50612 18788 50660 18844
rect 50716 18788 50764 18844
rect 50820 18788 50848 18844
rect 43036 14578 43092 14588
rect 50528 17276 50848 18788
rect 50528 17220 50556 17276
rect 50612 17220 50660 17276
rect 50716 17220 50764 17276
rect 50820 17220 50848 17276
rect 50528 15708 50848 17220
rect 50528 15652 50556 15708
rect 50612 15652 50660 15708
rect 50716 15652 50764 15708
rect 50820 15652 50848 15708
rect 36764 13794 36820 13804
rect 50528 14140 50848 15652
rect 50528 14084 50556 14140
rect 50612 14084 50660 14140
rect 50716 14084 50764 14140
rect 50820 14084 50848 14140
rect 36316 3378 36372 3388
rect 50528 12572 50848 14084
rect 50528 12516 50556 12572
rect 50612 12516 50660 12572
rect 50716 12516 50764 12572
rect 50820 12516 50848 12572
rect 50528 11004 50848 12516
rect 50528 10948 50556 11004
rect 50612 10948 50660 11004
rect 50716 10948 50764 11004
rect 50820 10948 50848 11004
rect 50528 9436 50848 10948
rect 50528 9380 50556 9436
rect 50612 9380 50660 9436
rect 50716 9380 50764 9436
rect 50820 9380 50848 9436
rect 50528 7868 50848 9380
rect 50528 7812 50556 7868
rect 50612 7812 50660 7868
rect 50716 7812 50764 7868
rect 50820 7812 50848 7868
rect 50528 6300 50848 7812
rect 50528 6244 50556 6300
rect 50612 6244 50660 6300
rect 50716 6244 50764 6300
rect 50820 6244 50848 6300
rect 50528 4732 50848 6244
rect 50528 4676 50556 4732
rect 50612 4676 50660 4732
rect 50716 4676 50764 4732
rect 50820 4676 50848 4732
rect 50528 3164 50848 4676
rect 50528 3108 50556 3164
rect 50612 3108 50660 3164
rect 50716 3108 50764 3164
rect 50820 3108 50848 3164
rect 50528 3076 50848 3108
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _1440_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 17584 0 1 42336
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1441_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 22288 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1442_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 23184 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1443_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 15344 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1444_
timestamp 1698431365
transform -1 0 16912 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1445_
timestamp 1698431365
transform -1 0 23632 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1446_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 24192 0 -1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1447_
timestamp 1698431365
transform 1 0 29680 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1448_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 31136 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1449_
timestamp 1698431365
transform 1 0 11760 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1450_
timestamp 1698431365
transform -1 0 14224 0 1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1451_
timestamp 1698431365
transform 1 0 11312 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1452_
timestamp 1698431365
transform 1 0 9632 0 -1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1453_
timestamp 1698431365
transform -1 0 19600 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _1454_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 11424 0 1 40768
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _1455_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 11424 0 1 40768
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _1456_
timestamp 1698431365
transform 1 0 10192 0 -1 42336
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1457_
timestamp 1698431365
transform -1 0 10640 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _1458_
timestamp 1698431365
transform -1 0 10528 0 1 42336
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1459_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 10528 0 1 42336
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1460_
timestamp 1698431365
transform 1 0 11536 0 -1 43904
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1461_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 12432 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1462_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 12656 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1463_
timestamp 1698431365
transform -1 0 21616 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1464_
timestamp 1698431365
transform -1 0 19376 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _1465_
timestamp 1698431365
transform 1 0 15232 0 1 31360
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  _1466_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 19264 0 -1 36064
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1467_
timestamp 1698431365
transform 1 0 16352 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1468_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 18256 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1469_
timestamp 1698431365
transform 1 0 21728 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1470_
timestamp 1698431365
transform 1 0 24192 0 -1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1471_
timestamp 1698431365
transform 1 0 25312 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1472_
timestamp 1698431365
transform 1 0 33488 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1473_
timestamp 1698431365
transform -1 0 21392 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1474_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 18256 0 -1 37632
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1475_
timestamp 1698431365
transform 1 0 19264 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1476_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 24864 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1477_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 20048 0 -1 39200
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1478_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 23184 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1479_
timestamp 1698431365
transform -1 0 23184 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1480_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 20048 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1481_
timestamp 1698431365
transform 1 0 21616 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1482_
timestamp 1698431365
transform 1 0 12096 0 -1 43904
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1483_
timestamp 1698431365
transform 1 0 12208 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1484_
timestamp 1698431365
transform 1 0 19824 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1485_
timestamp 1698431365
transform -1 0 20048 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1486_
timestamp 1698431365
transform 1 0 18704 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1487_
timestamp 1698431365
transform 1 0 17472 0 -1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1488_
timestamp 1698431365
transform -1 0 18928 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1489_
timestamp 1698431365
transform 1 0 14336 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1490_
timestamp 1698431365
transform -1 0 17808 0 -1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1491_
timestamp 1698431365
transform -1 0 16800 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1492_
timestamp 1698431365
transform -1 0 20160 0 1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1493_
timestamp 1698431365
transform 1 0 14784 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1494_
timestamp 1698431365
transform -1 0 17024 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1495_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 15680 0 -1 29792
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1496_
timestamp 1698431365
transform -1 0 20944 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1497_
timestamp 1698431365
transform -1 0 16912 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1498_
timestamp 1698431365
transform -1 0 14336 0 1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1499_
timestamp 1698431365
transform 1 0 14560 0 -1 32928
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1500_
timestamp 1698431365
transform -1 0 16464 0 -1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1501_
timestamp 1698431365
transform -1 0 15904 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1502_
timestamp 1698431365
transform -1 0 15344 0 1 32928
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1503_
timestamp 1698431365
transform 1 0 16576 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1504_
timestamp 1698431365
transform 1 0 23408 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1505_
timestamp 1698431365
transform 1 0 23968 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1506_
timestamp 1698431365
transform 1 0 18256 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1507_
timestamp 1698431365
transform 1 0 17136 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1508_
timestamp 1698431365
transform 1 0 16576 0 1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1509_
timestamp 1698431365
transform -1 0 15904 0 1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1510_
timestamp 1698431365
transform 1 0 13104 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1511_
timestamp 1698431365
transform 1 0 19600 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1512_
timestamp 1698431365
transform 1 0 23408 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1513_
timestamp 1698431365
transform 1 0 25872 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1514_
timestamp 1698431365
transform -1 0 24304 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1515_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 22512 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1516_
timestamp 1698431365
transform 1 0 15904 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai222_2  _1517_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 17248 0 1 26656
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1518_
timestamp 1698431365
transform -1 0 18592 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai222_2  _1519_
timestamp 1698431365
transform 1 0 17248 0 -1 26656
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1520_
timestamp 1698431365
transform -1 0 17248 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1521_
timestamp 1698431365
transform 1 0 19152 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai222_2  _1522_
timestamp 1698431365
transform 1 0 20272 0 -1 26656
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1523_
timestamp 1698431365
transform 1 0 17920 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1524_
timestamp 1698431365
transform 1 0 22512 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1525_
timestamp 1698431365
transform 1 0 15120 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1526_
timestamp 1698431365
transform 1 0 20496 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1527_
timestamp 1698431365
transform -1 0 21616 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai222_2  _1528_
timestamp 1698431365
transform 1 0 21168 0 -1 12544
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1529_
timestamp 1698431365
transform -1 0 21616 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1530_
timestamp 1698431365
transform 1 0 23184 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai222_2  _1531_
timestamp 1698431365
transform -1 0 20944 0 1 10976
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1532_
timestamp 1698431365
transform -1 0 23184 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai222_2  _1533_
timestamp 1698431365
transform 1 0 23184 0 1 12544
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1534_
timestamp 1698431365
transform -1 0 24752 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1535_
timestamp 1698431365
transform 1 0 32704 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1536_
timestamp 1698431365
transform -1 0 32704 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai222_2  _1537_
timestamp 1698431365
transform 1 0 25200 0 -1 9408
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1538_
timestamp 1698431365
transform -1 0 26768 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1539_
timestamp 1698431365
transform 1 0 30128 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1540_
timestamp 1698431365
transform 1 0 30128 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai222_2  _1541_
timestamp 1698431365
transform 1 0 27104 0 -1 12544
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1542_
timestamp 1698431365
transform -1 0 28336 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1543_
timestamp 1698431365
transform -1 0 34272 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai222_2  _1544_
timestamp 1698431365
transform 1 0 29232 0 1 10976
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1545_
timestamp 1698431365
transform -1 0 32704 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai222_2  _1546_
timestamp 1698431365
transform 1 0 29904 0 1 9408
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1547_
timestamp 1698431365
transform -1 0 31808 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1548_
timestamp 1698431365
transform 1 0 34608 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai222_2  _1549_
timestamp 1698431365
transform 1 0 32928 0 -1 10976
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1550_
timestamp 1698431365
transform -1 0 34272 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1551_
timestamp 1698431365
transform -1 0 36624 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1552_
timestamp 1698431365
transform -1 0 39200 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai222_2  _1553_
timestamp 1698431365
transform -1 0 38976 0 -1 10976
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1554_
timestamp 1698431365
transform -1 0 34944 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1555_
timestamp 1698431365
transform 1 0 36848 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai222_2  _1556_
timestamp 1698431365
transform -1 0 38528 0 -1 12544
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1557_
timestamp 1698431365
transform 1 0 36176 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai222_2  _1558_
timestamp 1698431365
transform -1 0 39872 0 1 10976
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1559_
timestamp 1698431365
transform -1 0 39872 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1560_
timestamp 1698431365
transform 1 0 42448 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai222_2  _1561_
timestamp 1698431365
transform 1 0 40768 0 1 10976
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1562_
timestamp 1698431365
transform -1 0 40544 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1563_
timestamp 1698431365
transform -1 0 44688 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1564_
timestamp 1698431365
transform 1 0 40768 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai222_2  _1565_
timestamp 1698431365
transform 1 0 41440 0 1 7840
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1566_
timestamp 1698431365
transform -1 0 42560 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1567_
timestamp 1698431365
transform 1 0 27328 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1568_
timestamp 1698431365
transform 1 0 42112 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai222_2  _1569_
timestamp 1698431365
transform 1 0 42448 0 -1 7840
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1570_
timestamp 1698431365
transform 1 0 42000 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai222_2  _1571_
timestamp 1698431365
transform 1 0 42784 0 -1 6272
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1572_
timestamp 1698431365
transform -1 0 46256 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1573_
timestamp 1698431365
transform 1 0 42672 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai222_2  _1574_
timestamp 1698431365
transform 1 0 44688 0 -1 12544
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1575_
timestamp 1698431365
transform 1 0 45360 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1576_
timestamp 1698431365
transform -1 0 47040 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1577_
timestamp 1698431365
transform 1 0 20496 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1578_
timestamp 1698431365
transform 1 0 42448 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai222_2  _1579_
timestamp 1698431365
transform 1 0 42784 0 -1 20384
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1580_
timestamp 1698431365
transform -1 0 44352 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1581_
timestamp 1698431365
transform 1 0 42448 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai222_2  _1582_
timestamp 1698431365
transform -1 0 46816 0 -1 23520
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1583_
timestamp 1698431365
transform 1 0 43344 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai222_2  _1584_
timestamp 1698431365
transform -1 0 45808 0 -1 26656
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1585_
timestamp 1698431365
transform 1 0 44688 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1586_
timestamp 1698431365
transform -1 0 19600 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1587_
timestamp 1698431365
transform 1 0 39088 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai222_2  _1588_
timestamp 1698431365
transform -1 0 43792 0 -1 25088
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1589_
timestamp 1698431365
transform -1 0 43792 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1590_
timestamp 1698431365
transform 1 0 41552 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1591_
timestamp 1698431365
transform 1 0 40656 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai222_2  _1592_
timestamp 1698431365
transform 1 0 40768 0 -1 23520
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1593_
timestamp 1698431365
transform -1 0 44240 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1594_
timestamp 1698431365
transform -1 0 36624 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai222_2  _1595_
timestamp 1698431365
transform 1 0 37408 0 1 20384
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1596_
timestamp 1698431365
transform -1 0 40432 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai222_2  _1597_
timestamp 1698431365
transform 1 0 36960 0 -1 21952
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1598_
timestamp 1698431365
transform 1 0 37184 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1599_
timestamp 1698431365
transform -1 0 37744 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai222_2  _1600_
timestamp 1698431365
transform -1 0 36624 0 -1 26656
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1601_
timestamp 1698431365
transform -1 0 37072 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1602_
timestamp 1698431365
transform 1 0 34608 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1603_
timestamp 1698431365
transform -1 0 24864 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai222_2  _1604_
timestamp 1698431365
transform 1 0 31584 0 1 25088
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1605_
timestamp 1698431365
transform -1 0 33600 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1606_
timestamp 1698431365
transform -1 0 27328 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai222_2  _1607_
timestamp 1698431365
transform 1 0 30128 0 1 21952
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1608_
timestamp 1698431365
transform 1 0 30800 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai222_2  _1609_
timestamp 1698431365
transform 1 0 29232 0 1 20384
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1610_
timestamp 1698431365
transform 1 0 29008 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1611_
timestamp 1698431365
transform -1 0 24528 0 1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1612_
timestamp 1698431365
transform 1 0 20496 0 -1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1613_
timestamp 1698431365
transform -1 0 21840 0 1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1614_
timestamp 1698431365
transform -1 0 20160 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1615_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 20384 0 1 43904
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1616_
timestamp 1698431365
transform -1 0 20944 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1617_
timestamp 1698431365
transform 1 0 21168 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1618_
timestamp 1698431365
transform 1 0 18144 0 -1 62720
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1619_
timestamp 1698431365
transform -1 0 22848 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1620_
timestamp 1698431365
transform 1 0 30016 0 -1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1621_
timestamp 1698431365
transform -1 0 32480 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1622_
timestamp 1698431365
transform -1 0 19264 0 -1 45472
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1623_
timestamp 1698431365
transform 1 0 18928 0 -1 59584
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1624_
timestamp 1698431365
transform 1 0 20272 0 1 59584
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1625_
timestamp 1698431365
transform 1 0 18144 0 1 51744
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1626_
timestamp 1698431365
transform 1 0 19376 0 -1 51744
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1627_
timestamp 1698431365
transform -1 0 20384 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1628_
timestamp 1698431365
transform -1 0 20608 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1629_
timestamp 1698431365
transform -1 0 20832 0 1 54880
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1630_
timestamp 1698431365
transform -1 0 19488 0 1 51744
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1631_
timestamp 1698431365
transform -1 0 22064 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1632_
timestamp 1698431365
transform -1 0 20832 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1633_
timestamp 1698431365
transform 1 0 23744 0 1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1634_
timestamp 1698431365
transform -1 0 22400 0 1 59584
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1635_
timestamp 1698431365
transform -1 0 20160 0 1 54880
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1636_
timestamp 1698431365
transform 1 0 20272 0 -1 61152
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1637_
timestamp 1698431365
transform 1 0 19376 0 -1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1638_
timestamp 1698431365
transform -1 0 19152 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1639_
timestamp 1698431365
transform 1 0 19712 0 1 65856
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1640_
timestamp 1698431365
transform 1 0 20048 0 -1 64288
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1641_
timestamp 1698431365
transform 1 0 21168 0 -1 61152
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1642_
timestamp 1698431365
transform 1 0 19600 0 1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1643_
timestamp 1698431365
transform -1 0 19600 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1644_
timestamp 1698431365
transform 1 0 23296 0 1 67424
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1645_
timestamp 1698431365
transform -1 0 23744 0 -1 65856
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1646_
timestamp 1698431365
transform 1 0 22624 0 1 67424
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1647_
timestamp 1698431365
transform 1 0 21168 0 1 64288
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1648_
timestamp 1698431365
transform 1 0 21616 0 1 65856
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1649_
timestamp 1698431365
transform 1 0 21616 0 -1 67424
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1650_
timestamp 1698431365
transform -1 0 21616 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1651_
timestamp 1698431365
transform -1 0 21616 0 -1 67424
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1652_
timestamp 1698431365
transform -1 0 23296 0 -1 67424
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1653_
timestamp 1698431365
transform 1 0 21728 0 1 67424
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1654_
timestamp 1698431365
transform 1 0 21168 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1655_
timestamp 1698431365
transform 1 0 30128 0 1 65856
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1656_
timestamp 1698431365
transform -1 0 30240 0 -1 67424
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1657_
timestamp 1698431365
transform -1 0 24528 0 -1 67424
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1658_
timestamp 1698431365
transform 1 0 23184 0 -1 68992
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1659_
timestamp 1698431365
transform -1 0 24864 0 -1 68992
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1660_
timestamp 1698431365
transform -1 0 24192 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1661_
timestamp 1698431365
transform 1 0 20048 0 -1 67424
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1662_
timestamp 1698431365
transform 1 0 25984 0 1 67424
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1663_
timestamp 1698431365
transform -1 0 25088 0 1 67424
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1664_
timestamp 1698431365
transform -1 0 25984 0 1 67424
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1665_
timestamp 1698431365
transform 1 0 25648 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1666_
timestamp 1698431365
transform 1 0 28112 0 1 67424
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1667_
timestamp 1698431365
transform -1 0 33600 0 1 67424
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1668_
timestamp 1698431365
transform -1 0 31808 0 -1 67424
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1669_
timestamp 1698431365
transform 1 0 29008 0 -1 67424
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1670_
timestamp 1698431365
transform 1 0 30464 0 1 68992
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1671_
timestamp 1698431365
transform 1 0 30240 0 -1 67424
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1672_
timestamp 1698431365
transform -1 0 31360 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1673_
timestamp 1698431365
transform -1 0 29568 0 1 68992
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1674_
timestamp 1698431365
transform -1 0 32032 0 1 68992
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1675_
timestamp 1698431365
transform 1 0 29568 0 1 68992
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1676_
timestamp 1698431365
transform -1 0 29456 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1677_
timestamp 1698431365
transform -1 0 34944 0 -1 68992
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1678_
timestamp 1698431365
transform 1 0 30800 0 1 65856
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1679_
timestamp 1698431365
transform 1 0 32928 0 -1 68992
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1680_
timestamp 1698431365
transform 1 0 32704 0 1 68992
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1681_
timestamp 1698431365
transform -1 0 32704 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1682_
timestamp 1698431365
transform 1 0 26208 0 -1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1683_
timestamp 1698431365
transform 1 0 35728 0 1 67424
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1684_
timestamp 1698431365
transform 1 0 35392 0 1 68992
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1685_
timestamp 1698431365
transform -1 0 35392 0 1 68992
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1686_
timestamp 1698431365
transform -1 0 34608 0 1 68992
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1687_
timestamp 1698431365
transform -1 0 35056 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1688_
timestamp 1698431365
transform 1 0 33376 0 1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1689_
timestamp 1698431365
transform -1 0 38976 0 1 67424
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1690_
timestamp 1698431365
transform 1 0 38304 0 -1 68992
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1691_
timestamp 1698431365
transform 1 0 35504 0 -1 68992
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1692_
timestamp 1698431365
transform 1 0 36176 0 -1 68992
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1693_
timestamp 1698431365
transform 1 0 36736 0 -1 68992
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1694_
timestamp 1698431365
transform -1 0 37856 0 1 68992
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1695_
timestamp 1698431365
transform 1 0 36176 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1696_
timestamp 1698431365
transform -1 0 37744 0 1 67424
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1697_
timestamp 1698431365
transform 1 0 37520 0 -1 68992
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1698_
timestamp 1698431365
transform -1 0 38752 0 1 68992
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1699_
timestamp 1698431365
transform -1 0 40544 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1700_
timestamp 1698431365
transform 1 0 40992 0 -1 67424
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1701_
timestamp 1698431365
transform 1 0 38976 0 -1 68992
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1702_
timestamp 1698431365
transform 1 0 39760 0 -1 68992
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1703_
timestamp 1698431365
transform -1 0 40544 0 -1 70560
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1704_
timestamp 1698431365
transform 1 0 40768 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1705_
timestamp 1698431365
transform -1 0 42336 0 -1 67424
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1706_
timestamp 1698431365
transform -1 0 41440 0 1 65856
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1707_
timestamp 1698431365
transform -1 0 41216 0 1 67424
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1708_
timestamp 1698431365
transform -1 0 41664 0 -1 68992
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1709_
timestamp 1698431365
transform 1 0 39088 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1710_
timestamp 1698431365
transform 1 0 42784 0 1 68992
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1711_
timestamp 1698431365
transform -1 0 48048 0 -1 65856
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1712_
timestamp 1698431365
transform 1 0 29008 0 1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1713_
timestamp 1698431365
transform 1 0 42448 0 1 58016
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1714_
timestamp 1698431365
transform 1 0 41440 0 1 65856
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1715_
timestamp 1698431365
transform 1 0 42672 0 1 65856
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1716_
timestamp 1698431365
transform -1 0 44912 0 -1 67424
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1717_
timestamp 1698431365
transform 1 0 45136 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1718_
timestamp 1698431365
transform -1 0 44128 0 -1 65856
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1719_
timestamp 1698431365
transform -1 0 43120 0 -1 67424
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1720_
timestamp 1698431365
transform -1 0 45808 0 -1 67424
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1721_
timestamp 1698431365
transform 1 0 45136 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1722_
timestamp 1698431365
transform 1 0 42000 0 1 65856
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1723_
timestamp 1698431365
transform -1 0 44688 0 -1 65856
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1724_
timestamp 1698431365
transform -1 0 44240 0 1 65856
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1725_
timestamp 1698431365
transform 1 0 43120 0 -1 67424
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1726_
timestamp 1698431365
transform -1 0 43904 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1727_
timestamp 1698431365
transform 1 0 43120 0 -1 62720
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1728_
timestamp 1698431365
transform -1 0 44352 0 -1 62720
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1729_
timestamp 1698431365
transform 1 0 43680 0 1 62720
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1730_
timestamp 1698431365
transform -1 0 45584 0 1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1731_
timestamp 1698431365
transform -1 0 44240 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1732_
timestamp 1698431365
transform -1 0 43568 0 1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1733_
timestamp 1698431365
transform -1 0 48496 0 1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1734_
timestamp 1698431365
transform 1 0 41328 0 1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1735_
timestamp 1698431365
transform -1 0 45696 0 -1 56448
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1736_
timestamp 1698431365
transform -1 0 45136 0 -1 56448
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1737_
timestamp 1698431365
transform 1 0 43568 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1738_
timestamp 1698431365
transform 1 0 45696 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1739_
timestamp 1698431365
transform -1 0 44240 0 1 56448
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1740_
timestamp 1698431365
transform 1 0 43568 0 -1 56448
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1741_
timestamp 1698431365
transform 1 0 43568 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1742_
timestamp 1698431365
transform 1 0 44688 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1743_
timestamp 1698431365
transform 1 0 32928 0 -1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1744_
timestamp 1698431365
transform -1 0 43568 0 1 53312
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1745_
timestamp 1698431365
transform -1 0 43344 0 -1 56448
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1746_
timestamp 1698431365
transform 1 0 42000 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1747_
timestamp 1698431365
transform 1 0 40880 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1748_
timestamp 1698431365
transform -1 0 40992 0 1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1749_
timestamp 1698431365
transform 1 0 41552 0 1 53312
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1750_
timestamp 1698431365
transform 1 0 42224 0 -1 53312
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1751_
timestamp 1698431365
transform 1 0 42112 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1752_
timestamp 1698431365
transform 1 0 43008 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1753_
timestamp 1698431365
transform 1 0 34272 0 -1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1754_
timestamp 1698431365
transform -1 0 36960 0 -1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1755_
timestamp 1698431365
transform -1 0 35840 0 1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1756_
timestamp 1698431365
transform -1 0 41552 0 1 53312
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1757_
timestamp 1698431365
transform -1 0 37184 0 -1 53312
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1758_
timestamp 1698431365
transform 1 0 35616 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1759_
timestamp 1698431365
transform -1 0 35056 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1760_
timestamp 1698431365
transform 1 0 37744 0 1 53312
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1761_
timestamp 1698431365
transform -1 0 36624 0 1 54880
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1762_
timestamp 1698431365
transform -1 0 37744 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1763_
timestamp 1698431365
transform 1 0 37296 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1764_
timestamp 1698431365
transform -1 0 32368 0 -1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1765_
timestamp 1698431365
transform -1 0 37744 0 -1 53312
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1766_
timestamp 1698431365
transform -1 0 35728 0 -1 54880
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1767_
timestamp 1698431365
transform -1 0 36624 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1768_
timestamp 1698431365
transform 1 0 36848 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1769_
timestamp 1698431365
transform 1 0 25536 0 -1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1770_
timestamp 1698431365
transform -1 0 34832 0 -1 53312
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1771_
timestamp 1698431365
transform 1 0 34832 0 -1 53312
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1772_
timestamp 1698431365
transform 1 0 34720 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1773_
timestamp 1698431365
transform 1 0 33152 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1774_
timestamp 1698431365
transform 1 0 19712 0 1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1775_
timestamp 1698431365
transform -1 0 31472 0 1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1776_
timestamp 1698431365
transform -1 0 30016 0 -1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1777_
timestamp 1698431365
transform -1 0 32928 0 1 51744
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1778_
timestamp 1698431365
transform -1 0 31472 0 -1 53312
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1779_
timestamp 1698431365
transform 1 0 29792 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1780_
timestamp 1698431365
transform -1 0 30240 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1781_
timestamp 1698431365
transform -1 0 31248 0 1 51744
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1782_
timestamp 1698431365
transform -1 0 30688 0 -1 53312
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1783_
timestamp 1698431365
transform 1 0 28672 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1784_
timestamp 1698431365
transform -1 0 28784 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1785_
timestamp 1698431365
transform 1 0 30688 0 -1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1786_
timestamp 1698431365
transform -1 0 28672 0 -1 53312
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1787_
timestamp 1698431365
transform 1 0 29008 0 1 51744
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1788_
timestamp 1698431365
transform 1 0 27104 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1789_
timestamp 1698431365
transform 1 0 25088 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1790_
timestamp 1698431365
transform -1 0 17024 0 -1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1791_
timestamp 1698431365
transform 1 0 26992 0 1 53312
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1792_
timestamp 1698431365
transform 1 0 27664 0 1 53312
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1793_
timestamp 1698431365
transform 1 0 26208 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1794_
timestamp 1698431365
transform -1 0 25536 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1795_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 18704 0 -1 45472
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1796_
timestamp 1698431365
transform -1 0 18256 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1797_
timestamp 1698431365
transform 1 0 11984 0 1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1798_
timestamp 1698431365
transform 1 0 13440 0 -1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1799_
timestamp 1698431365
transform 1 0 15568 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1800_
timestamp 1698431365
transform -1 0 14672 0 1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1801_
timestamp 1698431365
transform -1 0 16912 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1802_
timestamp 1698431365
transform 1 0 26096 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1803_
timestamp 1698431365
transform 1 0 25984 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1804_
timestamp 1698431365
transform -1 0 17024 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1805_
timestamp 1698431365
transform 1 0 15568 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1806_
timestamp 1698431365
transform 1 0 28448 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1807_
timestamp 1698431365
transform 1 0 29456 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1808_
timestamp 1698431365
transform 1 0 31248 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1809_
timestamp 1698431365
transform -1 0 32144 0 1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1810_
timestamp 1698431365
transform 1 0 26768 0 1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1811_
timestamp 1698431365
transform 1 0 25648 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1812_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 22064 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1813_
timestamp 1698431365
transform 1 0 31360 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1814_
timestamp 1698431365
transform 1 0 31808 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1815_
timestamp 1698431365
transform 1 0 30128 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1816_
timestamp 1698431365
transform -1 0 27888 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _1817_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 23184 0 -1 31360
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1818_
timestamp 1698431365
transform -1 0 23184 0 -1 32928
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1819_
timestamp 1698431365
transform -1 0 22176 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1820_
timestamp 1698431365
transform 1 0 26880 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1821_
timestamp 1698431365
transform 1 0 22176 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1822_
timestamp 1698431365
transform -1 0 22960 0 1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1823_
timestamp 1698431365
transform 1 0 21168 0 1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1824_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 20944 0 -1 36064
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1825_
timestamp 1698431365
transform 1 0 27328 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1826_
timestamp 1698431365
transform 1 0 22288 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1827_
timestamp 1698431365
transform 1 0 21504 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1828_
timestamp 1698431365
transform -1 0 20944 0 1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1829_
timestamp 1698431365
transform 1 0 27888 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1830_
timestamp 1698431365
transform 1 0 29456 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1831_
timestamp 1698431365
transform 1 0 30912 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1832_
timestamp 1698431365
transform 1 0 21392 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1833_
timestamp 1698431365
transform -1 0 28112 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1834_
timestamp 1698431365
transform 1 0 24976 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1835_
timestamp 1698431365
transform -1 0 23632 0 1 28224
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1836_
timestamp 1698431365
transform 1 0 21168 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1837_
timestamp 1698431365
transform -1 0 24416 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1838_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 23296 0 1 26656
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1839_
timestamp 1698431365
transform 1 0 23072 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1840_
timestamp 1698431365
transform -1 0 21840 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1841_
timestamp 1698431365
transform -1 0 24752 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1842_
timestamp 1698431365
transform 1 0 25088 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1843_
timestamp 1698431365
transform 1 0 22176 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1844_
timestamp 1698431365
transform 1 0 33264 0 1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1845_
timestamp 1698431365
transform 1 0 33600 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1846_
timestamp 1698431365
transform -1 0 25872 0 -1 26656
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1847_
timestamp 1698431365
transform -1 0 31584 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1848_
timestamp 1698431365
transform -1 0 25648 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1849_
timestamp 1698431365
transform 1 0 22064 0 1 23520
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1850_
timestamp 1698431365
transform -1 0 24192 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1851_
timestamp 1698431365
transform 1 0 24192 0 1 26656
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1852_
timestamp 1698431365
transform -1 0 24864 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1853_
timestamp 1698431365
transform -1 0 20944 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1854_
timestamp 1698431365
transform -1 0 24192 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1855_
timestamp 1698431365
transform -1 0 25088 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1856_
timestamp 1698431365
transform 1 0 22960 0 -1 18816
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1857_
timestamp 1698431365
transform 1 0 22064 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1858_
timestamp 1698431365
transform 1 0 26320 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1859_
timestamp 1698431365
transform 1 0 26992 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1860_
timestamp 1698431365
transform -1 0 24304 0 1 18816
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1861_
timestamp 1698431365
transform -1 0 22624 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1862_
timestamp 1698431365
transform -1 0 26320 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1863_
timestamp 1698431365
transform -1 0 24864 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1864_
timestamp 1698431365
transform 1 0 22624 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1865_
timestamp 1698431365
transform 1 0 23408 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1866_
timestamp 1698431365
transform 1 0 22512 0 -1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1867_
timestamp 1698431365
transform -1 0 24640 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1868_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 25088 0 1 15680
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1869_
timestamp 1698431365
transform 1 0 28112 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1870_
timestamp 1698431365
transform -1 0 26768 0 1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1871_
timestamp 1698431365
transform -1 0 26544 0 -1 14112
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1872_
timestamp 1698431365
transform -1 0 23968 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1873_
timestamp 1698431365
transform 1 0 23968 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1874_
timestamp 1698431365
transform -1 0 25648 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1875_
timestamp 1698431365
transform 1 0 23968 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1876_
timestamp 1698431365
transform -1 0 27440 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1877_
timestamp 1698431365
transform -1 0 25872 0 -1 12544
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1878_
timestamp 1698431365
transform -1 0 26768 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1879_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 26320 0 1 14112
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1880_
timestamp 1698431365
transform 1 0 28448 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1881_
timestamp 1698431365
transform -1 0 29568 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1882_
timestamp 1698431365
transform -1 0 28000 0 -1 15680
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1883_
timestamp 1698431365
transform -1 0 26656 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1884_
timestamp 1698431365
transform 1 0 33152 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1885_
timestamp 1698431365
transform -1 0 33600 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1886_
timestamp 1698431365
transform 1 0 27552 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1887_
timestamp 1698431365
transform 1 0 25088 0 -1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1888_
timestamp 1698431365
transform -1 0 26656 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1889_
timestamp 1698431365
transform -1 0 34496 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1890_
timestamp 1698431365
transform -1 0 28784 0 -1 15680
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1891_
timestamp 1698431365
transform 1 0 26656 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1892_
timestamp 1698431365
transform 1 0 25872 0 -1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1893_
timestamp 1698431365
transform -1 0 26432 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1894_
timestamp 1698431365
transform 1 0 26768 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1895_
timestamp 1698431365
transform -1 0 27664 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1896_
timestamp 1698431365
transform 1 0 25872 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1897_
timestamp 1698431365
transform -1 0 25648 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1898_
timestamp 1698431365
transform -1 0 25872 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1899_
timestamp 1698431365
transform 1 0 31808 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1900_
timestamp 1698431365
transform 1 0 29680 0 1 17248
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1901_
timestamp 1698431365
transform 1 0 29232 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1902_
timestamp 1698431365
transform -1 0 32704 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1903_
timestamp 1698431365
transform 1 0 31024 0 1 17248
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1904_
timestamp 1698431365
transform -1 0 31696 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1905_
timestamp 1698431365
transform 1 0 32032 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1906_
timestamp 1698431365
transform -1 0 33376 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1907_
timestamp 1698431365
transform -1 0 31696 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1908_
timestamp 1698431365
transform 1 0 30128 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1909_
timestamp 1698431365
transform 1 0 30464 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1910_
timestamp 1698431365
transform 1 0 29680 0 -1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1911_
timestamp 1698431365
transform 1 0 31808 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1912_
timestamp 1698431365
transform -1 0 31920 0 -1 15680
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1913_
timestamp 1698431365
transform -1 0 31584 0 -1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1914_
timestamp 1698431365
transform -1 0 31920 0 1 12544
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1915_
timestamp 1698431365
transform -1 0 30128 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1916_
timestamp 1698431365
transform -1 0 31024 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1917_
timestamp 1698431365
transform 1 0 32032 0 -1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1918_
timestamp 1698431365
transform 1 0 32928 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1919_
timestamp 1698431365
transform 1 0 31920 0 1 12544
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1920_
timestamp 1698431365
transform -1 0 32592 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1921_
timestamp 1698431365
transform -1 0 32480 0 1 14112
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1922_
timestamp 1698431365
transform 1 0 35056 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1923_
timestamp 1698431365
transform -1 0 35392 0 -1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1924_
timestamp 1698431365
transform -1 0 34832 0 -1 14112
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1925_
timestamp 1698431365
transform 1 0 33040 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1926_
timestamp 1698431365
transform -1 0 35616 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1927_
timestamp 1698431365
transform -1 0 35504 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1928_
timestamp 1698431365
transform 1 0 33824 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1929_
timestamp 1698431365
transform -1 0 37632 0 1 14112
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1930_
timestamp 1698431365
transform 1 0 35616 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1931_
timestamp 1698431365
transform 1 0 35056 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1932_
timestamp 1698431365
transform -1 0 36288 0 1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1933_
timestamp 1698431365
transform 1 0 34496 0 1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1934_
timestamp 1698431365
transform 1 0 35952 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1935_
timestamp 1698431365
transform 1 0 34608 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1936_
timestamp 1698431365
transform -1 0 35168 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1937_
timestamp 1698431365
transform -1 0 35280 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1938_
timestamp 1698431365
transform 1 0 39536 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1939_
timestamp 1698431365
transform 1 0 34048 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1940_
timestamp 1698431365
transform 1 0 33824 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1941_
timestamp 1698431365
transform 1 0 33488 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1942_
timestamp 1698431365
transform 1 0 27328 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1943_
timestamp 1698431365
transform -1 0 38976 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1944_
timestamp 1698431365
transform -1 0 38192 0 -1 17248
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1945_
timestamp 1698431365
transform 1 0 35728 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1946_
timestamp 1698431365
transform -1 0 36960 0 -1 18816
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1947_
timestamp 1698431365
transform 1 0 36288 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1948_
timestamp 1698431365
transform 1 0 38976 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1949_
timestamp 1698431365
transform -1 0 39424 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1950_
timestamp 1698431365
transform 1 0 36960 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1951_
timestamp 1698431365
transform 1 0 38192 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1952_
timestamp 1698431365
transform 1 0 36064 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1953_
timestamp 1698431365
transform -1 0 38192 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1954_
timestamp 1698431365
transform 1 0 37184 0 -1 15680
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1955_
timestamp 1698431365
transform 1 0 37184 0 -1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1956_
timestamp 1698431365
transform -1 0 39984 0 -1 12544
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1957_
timestamp 1698431365
transform 1 0 37744 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1958_
timestamp 1698431365
transform -1 0 38528 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1959_
timestamp 1698431365
transform 1 0 38864 0 -1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1960_
timestamp 1698431365
transform 1 0 38640 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1961_
timestamp 1698431365
transform 1 0 39872 0 1 10976
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1962_
timestamp 1698431365
transform -1 0 40656 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1963_
timestamp 1698431365
transform -1 0 39984 0 1 14112
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1964_
timestamp 1698431365
transform 1 0 40656 0 1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1965_
timestamp 1698431365
transform 1 0 40768 0 -1 14112
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1966_
timestamp 1698431365
transform 1 0 39648 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1967_
timestamp 1698431365
transform -1 0 40544 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1968_
timestamp 1698431365
transform -1 0 42672 0 -1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1969_
timestamp 1698431365
transform 1 0 41664 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1970_
timestamp 1698431365
transform 1 0 37072 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1971_
timestamp 1698431365
transform 1 0 40768 0 -1 17248
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1972_
timestamp 1698431365
transform 1 0 40768 0 -1 15680
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1973_
timestamp 1698431365
transform -1 0 42224 0 -1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1974_
timestamp 1698431365
transform 1 0 42448 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1975_
timestamp 1698431365
transform -1 0 41888 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1976_
timestamp 1698431365
transform 1 0 40544 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1977_
timestamp 1698431365
transform -1 0 40544 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1978_
timestamp 1698431365
transform -1 0 42000 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1979_
timestamp 1698431365
transform 1 0 40768 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1980_
timestamp 1698431365
transform 1 0 45584 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1981_
timestamp 1698431365
transform -1 0 45472 0 -1 17248
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1982_
timestamp 1698431365
transform 1 0 43232 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1983_
timestamp 1698431365
transform 1 0 34048 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1984_
timestamp 1698431365
transform 1 0 44688 0 1 17248
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1985_
timestamp 1698431365
transform 1 0 46144 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1986_
timestamp 1698431365
transform 1 0 45472 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1987_
timestamp 1698431365
transform -1 0 46032 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1988_
timestamp 1698431365
transform 1 0 44688 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1989_
timestamp 1698431365
transform 1 0 45472 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1990_
timestamp 1698431365
transform -1 0 34720 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1991_
timestamp 1698431365
transform 1 0 44688 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1992_
timestamp 1698431365
transform 1 0 46480 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1993_
timestamp 1698431365
transform -1 0 47824 0 -1 15680
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1994_
timestamp 1698431365
transform 1 0 44128 0 -1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1995_
timestamp 1698431365
transform 1 0 45024 0 1 12544
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1996_
timestamp 1698431365
transform 1 0 46480 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1997_
timestamp 1698431365
transform 1 0 46704 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1998_
timestamp 1698431365
transform 1 0 47264 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1999_
timestamp 1698431365
transform 1 0 47712 0 -1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2000_
timestamp 1698431365
transform 1 0 47376 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2001_
timestamp 1698431365
transform 1 0 44800 0 1 10976
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2002_
timestamp 1698431365
transform 1 0 45920 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2003_
timestamp 1698431365
transform 1 0 45808 0 -1 14112
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2004_
timestamp 1698431365
transform 1 0 45808 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2005_
timestamp 1698431365
transform 1 0 46368 0 1 14112
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2006_
timestamp 1698431365
transform 1 0 47488 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2007_
timestamp 1698431365
transform 1 0 48608 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2008_
timestamp 1698431365
transform -1 0 49728 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2009_
timestamp 1698431365
transform 1 0 48272 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2010_
timestamp 1698431365
transform 1 0 48384 0 1 15680
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2011_
timestamp 1698431365
transform 1 0 48608 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2012_
timestamp 1698431365
transform 1 0 45920 0 1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2013_
timestamp 1698431365
transform -1 0 47040 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2014_
timestamp 1698431365
transform 1 0 46480 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2015_
timestamp 1698431365
transform 1 0 48608 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2016_
timestamp 1698431365
transform -1 0 48608 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2017_
timestamp 1698431365
transform 1 0 47152 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2018_
timestamp 1698431365
transform -1 0 49504 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2019_
timestamp 1698431365
transform -1 0 50960 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2020_
timestamp 1698431365
transform -1 0 49952 0 -1 23520
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2021_
timestamp 1698431365
transform 1 0 45472 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2022_
timestamp 1698431365
transform 1 0 44688 0 1 21952
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2023_
timestamp 1698431365
transform 1 0 47712 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2024_
timestamp 1698431365
transform 1 0 46816 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2025_
timestamp 1698431365
transform -1 0 48384 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2026_
timestamp 1698431365
transform -1 0 47712 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2027_
timestamp 1698431365
transform 1 0 50288 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2028_
timestamp 1698431365
transform 1 0 47040 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2029_
timestamp 1698431365
transform -1 0 50512 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2030_
timestamp 1698431365
transform -1 0 50288 0 -1 25088
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2031_
timestamp 1698431365
transform 1 0 45584 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2032_
timestamp 1698431365
transform 1 0 46928 0 1 26656
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2033_
timestamp 1698431365
transform 1 0 48608 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2034_
timestamp 1698431365
transform -1 0 48384 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2035_
timestamp 1698431365
transform -1 0 50624 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2036_
timestamp 1698431365
transform 1 0 49504 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2037_
timestamp 1698431365
transform 1 0 46144 0 1 26656
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2038_
timestamp 1698431365
transform 1 0 47824 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2039_
timestamp 1698431365
transform 1 0 48608 0 -1 28224
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2040_
timestamp 1698431365
transform 1 0 47040 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2041_
timestamp 1698431365
transform 1 0 47264 0 1 29792
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2042_
timestamp 1698431365
transform 1 0 49504 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2043_
timestamp 1698431365
transform -1 0 46816 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2044_
timestamp 1698431365
transform -1 0 48272 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2045_
timestamp 1698431365
transform -1 0 50960 0 1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2046_
timestamp 1698431365
transform 1 0 48608 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2047_
timestamp 1698431365
transform 1 0 47264 0 -1 29792
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2048_
timestamp 1698431365
transform 1 0 46368 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2049_
timestamp 1698431365
transform 1 0 44688 0 1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2050_
timestamp 1698431365
transform -1 0 45584 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2051_
timestamp 1698431365
transform 1 0 45808 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2052_
timestamp 1698431365
transform -1 0 46928 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2053_
timestamp 1698431365
transform -1 0 46032 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2054_
timestamp 1698431365
transform -1 0 47040 0 1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2055_
timestamp 1698431365
transform 1 0 45248 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2056_
timestamp 1698431365
transform -1 0 41440 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2057_
timestamp 1698431365
transform -1 0 40656 0 1 26656
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2058_
timestamp 1698431365
transform 1 0 38528 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2059_
timestamp 1698431365
transform 1 0 32256 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2060_
timestamp 1698431365
transform 1 0 37408 0 1 26656
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2061_
timestamp 1698431365
transform 1 0 37856 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2062_
timestamp 1698431365
transform 1 0 31696 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2063_
timestamp 1698431365
transform 1 0 34272 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2064_
timestamp 1698431365
transform -1 0 39648 0 -1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2065_
timestamp 1698431365
transform 1 0 38192 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2066_
timestamp 1698431365
transform -1 0 42112 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2067_
timestamp 1698431365
transform 1 0 40096 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2068_
timestamp 1698431365
transform -1 0 42336 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2069_
timestamp 1698431365
transform -1 0 42224 0 1 28224
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2070_
timestamp 1698431365
transform 1 0 39984 0 -1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2071_
timestamp 1698431365
transform 1 0 41664 0 1 29792
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2072_
timestamp 1698431365
transform -1 0 43120 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2073_
timestamp 1698431365
transform 1 0 42448 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2074_
timestamp 1698431365
transform -1 0 41552 0 -1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2075_
timestamp 1698431365
transform -1 0 42448 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2076_
timestamp 1698431365
transform 1 0 42336 0 1 26656
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2077_
timestamp 1698431365
transform -1 0 43568 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2078_
timestamp 1698431365
transform 1 0 40208 0 1 29792
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2079_
timestamp 1698431365
transform 1 0 36848 0 1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2080_
timestamp 1698431365
transform 1 0 37632 0 1 29792
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2081_
timestamp 1698431365
transform -1 0 39760 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2082_
timestamp 1698431365
transform 1 0 38976 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2083_
timestamp 1698431365
transform -1 0 40208 0 1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2084_
timestamp 1698431365
transform 1 0 38752 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2085_
timestamp 1698431365
transform 1 0 38192 0 -1 29792
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2086_
timestamp 1698431365
transform 1 0 37968 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2087_
timestamp 1698431365
transform 1 0 34160 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2088_
timestamp 1698431365
transform 1 0 34608 0 1 32928
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2089_
timestamp 1698431365
transform -1 0 35056 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2090_
timestamp 1698431365
transform 1 0 34384 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2091_
timestamp 1698431365
transform -1 0 34608 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2092_
timestamp 1698431365
transform -1 0 37744 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2093_
timestamp 1698431365
transform 1 0 30800 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2094_
timestamp 1698431365
transform -1 0 31696 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2095_
timestamp 1698431365
transform -1 0 35840 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2096_
timestamp 1698431365
transform -1 0 37408 0 1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2097_
timestamp 1698431365
transform 1 0 35728 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2098_
timestamp 1698431365
transform 1 0 36848 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2099_
timestamp 1698431365
transform 1 0 34048 0 1 28224
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2100_
timestamp 1698431365
transform 1 0 34272 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2101_
timestamp 1698431365
transform -1 0 35952 0 1 26656
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2102_
timestamp 1698431365
transform -1 0 34048 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2103_
timestamp 1698431365
transform 1 0 30800 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2104_
timestamp 1698431365
transform 1 0 32592 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2105_
timestamp 1698431365
transform -1 0 34272 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2106_
timestamp 1698431365
transform 1 0 35392 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2107_
timestamp 1698431365
transform 1 0 33712 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2108_
timestamp 1698431365
transform -1 0 36624 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2109_
timestamp 1698431365
transform -1 0 35952 0 -1 29792
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2110_
timestamp 1698431365
transform 1 0 29568 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2111_
timestamp 1698431365
transform 1 0 30688 0 1 28224
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2112_
timestamp 1698431365
transform -1 0 31920 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2113_
timestamp 1698431365
transform 1 0 31136 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2114_
timestamp 1698431365
transform 1 0 32032 0 -1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2115_
timestamp 1698431365
transform 1 0 29792 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2116_
timestamp 1698431365
transform -1 0 32704 0 -1 28224
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2117_
timestamp 1698431365
transform -1 0 32592 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2118_
timestamp 1698431365
transform -1 0 32256 0 1 29792
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2119_
timestamp 1698431365
transform 1 0 29008 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2120_
timestamp 1698431365
transform -1 0 31024 0 -1 29792
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2121_
timestamp 1698431365
transform -1 0 28784 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2122_
timestamp 1698431365
transform -1 0 27888 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2123_
timestamp 1698431365
transform 1 0 30688 0 -1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2124_
timestamp 1698431365
transform 1 0 27888 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2125_
timestamp 1698431365
transform 1 0 27104 0 1 31360
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2126_
timestamp 1698431365
transform 1 0 29120 0 1 29792
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2127_
timestamp 1698431365
transform 1 0 27552 0 1 34496
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2128_
timestamp 1698431365
transform -1 0 27552 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2129_
timestamp 1698431365
transform -1 0 30464 0 -1 34496
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2130_
timestamp 1698431365
transform -1 0 27888 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2131_
timestamp 1698431365
transform -1 0 28784 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2132_
timestamp 1698431365
transform 1 0 29904 0 1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2133_
timestamp 1698431365
transform 1 0 29008 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _2134_
timestamp 1698431365
transform -1 0 29456 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2135_
timestamp 1698431365
transform -1 0 26656 0 -1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2136_
timestamp 1698431365
transform 1 0 23744 0 -1 53312
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2137_
timestamp 1698431365
transform 1 0 31920 0 1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2138_
timestamp 1698431365
transform -1 0 33824 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2139_
timestamp 1698431365
transform -1 0 24752 0 -1 56448
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2140_
timestamp 1698431365
transform 1 0 25088 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2141_
timestamp 1698431365
transform 1 0 25088 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2142_
timestamp 1698431365
transform 1 0 26656 0 -1 54880
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2143_
timestamp 1698431365
transform -1 0 30688 0 1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2144_
timestamp 1698431365
transform 1 0 24304 0 -1 54880
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2145_
timestamp 1698431365
transform -1 0 26992 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2146_
timestamp 1698431365
transform -1 0 20944 0 1 50176
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2147_
timestamp 1698431365
transform 1 0 22624 0 -1 53312
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2148_
timestamp 1698431365
transform 1 0 24416 0 1 53312
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2149_
timestamp 1698431365
transform 1 0 29904 0 1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2150_
timestamp 1698431365
transform 1 0 33152 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2151_
timestamp 1698431365
transform 1 0 21840 0 1 50176
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2152_
timestamp 1698431365
transform -1 0 34720 0 1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2153_
timestamp 1698431365
transform 1 0 20160 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2154_
timestamp 1698431365
transform 1 0 21952 0 -1 51744
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2155_
timestamp 1698431365
transform 1 0 23072 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2156_
timestamp 1698431365
transform 1 0 21056 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2157_
timestamp 1698431365
transform -1 0 20944 0 1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2158_
timestamp 1698431365
transform 1 0 17248 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2159_
timestamp 1698431365
transform -1 0 20608 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2160_
timestamp 1698431365
transform -1 0 18704 0 1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2161_
timestamp 1698431365
transform 1 0 21840 0 1 51744
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2162_
timestamp 1698431365
transform 1 0 32144 0 1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2163_
timestamp 1698431365
transform 1 0 19600 0 -1 59584
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2164_
timestamp 1698431365
transform -1 0 21280 0 -1 58016
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2165_
timestamp 1698431365
transform -1 0 20048 0 1 58016
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2166_
timestamp 1698431365
transform 1 0 21168 0 1 56448
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2167_
timestamp 1698431365
transform -1 0 31696 0 1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2168_
timestamp 1698431365
transform 1 0 21280 0 -1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2169_
timestamp 1698431365
transform 1 0 20048 0 1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2170_
timestamp 1698431365
transform -1 0 19600 0 1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2171_
timestamp 1698431365
transform -1 0 19152 0 1 58016
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2172_
timestamp 1698431365
transform 1 0 20384 0 -1 59584
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2173_
timestamp 1698431365
transform 1 0 26768 0 1 59584
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2174_
timestamp 1698431365
transform -1 0 28448 0 1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2175_
timestamp 1698431365
transform -1 0 28560 0 1 59584
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2176_
timestamp 1698431365
transform 1 0 25872 0 1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2177_
timestamp 1698431365
transform -1 0 31472 0 1 59584
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2178_
timestamp 1698431365
transform 1 0 26656 0 1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2179_
timestamp 1698431365
transform 1 0 26096 0 1 61152
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2180_
timestamp 1698431365
transform 1 0 28336 0 -1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _2181_
timestamp 1698431365
transform -1 0 31136 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2182_
timestamp 1698431365
transform -1 0 27216 0 1 58016
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2183_
timestamp 1698431365
transform 1 0 23968 0 1 56448
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2184_
timestamp 1698431365
transform -1 0 24864 0 -1 58016
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2185_
timestamp 1698431365
transform -1 0 25984 0 -1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2186_
timestamp 1698431365
transform -1 0 23968 0 1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2187_
timestamp 1698431365
transform 1 0 25984 0 -1 59584
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2188_
timestamp 1698431365
transform -1 0 24864 0 -1 59584
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2189_
timestamp 1698431365
transform 1 0 22512 0 -1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2190_
timestamp 1698431365
transform 1 0 21952 0 -1 61152
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2191_
timestamp 1698431365
transform 1 0 22288 0 1 56448
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2192_
timestamp 1698431365
transform 1 0 24864 0 1 58016
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2193_
timestamp 1698431365
transform 1 0 22624 0 1 62720
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2194_
timestamp 1698431365
transform -1 0 22624 0 1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2195_
timestamp 1698431365
transform 1 0 23744 0 1 62720
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2196_
timestamp 1698431365
transform -1 0 23408 0 -1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2197_
timestamp 1698431365
transform -1 0 24640 0 -1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2198_
timestamp 1698431365
transform -1 0 22848 0 -1 64288
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2199_
timestamp 1698431365
transform 1 0 24192 0 -1 61152
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2200_
timestamp 1698431365
transform 1 0 25984 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2201_
timestamp 1698431365
transform -1 0 26768 0 1 64288
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2202_
timestamp 1698431365
transform 1 0 24416 0 1 61152
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2203_
timestamp 1698431365
transform -1 0 25872 0 1 65856
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2204_
timestamp 1698431365
transform -1 0 33824 0 -1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2205_
timestamp 1698431365
transform -1 0 26432 0 1 65856
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2206_
timestamp 1698431365
transform -1 0 26880 0 -1 64288
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2207_
timestamp 1698431365
transform 1 0 24528 0 1 65856
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2208_
timestamp 1698431365
transform -1 0 25984 0 -1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2209_
timestamp 1698431365
transform 1 0 24864 0 1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2210_
timestamp 1698431365
transform -1 0 23744 0 -1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2211_
timestamp 1698431365
transform -1 0 24752 0 -1 65856
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2212_
timestamp 1698431365
transform -1 0 26320 0 -1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2213_
timestamp 1698431365
transform 1 0 27664 0 1 64288
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2214_
timestamp 1698431365
transform 1 0 27664 0 1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2215_
timestamp 1698431365
transform 1 0 27888 0 -1 64288
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2216_
timestamp 1698431365
transform -1 0 27664 0 1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2217_
timestamp 1698431365
transform 1 0 29904 0 -1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2218_
timestamp 1698431365
transform -1 0 29120 0 -1 64288
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2219_
timestamp 1698431365
transform -1 0 27664 0 1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _2220_
timestamp 1698431365
transform 1 0 32144 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2221_
timestamp 1698431365
transform 1 0 34832 0 1 61152
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2222_
timestamp 1698431365
transform 1 0 33040 0 1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2223_
timestamp 1698431365
transform -1 0 34048 0 -1 59584
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2224_
timestamp 1698431365
transform 1 0 33824 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2225_
timestamp 1698431365
transform -1 0 34832 0 1 61152
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2226_
timestamp 1698431365
transform 1 0 32816 0 1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2227_
timestamp 1698431365
transform 1 0 32928 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2228_
timestamp 1698431365
transform -1 0 32704 0 -1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2229_
timestamp 1698431365
transform 1 0 34048 0 -1 59584
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2230_
timestamp 1698431365
transform 1 0 34720 0 1 58016
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2231_
timestamp 1698431365
transform 1 0 34048 0 1 58016
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2232_
timestamp 1698431365
transform 1 0 34608 0 -1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2233_
timestamp 1698431365
transform -1 0 29568 0 1 61152
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2234_
timestamp 1698431365
transform 1 0 34720 0 1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2235_
timestamp 1698431365
transform -1 0 33712 0 -1 62720
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2236_
timestamp 1698431365
transform 1 0 32928 0 -1 61152
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2237_
timestamp 1698431365
transform 1 0 29568 0 1 61152
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2238_
timestamp 1698431365
transform -1 0 30800 0 -1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2239_
timestamp 1698431365
transform 1 0 30128 0 -1 64288
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2240_
timestamp 1698431365
transform 1 0 32144 0 1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2241_
timestamp 1698431365
transform 1 0 29232 0 -1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2242_
timestamp 1698431365
transform 1 0 28000 0 -1 62720
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2243_
timestamp 1698431365
transform -1 0 34272 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2244_
timestamp 1698431365
transform -1 0 32704 0 -1 64288
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2245_
timestamp 1698431365
transform 1 0 30688 0 1 61152
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2246_
timestamp 1698431365
transform 1 0 33712 0 -1 62720
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2247_
timestamp 1698431365
transform -1 0 34384 0 -1 64288
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2248_
timestamp 1698431365
transform -1 0 33824 0 1 65856
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2249_
timestamp 1698431365
transform 1 0 31472 0 -1 64288
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2250_
timestamp 1698431365
transform -1 0 33824 0 -1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2251_
timestamp 1698431365
transform -1 0 33824 0 -1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2252_
timestamp 1698431365
transform 1 0 34272 0 1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2253_
timestamp 1698431365
transform -1 0 32704 0 -1 65856
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2254_
timestamp 1698431365
transform 1 0 33824 0 -1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2255_
timestamp 1698431365
transform 1 0 35504 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2256_
timestamp 1698431365
transform 1 0 35504 0 1 64288
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2257_
timestamp 1698431365
transform 1 0 36848 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2258_
timestamp 1698431365
transform -1 0 38640 0 1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2259_
timestamp 1698431365
transform -1 0 36624 0 1 65856
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2260_
timestamp 1698431365
transform 1 0 35056 0 1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2261_
timestamp 1698431365
transform 1 0 37632 0 -1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2262_
timestamp 1698431365
transform -1 0 37408 0 1 62720
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2263_
timestamp 1698431365
transform -1 0 36288 0 1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _2264_
timestamp 1698431365
transform -1 0 36624 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2265_
timestamp 1698431365
transform 1 0 38864 0 1 61152
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2266_
timestamp 1698431365
transform -1 0 38976 0 -1 59584
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2267_
timestamp 1698431365
transform -1 0 38864 0 1 61152
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2268_
timestamp 1698431365
transform -1 0 37744 0 1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2269_
timestamp 1698431365
transform -1 0 37968 0 1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2270_
timestamp 1698431365
transform 1 0 37968 0 1 58016
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2271_
timestamp 1698431365
transform -1 0 40208 0 -1 59584
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2272_
timestamp 1698431365
transform 1 0 38752 0 -1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2273_
timestamp 1698431365
transform 1 0 38304 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2274_
timestamp 1698431365
transform 1 0 39088 0 -1 59584
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2275_
timestamp 1698431365
transform -1 0 40208 0 1 59584
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2276_
timestamp 1698431365
transform -1 0 39424 0 1 59584
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2277_
timestamp 1698431365
transform 1 0 38528 0 1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2278_
timestamp 1698431365
transform 1 0 39872 0 1 58016
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2279_
timestamp 1698431365
transform 1 0 33824 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2280_
timestamp 1698431365
transform -1 0 39872 0 1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2281_
timestamp 1698431365
transform 1 0 40992 0 1 58016
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2282_
timestamp 1698431365
transform 1 0 38192 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2283_
timestamp 1698431365
transform -1 0 41664 0 -1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2284_
timestamp 1698431365
transform 1 0 41664 0 -1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2285_
timestamp 1698431365
transform -1 0 40768 0 1 59584
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2286_
timestamp 1698431365
transform -1 0 42448 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2287_
timestamp 1698431365
transform -1 0 42000 0 1 61152
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2288_
timestamp 1698431365
transform 1 0 40768 0 -1 59584
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2289_
timestamp 1698431365
transform 1 0 37856 0 1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2290_
timestamp 1698431365
transform -1 0 42448 0 -1 62720
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2291_
timestamp 1698431365
transform -1 0 42784 0 -1 64288
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2292_
timestamp 1698431365
transform -1 0 42224 0 -1 64288
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2293_
timestamp 1698431365
transform -1 0 40432 0 1 61152
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2294_
timestamp 1698431365
transform 1 0 40768 0 -1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2295_
timestamp 1698431365
transform 1 0 39648 0 -1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2296_
timestamp 1698431365
transform 1 0 40432 0 1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2297_
timestamp 1698431365
transform -1 0 43120 0 -1 62720
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2298_
timestamp 1698431365
transform 1 0 39200 0 1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2299_
timestamp 1698431365
transform 1 0 40768 0 1 64288
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2300_
timestamp 1698431365
transform 1 0 40768 0 -1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2301_
timestamp 1698431365
transform 1 0 40768 0 -1 65856
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2302_
timestamp 1698431365
transform -1 0 40320 0 -1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2303_
timestamp 1698431365
transform -1 0 39536 0 1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2304_
timestamp 1698431365
transform -1 0 40096 0 1 65856
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2305_
timestamp 1698431365
transform 1 0 38528 0 -1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _2306_
timestamp 1698431365
transform -1 0 49168 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2307_
timestamp 1698431365
transform -1 0 51072 0 1 61152
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2308_
timestamp 1698431365
transform 1 0 47152 0 1 59584
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2309_
timestamp 1698431365
transform -1 0 50064 0 -1 61152
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2310_
timestamp 1698431365
transform -1 0 49504 0 1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2311_
timestamp 1698431365
transform -1 0 45584 0 1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2312_
timestamp 1698431365
transform 1 0 46928 0 -1 64288
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2313_
timestamp 1698431365
transform 1 0 23408 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2314_
timestamp 1698431365
transform 1 0 44912 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2315_
timestamp 1698431365
transform -1 0 49168 0 -1 59584
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2316_
timestamp 1698431365
transform 1 0 47488 0 -1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2317_
timestamp 1698431365
transform -1 0 48384 0 -1 58016
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2318_
timestamp 1698431365
transform 1 0 46368 0 1 59584
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2319_
timestamp 1698431365
transform 1 0 46704 0 -1 61152
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2320_
timestamp 1698431365
transform 1 0 45808 0 -1 58016
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2321_
timestamp 1698431365
transform 1 0 44912 0 -1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2322_
timestamp 1698431365
transform 1 0 46032 0 -1 59584
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2323_
timestamp 1698431365
transform 1 0 46928 0 -1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2324_
timestamp 1698431365
transform 1 0 47152 0 -1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2325_
timestamp 1698431365
transform 1 0 47152 0 1 56448
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2326_
timestamp 1698431365
transform -1 0 45808 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2327_
timestamp 1698431365
transform -1 0 42560 0 1 59584
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2328_
timestamp 1698431365
transform 1 0 45584 0 1 58016
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2329_
timestamp 1698431365
transform 1 0 42560 0 1 59584
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2330_
timestamp 1698431365
transform 1 0 42336 0 -1 59584
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2331_
timestamp 1698431365
transform 1 0 43456 0 1 58016
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2332_
timestamp 1698431365
transform -1 0 44016 0 -1 58016
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2333_
timestamp 1698431365
transform -1 0 45584 0 1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2334_
timestamp 1698431365
transform 1 0 43344 0 -1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2335_
timestamp 1698431365
transform 1 0 43344 0 1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2336_
timestamp 1698431365
transform 1 0 44688 0 1 59584
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2337_
timestamp 1698431365
transform 1 0 44240 0 -1 59584
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2338_
timestamp 1698431365
transform 1 0 44800 0 1 47040
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2339_
timestamp 1698431365
transform 1 0 43568 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2340_
timestamp 1698431365
transform 1 0 46816 0 1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2341_
timestamp 1698431365
transform 1 0 46368 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2342_
timestamp 1698431365
transform 1 0 31808 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2343_
timestamp 1698431365
transform -1 0 46368 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2344_
timestamp 1698431365
transform 1 0 47488 0 1 47040
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2345_
timestamp 1698431365
transform 1 0 47264 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _2346_
timestamp 1698431365
transform -1 0 50624 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2347_
timestamp 1698431365
transform -1 0 49616 0 -1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2348_
timestamp 1698431365
transform 1 0 48608 0 -1 56448
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2349_
timestamp 1698431365
transform -1 0 49728 0 1 54880
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2350_
timestamp 1698431365
transform 1 0 49168 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2351_
timestamp 1698431365
transform -1 0 48384 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2352_
timestamp 1698431365
transform 1 0 47824 0 -1 53312
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2353_
timestamp 1698431365
transform 1 0 50064 0 1 53312
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2354_
timestamp 1698431365
transform 1 0 49728 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2355_
timestamp 1698431365
transform 1 0 47264 0 -1 51744
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2356_
timestamp 1698431365
transform 1 0 47488 0 -1 56448
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2357_
timestamp 1698431365
transform 1 0 47488 0 1 53312
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2358_
timestamp 1698431365
transform 1 0 45584 0 -1 53312
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2359_
timestamp 1698431365
transform 1 0 44688 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2360_
timestamp 1698431365
transform 1 0 46704 0 -1 53312
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2361_
timestamp 1698431365
transform 1 0 48608 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2362_
timestamp 1698431365
transform 1 0 46368 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2363_
timestamp 1698431365
transform 1 0 47824 0 -1 51744
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2364_
timestamp 1698431365
transform -1 0 44128 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2365_
timestamp 1698431365
transform -1 0 42560 0 1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2366_
timestamp 1698431365
transform 1 0 45808 0 -1 51744
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2367_
timestamp 1698431365
transform 1 0 42560 0 1 48608
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2368_
timestamp 1698431365
transform 1 0 41328 0 1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2369_
timestamp 1698431365
transform 1 0 42000 0 -1 50176
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2370_
timestamp 1698431365
transform 1 0 43120 0 -1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2371_
timestamp 1698431365
transform -1 0 44240 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2372_
timestamp 1698431365
transform 1 0 43904 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2373_
timestamp 1698431365
transform 1 0 43456 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2374_
timestamp 1698431365
transform 1 0 45136 0 1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2375_
timestamp 1698431365
transform -1 0 43904 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2376_
timestamp 1698431365
transform -1 0 44240 0 1 45472
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2377_
timestamp 1698431365
transform 1 0 44240 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2378_
timestamp 1698431365
transform -1 0 43120 0 1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2379_
timestamp 1698431365
transform 1 0 43344 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2380_
timestamp 1698431365
transform 1 0 44688 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2381_
timestamp 1698431365
transform -1 0 46144 0 -1 45472
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2382_
timestamp 1698431365
transform 1 0 44016 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _2383_
timestamp 1698431365
transform -1 0 43568 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2384_
timestamp 1698431365
transform -1 0 36736 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2385_
timestamp 1698431365
transform 1 0 35504 0 1 48608
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2386_
timestamp 1698431365
transform -1 0 38304 0 1 50176
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2387_
timestamp 1698431365
transform 1 0 37744 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2388_
timestamp 1698431365
transform 1 0 36848 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2389_
timestamp 1698431365
transform -1 0 35504 0 -1 50176
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2390_
timestamp 1698431365
transform -1 0 35616 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2391_
timestamp 1698431365
transform -1 0 38304 0 1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2392_
timestamp 1698431365
transform -1 0 35392 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2393_
timestamp 1698431365
transform 1 0 41552 0 1 50176
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2394_
timestamp 1698431365
transform 1 0 35840 0 1 50176
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2395_
timestamp 1698431365
transform 1 0 36736 0 -1 50176
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2396_
timestamp 1698431365
transform -1 0 40320 0 1 51744
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2397_
timestamp 1698431365
transform 1 0 38976 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2398_
timestamp 1698431365
transform -1 0 40320 0 -1 51744
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2399_
timestamp 1698431365
transform -1 0 39200 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2400_
timestamp 1698431365
transform -1 0 39200 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2401_
timestamp 1698431365
transform 1 0 37744 0 -1 51744
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2402_
timestamp 1698431365
transform 1 0 40768 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2403_
timestamp 1698431365
transform 1 0 40880 0 1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2404_
timestamp 1698431365
transform -1 0 40432 0 -1 50176
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2405_
timestamp 1698431365
transform 1 0 37856 0 -1 48608
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2406_
timestamp 1698431365
transform -1 0 39984 0 1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2407_
timestamp 1698431365
transform 1 0 38864 0 1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2408_
timestamp 1698431365
transform -1 0 41328 0 -1 47040
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2409_
timestamp 1698431365
transform -1 0 40432 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2410_
timestamp 1698431365
transform -1 0 40880 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2411_
timestamp 1698431365
transform -1 0 39984 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2412_
timestamp 1698431365
transform -1 0 39088 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2413_
timestamp 1698431365
transform -1 0 39536 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2414_
timestamp 1698431365
transform -1 0 34496 0 -1 47040
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2415_
timestamp 1698431365
transform 1 0 34496 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2416_
timestamp 1698431365
transform -1 0 33824 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2417_
timestamp 1698431365
transform -1 0 36624 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2418_
timestamp 1698431365
transform 1 0 35392 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2419_
timestamp 1698431365
transform -1 0 37408 0 1 45472
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2420_
timestamp 1698431365
transform 1 0 35616 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _2421_
timestamp 1698431365
transform -1 0 34272 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2422_
timestamp 1698431365
transform -1 0 33600 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2423_
timestamp 1698431365
transform -1 0 31472 0 1 47040
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2424_
timestamp 1698431365
transform -1 0 32256 0 -1 48608
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2425_
timestamp 1698431365
transform 1 0 31472 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2426_
timestamp 1698431365
transform 1 0 29456 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2427_
timestamp 1698431365
transform -1 0 29568 0 1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2428_
timestamp 1698431365
transform 1 0 32144 0 -1 45472
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2429_
timestamp 1698431365
transform 1 0 32368 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2430_
timestamp 1698431365
transform -1 0 27440 0 -1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2431_
timestamp 1698431365
transform 1 0 30016 0 -1 50176
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2432_
timestamp 1698431365
transform 1 0 30128 0 -1 47040
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2433_
timestamp 1698431365
transform -1 0 29008 0 -1 45472
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2434_
timestamp 1698431365
transform -1 0 29904 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2435_
timestamp 1698431365
transform -1 0 28560 0 1 43904
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2436_
timestamp 1698431365
transform -1 0 15344 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2437_
timestamp 1698431365
transform -1 0 27440 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2438_
timestamp 1698431365
transform -1 0 27776 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2439_
timestamp 1698431365
transform -1 0 27328 0 1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2440_
timestamp 1698431365
transform 1 0 27328 0 1 45472
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2441_
timestamp 1698431365
transform -1 0 28448 0 -1 50176
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2442_
timestamp 1698431365
transform -1 0 28448 0 1 48608
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2443_
timestamp 1698431365
transform 1 0 26432 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2444_
timestamp 1698431365
transform 1 0 27888 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2445_
timestamp 1698431365
transform -1 0 28896 0 -1 47040
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2446_
timestamp 1698431365
transform 1 0 27328 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2447_
timestamp 1698431365
transform 1 0 27104 0 -1 50176
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2448_
timestamp 1698431365
transform 1 0 26208 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2449_
timestamp 1698431365
transform -1 0 28672 0 1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2450_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 25088 0 1 36064
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2451_
timestamp 1698431365
transform 1 0 31472 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2452_
timestamp 1698431365
transform -1 0 25648 0 -1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2453_
timestamp 1698431365
transform -1 0 26544 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2454_
timestamp 1698431365
transform -1 0 23856 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2455_
timestamp 1698431365
transform 1 0 23408 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2456_
timestamp 1698431365
transform -1 0 24864 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2457_
timestamp 1698431365
transform 1 0 22736 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2458_
timestamp 1698431365
transform 1 0 27664 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2459_
timestamp 1698431365
transform -1 0 30800 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2460_
timestamp 1698431365
transform 1 0 27888 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2461_
timestamp 1698431365
transform 1 0 32928 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2462_
timestamp 1698431365
transform 1 0 35280 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2463_
timestamp 1698431365
transform -1 0 37408 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2464_
timestamp 1698431365
transform 1 0 35392 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2465_
timestamp 1698431365
transform -1 0 43120 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2466_
timestamp 1698431365
transform -1 0 44016 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2467_
timestamp 1698431365
transform -1 0 45248 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2468_
timestamp 1698431365
transform 1 0 43344 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2469_
timestamp 1698431365
transform -1 0 48160 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2470_
timestamp 1698431365
transform -1 0 48048 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2471_
timestamp 1698431365
transform -1 0 48048 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2472_
timestamp 1698431365
transform 1 0 45584 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2473_
timestamp 1698431365
transform 1 0 43120 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2474_
timestamp 1698431365
transform -1 0 44464 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2475_
timestamp 1698431365
transform 1 0 33264 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2476_
timestamp 1698431365
transform -1 0 36736 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2477_
timestamp 1698431365
transform 1 0 36176 0 -1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2478_
timestamp 1698431365
transform 1 0 35168 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2479_
timestamp 1698431365
transform 1 0 29792 0 1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2480_
timestamp 1698431365
transform -1 0 29344 0 -1 34496
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _2481_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 28784 0 1 54880
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2482_
timestamp 1698431365
transform 1 0 26768 0 -1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _2483_
timestamp 1698431365
transform 1 0 27552 0 1 58016
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2484_
timestamp 1698431365
transform -1 0 29904 0 1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _2485_
timestamp 1698431365
transform 1 0 29344 0 1 58016
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2486_
timestamp 1698431365
transform 1 0 34608 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2487_
timestamp 1698431365
transform -1 0 37744 0 1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _2488_
timestamp 1698431365
transform -1 0 36400 0 1 59584
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2489_
timestamp 1698431365
transform 1 0 31024 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2490_
timestamp 1698431365
transform -1 0 42784 0 1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _2491_
timestamp 1698431365
transform 1 0 45584 0 1 61152
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2492_
timestamp 1698431365
transform 1 0 45920 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _2493_
timestamp 1698431365
transform 1 0 45808 0 1 48608
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2494_
timestamp 1698431365
transform 1 0 42448 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _2495_
timestamp 1698431365
transform -1 0 42448 0 -1 47040
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2496_
timestamp 1698431365
transform 1 0 29680 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2497_
timestamp 1698431365
transform -1 0 35728 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _2498_
timestamp 1698431365
transform -1 0 32144 0 -1 45472
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2499_
timestamp 1698431365
transform 1 0 17248 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _2500_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 19152 0 1 39200
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2501_
timestamp 1698431365
transform -1 0 18928 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2502_
timestamp 1698431365
transform -1 0 22064 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai222_2  _2503_
timestamp 1698431365
transform -1 0 24192 0 1 20384
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2504_
timestamp 1698431365
transform 1 0 24192 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2505_
timestamp 1698431365
transform 1 0 18368 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai222_2  _2506_
timestamp 1698431365
transform 1 0 17920 0 1 21952
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2507_
timestamp 1698431365
transform -1 0 20608 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai222_2  _2508_
timestamp 1698431365
transform 1 0 18592 0 -1 20384
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2509_
timestamp 1698431365
transform 1 0 16576 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2510_
timestamp 1698431365
transform 1 0 17472 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai222_2  _2511_
timestamp 1698431365
transform 1 0 18816 0 -1 18816
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2512_
timestamp 1698431365
transform -1 0 19824 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2513_
timestamp 1698431365
transform -1 0 18368 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai222_2  _2514_
timestamp 1698431365
transform 1 0 17808 0 1 14112
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2515_
timestamp 1698431365
transform -1 0 18816 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2516_
timestamp 1698431365
transform -1 0 14448 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2517_
timestamp 1698431365
transform 1 0 13776 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai222_2  _2518_
timestamp 1698431365
transform 1 0 16352 0 1 17248
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2519_
timestamp 1698431365
transform -1 0 17024 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai222_1  _2520_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 15232 0 -1 18816
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2521_
timestamp 1698431365
transform -1 0 17696 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2522_
timestamp 1698431365
transform 1 0 15904 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai222_2  _2523_
timestamp 1698431365
transform 1 0 13888 0 1 20384
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2524_
timestamp 1698431365
transform 1 0 16576 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2525_
timestamp 1698431365
transform -1 0 14000 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2526_
timestamp 1698431365
transform 1 0 12208 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai222_2  _2527_
timestamp 1698431365
transform 1 0 13552 0 1 18816
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2528_
timestamp 1698431365
transform -1 0 14896 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2529_
timestamp 1698431365
transform 1 0 15008 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai222_2  _2530_
timestamp 1698431365
transform 1 0 13328 0 1 17248
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2531_
timestamp 1698431365
transform -1 0 13776 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai222_2  _2532_
timestamp 1698431365
transform -1 0 19600 0 1 18816
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2533_
timestamp 1698431365
transform -1 0 13664 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2534_
timestamp 1698431365
transform -1 0 13104 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai222_2  _2535_
timestamp 1698431365
transform 1 0 10080 0 1 18816
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2536_
timestamp 1698431365
transform 1 0 12544 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2537_
timestamp 1698431365
transform -1 0 11984 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai222_2  _2538_
timestamp 1698431365
transform 1 0 7056 0 1 18816
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2539_
timestamp 1698431365
transform -1 0 11312 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2540_
timestamp 1698431365
transform -1 0 10304 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai222_2  _2541_
timestamp 1698431365
transform 1 0 9408 0 1 14112
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2542_
timestamp 1698431365
transform 1 0 8736 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai222_2  _2543_
timestamp 1698431365
transform 1 0 6160 0 -1 18816
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2544_
timestamp 1698431365
transform -1 0 10752 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2545_
timestamp 1698431365
transform -1 0 15120 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2546_
timestamp 1698431365
transform -1 0 10416 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai222_2  _2547_
timestamp 1698431365
transform 1 0 9184 0 1 20384
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2548_
timestamp 1698431365
transform 1 0 6608 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2549_
timestamp 1698431365
transform -1 0 12432 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai222_2  _2550_
timestamp 1698431365
transform 1 0 6160 0 -1 21952
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2551_
timestamp 1698431365
transform -1 0 9856 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2552_
timestamp 1698431365
transform -1 0 11536 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai222_2  _2553_
timestamp 1698431365
transform -1 0 10640 0 1 21952
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2554_
timestamp 1698431365
transform -1 0 7280 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai222_1  _2555_
timestamp 1698431365
transform 1 0 6832 0 1 23520
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2556_
timestamp 1698431365
transform -1 0 9072 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2557_
timestamp 1698431365
transform 1 0 10976 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai222_2  _2558_
timestamp 1698431365
transform 1 0 9408 0 -1 23520
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2559_
timestamp 1698431365
transform -1 0 8512 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2560_
timestamp 1698431365
transform -1 0 13328 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai222_2  _2561_
timestamp 1698431365
transform 1 0 10080 0 1 25088
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2562_
timestamp 1698431365
transform 1 0 10976 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2563_
timestamp 1698431365
transform -1 0 12096 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai222_2  _2564_
timestamp 1698431365
transform 1 0 13328 0 1 26656
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2565_
timestamp 1698431365
transform -1 0 13776 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai222_2  _2566_
timestamp 1698431365
transform 1 0 11424 0 -1 25088
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2567_
timestamp 1698431365
transform -1 0 13776 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2568_
timestamp 1698431365
transform 1 0 11088 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai222_2  _2569_
timestamp 1698431365
transform 1 0 12656 0 -1 29792
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2570_
timestamp 1698431365
transform -1 0 10192 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2571_
timestamp 1698431365
transform -1 0 13104 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai222_2  _2572_
timestamp 1698431365
transform 1 0 9632 0 -1 29792
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2573_
timestamp 1698431365
transform -1 0 9184 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2574_
timestamp 1698431365
transform -1 0 12880 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai222_2  _2575_
timestamp 1698431365
transform 1 0 9632 0 -1 31360
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2576_
timestamp 1698431365
transform -1 0 9184 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai222_2  _2577_
timestamp 1698431365
transform 1 0 11312 0 -1 32928
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2578_
timestamp 1698431365
transform -1 0 10192 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2579_
timestamp 1698431365
transform -1 0 14336 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai222_2  _2580_
timestamp 1698431365
transform 1 0 10416 0 -1 34496
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2581_
timestamp 1698431365
transform -1 0 10416 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai222_2  _2582_
timestamp 1698431365
transform 1 0 10416 0 -1 36064
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2583_
timestamp 1698431365
transform -1 0 10528 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai222_2  _2584_
timestamp 1698431365
transform -1 0 16352 0 1 37632
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2585_
timestamp 1698431365
transform -1 0 10976 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai222_2  _2586_
timestamp 1698431365
transform 1 0 10080 0 1 39200
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2587_
timestamp 1698431365
transform -1 0 13776 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2588_
timestamp 1698431365
transform -1 0 14000 0 1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2589_
timestamp 1698431365
transform 1 0 13664 0 1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2590_
timestamp 1698431365
transform 1 0 17808 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2591_
timestamp 1698431365
transform -1 0 18592 0 -1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2592_
timestamp 1698431365
transform 1 0 17248 0 -1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2593_
timestamp 1698431365
transform 1 0 17472 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2594_
timestamp 1698431365
transform 1 0 17696 0 1 48608
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2595_
timestamp 1698431365
transform -1 0 17024 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2596_
timestamp 1698431365
transform 1 0 16016 0 -1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2597_
timestamp 1698431365
transform -1 0 16576 0 -1 51744
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2598_
timestamp 1698431365
transform 1 0 15904 0 -1 50176
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2599_
timestamp 1698431365
transform -1 0 17024 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2600_
timestamp 1698431365
transform 1 0 16128 0 1 53312
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2601_
timestamp 1698431365
transform -1 0 16128 0 -1 53312
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2602_
timestamp 1698431365
transform -1 0 14784 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2603_
timestamp 1698431365
transform -1 0 15456 0 -1 54880
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2604_
timestamp 1698431365
transform -1 0 15120 0 -1 53312
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2605_
timestamp 1698431365
transform 1 0 14000 0 1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2606_
timestamp 1698431365
transform -1 0 15904 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2607_
timestamp 1698431365
transform 1 0 13888 0 1 58016
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2608_
timestamp 1698431365
transform -1 0 16912 0 -1 56448
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2609_
timestamp 1698431365
transform -1 0 16352 0 -1 56448
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2610_
timestamp 1698431365
transform 1 0 13552 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2611_
timestamp 1698431365
transform 1 0 16352 0 -1 61152
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2612_
timestamp 1698431365
transform -1 0 18144 0 1 58016
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2613_
timestamp 1698431365
transform -1 0 15680 0 1 58016
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2614_
timestamp 1698431365
transform -1 0 17696 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2615_
timestamp 1698431365
transform 1 0 17024 0 1 58016
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2616_
timestamp 1698431365
transform -1 0 16688 0 1 58016
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2617_
timestamp 1698431365
transform -1 0 16688 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2618_
timestamp 1698431365
transform -1 0 16352 0 -1 61152
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2619_
timestamp 1698431365
transform -1 0 16240 0 1 59584
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2620_
timestamp 1698431365
transform 1 0 14336 0 -1 61152
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2621_
timestamp 1698431365
transform -1 0 17696 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2622_
timestamp 1698431365
transform 1 0 13440 0 1 61152
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2623_
timestamp 1698431365
transform -1 0 17024 0 -1 62720
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2624_
timestamp 1698431365
transform -1 0 16464 0 -1 62720
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2625_
timestamp 1698431365
transform -1 0 17696 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2626_
timestamp 1698431365
transform -1 0 15792 0 -1 64288
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2627_
timestamp 1698431365
transform -1 0 16688 0 -1 65856
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2628_
timestamp 1698431365
transform 1 0 15792 0 -1 64288
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2629_
timestamp 1698431365
transform -1 0 18704 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2630_
timestamp 1698431365
transform -1 0 15120 0 -1 64288
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2631_
timestamp 1698431365
transform 1 0 17248 0 -1 65856
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2632_
timestamp 1698431365
transform -1 0 15568 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2633_
timestamp 1698431365
transform 1 0 13776 0 1 65856
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2634_
timestamp 1698431365
transform 1 0 13440 0 1 64288
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2635_
timestamp 1698431365
transform -1 0 13104 0 1 61152
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2636_
timestamp 1698431365
transform -1 0 14224 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2637_
timestamp 1698431365
transform -1 0 13328 0 -1 61152
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2638_
timestamp 1698431365
transform 1 0 13216 0 -1 64288
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2639_
timestamp 1698431365
transform -1 0 13216 0 -1 64288
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2640_
timestamp 1698431365
transform -1 0 12880 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2641_
timestamp 1698431365
transform -1 0 12208 0 -1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2642_
timestamp 1698431365
transform 1 0 11088 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2643_
timestamp 1698431365
transform -1 0 13216 0 -1 62720
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2644_
timestamp 1698431365
transform -1 0 12208 0 -1 64288
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2645_
timestamp 1698431365
transform 1 0 9856 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2646_
timestamp 1698431365
transform -1 0 11984 0 1 62720
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2647_
timestamp 1698431365
transform -1 0 11312 0 1 61152
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2648_
timestamp 1698431365
transform -1 0 12432 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2649_
timestamp 1698431365
transform -1 0 11984 0 1 59584
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2650_
timestamp 1698431365
transform 1 0 11312 0 1 61152
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2651_
timestamp 1698431365
transform -1 0 11648 0 1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2652_
timestamp 1698431365
transform -1 0 9968 0 1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2653_
timestamp 1698431365
transform -1 0 11984 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2654_
timestamp 1698431365
transform -1 0 10416 0 -1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2655_
timestamp 1698431365
transform 1 0 9520 0 -1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2656_
timestamp 1698431365
transform -1 0 11536 0 1 56448
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2657_
timestamp 1698431365
transform -1 0 11200 0 -1 58016
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2658_
timestamp 1698431365
transform -1 0 11424 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2659_
timestamp 1698431365
transform -1 0 9184 0 -1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2660_
timestamp 1698431365
transform -1 0 10528 0 1 56448
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2661_
timestamp 1698431365
transform 1 0 9968 0 1 53312
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2662_
timestamp 1698431365
transform -1 0 10976 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2663_
timestamp 1698431365
transform 1 0 9408 0 -1 58016
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2664_
timestamp 1698431365
transform 1 0 9744 0 -1 56448
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2665_
timestamp 1698431365
transform -1 0 9184 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2666_
timestamp 1698431365
transform 1 0 8624 0 -1 56448
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2667_
timestamp 1698431365
transform -1 0 9744 0 1 56448
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2668_
timestamp 1698431365
transform -1 0 8288 0 -1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2669_
timestamp 1698431365
transform -1 0 8624 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2670_
timestamp 1698431365
transform -1 0 8960 0 -1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2671_
timestamp 1698431365
transform -1 0 7952 0 -1 54880
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2672_
timestamp 1698431365
transform -1 0 7728 0 -1 56448
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2673_
timestamp 1698431365
transform -1 0 8176 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2674_
timestamp 1698431365
transform -1 0 8736 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2675_
timestamp 1698431365
transform -1 0 7952 0 1 53312
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2676_
timestamp 1698431365
transform -1 0 7392 0 -1 54880
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2677_
timestamp 1698431365
transform -1 0 8400 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2678_
timestamp 1698431365
transform -1 0 7952 0 1 51744
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2679_
timestamp 1698431365
transform -1 0 7392 0 1 53312
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2680_
timestamp 1698431365
transform -1 0 8400 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2681_
timestamp 1698431365
transform -1 0 7392 0 1 50176
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2682_
timestamp 1698431365
transform -1 0 7392 0 1 51744
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2683_
timestamp 1698431365
transform -1 0 8288 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2684_
timestamp 1698431365
transform -1 0 9184 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2685_
timestamp 1698431365
transform -1 0 8064 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2686_
timestamp 1698431365
transform -1 0 7392 0 -1 50176
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2687_
timestamp 1698431365
transform 1 0 6608 0 -1 48608
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2688_
timestamp 1698431365
transform 1 0 6160 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2689_
timestamp 1698431365
transform -1 0 9184 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2690_
timestamp 1698431365
transform 1 0 8736 0 1 45472
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2691_
timestamp 1698431365
transform -1 0 8624 0 -1 47040
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2692_
timestamp 1698431365
transform -1 0 7952 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2693_
timestamp 1698431365
transform -1 0 8736 0 1 45472
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2694_
timestamp 1698431365
transform -1 0 7168 0 1 45472
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2695_
timestamp 1698431365
transform -1 0 9296 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2696_
timestamp 1698431365
transform -1 0 9184 0 -1 45472
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2697_
timestamp 1698431365
transform -1 0 8176 0 1 45472
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2698_
timestamp 1698431365
transform 1 0 9968 0 1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2699_
timestamp 1698431365
transform -1 0 11424 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2700_
timestamp 1698431365
transform 1 0 9296 0 1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2701_
timestamp 1698431365
transform -1 0 10416 0 -1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2702_
timestamp 1698431365
transform 1 0 9968 0 1 45472
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2703_
timestamp 1698431365
transform 1 0 11424 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2704_
timestamp 1698431365
transform -1 0 11984 0 -1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2705_
timestamp 1698431365
transform 1 0 11088 0 1 47040
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2706_
timestamp 1698431365
transform 1 0 12544 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2707_
timestamp 1698431365
transform -1 0 12208 0 1 51744
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2708_
timestamp 1698431365
transform -1 0 14336 0 1 48608
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2709_
timestamp 1698431365
transform -1 0 13104 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2710_
timestamp 1698431365
transform -1 0 13104 0 1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2711_
timestamp 1698431365
transform -1 0 11648 0 1 50176
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2712_
timestamp 1698431365
transform -1 0 25536 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2713_
timestamp 1698431365
transform 1 0 30352 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2714_
timestamp 1698431365
transform -1 0 32144 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2715_
timestamp 1698431365
transform -1 0 25424 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _2716_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 19264 0 -1 43904
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2717_
timestamp 1698431365
transform 1 0 19264 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2718_
timestamp 1698431365
transform 1 0 21728 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2719_
timestamp 1698431365
transform 1 0 22512 0 -1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2720_
timestamp 1698431365
transform -1 0 25312 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2721_
timestamp 1698431365
transform -1 0 24752 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2722_
timestamp 1698431365
transform 1 0 22960 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2723_
timestamp 1698431365
transform 1 0 22960 0 1 45472
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2724_
timestamp 1698431365
transform -1 0 22848 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2725_
timestamp 1698431365
transform -1 0 22400 0 -1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2726_
timestamp 1698431365
transform 1 0 21728 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2727_
timestamp 1698431365
transform 1 0 21728 0 1 45472
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2728_
timestamp 1698431365
transform 1 0 21280 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2729_
timestamp 1698431365
transform -1 0 22400 0 1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2730_
timestamp 1698431365
transform 1 0 20832 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2731_
timestamp 1698431365
transform 1 0 21392 0 1 47040
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2732_
timestamp 1698431365
transform 1 0 21840 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2733_
timestamp 1698431365
transform -1 0 24864 0 -1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2734_
timestamp 1698431365
transform 1 0 22960 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2735_
timestamp 1698431365
transform 1 0 23632 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2736_
timestamp 1698431365
transform -1 0 23520 0 -1 43904
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2737_
timestamp 1698431365
transform -1 0 27216 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2738_
timestamp 1698431365
transform 1 0 25536 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2739_
timestamp 1698431365
transform -1 0 26432 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2740_
timestamp 1698431365
transform -1 0 26768 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2741_
timestamp 1698431365
transform 1 0 24304 0 -1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2742_
timestamp 1698431365
transform -1 0 25760 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2743_
timestamp 1698431365
transform 1 0 23632 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2744_
timestamp 1698431365
transform 1 0 25088 0 -1 34496
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2745_
timestamp 1698431365
transform 1 0 23408 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2746_
timestamp 1698431365
transform -1 0 25648 0 -1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2747_
timestamp 1698431365
transform 1 0 23856 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2748_
timestamp 1698431365
transform 1 0 23856 0 -1 34496
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2749_
timestamp 1698431365
transform -1 0 26544 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2750_
timestamp 1698431365
transform -1 0 22848 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2751_
timestamp 1698431365
transform 1 0 24528 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2752_
timestamp 1698431365
transform 1 0 25088 0 1 31360
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2753_
timestamp 1698431365
transform -1 0 27104 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2754_
timestamp 1698431365
transform 1 0 24304 0 -1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2755_
timestamp 1698431365
transform 1 0 26208 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2756_
timestamp 1698431365
transform -1 0 26768 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2757_
timestamp 1698431365
transform -1 0 26208 0 -1 29792
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2758_
timestamp 1698431365
transform -1 0 36064 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2759_
timestamp 1698431365
transform 1 0 34384 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2760_
timestamp 1698431365
transform 1 0 31136 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2761_
timestamp 1698431365
transform 1 0 31808 0 1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2762_
timestamp 1698431365
transform -1 0 35952 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2763_
timestamp 1698431365
transform 1 0 33600 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2764_
timestamp 1698431365
transform 1 0 33600 0 -1 40768
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2765_
timestamp 1698431365
transform -1 0 34720 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2766_
timestamp 1698431365
transform 1 0 33040 0 1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2767_
timestamp 1698431365
transform 1 0 32704 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2768_
timestamp 1698431365
transform 1 0 33040 0 -1 36064
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2769_
timestamp 1698431365
transform -1 0 36512 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2770_
timestamp 1698431365
transform -1 0 35616 0 1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2771_
timestamp 1698431365
transform 1 0 34496 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2772_
timestamp 1698431365
transform 1 0 34608 0 -1 40768
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2773_
timestamp 1698431365
transform -1 0 37408 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2774_
timestamp 1698431365
transform 1 0 35616 0 1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2775_
timestamp 1698431365
transform 1 0 37408 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2776_
timestamp 1698431365
transform -1 0 39312 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2777_
timestamp 1698431365
transform -1 0 36624 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2778_
timestamp 1698431365
transform -1 0 36512 0 1 36064
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2779_
timestamp 1698431365
transform -1 0 41216 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2780_
timestamp 1698431365
transform -1 0 43120 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2781_
timestamp 1698431365
transform 1 0 38304 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2782_
timestamp 1698431365
transform 1 0 39984 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2783_
timestamp 1698431365
transform -1 0 40320 0 -1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2784_
timestamp 1698431365
transform 1 0 37520 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2785_
timestamp 1698431365
transform -1 0 39424 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2786_
timestamp 1698431365
transform 1 0 39312 0 -1 36064
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2787_
timestamp 1698431365
transform -1 0 43680 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2788_
timestamp 1698431365
transform 1 0 40768 0 1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2789_
timestamp 1698431365
transform 1 0 40880 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2790_
timestamp 1698431365
transform 1 0 40992 0 1 34496
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2791_
timestamp 1698431365
transform -1 0 44016 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2792_
timestamp 1698431365
transform 1 0 44688 0 1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2793_
timestamp 1698431365
transform 1 0 42112 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2794_
timestamp 1698431365
transform 1 0 42000 0 1 37632
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2795_
timestamp 1698431365
transform -1 0 44464 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2796_
timestamp 1698431365
transform -1 0 44128 0 1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2797_
timestamp 1698431365
transform -1 0 46368 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2798_
timestamp 1698431365
transform -1 0 42672 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2799_
timestamp 1698431365
transform 1 0 42000 0 1 34496
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2800_
timestamp 1698431365
transform -1 0 47040 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2801_
timestamp 1698431365
transform 1 0 45360 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2802_
timestamp 1698431365
transform 1 0 45472 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2803_
timestamp 1698431365
transform -1 0 47040 0 -1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2804_
timestamp 1698431365
transform 1 0 47040 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2805_
timestamp 1698431365
transform 1 0 47152 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2806_
timestamp 1698431365
transform -1 0 47040 0 -1 36064
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2807_
timestamp 1698431365
transform -1 0 50736 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2808_
timestamp 1698431365
transform 1 0 47824 0 1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2809_
timestamp 1698431365
transform -1 0 48944 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2810_
timestamp 1698431365
transform 1 0 48608 0 -1 37632
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2811_
timestamp 1698431365
transform -1 0 48720 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2812_
timestamp 1698431365
transform -1 0 47936 0 -1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2813_
timestamp 1698431365
transform 1 0 46256 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2814_
timestamp 1698431365
transform 1 0 47040 0 1 37632
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2815_
timestamp 1698431365
transform -1 0 51184 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2816_
timestamp 1698431365
transform 1 0 48608 0 1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2817_
timestamp 1698431365
transform 1 0 46816 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2818_
timestamp 1698431365
transform 1 0 47488 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2819_
timestamp 1698431365
transform 1 0 47376 0 -1 36064
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2820_
timestamp 1698431365
transform -1 0 51744 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2821_
timestamp 1698431365
transform 1 0 45136 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2822_
timestamp 1698431365
transform 1 0 45808 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2823_
timestamp 1698431365
transform -1 0 50288 0 1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2824_
timestamp 1698431365
transform -1 0 47040 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2825_
timestamp 1698431365
transform 1 0 49056 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2826_
timestamp 1698431365
transform -1 0 49840 0 -1 39200
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2827_
timestamp 1698431365
transform -1 0 51296 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2828_
timestamp 1698431365
transform -1 0 50848 0 1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2829_
timestamp 1698431365
transform -1 0 47488 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2830_
timestamp 1698431365
transform 1 0 48944 0 -1 42336
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2831_
timestamp 1698431365
transform -1 0 50848 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2832_
timestamp 1698431365
transform -1 0 49728 0 1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2833_
timestamp 1698431365
transform -1 0 49056 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2834_
timestamp 1698431365
transform 1 0 48944 0 1 42336
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2835_
timestamp 1698431365
transform -1 0 47936 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2836_
timestamp 1698431365
transform -1 0 46592 0 1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2837_
timestamp 1698431365
transform -1 0 45360 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2838_
timestamp 1698431365
transform 1 0 45360 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2839_
timestamp 1698431365
transform 1 0 45808 0 1 39200
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2840_
timestamp 1698431365
transform -1 0 41216 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2841_
timestamp 1698431365
transform 1 0 40432 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2842_
timestamp 1698431365
transform -1 0 39872 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2843_
timestamp 1698431365
transform 1 0 39200 0 -1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2844_
timestamp 1698431365
transform -1 0 39872 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2845_
timestamp 1698431365
transform -1 0 40320 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2846_
timestamp 1698431365
transform -1 0 40320 0 -1 40768
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2847_
timestamp 1698431365
transform -1 0 43680 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2848_
timestamp 1698431365
transform 1 0 43008 0 1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2849_
timestamp 1698431365
transform -1 0 42112 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2850_
timestamp 1698431365
transform -1 0 42112 0 1 39200
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2851_
timestamp 1698431365
transform -1 0 43232 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2852_
timestamp 1698431365
transform 1 0 40768 0 -1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2853_
timestamp 1698431365
transform -1 0 41216 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2854_
timestamp 1698431365
transform 1 0 40880 0 -1 42336
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2855_
timestamp 1698431365
transform -1 0 39648 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2856_
timestamp 1698431365
transform -1 0 38976 0 1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2857_
timestamp 1698431365
transform 1 0 36848 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2858_
timestamp 1698431365
transform 1 0 37632 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2859_
timestamp 1698431365
transform 1 0 38304 0 -1 40768
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2860_
timestamp 1698431365
transform -1 0 34160 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2861_
timestamp 1698431365
transform -1 0 32704 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2862_
timestamp 1698431365
transform 1 0 29904 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2863_
timestamp 1698431365
transform 1 0 31248 0 -1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2864_
timestamp 1698431365
transform -1 0 31472 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2865_
timestamp 1698431365
transform 1 0 31024 0 -1 39200
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2866_
timestamp 1698431365
transform -1 0 32032 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2867_
timestamp 1698431365
transform 1 0 30576 0 1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2868_
timestamp 1698431365
transform -1 0 30240 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2869_
timestamp 1698431365
transform 1 0 30576 0 1 39200
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2870_
timestamp 1698431365
transform 1 0 29008 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2871_
timestamp 1698431365
transform -1 0 30688 0 -1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2872_
timestamp 1698431365
transform -1 0 29680 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2873_
timestamp 1698431365
transform 1 0 28896 0 -1 42336
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2874_
timestamp 1698431365
transform 1 0 27440 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2875_
timestamp 1698431365
transform 1 0 29008 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2876_
timestamp 1698431365
transform -1 0 30464 0 1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2877_
timestamp 1698431365
transform 1 0 29008 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2878_
timestamp 1698431365
transform -1 0 18816 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2879_
timestamp 1698431365
transform 1 0 18032 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2880_
timestamp 1698431365
transform -1 0 15904 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2881_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 13552 0 -1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2882_
timestamp 1698431365
transform 1 0 12320 0 -1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2883_
timestamp 1698431365
transform -1 0 20608 0 1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2884_
timestamp 1698431365
transform 1 0 21168 0 -1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2885_
timestamp 1698431365
transform 1 0 15904 0 1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2886_
timestamp 1698431365
transform 1 0 13552 0 1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2887_
timestamp 1698431365
transform -1 0 19824 0 1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2888_
timestamp 1698431365
transform 1 0 13328 0 1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2889_
timestamp 1698431365
transform -1 0 15904 0 -1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2890_
timestamp 1698431365
transform 1 0 13328 0 1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2891_
timestamp 1698431365
transform 1 0 13440 0 -1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2892_
timestamp 1698431365
transform -1 0 17024 0 -1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2893_
timestamp 1698431365
transform 1 0 29456 0 -1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2894_
timestamp 1698431365
transform 1 0 13776 0 -1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2895_
timestamp 1698431365
transform 1 0 17360 0 1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2896_
timestamp 1698431365
transform 1 0 15344 0 1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2897_
timestamp 1698431365
transform 1 0 17248 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2898_
timestamp 1698431365
transform 1 0 18368 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2899_
timestamp 1698431365
transform 1 0 21616 0 -1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2900_
timestamp 1698431365
transform 1 0 22064 0 1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2901_
timestamp 1698431365
transform 1 0 25312 0 1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2902_
timestamp 1698431365
transform 1 0 26880 0 -1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2903_
timestamp 1698431365
transform -1 0 31808 0 -1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2904_
timestamp 1698431365
transform 1 0 30576 0 1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2905_
timestamp 1698431365
transform 1 0 32928 0 1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2906_
timestamp 1698431365
transform 1 0 33376 0 1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2907_
timestamp 1698431365
transform 1 0 36848 0 1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2908_
timestamp 1698431365
transform -1 0 40544 0 -1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2909_
timestamp 1698431365
transform 1 0 39200 0 1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2910_
timestamp 1698431365
transform 1 0 41216 0 1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2911_
timestamp 1698431365
transform 1 0 42112 0 -1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2912_
timestamp 1698431365
transform 1 0 44800 0 1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2913_
timestamp 1698431365
transform 1 0 44688 0 1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2914_
timestamp 1698431365
transform 1 0 43120 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2915_
timestamp 1698431365
transform 1 0 43792 0 -1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2916_
timestamp 1698431365
transform 1 0 44688 0 1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2917_
timestamp 1698431365
transform -1 0 44352 0 1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2918_
timestamp 1698431365
transform -1 0 42224 0 1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2919_
timestamp 1698431365
transform 1 0 37408 0 1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2920_
timestamp 1698431365
transform 1 0 36848 0 1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2921_
timestamp 1698431365
transform -1 0 36624 0 1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2922_
timestamp 1698431365
transform 1 0 31808 0 1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2923_
timestamp 1698431365
transform -1 0 32032 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _2924_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 30464 0 -1 25088
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2925_
timestamp 1698431365
transform -1 0 20272 0 1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2926_
timestamp 1698431365
transform 1 0 17696 0 1 53312
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2927_
timestamp 1698431365
transform 1 0 17248 0 -1 53312
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2928_
timestamp 1698431365
transform 1 0 17360 0 1 61152
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2929_
timestamp 1698431365
transform 1 0 17696 0 1 64288
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2930_
timestamp 1698431365
transform 1 0 19824 0 -1 65856
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2931_
timestamp 1698431365
transform -1 0 22960 0 -1 68992
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2932_
timestamp 1698431365
transform 1 0 21952 0 1 68992
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2933_
timestamp 1698431365
transform 1 0 25200 0 1 68992
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2934_
timestamp 1698431365
transform 1 0 29456 0 1 67424
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2935_
timestamp 1698431365
transform 1 0 27664 0 -1 70560
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2936_
timestamp 1698431365
transform 1 0 31360 0 1 70560
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2937_
timestamp 1698431365
transform 1 0 33040 0 -1 70560
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2938_
timestamp 1698431365
transform 1 0 36288 0 -1 70560
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2939_
timestamp 1698431365
transform -1 0 40096 0 -1 72128
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2940_
timestamp 1698431365
transform 1 0 40768 0 -1 70560
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2941_
timestamp 1698431365
transform 1 0 39536 0 1 68992
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2942_
timestamp 1698431365
transform 1 0 45024 0 1 65856
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2943_
timestamp 1698431365
transform -1 0 47936 0 1 67424
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2944_
timestamp 1698431365
transform -1 0 44464 0 1 67424
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2945_
timestamp 1698431365
transform 1 0 42896 0 -1 64288
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2946_
timestamp 1698431365
transform 1 0 45024 0 1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2947_
timestamp 1698431365
transform 1 0 44016 0 -1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2948_
timestamp 1698431365
transform 1 0 40768 0 -1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2949_
timestamp 1698431365
transform -1 0 44352 0 -1 51744
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2950_
timestamp 1698431365
transform 1 0 33040 0 -1 51744
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2951_
timestamp 1698431365
transform 1 0 36624 0 -1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2952_
timestamp 1698431365
transform 1 0 36848 0 1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2953_
timestamp 1698431365
transform -1 0 34720 0 1 53312
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2954_
timestamp 1698431365
transform 1 0 28784 0 -1 51744
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2955_
timestamp 1698431365
transform 1 0 25536 0 1 51744
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2956_
timestamp 1698431365
transform 1 0 25088 0 -1 51744
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2957_
timestamp 1698431365
transform 1 0 23408 0 1 48608
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2958_
timestamp 1698431365
transform -1 0 15568 0 -1 48608
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2959_
timestamp 1698431365
transform 1 0 14112 0 1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2960_
timestamp 1698431365
transform 1 0 19936 0 -1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2961_
timestamp 1698431365
transform 1 0 18928 0 -1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2962_
timestamp 1698431365
transform 1 0 18928 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2963_
timestamp 1698431365
transform -1 0 23408 0 -1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2964_
timestamp 1698431365
transform 1 0 21168 0 1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2965_
timestamp 1698431365
transform 1 0 21616 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2966_
timestamp 1698431365
transform 1 0 25536 0 1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2967_
timestamp 1698431365
transform -1 0 27440 0 1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2968_
timestamp 1698431365
transform 1 0 28784 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2969_
timestamp 1698431365
transform -1 0 32144 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2970_
timestamp 1698431365
transform 1 0 32480 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2971_
timestamp 1698431365
transform 1 0 31920 0 1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2972_
timestamp 1698431365
transform 1 0 36848 0 1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2973_
timestamp 1698431365
transform 1 0 36960 0 1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2974_
timestamp 1698431365
transform 1 0 39984 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2975_
timestamp 1698431365
transform 1 0 39200 0 1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2976_
timestamp 1698431365
transform 1 0 42896 0 -1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2977_
timestamp 1698431365
transform -1 0 49616 0 1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2978_
timestamp 1698431365
transform 1 0 47712 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2979_
timestamp 1698431365
transform -1 0 51856 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2980_
timestamp 1698431365
transform 1 0 46928 0 1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2981_
timestamp 1698431365
transform -1 0 51632 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2982_
timestamp 1698431365
transform 1 0 47488 0 1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2983_
timestamp 1698431365
transform -1 0 47264 0 -1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2984_
timestamp 1698431365
transform 1 0 37296 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2985_
timestamp 1698431365
transform 1 0 40992 0 1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2986_
timestamp 1698431365
transform 1 0 37296 0 -1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2987_
timestamp 1698431365
transform 1 0 35280 0 -1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2988_
timestamp 1698431365
transform 1 0 32928 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2989_
timestamp 1698431365
transform 1 0 29008 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2990_
timestamp 1698431365
transform 1 0 26432 0 -1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2991_
timestamp 1698431365
transform -1 0 30016 0 -1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2992_
timestamp 1698431365
transform 1 0 21168 0 1 53312
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2993_
timestamp 1698431365
transform 1 0 19152 0 -1 50176
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2994_
timestamp 1698431365
transform 1 0 17472 0 -1 58016
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2995_
timestamp 1698431365
transform -1 0 28336 0 -1 61152
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2996_
timestamp 1698431365
transform 1 0 21616 0 1 58016
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2997_
timestamp 1698431365
transform 1 0 21168 0 1 61152
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2998_
timestamp 1698431365
transform 1 0 22848 0 1 64288
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _2999_
timestamp 1698431365
transform 1 0 26432 0 -1 65856
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3000_
timestamp 1698431365
transform 1 0 31920 0 1 59584
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _3001_
timestamp 1698431365
transform 1 0 28560 0 -1 62720
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3002_
timestamp 1698431365
transform 1 0 31024 0 1 64288
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3003_
timestamp 1698431365
transform -1 0 37632 0 -1 64288
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3004_
timestamp 1698431365
transform 1 0 35504 0 -1 61152
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3005_
timestamp 1698431365
transform -1 0 42448 0 1 56448
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3006_
timestamp 1698431365
transform -1 0 43344 0 1 62720
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _3007_
timestamp 1698431365
transform 1 0 37296 0 1 64288
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3008_
timestamp 1698431365
transform 1 0 47152 0 1 61152
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3009_
timestamp 1698431365
transform 1 0 47040 0 1 58016
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3010_
timestamp 1698431365
transform -1 0 46368 0 -1 61152
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3011_
timestamp 1698431365
transform -1 0 49504 0 1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3012_
timestamp 1698431365
transform -1 0 51856 0 -1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3013_
timestamp 1698431365
transform -1 0 50176 0 1 50176
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3014_
timestamp 1698431365
transform 1 0 45136 0 -1 48608
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3015_
timestamp 1698431365
transform 1 0 42896 0 -1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3016_
timestamp 1698431365
transform 1 0 34496 0 -1 48608
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3017_
timestamp 1698431365
transform 1 0 38304 0 1 50176
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3018_
timestamp 1698431365
transform 1 0 37296 0 -1 47040
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3019_
timestamp 1698431365
transform 1 0 34720 0 -1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3020_
timestamp 1698431365
transform 1 0 29568 0 1 48608
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3021_
timestamp 1698431365
transform 1 0 25424 0 -1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3022_
timestamp 1698431365
transform 1 0 24640 0 1 47040
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3023_
timestamp 1698431365
transform 1 0 24080 0 1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3024_
timestamp 1698431365
transform 1 0 21616 0 -1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3025_
timestamp 1698431365
transform 1 0 26992 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3026_
timestamp 1698431365
transform 1 0 35168 0 -1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3027_
timestamp 1698431365
transform 1 0 42000 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3028_
timestamp 1698431365
transform 1 0 47040 0 1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3029_
timestamp 1698431365
transform -1 0 45472 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3030_
timestamp 1698431365
transform 1 0 32928 0 -1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3031_
timestamp 1698431365
transform 1 0 26432 0 -1 56448
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3032_
timestamp 1698431365
transform 1 0 25536 0 1 56448
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3033_
timestamp 1698431365
transform 1 0 28896 0 -1 59584
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3034_
timestamp 1698431365
transform 1 0 34608 0 -1 59584
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3035_
timestamp 1698431365
transform 1 0 45136 0 -1 62720
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3036_
timestamp 1698431365
transform 1 0 46928 0 1 48608
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3037_
timestamp 1698431365
transform 1 0 40768 0 -1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3038_
timestamp 1698431365
transform 1 0 30352 0 1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3039_
timestamp 1698431365
transform 1 0 17696 0 -1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3040_
timestamp 1698431365
transform 1 0 24640 0 1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3041_
timestamp 1698431365
transform 1 0 19264 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3042_
timestamp 1698431365
transform 1 0 16912 0 1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3043_
timestamp 1698431365
transform 1 0 17696 0 1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3044_
timestamp 1698431365
transform 1 0 17472 0 -1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3045_
timestamp 1698431365
transform 1 0 14224 0 1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3046_
timestamp 1698431365
transform 1 0 13776 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3047_
timestamp 1698431365
transform -1 0 17920 0 1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3048_
timestamp 1698431365
transform 1 0 13328 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3049_
timestamp 1698431365
transform 1 0 10080 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3050_
timestamp 1698431365
transform 1 0 11984 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3051_
timestamp 1698431365
transform -1 0 14672 0 -1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3052_
timestamp 1698431365
transform 1 0 9632 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3053_
timestamp 1698431365
transform 1 0 8176 0 1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3054_
timestamp 1698431365
transform 1 0 6944 0 1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3055_
timestamp 1698431365
transform 1 0 5936 0 -1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3056_
timestamp 1698431365
transform 1 0 5936 0 1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3057_
timestamp 1698431365
transform 1 0 5152 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3058_
timestamp 1698431365
transform 1 0 5376 0 -1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3059_
timestamp 1698431365
transform 1 0 6272 0 1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3060_
timestamp 1698431365
transform -1 0 13104 0 1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3061_
timestamp 1698431365
transform 1 0 11872 0 -1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3062_
timestamp 1698431365
transform 1 0 10864 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3063_
timestamp 1698431365
transform 1 0 8176 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3064_
timestamp 1698431365
transform 1 0 7728 0 1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3065_
timestamp 1698431365
transform 1 0 7728 0 1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3066_
timestamp 1698431365
transform 1 0 8064 0 1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3067_
timestamp 1698431365
transform 1 0 8176 0 1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3068_
timestamp 1698431365
transform 1 0 8288 0 1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3069_
timestamp 1698431365
transform 1 0 8848 0 1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3070_
timestamp 1698431365
transform 1 0 10976 0 -1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3071_
timestamp 1698431365
transform -1 0 19376 0 1 47040
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3072_
timestamp 1698431365
transform 1 0 14448 0 1 48608
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3073_
timestamp 1698431365
transform 1 0 14336 0 1 51744
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3074_
timestamp 1698431365
transform 1 0 12656 0 -1 50176
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3075_
timestamp 1698431365
transform -1 0 16576 0 1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3076_
timestamp 1698431365
transform 1 0 12096 0 -1 56448
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3077_
timestamp 1698431365
transform 1 0 14784 0 1 56448
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3078_
timestamp 1698431365
transform 1 0 13776 0 -1 59584
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3079_
timestamp 1698431365
transform 1 0 14112 0 1 61152
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3080_
timestamp 1698431365
transform 1 0 14448 0 1 64288
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3081_
timestamp 1698431365
transform 1 0 14336 0 1 65856
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3082_
timestamp 1698431365
transform 1 0 12880 0 -1 65856
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3083_
timestamp 1698431365
transform 1 0 9632 0 -1 65856
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3084_
timestamp 1698431365
transform 1 0 9856 0 1 64288
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3085_
timestamp 1698431365
transform 1 0 9408 0 -1 62720
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3086_
timestamp 1698431365
transform 1 0 9408 0 -1 61152
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3087_
timestamp 1698431365
transform 1 0 9408 0 -1 59584
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3088_
timestamp 1698431365
transform 1 0 9408 0 -1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3089_
timestamp 1698431365
transform -1 0 12432 0 1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3090_
timestamp 1698431365
transform 1 0 5936 0 -1 58016
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3091_
timestamp 1698431365
transform 1 0 5488 0 1 56448
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3092_
timestamp 1698431365
transform 1 0 5488 0 1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3093_
timestamp 1698431365
transform 1 0 4368 0 -1 53312
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3094_
timestamp 1698431365
transform 1 0 4368 0 -1 51744
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3095_
timestamp 1698431365
transform 1 0 5488 0 1 48608
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3096_
timestamp 1698431365
transform 1 0 4368 0 -1 47040
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3097_
timestamp 1698431365
transform 1 0 5040 0 -1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3098_
timestamp 1698431365
transform 1 0 5600 0 1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3099_
timestamp 1698431365
transform -1 0 12656 0 -1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3100_
timestamp 1698431365
transform -1 0 12656 0 -1 47040
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3101_
timestamp 1698431365
transform 1 0 9408 0 -1 50176
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3102_
timestamp 1698431365
transform 1 0 9296 0 1 48608
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3103_
timestamp 1698431365
transform -1 0 24864 0 -1 47040
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3104_
timestamp 1698431365
transform -1 0 21616 0 -1 47040
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3105_
timestamp 1698431365
transform -1 0 22512 0 -1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3106_
timestamp 1698431365
transform -1 0 23296 0 -1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3107_
timestamp 1698431365
transform -1 0 26208 0 1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3108_
timestamp 1698431365
transform -1 0 25760 0 1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _3109_
timestamp 1698431365
transform -1 0 26880 0 1 29792
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3110_
timestamp 1698431365
transform 1 0 23744 0 1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3111_
timestamp 1698431365
transform 1 0 33040 0 1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3112_
timestamp 1698431365
transform 1 0 32032 0 1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3113_
timestamp 1698431365
transform 1 0 34048 0 -1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3114_
timestamp 1698431365
transform 1 0 35056 0 -1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3115_
timestamp 1698431365
transform 1 0 37296 0 -1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3116_
timestamp 1698431365
transform 1 0 41328 0 -1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3117_
timestamp 1698431365
transform 1 0 41664 0 -1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3118_
timestamp 1698431365
transform 1 0 41216 0 -1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3119_
timestamp 1698431365
transform 1 0 44912 0 -1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3120_
timestamp 1698431365
transform 1 0 48608 0 -1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3121_
timestamp 1698431365
transform 1 0 46144 0 1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3122_
timestamp 1698431365
transform 1 0 48608 0 -1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3123_
timestamp 1698431365
transform 1 0 48384 0 1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3124_
timestamp 1698431365
transform 1 0 48608 0 -1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3125_
timestamp 1698431365
transform 1 0 48608 0 -1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3126_
timestamp 1698431365
transform 1 0 44688 0 -1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3127_
timestamp 1698431365
transform 1 0 37296 0 1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3128_
timestamp 1698431365
transform 1 0 41104 0 -1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3129_
timestamp 1698431365
transform 1 0 40880 0 1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3130_
timestamp 1698431365
transform 1 0 36960 0 1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3131_
timestamp 1698431365
transform 1 0 30464 0 1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3132_
timestamp 1698431365
transform 1 0 29456 0 1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3133_
timestamp 1698431365
transform -1 0 30576 0 -1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3134_
timestamp 1698431365
transform -1 0 30128 0 -1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _3135_
timestamp 1698431365
transform 1 0 13328 0 1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _3136_
timestamp 1698431365
transform 1 0 32368 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1441__I dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 21616 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1445__I
timestamp 1698431365
transform 1 0 25760 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1451__I
timestamp 1698431365
transform 1 0 11088 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1454__A1
timestamp 1698431365
transform 1 0 12656 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1454__A3
timestamp 1698431365
transform 1 0 11200 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1456__A4
timestamp 1698431365
transform -1 0 10192 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1458__A4
timestamp 1698431365
transform -1 0 9408 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1467__I
timestamp 1698431365
transform 1 0 16128 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1468__B
timestamp 1698431365
transform 1 0 17472 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1473__A2
timestamp 1698431365
transform 1 0 21392 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1476__I
timestamp 1698431365
transform -1 0 25536 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1478__I
timestamp 1698431365
transform 1 0 23184 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1479__I
timestamp 1698431365
transform -1 0 21840 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1480__A2
timestamp 1698431365
transform 1 0 21616 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1482__A1
timestamp 1698431365
transform -1 0 11536 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1484__I
timestamp 1698431365
transform -1 0 19376 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1486__I
timestamp 1698431365
transform 1 0 19600 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1487__A2
timestamp 1698431365
transform 1 0 18032 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1488__A2
timestamp 1698431365
transform 1 0 18480 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1489__A2
timestamp 1698431365
transform 1 0 15568 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1493__I
timestamp 1698431365
transform 1 0 14560 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1497__A1
timestamp 1698431365
transform 1 0 16912 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1504__I
timestamp 1698431365
transform 1 0 22736 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1505__I
timestamp 1698431365
transform 1 0 23744 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1506__I
timestamp 1698431365
transform 1 0 19040 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1507__B
timestamp 1698431365
transform 1 0 18032 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1511__I
timestamp 1698431365
transform 1 0 19376 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1515__I
timestamp 1698431365
transform 1 0 21840 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1517__A1
timestamp 1698431365
transform 1 0 18256 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1517__B1
timestamp 1698431365
transform -1 0 18928 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1519__A1
timestamp 1698431365
transform -1 0 19152 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1519__B1
timestamp 1698431365
transform 1 0 19936 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1521__I
timestamp 1698431365
transform -1 0 18816 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1522__A1
timestamp 1698431365
transform -1 0 19712 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1522__A2
timestamp 1698431365
transform 1 0 23520 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1522__B1
timestamp 1698431365
transform 1 0 23072 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1522__C2
timestamp 1698431365
transform -1 0 19264 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1525__I
timestamp 1698431365
transform 1 0 16576 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1526__I
timestamp 1698431365
transform -1 0 20048 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1527__I
timestamp 1698431365
transform 1 0 21616 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1528__A1
timestamp 1698431365
transform 1 0 20272 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1528__B1
timestamp 1698431365
transform -1 0 23184 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1528__B2
timestamp 1698431365
transform 1 0 20720 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1530__I
timestamp 1698431365
transform -1 0 24304 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1531__A1
timestamp 1698431365
transform -1 0 21616 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1533__A1
timestamp 1698431365
transform 1 0 22960 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1535__I
timestamp 1698431365
transform -1 0 32704 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1540__I
timestamp 1698431365
transform 1 0 29680 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1543__I
timestamp 1698431365
transform 1 0 34160 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1552__I
timestamp 1698431365
transform 1 0 38752 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1555__I
timestamp 1698431365
transform 1 0 36400 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1564__I
timestamp 1698431365
transform -1 0 40768 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1569__B1
timestamp 1698431365
transform 1 0 45696 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1571__B1
timestamp 1698431365
transform 1 0 42560 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1574__A1
timestamp 1698431365
transform -1 0 44464 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1574__B1
timestamp 1698431365
transform -1 0 42672 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1577__I
timestamp 1698431365
transform 1 0 20272 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1578__I
timestamp 1698431365
transform 1 0 41888 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1579__A1
timestamp 1698431365
transform 1 0 45808 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1579__B1
timestamp 1698431365
transform 1 0 42560 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1582__A1
timestamp 1698431365
transform 1 0 43568 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1584__A1
timestamp 1698431365
transform -1 0 46704 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1586__I
timestamp 1698431365
transform 1 0 19824 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1587__I
timestamp 1698431365
transform 1 0 40208 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1591__I
timestamp 1698431365
transform 1 0 40992 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1592__C2
timestamp 1698431365
transform 1 0 44016 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1597__C2
timestamp 1698431365
transform 1 0 40656 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1599__I
timestamp 1698431365
transform 1 0 37968 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1600__C2
timestamp 1698431365
transform 1 0 37856 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1603__I
timestamp 1698431365
transform 1 0 22624 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1604__C2
timestamp 1698431365
transform 1 0 34608 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1607__C2
timestamp 1698431365
transform 1 0 33152 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1609__A2
timestamp 1698431365
transform -1 0 27888 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1613__I
timestamp 1698431365
transform 1 0 21392 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1614__A2
timestamp 1698431365
transform -1 0 19264 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1615__A2
timestamp 1698431365
transform -1 0 20832 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1615__C
timestamp 1698431365
transform 1 0 17472 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1616__A1
timestamp 1698431365
transform 1 0 20048 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1616__A2
timestamp 1698431365
transform 1 0 20496 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1618__I
timestamp 1698431365
transform 1 0 17920 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1620__I
timestamp 1698431365
transform 1 0 29120 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1623__I
timestamp 1698431365
transform -1 0 18928 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1624__I
timestamp 1698431365
transform 1 0 19600 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1625__A2
timestamp 1698431365
transform -1 0 18144 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1626__A1
timestamp 1698431365
transform -1 0 17920 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1630__A1
timestamp 1698431365
transform 1 0 17920 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1633__I
timestamp 1698431365
transform -1 0 23744 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1634__I
timestamp 1698431365
transform 1 0 22624 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1639__I
timestamp 1698431365
transform 1 0 20608 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1644__I
timestamp 1698431365
transform 1 0 23520 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1646__I
timestamp 1698431365
transform 1 0 20720 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1655__I
timestamp 1698431365
transform -1 0 30128 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1661__I
timestamp 1698431365
transform 1 0 19824 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1666__I
timestamp 1698431365
transform -1 0 28112 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1668__I
timestamp 1698431365
transform 1 0 32032 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1683__I
timestamp 1698431365
transform -1 0 35728 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1688__I
timestamp 1698431365
transform -1 0 33376 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1689__I
timestamp 1698431365
transform 1 0 38080 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1691__I
timestamp 1698431365
transform 1 0 35280 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1705__I
timestamp 1698431365
transform 1 0 39648 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1710__I
timestamp 1698431365
transform 1 0 44128 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1712__I
timestamp 1698431365
transform 1 0 30352 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1727__I
timestamp 1698431365
transform 1 0 44576 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1730__A2
timestamp 1698431365
transform -1 0 46032 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1732__I
timestamp 1698431365
transform 1 0 42336 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1735__A2
timestamp 1698431365
transform 1 0 46368 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1748__I
timestamp 1698431365
transform 1 0 40096 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1753__I
timestamp 1698431365
transform 1 0 34048 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1774__I
timestamp 1698431365
transform -1 0 19712 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1791__A1
timestamp 1698431365
transform 1 0 27440 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1796__A1
timestamp 1698431365
transform 1 0 18480 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1799__A1
timestamp 1698431365
transform -1 0 16128 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1802__I
timestamp 1698431365
transform 1 0 24864 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1803__I
timestamp 1698431365
transform 1 0 26880 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1804__A1
timestamp 1698431365
transform 1 0 17472 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1807__I
timestamp 1698431365
transform 1 0 29232 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1810__I
timestamp 1698431365
transform 1 0 28336 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1811__I
timestamp 1698431365
transform 1 0 26768 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1812__A2
timestamp 1698431365
transform -1 0 23408 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1813__I
timestamp 1698431365
transform 1 0 29344 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1815__I
timestamp 1698431365
transform -1 0 29120 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1816__I
timestamp 1698431365
transform 1 0 27888 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1817__A3
timestamp 1698431365
transform 1 0 23520 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1818__A1
timestamp 1698431365
transform 1 0 21952 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1818__B1
timestamp 1698431365
transform 1 0 23408 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1820__I
timestamp 1698431365
transform 1 0 28000 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1822__A1
timestamp 1698431365
transform 1 0 23632 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1823__A2
timestamp 1698431365
transform -1 0 24080 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1826__B
timestamp 1698431365
transform -1 0 23632 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1830__I
timestamp 1698431365
transform 1 0 28560 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1832__A2
timestamp 1698431365
transform -1 0 20944 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1833__I
timestamp 1698431365
transform -1 0 28336 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1834__I
timestamp 1698431365
transform 1 0 25872 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1835__A3
timestamp 1698431365
transform -1 0 23408 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1837__A2
timestamp 1698431365
transform 1 0 26320 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1841__A1
timestamp 1698431365
transform 1 0 28112 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1842__A1
timestamp 1698431365
transform 1 0 24640 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1846__A3
timestamp 1698431365
transform 1 0 27664 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1848__A1
timestamp 1698431365
transform 1 0 25312 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1852__A1
timestamp 1698431365
transform 1 0 21840 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1853__A1
timestamp 1698431365
transform -1 0 21616 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1857__A2
timestamp 1698431365
transform -1 0 23296 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1859__I
timestamp 1698431365
transform 1 0 26768 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1860__A2
timestamp 1698431365
transform 1 0 25312 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1861__A1
timestamp 1698431365
transform 1 0 20720 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1862__I
timestamp 1698431365
transform -1 0 28336 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1866__A2
timestamp 1698431365
transform 1 0 22288 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1869__I
timestamp 1698431365
transform -1 0 29456 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1870__A2
timestamp 1698431365
transform 1 0 26992 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1871__A1
timestamp 1698431365
transform -1 0 24864 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1873__B
timestamp 1698431365
transform -1 0 23968 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1874__A2
timestamp 1698431365
transform 1 0 25312 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1876__I
timestamp 1698431365
transform -1 0 27664 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1877__A1
timestamp 1698431365
transform 1 0 26544 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1877__A3
timestamp 1698431365
transform 1 0 26096 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1880__I
timestamp 1698431365
transform 1 0 28224 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1881__A2
timestamp 1698431365
transform -1 0 29232 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1882__A1
timestamp 1698431365
transform -1 0 27888 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1884__I
timestamp 1698431365
transform 1 0 34048 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1885__I
timestamp 1698431365
transform -1 0 34048 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1887__A2
timestamp 1698431365
transform -1 0 27216 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1890__A1
timestamp 1698431365
transform 1 0 28560 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1890__A3
timestamp 1698431365
transform 1 0 28112 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1892__A3
timestamp 1698431365
transform 1 0 28112 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1893__A2
timestamp 1698431365
transform -1 0 28448 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1900__A1
timestamp 1698431365
transform -1 0 31584 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1901__A2
timestamp 1698431365
transform 1 0 28560 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1903__A2
timestamp 1698431365
transform 1 0 30240 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1904__A1
timestamp 1698431365
transform 1 0 31920 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1905__I
timestamp 1698431365
transform 1 0 33152 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1906__I
timestamp 1698431365
transform 1 0 33600 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1907__A2
timestamp 1698431365
transform 1 0 32256 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1910__A2
timestamp 1698431365
transform 1 0 30016 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1911__A1
timestamp 1698431365
transform 1 0 33152 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1913__A2
timestamp 1698431365
transform 1 0 30240 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1914__A1
timestamp 1698431365
transform -1 0 32480 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1917__A2
timestamp 1698431365
transform -1 0 29680 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1919__A1
timestamp 1698431365
transform -1 0 33376 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1919__A3
timestamp 1698431365
transform 1 0 31808 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1923__A2
timestamp 1698431365
transform 1 0 36736 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1924__A1
timestamp 1698431365
transform -1 0 35392 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1927__A2
timestamp 1698431365
transform 1 0 38416 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1929__A1
timestamp 1698431365
transform -1 0 33488 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1929__A3
timestamp 1698431365
transform 1 0 40208 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1931__I
timestamp 1698431365
transform 1 0 34272 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1932__A1
timestamp 1698431365
transform 1 0 37632 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1932__A3
timestamp 1698431365
transform 1 0 38080 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1934__I
timestamp 1698431365
transform 1 0 35728 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1935__A2
timestamp 1698431365
transform -1 0 33488 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1935__B
timestamp 1698431365
transform -1 0 36960 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1938__I
timestamp 1698431365
transform -1 0 39536 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1940__A2
timestamp 1698431365
transform -1 0 34048 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1942__I
timestamp 1698431365
transform 1 0 27104 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1944__A1
timestamp 1698431365
transform 1 0 40096 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1945__A2
timestamp 1698431365
transform 1 0 37072 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1946__A2
timestamp 1698431365
transform -1 0 36288 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1947__A1
timestamp 1698431365
transform 1 0 39648 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1948__I
timestamp 1698431365
transform 1 0 38976 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1949__A2
timestamp 1698431365
transform 1 0 40320 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1952__A2
timestamp 1698431365
transform 1 0 36288 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1953__A1
timestamp 1698431365
transform 1 0 38640 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1955__A2
timestamp 1698431365
transform -1 0 38192 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1956__A1
timestamp 1698431365
transform 1 0 41440 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1959__A2
timestamp 1698431365
transform 1 0 43456 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1961__A1
timestamp 1698431365
transform -1 0 41216 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1961__A3
timestamp 1698431365
transform 1 0 39648 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1964__A2
timestamp 1698431365
transform -1 0 41216 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1965__A1
timestamp 1698431365
transform -1 0 43120 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1968__A2
timestamp 1698431365
transform -1 0 43568 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1970__I
timestamp 1698431365
transform -1 0 38192 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1971__A1
timestamp 1698431365
transform 1 0 46928 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1971__A3
timestamp 1698431365
transform 1 0 42784 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1973__A1
timestamp 1698431365
transform 1 0 41440 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1973__A3
timestamp 1698431365
transform 1 0 42448 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1974__A2
timestamp 1698431365
transform 1 0 45472 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1974__B
timestamp 1698431365
transform 1 0 43008 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1978__A2
timestamp 1698431365
transform 1 0 43904 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1981__A1
timestamp 1698431365
transform 1 0 47264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1982__A2
timestamp 1698431365
transform -1 0 44128 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1983__I
timestamp 1698431365
transform 1 0 35728 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1984__A2
timestamp 1698431365
transform 1 0 46704 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1985__A1
timestamp 1698431365
transform 1 0 48048 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1986__I
timestamp 1698431365
transform 1 0 46256 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1987__A2
timestamp 1698431365
transform 1 0 47824 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1991__A2
timestamp 1698431365
transform 1 0 45472 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1992__A1
timestamp 1698431365
transform 1 0 49952 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1994__A2
timestamp 1698431365
transform 1 0 43904 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1995__A1
timestamp 1698431365
transform 1 0 49392 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1997__I
timestamp 1698431365
transform 1 0 46480 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1999__A2
timestamp 1698431365
transform 1 0 48832 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2001__A1
timestamp 1698431365
transform -1 0 46704 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2001__A3
timestamp 1698431365
transform -1 0 44464 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2004__A2
timestamp 1698431365
transform 1 0 45584 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2005__A1
timestamp 1698431365
transform -1 0 49952 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2008__A2
timestamp 1698431365
transform 1 0 49728 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2010__A1
timestamp 1698431365
transform 1 0 50400 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2010__A3
timestamp 1698431365
transform 1 0 49728 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2012__A1
timestamp 1698431365
transform 1 0 48272 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2012__A3
timestamp 1698431365
transform -1 0 46480 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2013__A2
timestamp 1698431365
transform 1 0 47376 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2013__B
timestamp 1698431365
transform 1 0 49728 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2017__A2
timestamp 1698431365
transform 1 0 50176 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2021__A2
timestamp 1698431365
transform 1 0 45248 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2022__A2
timestamp 1698431365
transform 1 0 46592 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2023__A1
timestamp 1698431365
transform 1 0 47824 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2024__I
timestamp 1698431365
transform 1 0 47152 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2028__A2
timestamp 1698431365
transform 1 0 46816 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2031__A2
timestamp 1698431365
transform 1 0 45360 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2037__A3
timestamp 1698431365
transform -1 0 46256 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2040__A2
timestamp 1698431365
transform -1 0 47040 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2043__I
timestamp 1698431365
transform -1 0 45248 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2047__A3
timestamp 1698431365
transform 1 0 47824 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2049__A3
timestamp 1698431365
transform 1 0 45696 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2050__A2
timestamp 1698431365
transform -1 0 44464 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2058__A2
timestamp 1698431365
transform 1 0 38304 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2060__A2
timestamp 1698431365
transform -1 0 37408 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2061__A1
timestamp 1698431365
transform 1 0 39088 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2062__I
timestamp 1698431365
transform 1 0 30800 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2063__I
timestamp 1698431365
transform -1 0 34272 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2067__A2
timestamp 1698431365
transform -1 0 41104 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2070__A2
timestamp 1698431365
transform 1 0 39760 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2076__A3
timestamp 1698431365
transform 1 0 41552 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2085__A3
timestamp 1698431365
transform 1 0 38640 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2087__I
timestamp 1698431365
transform 1 0 34720 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2088__A3
timestamp 1698431365
transform 1 0 37632 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2089__I
timestamp 1698431365
transform -1 0 34384 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2090__A2
timestamp 1698431365
transform -1 0 33936 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2093__I
timestamp 1698431365
transform 1 0 30576 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2094__I
timestamp 1698431365
transform 1 0 32592 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2100__A2
timestamp 1698431365
transform -1 0 33376 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2101__A2
timestamp 1698431365
transform -1 0 36400 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2102__A1
timestamp 1698431365
transform 1 0 33600 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2103__I
timestamp 1698431365
transform 1 0 31696 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2107__A2
timestamp 1698431365
transform -1 0 35952 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2110__A2
timestamp 1698431365
transform 1 0 29344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2116__A3
timestamp 1698431365
transform 1 0 32480 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2119__A1
timestamp 1698431365
transform 1 0 28448 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2125__A2
timestamp 1698431365
transform 1 0 28112 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2125__A3
timestamp 1698431365
transform -1 0 26096 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2127__A2
timestamp 1698431365
transform 1 0 27328 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2127__A3
timestamp 1698431365
transform 1 0 29232 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2128__A1
timestamp 1698431365
transform 1 0 26432 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2128__A2
timestamp 1698431365
transform -1 0 27776 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2136__A3
timestamp 1698431365
transform 1 0 25312 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2137__I
timestamp 1698431365
transform -1 0 31920 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2142__A1
timestamp 1698431365
transform 1 0 27888 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2143__I
timestamp 1698431365
transform 1 0 30912 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2146__A1
timestamp 1698431365
transform 1 0 21392 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2147__A3
timestamp 1698431365
transform 1 0 23520 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2149__I
timestamp 1698431365
transform 1 0 29680 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2151__A3
timestamp 1698431365
transform -1 0 23408 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2153__A2
timestamp 1698431365
transform -1 0 19376 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2155__B
timestamp 1698431365
transform 1 0 24192 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2158__I
timestamp 1698431365
transform 1 0 18368 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2160__A1
timestamp 1698431365
transform 1 0 17920 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2163__A3
timestamp 1698431365
transform 1 0 20048 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2164__A2
timestamp 1698431365
transform -1 0 22512 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2167__I
timestamp 1698431365
transform 1 0 31920 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2168__B
timestamp 1698431365
transform -1 0 21616 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2173__A1
timestamp 1698431365
transform 1 0 25200 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2173__A3
timestamp 1698431365
transform 1 0 27888 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2174__A2
timestamp 1698431365
transform 1 0 28448 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2174__B
timestamp 1698431365
transform -1 0 27552 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2177__I
timestamp 1698431365
transform -1 0 31920 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2179__A2
timestamp 1698431365
transform -1 0 26096 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2183__A1
timestamp 1698431365
transform 1 0 22064 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2183__A3
timestamp 1698431365
transform 1 0 25312 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2187__A1
timestamp 1698431365
transform -1 0 25872 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2188__A2
timestamp 1698431365
transform 1 0 23632 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2190__A1
timestamp 1698431365
transform 1 0 21504 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2190__A2
timestamp 1698431365
transform 1 0 22736 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2191__A1
timestamp 1698431365
transform -1 0 21728 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2191__A3
timestamp 1698431365
transform -1 0 22176 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2193__A1
timestamp 1698431365
transform 1 0 25312 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2193__A3
timestamp 1698431365
transform -1 0 21728 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2194__A2
timestamp 1698431365
transform -1 0 22848 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2194__B
timestamp 1698431365
transform -1 0 22288 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2196__B
timestamp 1698431365
transform 1 0 23072 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2199__I
timestamp 1698431365
transform 1 0 23968 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2200__I
timestamp 1698431365
transform 1 0 26432 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2201__A1
timestamp 1698431365
transform 1 0 25984 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2203__A1
timestamp 1698431365
transform -1 0 25760 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2203__A3
timestamp 1698431365
transform -1 0 24528 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2205__A2
timestamp 1698431365
transform -1 0 27104 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2208__B
timestamp 1698431365
transform -1 0 26208 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2213__A1
timestamp 1698431365
transform 1 0 30576 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2213__A3
timestamp 1698431365
transform 1 0 27664 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2214__A2
timestamp 1698431365
transform -1 0 28784 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2214__B
timestamp 1698431365
transform -1 0 29456 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2218__A2
timestamp 1698431365
transform 1 0 30128 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2222__I
timestamp 1698431365
transform 1 0 32480 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2223__A1
timestamp 1698431365
transform -1 0 32816 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2223__A3
timestamp 1698431365
transform -1 0 32704 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2225__A2
timestamp 1698431365
transform 1 0 36176 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2229__A1
timestamp 1698431365
transform 1 0 34048 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2230__I
timestamp 1698431365
transform 1 0 35616 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2231__A2
timestamp 1698431365
transform 1 0 36064 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2233__A1
timestamp 1698431365
transform -1 0 28000 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2233__A2
timestamp 1698431365
transform 1 0 29568 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2235__A1
timestamp 1698431365
transform 1 0 35616 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2235__A3
timestamp 1698431365
transform 1 0 36064 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2237__A1
timestamp 1698431365
transform 1 0 32256 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2237__A3
timestamp 1698431365
transform 1 0 29680 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2238__A2
timestamp 1698431365
transform 1 0 31472 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2238__B
timestamp 1698431365
transform 1 0 31024 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2240__B
timestamp 1698431365
transform 1 0 34720 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2243__I
timestamp 1698431365
transform -1 0 34496 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2244__A1
timestamp 1698431365
transform -1 0 32032 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2246__A1
timestamp 1698431365
transform 1 0 35168 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2246__A3
timestamp 1698431365
transform 1 0 35168 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2247__A2
timestamp 1698431365
transform 1 0 34496 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2250__B
timestamp 1698431365
transform 1 0 32704 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2255__I
timestamp 1698431365
transform 1 0 36400 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2256__A1
timestamp 1698431365
transform -1 0 37296 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2256__A3
timestamp 1698431365
transform -1 0 36848 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2257__I
timestamp 1698431365
transform 1 0 38864 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2258__A2
timestamp 1698431365
transform 1 0 38864 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2258__B
timestamp 1698431365
transform 1 0 38080 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2262__A2
timestamp 1698431365
transform 1 0 37632 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2266__A1
timestamp 1698431365
transform 1 0 40992 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2266__A3
timestamp 1698431365
transform -1 0 37408 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2267__A2
timestamp 1698431365
transform -1 0 37408 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2270__A1
timestamp 1698431365
transform 1 0 38752 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2271__A2
timestamp 1698431365
transform 1 0 40320 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2273__I
timestamp 1698431365
transform 1 0 38080 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2274__A1
timestamp 1698431365
transform -1 0 40096 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2275__A1
timestamp 1698431365
transform 1 0 41440 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2275__A3
timestamp 1698431365
transform 1 0 40992 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2283__B
timestamp 1698431365
transform 1 0 40992 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2286__I
timestamp 1698431365
transform 1 0 43120 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2287__A1
timestamp 1698431365
transform 1 0 42672 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2290__A1
timestamp 1698431365
transform -1 0 39200 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2290__A3
timestamp 1698431365
transform 1 0 43568 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2291__A2
timestamp 1698431365
transform 1 0 42560 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2294__B
timestamp 1698431365
transform 1 0 39424 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2299__A1
timestamp 1698431365
transform 1 0 42112 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2299__A3
timestamp 1698431365
transform 1 0 43008 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2300__A2
timestamp 1698431365
transform -1 0 41888 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2300__B
timestamp 1698431365
transform 1 0 40320 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2304__A2
timestamp 1698431365
transform -1 0 40320 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2308__A1
timestamp 1698431365
transform 1 0 49840 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2308__A3
timestamp 1698431365
transform 1 0 49728 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2309__A2
timestamp 1698431365
transform 1 0 50288 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2312__A1
timestamp 1698431365
transform -1 0 46928 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2314__I
timestamp 1698431365
transform 1 0 44912 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2315__A1
timestamp 1698431365
transform 1 0 49392 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2315__A2
timestamp 1698431365
transform 1 0 50288 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2317__A1
timestamp 1698431365
transform 1 0 49728 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2317__A2
timestamp 1698431365
transform 1 0 49280 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2318__A1
timestamp 1698431365
transform 1 0 50176 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2318__A3
timestamp 1698431365
transform 1 0 46928 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2320__A1
timestamp 1698431365
transform 1 0 48832 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2321__B
timestamp 1698431365
transform 1 0 45808 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2323__B
timestamp 1698431365
transform 1 0 46704 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2326__I
timestamp 1698431365
transform 1 0 46032 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2327__A1
timestamp 1698431365
transform 1 0 41664 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2329__A1
timestamp 1698431365
transform -1 0 43120 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2329__A3
timestamp 1698431365
transform 1 0 42336 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2330__A2
timestamp 1698431365
transform 1 0 43120 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2333__B
timestamp 1698431365
transform -1 0 44464 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2338__A2
timestamp 1698431365
transform 1 0 48272 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2338__A3
timestamp 1698431365
transform 1 0 44912 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2339__A1
timestamp 1698431365
transform 1 0 44800 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2339__A2
timestamp 1698431365
transform 1 0 42896 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2342__I
timestamp 1698431365
transform 1 0 33152 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2343__B
timestamp 1698431365
transform -1 0 45584 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2344__A1
timestamp 1698431365
transform 1 0 48720 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2348__A3
timestamp 1698431365
transform 1 0 48720 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2349__A2
timestamp 1698431365
transform 1 0 47264 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2352__A1
timestamp 1698431365
transform 1 0 45360 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2353__A1
timestamp 1698431365
transform 1 0 50848 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2355__A1
timestamp 1698431365
transform 1 0 46704 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2356__A3
timestamp 1698431365
transform -1 0 47040 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2361__B
timestamp 1698431365
transform 1 0 49728 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2365__A1
timestamp 1698431365
transform 1 0 41104 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2367__A3
timestamp 1698431365
transform -1 0 42560 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2371__B
timestamp 1698431365
transform 1 0 43120 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2376__A3
timestamp 1698431365
transform 1 0 42896 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2377__A2
timestamp 1698431365
transform 1 0 44352 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2380__B
timestamp 1698431365
transform 1 0 45808 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2381__A1
timestamp 1698431365
transform 1 0 46368 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2385__A3
timestamp 1698431365
transform -1 0 35952 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2386__A2
timestamp 1698431365
transform 1 0 37184 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2389__A1
timestamp 1698431365
transform 1 0 34720 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2390__I
timestamp 1698431365
transform 1 0 34048 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2393__A1
timestamp 1698431365
transform 1 0 42336 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2394__A3
timestamp 1698431365
transform 1 0 35616 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2399__B
timestamp 1698431365
transform -1 0 38304 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2403__A1
timestamp 1698431365
transform 1 0 42224 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2405__A3
timestamp 1698431365
transform 1 0 38640 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2409__B
timestamp 1698431365
transform 1 0 40208 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2414__A3
timestamp 1698431365
transform -1 0 34720 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2415__A2
timestamp 1698431365
transform 1 0 36736 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2418__B
timestamp 1698431365
transform -1 0 34496 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2423__A3
timestamp 1698431365
transform 1 0 32480 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2427__A1
timestamp 1698431365
transform 1 0 29568 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2430__A1
timestamp 1698431365
transform 1 0 27664 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2433__A3
timestamp 1698431365
transform 1 0 29232 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2437__B
timestamp 1698431365
transform -1 0 26544 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2444__B
timestamp 1698431365
transform 1 0 29232 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2447__A3
timestamp 1698431365
transform 1 0 28672 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2449__A1
timestamp 1698431365
transform -1 0 27328 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2451__I
timestamp 1698431365
transform -1 0 30800 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2452__A1
timestamp 1698431365
transform 1 0 24864 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2453__A1
timestamp 1698431365
transform 1 0 24416 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2456__A1
timestamp 1698431365
transform 1 0 25312 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2457__A1
timestamp 1698431365
transform 1 0 22176 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2459__A1
timestamp 1698431365
transform 1 0 31472 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2460__A1
timestamp 1698431365
transform 1 0 28560 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2463__A1
timestamp 1698431365
transform 1 0 38528 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2464__A1
timestamp 1698431365
transform 1 0 37072 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2466__I
timestamp 1698431365
transform -1 0 43120 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2467__A1
timestamp 1698431365
transform 1 0 46032 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2468__A1
timestamp 1698431365
transform -1 0 43680 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2470__A1
timestamp 1698431365
transform 1 0 47264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2471__A1
timestamp 1698431365
transform 1 0 48832 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2473__A1
timestamp 1698431365
transform 1 0 43904 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2474__A1
timestamp 1698431365
transform -1 0 43568 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2475__I
timestamp 1698431365
transform 1 0 35168 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2477__A1
timestamp 1698431365
transform 1 0 36960 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2478__A1
timestamp 1698431365
transform 1 0 36288 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2481__B1
timestamp 1698431365
transform 1 0 30688 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2481__B2
timestamp 1698431365
transform 1 0 29904 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2483__B1
timestamp 1698431365
transform -1 0 28896 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2485__B1
timestamp 1698431365
transform 1 0 31360 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2486__I
timestamp 1698431365
transform 1 0 34384 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2488__B1
timestamp 1698431365
transform 1 0 35728 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2491__A1
timestamp 1698431365
transform -1 0 44464 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2491__B1
timestamp 1698431365
transform 1 0 46368 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2493__A1
timestamp 1698431365
transform 1 0 45360 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2493__B1
timestamp 1698431365
transform 1 0 45808 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2495__A1
timestamp 1698431365
transform 1 0 41776 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2495__B1
timestamp 1698431365
transform 1 0 41440 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2498__A1
timestamp 1698431365
transform -1 0 32368 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2498__B1
timestamp 1698431365
transform -1 0 31024 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2500__B1
timestamp 1698431365
transform 1 0 20720 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2502__I
timestamp 1698431365
transform 1 0 19824 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2503__A2
timestamp 1698431365
transform 1 0 25760 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2503__C2
timestamp 1698431365
transform 1 0 25312 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2505__I
timestamp 1698431365
transform -1 0 18592 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2506__B2
timestamp 1698431365
transform 1 0 20720 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2506__C2
timestamp 1698431365
transform 1 0 21392 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2508__B2
timestamp 1698431365
transform -1 0 20496 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2510__I
timestamp 1698431365
transform 1 0 20048 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2513__I
timestamp 1698431365
transform 1 0 17920 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2516__I
timestamp 1698431365
transform -1 0 15568 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2522__I
timestamp 1698431365
transform 1 0 13664 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2525__I
timestamp 1698431365
transform -1 0 14448 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2532__C2
timestamp 1698431365
transform 1 0 16352 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2534__I
timestamp 1698431365
transform -1 0 12208 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2563__I
timestamp 1698431365
transform 1 0 12320 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2571__I
timestamp 1698431365
transform -1 0 12208 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2574__I
timestamp 1698431365
transform -1 0 13776 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2582__A1
timestamp 1698431365
transform 1 0 12880 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2584__A1
timestamp 1698431365
transform 1 0 18480 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2586__A1
timestamp 1698431365
transform 1 0 14000 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2588__I
timestamp 1698431365
transform -1 0 13104 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2591__I
timestamp 1698431365
transform -1 0 17696 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2593__B
timestamp 1698431365
transform -1 0 17024 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2596__I
timestamp 1698431365
transform 1 0 17472 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2611__I
timestamp 1698431365
transform 1 0 17920 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2626__I
timestamp 1698431365
transform 1 0 17920 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2651__I
timestamp 1698431365
transform -1 0 12656 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2712__I
timestamp 1698431365
transform 1 0 25760 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2717__I
timestamp 1698431365
transform 1 0 19040 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2724__I
timestamp 1698431365
transform 1 0 22848 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2728__I
timestamp 1698431365
transform 1 0 22064 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2732__I
timestamp 1698431365
transform 1 0 20720 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2735__A1
timestamp 1698431365
transform -1 0 24080 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2737__I
timestamp 1698431365
transform 1 0 26544 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2739__I
timestamp 1698431365
transform 1 0 26880 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2743__A1
timestamp 1698431365
transform -1 0 23856 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2745__I
timestamp 1698431365
transform 1 0 23184 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2746__A1
timestamp 1698431365
transform -1 0 24304 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2747__A1
timestamp 1698431365
transform 1 0 25312 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2749__I
timestamp 1698431365
transform -1 0 24640 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2750__A1
timestamp 1698431365
transform -1 0 20944 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2751__A1
timestamp 1698431365
transform -1 0 26208 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2753__I
timestamp 1698431365
transform 1 0 28560 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2756__A1
timestamp 1698431365
transform -1 0 25872 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2758__I
timestamp 1698431365
transform -1 0 36960 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2759__I
timestamp 1698431365
transform -1 0 35504 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2761__A1
timestamp 1698431365
transform 1 0 32368 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2763__A1
timestamp 1698431365
transform 1 0 34496 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2765__I
timestamp 1698431365
transform -1 0 36624 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2766__A1
timestamp 1698431365
transform 1 0 33824 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2767__A1
timestamp 1698431365
transform 1 0 32480 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2769__I
timestamp 1698431365
transform 1 0 37184 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2770__A1
timestamp 1698431365
transform -1 0 38304 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2771__A1
timestamp 1698431365
transform -1 0 34496 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2773__I
timestamp 1698431365
transform 1 0 38080 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2774__A1
timestamp 1698431365
transform 1 0 37632 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2775__I
timestamp 1698431365
transform -1 0 37408 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2777__A1
timestamp 1698431365
transform -1 0 36400 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2779__I
timestamp 1698431365
transform -1 0 41216 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2780__I
timestamp 1698431365
transform 1 0 41440 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2781__I
timestamp 1698431365
transform 1 0 38752 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2783__A1
timestamp 1698431365
transform 1 0 39536 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2785__A1
timestamp 1698431365
transform 1 0 39536 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2788__A1
timestamp 1698431365
transform -1 0 40768 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2792__A1
timestamp 1698431365
transform 1 0 44800 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2793__A1
timestamp 1698431365
transform -1 0 42336 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2796__A1
timestamp 1698431365
transform 1 0 43344 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2798__A1
timestamp 1698431365
transform 1 0 41552 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2801__I
timestamp 1698431365
transform 1 0 45136 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2803__A1
timestamp 1698431365
transform 1 0 45584 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2805__A1
timestamp 1698431365
transform 1 0 50176 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2808__A1
timestamp 1698431365
transform -1 0 47824 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2809__A1
timestamp 1698431365
transform -1 0 48160 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2812__A1
timestamp 1698431365
transform 1 0 48160 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2813__A1
timestamp 1698431365
transform 1 0 46368 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2816__A1
timestamp 1698431365
transform 1 0 49168 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2857__I
timestamp 1698431365
transform -1 0 36848 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2860__I
timestamp 1698431365
transform -1 0 33712 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2862__I
timestamp 1698431365
transform 1 0 28560 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2866__I
timestamp 1698431365
transform -1 0 32480 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2870__I
timestamp 1698431365
transform -1 0 28784 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2876__A1
timestamp 1698431365
transform 1 0 30800 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3005__CLK
timestamp 1698431365
transform 1 0 40320 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__3136__I
timestamp 1698431365
transform -1 0 33376 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_clk_I
timestamp 1698431365
transform 1 0 26432 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_2_0__f_clk_I
timestamp 1698431365
transform 1 0 27216 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_2_1__f_clk_I
timestamp 1698431365
transform 1 0 36176 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_2_2__f_clk_I
timestamp 1698431365
transform -1 0 26432 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_2_3__f_clk_I
timestamp 1698431365
transform 1 0 34944 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_0_clk_I
timestamp 1698431365
transform 1 0 15120 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_1_clk_I
timestamp 1698431365
transform 1 0 17696 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_2_clk_I
timestamp 1698431365
transform 1 0 14336 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_3_clk_I
timestamp 1698431365
transform 1 0 17696 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_4_clk_I
timestamp 1698431365
transform 1 0 23072 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_5_clk_I
timestamp 1698431365
transform 1 0 27440 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_6_clk_I
timestamp 1698431365
transform 1 0 25312 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_7_clk_I
timestamp 1698431365
transform 1 0 23632 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_8_clk_I
timestamp 1698431365
transform -1 0 22736 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_9_clk_I
timestamp 1698431365
transform 1 0 11088 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_10_clk_I
timestamp 1698431365
transform 1 0 16912 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_11_clk_I
timestamp 1698431365
transform 1 0 17472 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_12_clk_I
timestamp 1698431365
transform 1 0 12656 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_13_clk_I
timestamp 1698431365
transform 1 0 19152 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_14_clk_I
timestamp 1698431365
transform 1 0 24640 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_15_clk_I
timestamp 1698431365
transform -1 0 25536 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_16_clk_I
timestamp 1698431365
transform 1 0 24080 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_17_clk_I
timestamp 1698431365
transform 1 0 23072 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_18_clk_I
timestamp 1698431365
transform 1 0 24416 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_19_clk_I
timestamp 1698431365
transform 1 0 35840 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_20_clk_I
timestamp 1698431365
transform 1 0 40320 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_21_clk_I
timestamp 1698431365
transform 1 0 36512 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_22_clk_I
timestamp 1698431365
transform 1 0 42672 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_23_clk_I
timestamp 1698431365
transform 1 0 43008 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_25_clk_I
timestamp 1698431365
transform 1 0 43568 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_26_clk_I
timestamp 1698431365
transform 1 0 40208 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_27_clk_I
timestamp 1698431365
transform 1 0 49392 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_28_clk_I
timestamp 1698431365
transform 1 0 44240 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_29_clk_I
timestamp 1698431365
transform 1 0 49280 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_30_clk_I
timestamp 1698431365
transform -1 0 45248 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_31_clk_I
timestamp 1698431365
transform 1 0 43344 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_32_clk_I
timestamp 1698431365
transform -1 0 38976 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_33_clk_I
timestamp 1698431365
transform 1 0 43232 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_34_clk_I
timestamp 1698431365
transform 1 0 40320 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_35_clk_I
timestamp 1698431365
transform 1 0 44688 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_36_clk_I
timestamp 1698431365
transform 1 0 48832 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_37_clk_I
timestamp 1698431365
transform 1 0 47264 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_38_clk_I
timestamp 1698431365
transform 1 0 50400 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_39_clk_I
timestamp 1698431365
transform 1 0 41888 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_40_clk_I
timestamp 1698431365
transform 1 0 42672 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_41_clk_I
timestamp 1698431365
transform 1 0 39200 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_42_clk_I
timestamp 1698431365
transform 1 0 35840 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_43_clk_I
timestamp 1698431365
transform 1 0 38752 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_44_clk_I
timestamp 1698431365
transform 1 0 35168 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_45_clk_I
timestamp 1698431365
transform 1 0 23968 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_46_clk_I
timestamp 1698431365
transform 1 0 27664 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_47_clk_I
timestamp 1698431365
transform 1 0 24752 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_48_clk_I
timestamp 1698431365
transform -1 0 22736 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_leaf_49_clk_I
timestamp 1698431365
transform 1 0 22848 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input1_I
timestamp 1698431365
transform 1 0 2464 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input2_I
timestamp 1698431365
transform 1 0 2464 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input3_I
timestamp 1698431365
transform 1 0 2912 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input4_I
timestamp 1698431365
transform 1 0 3136 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input5_I
timestamp 1698431365
transform 1 0 2464 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input6_I
timestamp 1698431365
transform 1 0 2464 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input7_I
timestamp 1698431365
transform 1 0 3136 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input8_I
timestamp 1698431365
transform 1 0 2464 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input9_I
timestamp 1698431365
transform 1 0 2464 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input10_I
timestamp 1698431365
transform 1 0 2464 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input11_I
timestamp 1698431365
transform 1 0 2464 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input12_I
timestamp 1698431365
transform 1 0 2464 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input13_I
timestamp 1698431365
transform 1 0 2464 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input14_I
timestamp 1698431365
transform 1 0 2464 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input15_I
timestamp 1698431365
transform 1 0 2464 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input16_I
timestamp 1698431365
transform 1 0 3136 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input17_I
timestamp 1698431365
transform 1 0 2912 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input18_I
timestamp 1698431365
transform 1 0 2912 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input19_I
timestamp 1698431365
transform -1 0 24416 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input20_I
timestamp 1698431365
transform -1 0 12768 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input21_I
timestamp 1698431365
transform 1 0 1792 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input22_I
timestamp 1698431365
transform 1 0 3136 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input23_I
timestamp 1698431365
transform 1 0 2464 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input24_I
timestamp 1698431365
transform 1 0 2464 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input25_I
timestamp 1698431365
transform 1 0 2464 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input26_I
timestamp 1698431365
transform 1 0 2464 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input27_I
timestamp 1698431365
transform 1 0 2464 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input28_I
timestamp 1698431365
transform 1 0 2464 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input29_I
timestamp 1698431365
transform 1 0 2464 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input30_I
timestamp 1698431365
transform 1 0 21840 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input31_I
timestamp 1698431365
transform 1 0 2464 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input32_I
timestamp 1698431365
transform 1 0 3136 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input33_I
timestamp 1698431365
transform 1 0 2464 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input34_I
timestamp 1698431365
transform 1 0 2912 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input35_I
timestamp 1698431365
transform 1 0 3136 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input36_I
timestamp 1698431365
transform 1 0 2464 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input37_I
timestamp 1698431365
transform 1 0 2464 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input38_I
timestamp 1698431365
transform 1 0 2464 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input39_I
timestamp 1698431365
transform 1 0 2464 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input40_I
timestamp 1698431365
transform 1 0 2464 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input41_I
timestamp 1698431365
transform 1 0 19712 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input42_I
timestamp 1698431365
transform 1 0 3136 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input43_I
timestamp 1698431365
transform 1 0 2464 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input44_I
timestamp 1698431365
transform 1 0 19040 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input45_I
timestamp 1698431365
transform 1 0 18368 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input46_I
timestamp 1698431365
transform -1 0 16912 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input47_I
timestamp 1698431365
transform -1 0 15904 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input48_I
timestamp 1698431365
transform 1 0 2912 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input49_I
timestamp 1698431365
transform 1 0 3136 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input50_I
timestamp 1698431365
transform 1 0 2464 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input51_I
timestamp 1698431365
transform 1 0 2464 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input52_I
timestamp 1698431365
transform -1 0 31472 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input53_I
timestamp 1698431365
transform -1 0 33040 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input54_I
timestamp 1698431365
transform -1 0 34384 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input55_I
timestamp 1698431365
transform -1 0 36512 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input56_I
timestamp 1698431365
transform -1 0 38528 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input57_I
timestamp 1698431365
transform -1 0 39760 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input58_I
timestamp 1698431365
transform -1 0 41216 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input59_I
timestamp 1698431365
transform -1 0 42448 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input60_I
timestamp 1698431365
transform -1 0 43456 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input61_I
timestamp 1698431365
transform -1 0 44128 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input62_I
timestamp 1698431365
transform 1 0 2464 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input63_I
timestamp 1698431365
transform -1 0 57680 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input64_I
timestamp 1698431365
transform -1 0 57680 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input65_I
timestamp 1698431365
transform -1 0 57680 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input66_I
timestamp 1698431365
transform -1 0 57680 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input67_I
timestamp 1698431365
transform -1 0 40432 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input68_I
timestamp 1698431365
transform -1 0 37856 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input69_I
timestamp 1698431365
transform -1 0 37184 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input70_I
timestamp 1698431365
transform -1 0 35616 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input71_I
timestamp 1698431365
transform -1 0 33712 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input72_I
timestamp 1698431365
transform -1 0 30352 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input73_I
timestamp 1698431365
transform 1 0 2464 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input74_I
timestamp 1698431365
transform -1 0 28784 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input75_I
timestamp 1698431365
transform 1 0 2464 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input76_I
timestamp 1698431365
transform 1 0 2912 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input77_I
timestamp 1698431365
transform -1 0 20944 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input78_I
timestamp 1698431365
transform 1 0 23520 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input79_I
timestamp 1698431365
transform 1 0 24640 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input80_I
timestamp 1698431365
transform -1 0 25648 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input81_I
timestamp 1698431365
transform -1 0 26880 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input82_I
timestamp 1698431365
transform -1 0 29680 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input83_I
timestamp 1698431365
transform 1 0 2912 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output84_I
timestamp 1698431365
transform 1 0 4704 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output85_I
timestamp 1698431365
transform -1 0 53312 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output86_I
timestamp 1698431365
transform -1 0 53312 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output87_I
timestamp 1698431365
transform -1 0 55440 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output95_I
timestamp 1698431365
transform -1 0 4928 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output104_I
timestamp 1698431365
transform -1 0 53312 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output105_I
timestamp 1698431365
transform -1 0 55440 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output106_I
timestamp 1698431365
transform 1 0 4704 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output107_I
timestamp 1698431365
transform -1 0 53312 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output108_I
timestamp 1698431365
transform -1 0 4928 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output109_I
timestamp 1698431365
transform -1 0 4928 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output110_I
timestamp 1698431365
transform -1 0 4928 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output111_I
timestamp 1698431365
transform 1 0 4704 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output112_I
timestamp 1698431365
transform -1 0 27328 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output113_I
timestamp 1698431365
transform -1 0 26992 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output114_I
timestamp 1698431365
transform -1 0 55440 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output115_I
timestamp 1698431365
transform 1 0 52080 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output116_I
timestamp 1698431365
transform -1 0 53312 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output118_I
timestamp 1698431365
transform -1 0 55440 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_clk dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 27104 0 -1 40768
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_2_0__f_clk
timestamp 1698431365
transform -1 0 26768 0 1 25088
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_2_1__f_clk
timestamp 1698431365
transform 1 0 34944 0 -1 25088
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_2_2__f_clk
timestamp 1698431365
transform -1 0 26768 0 1 54880
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_2_3__f_clk
timestamp 1698431365
transform 1 0 34496 0 -1 56448
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_0_clk
timestamp 1698431365
transform -1 0 15008 0 -1 20384
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_1_clk
timestamp 1698431365
transform -1 0 18928 0 1 23520
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_2_clk
timestamp 1698431365
transform -1 0 12992 0 1 28224
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_3_clk
timestamp 1698431365
transform -1 0 17024 0 -1 37632
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_4_clk
timestamp 1698431365
transform -1 0 22848 0 -1 29792
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_5_clk
timestamp 1698431365
transform -1 0 27216 0 1 39200
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_6_clk
timestamp 1698431365
transform -1 0 24864 0 -1 45472
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_7_clk
timestamp 1698431365
transform -1 0 20384 0 1 50176
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_8_clk
timestamp 1698431365
transform -1 0 19264 0 1 43904
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_9_clk
timestamp 1698431365
transform -1 0 11088 0 1 47040
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_10_clk
timestamp 1698431365
transform -1 0 16016 0 -1 51744
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_11_clk
timestamp 1698431365
transform 1 0 11200 0 -1 58016
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_12_clk
timestamp 1698431365
transform -1 0 12432 0 1 58016
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_13_clk
timestamp 1698431365
transform -1 0 18928 0 1 62720
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_14_clk
timestamp 1698431365
transform -1 0 24416 0 -1 62720
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_15_clk
timestamp 1698431365
transform 1 0 25088 0 -1 68992
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_16_clk
timestamp 1698431365
transform 1 0 25088 0 -1 58016
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_17_clk
timestamp 1698431365
transform -1 0 24192 0 -1 54880
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_18_clk
timestamp 1698431365
transform 1 0 25088 0 -1 48608
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_19_clk
timestamp 1698431365
transform -1 0 34832 0 1 45472
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_20_clk
timestamp 1698431365
transform -1 0 40096 0 -1 58016
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_21_clk
timestamp 1698431365
transform -1 0 34944 0 1 62720
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_22_clk
timestamp 1698431365
transform -1 0 42448 0 1 70560
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_23_clk
timestamp 1698431365
transform -1 0 40544 0 -1 65856
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_25_clk
timestamp 1698431365
transform -1 0 50288 0 1 62720
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_26_clk
timestamp 1698431365
transform -1 0 47488 0 -1 68992
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_27_clk
timestamp 1698431365
transform 1 0 48608 0 -1 62720
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_28_clk
timestamp 1698431365
transform -1 0 50288 0 1 51744
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_29_clk
timestamp 1698431365
transform 1 0 49504 0 -1 50176
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_30_clk
timestamp 1698431365
transform -1 0 50848 0 1 40768
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_31_clk
timestamp 1698431365
transform -1 0 43008 0 1 45472
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_32_clk
timestamp 1698431365
transform -1 0 38528 0 -1 39200
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_33_clk
timestamp 1698431365
transform -1 0 42448 0 1 36064
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_34_clk
timestamp 1698431365
transform -1 0 46368 0 -1 29792
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_35_clk
timestamp 1698431365
transform 1 0 44688 0 1 36064
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_36_clk
timestamp 1698431365
transform 1 0 48608 0 -1 31360
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_37_clk
timestamp 1698431365
transform -1 0 50288 0 1 23520
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_38_clk
timestamp 1698431365
transform 1 0 50624 0 -1 15680
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_39_clk
timestamp 1698431365
transform -1 0 48160 0 -1 10976
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_40_clk
timestamp 1698431365
transform -1 0 44464 0 1 15680
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_41_clk
timestamp 1698431365
transform -1 0 38528 0 -1 9408
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_42_clk
timestamp 1698431365
transform -1 0 35840 0 1 15680
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_43_clk
timestamp 1698431365
transform 1 0 33376 0 -1 23520
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_44_clk
timestamp 1698431365
transform -1 0 35168 0 1 31360
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_45_clk
timestamp 1698431365
transform 1 0 25088 0 -1 31360
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_46_clk
timestamp 1698431365
transform -1 0 26768 0 1 21952
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_47_clk
timestamp 1698431365
transform 1 0 25536 0 -1 20384
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_48_clk
timestamp 1698431365
transform 1 0 23184 0 1 10976
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_leaf_49_clk
timestamp 1698431365
transform -1 0 22848 0 -1 17248
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1568 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_36
timestamp 1698431365
transform 1 0 5376 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_70 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 9184 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_86 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 10976 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_94 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 11872 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_98 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 12320 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_110
timestamp 1698431365
transform 1 0 13664 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_126
timestamp 1698431365
transform 1 0 15456 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_138 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 16800 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_145
timestamp 1698431365
transform 1 0 17584 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_172
timestamp 1698431365
transform 1 0 20608 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_174
timestamp 1698431365
transform 1 0 20832 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_181
timestamp 1698431365
transform 1 0 21616 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_185
timestamp 1698431365
transform 1 0 22064 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_189
timestamp 1698431365
transform 1 0 22512 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_191
timestamp 1698431365
transform 1 0 22736 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_212
timestamp 1698431365
transform 1 0 25088 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_214
timestamp 1698431365
transform 1 0 25312 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_223
timestamp 1698431365
transform 1 0 26320 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_225
timestamp 1698431365
transform 1 0 26544 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_228
timestamp 1698431365
transform 1 0 26880 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_274
timestamp 1698431365
transform 1 0 32032 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_278
timestamp 1698431365
transform 1 0 32480 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_280
timestamp 1698431365
transform 1 0 32704 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_301
timestamp 1698431365
transform 1 0 35056 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_303
timestamp 1698431365
transform 1 0 35280 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_338
timestamp 1698431365
transform 1 0 39200 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_342
timestamp 1698431365
transform 1 0 39648 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_361
timestamp 1698431365
transform 1 0 41776 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_373
timestamp 1698431365
transform 1 0 43120 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_388
timestamp 1698431365
transform 1 0 44800 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_404
timestamp 1698431365
transform 1 0 46592 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_410
timestamp 1698431365
transform 1 0 47264 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_444
timestamp 1698431365
transform 1 0 51072 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_478
timestamp 1698431365
transform 1 0 54880 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_494
timestamp 1698431365
transform 1 0 56672 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_502
timestamp 1698431365
transform 1 0 57568 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_506
timestamp 1698431365
transform 1 0 58016 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_508
timestamp 1698431365
transform 1 0 58240 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1568 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_66
timestamp 1698431365
transform 1 0 8736 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_72
timestamp 1698431365
transform 1 0 9408 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_136
timestamp 1698431365
transform 1 0 16576 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_139
timestamp 1698431365
transform 1 0 16912 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_142
timestamp 1698431365
transform 1 0 17248 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_150
timestamp 1698431365
transform 1 0 18144 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_154
timestamp 1698431365
transform 1 0 18592 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_160
timestamp 1698431365
transform 1 0 19264 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_166
timestamp 1698431365
transform 1 0 19936 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_170
timestamp 1698431365
transform 1 0 20384 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_172
timestamp 1698431365
transform 1 0 20608 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_175
timestamp 1698431365
transform 1 0 20944 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_191
timestamp 1698431365
transform 1 0 22736 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_195
timestamp 1698431365
transform 1 0 23184 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_197
timestamp 1698431365
transform 1 0 23408 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_200
timestamp 1698431365
transform 1 0 23744 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_206
timestamp 1698431365
transform 1 0 24416 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_212
timestamp 1698431365
transform 1 0 25088 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_220
timestamp 1698431365
transform 1 0 25984 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_224
timestamp 1698431365
transform 1 0 26432 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_226
timestamp 1698431365
transform 1 0 26656 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_255
timestamp 1698431365
transform 1 0 29904 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_265
timestamp 1698431365
transform 1 0 31024 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_269
timestamp 1698431365
transform 1 0 31472 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_277
timestamp 1698431365
transform 1 0 32368 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_279
timestamp 1698431365
transform 1 0 32592 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_282
timestamp 1698431365
transform 1 0 32928 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_286
timestamp 1698431365
transform 1 0 33376 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_289
timestamp 1698431365
transform 1 0 33712 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_295
timestamp 1698431365
transform 1 0 34384 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_311
timestamp 1698431365
transform 1 0 36176 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_314
timestamp 1698431365
transform 1 0 36512 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_320
timestamp 1698431365
transform 1 0 37184 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_326
timestamp 1698431365
transform 1 0 37856 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_332
timestamp 1698431365
transform 1 0 38528 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_340
timestamp 1698431365
transform 1 0 39424 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_343
timestamp 1698431365
transform 1 0 39760 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_349
timestamp 1698431365
transform 1 0 40432 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_352
timestamp 1698431365
transform 1 0 40768 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_356
timestamp 1698431365
transform 1 0 41216 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_372
timestamp 1698431365
transform 1 0 43008 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_376
timestamp 1698431365
transform 1 0 43456 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_1_382
timestamp 1698431365
transform 1 0 44128 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_414
timestamp 1698431365
transform 1 0 47712 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_418
timestamp 1698431365
transform 1 0 48160 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_422
timestamp 1698431365
transform 1 0 48608 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_486
timestamp 1698431365
transform 1 0 55776 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_492
timestamp 1698431365
transform 1 0 56448 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_508
timestamp 1698431365
transform 1 0 58240 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_2
timestamp 1698431365
transform 1 0 1568 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_34
timestamp 1698431365
transform 1 0 5152 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_37
timestamp 1698431365
transform 1 0 5488 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_101
timestamp 1698431365
transform 1 0 12656 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_107
timestamp 1698431365
transform 1 0 13328 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_171
timestamp 1698431365
transform 1 0 20496 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_177
timestamp 1698431365
transform 1 0 21168 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_241
timestamp 1698431365
transform 1 0 28336 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_259
timestamp 1698431365
transform 1 0 30352 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_291
timestamp 1698431365
transform 1 0 33936 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_307
timestamp 1698431365
transform 1 0 35728 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_317
timestamp 1698431365
transform 1 0 36848 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_381
timestamp 1698431365
transform 1 0 44016 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_387
timestamp 1698431365
transform 1 0 44688 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_451
timestamp 1698431365
transform 1 0 51856 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_457
timestamp 1698431365
transform 1 0 52528 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_489
timestamp 1698431365
transform 1 0 56112 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_505
timestamp 1698431365
transform 1 0 57904 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_2
timestamp 1698431365
transform 1 0 1568 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_66
timestamp 1698431365
transform 1 0 8736 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_72
timestamp 1698431365
transform 1 0 9408 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_136
timestamp 1698431365
transform 1 0 16576 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_142
timestamp 1698431365
transform 1 0 17248 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_206
timestamp 1698431365
transform 1 0 24416 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_3_212
timestamp 1698431365
transform 1 0 25088 0 -1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_244
timestamp 1698431365
transform 1 0 28672 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_248
timestamp 1698431365
transform 1 0 29120 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_250
timestamp 1698431365
transform 1 0 29344 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_253
timestamp 1698431365
transform 1 0 29680 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_269
timestamp 1698431365
transform 1 0 31472 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_277
timestamp 1698431365
transform 1 0 32368 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_279
timestamp 1698431365
transform 1 0 32592 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_282
timestamp 1698431365
transform 1 0 32928 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_346
timestamp 1698431365
transform 1 0 40096 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_352
timestamp 1698431365
transform 1 0 40768 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_397
timestamp 1698431365
transform 1 0 45808 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_413
timestamp 1698431365
transform 1 0 47600 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_417
timestamp 1698431365
transform 1 0 48048 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_419
timestamp 1698431365
transform 1 0 48272 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_422
timestamp 1698431365
transform 1 0 48608 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_486
timestamp 1698431365
transform 1 0 55776 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_492
timestamp 1698431365
transform 1 0 56448 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_508
timestamp 1698431365
transform 1 0 58240 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_2
timestamp 1698431365
transform 1 0 1568 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_34
timestamp 1698431365
transform 1 0 5152 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_37
timestamp 1698431365
transform 1 0 5488 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_101
timestamp 1698431365
transform 1 0 12656 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_107
timestamp 1698431365
transform 1 0 13328 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_171
timestamp 1698431365
transform 1 0 20496 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_177
timestamp 1698431365
transform 1 0 21168 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_241
timestamp 1698431365
transform 1 0 28336 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_247
timestamp 1698431365
transform 1 0 29008 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_311
timestamp 1698431365
transform 1 0 36176 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_317
timestamp 1698431365
transform 1 0 36848 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_381
timestamp 1698431365
transform 1 0 44016 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_387
timestamp 1698431365
transform 1 0 44688 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_451
timestamp 1698431365
transform 1 0 51856 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_457
timestamp 1698431365
transform 1 0 52528 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_4_489
timestamp 1698431365
transform 1 0 56112 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_505
timestamp 1698431365
transform 1 0 57904 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_2
timestamp 1698431365
transform 1 0 1568 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_66
timestamp 1698431365
transform 1 0 8736 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_72
timestamp 1698431365
transform 1 0 9408 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_136
timestamp 1698431365
transform 1 0 16576 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_142
timestamp 1698431365
transform 1 0 17248 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_206
timestamp 1698431365
transform 1 0 24416 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_212
timestamp 1698431365
transform 1 0 25088 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_276
timestamp 1698431365
transform 1 0 32256 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_5_282
timestamp 1698431365
transform 1 0 32928 0 -1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_314
timestamp 1698431365
transform 1 0 36512 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_318
timestamp 1698431365
transform 1 0 36960 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_320
timestamp 1698431365
transform 1 0 37184 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_352
timestamp 1698431365
transform 1 0 40768 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_360
timestamp 1698431365
transform 1 0 41664 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_362
timestamp 1698431365
transform 1 0 41888 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_394
timestamp 1698431365
transform 1 0 45472 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_5_398
timestamp 1698431365
transform 1 0 45920 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_414
timestamp 1698431365
transform 1 0 47712 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_418
timestamp 1698431365
transform 1 0 48160 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_422
timestamp 1698431365
transform 1 0 48608 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_486
timestamp 1698431365
transform 1 0 55776 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_5_492
timestamp 1698431365
transform 1 0 56448 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_508
timestamp 1698431365
transform 1 0 58240 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_2
timestamp 1698431365
transform 1 0 1568 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_34
timestamp 1698431365
transform 1 0 5152 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_37
timestamp 1698431365
transform 1 0 5488 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_101
timestamp 1698431365
transform 1 0 12656 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_107
timestamp 1698431365
transform 1 0 13328 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_171
timestamp 1698431365
transform 1 0 20496 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_177
timestamp 1698431365
transform 1 0 21168 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_193
timestamp 1698431365
transform 1 0 22960 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_201
timestamp 1698431365
transform 1 0 23856 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_205
timestamp 1698431365
transform 1 0 24304 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_221
timestamp 1698431365
transform 1 0 26096 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_227
timestamp 1698431365
transform 1 0 26768 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_235
timestamp 1698431365
transform 1 0 27664 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_241
timestamp 1698431365
transform 1 0 28336 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_247
timestamp 1698431365
transform 1 0 29008 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_255
timestamp 1698431365
transform 1 0 29904 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_259
timestamp 1698431365
transform 1 0 30352 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_294
timestamp 1698431365
transform 1 0 34272 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_310
timestamp 1698431365
transform 1 0 36064 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_346
timestamp 1698431365
transform 1 0 40096 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_352
timestamp 1698431365
transform 1 0 40768 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_356
timestamp 1698431365
transform 1 0 41216 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_387
timestamp 1698431365
transform 1 0 44688 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_417
timestamp 1698431365
transform 1 0 48048 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_449
timestamp 1698431365
transform 1 0 51632 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_453
timestamp 1698431365
transform 1 0 52080 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_457
timestamp 1698431365
transform 1 0 52528 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_489
timestamp 1698431365
transform 1 0 56112 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_505
timestamp 1698431365
transform 1 0 57904 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_2
timestamp 1698431365
transform 1 0 1568 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_66
timestamp 1698431365
transform 1 0 8736 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_72
timestamp 1698431365
transform 1 0 9408 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_136
timestamp 1698431365
transform 1 0 16576 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_7_142
timestamp 1698431365
transform 1 0 17248 0 -1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_174
timestamp 1698431365
transform 1 0 20832 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_190
timestamp 1698431365
transform 1 0 22624 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_203
timestamp 1698431365
transform 1 0 24080 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_209
timestamp 1698431365
transform 1 0 24752 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_212
timestamp 1698431365
transform 1 0 25088 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_240
timestamp 1698431365
transform 1 0 28224 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_242
timestamp 1698431365
transform 1 0 28448 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_272
timestamp 1698431365
transform 1 0 31808 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_276
timestamp 1698431365
transform 1 0 32256 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_332
timestamp 1698431365
transform 1 0 38528 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_336
timestamp 1698431365
transform 1 0 38976 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_344
timestamp 1698431365
transform 1 0 39872 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_360
timestamp 1698431365
transform 1 0 41664 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_401
timestamp 1698431365
transform 1 0 46256 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_405
timestamp 1698431365
transform 1 0 46704 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_413
timestamp 1698431365
transform 1 0 47600 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_417
timestamp 1698431365
transform 1 0 48048 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_419
timestamp 1698431365
transform 1 0 48272 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_422
timestamp 1698431365
transform 1 0 48608 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_486
timestamp 1698431365
transform 1 0 55776 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_492
timestamp 1698431365
transform 1 0 56448 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_508
timestamp 1698431365
transform 1 0 58240 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_2
timestamp 1698431365
transform 1 0 1568 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_34
timestamp 1698431365
transform 1 0 5152 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_37
timestamp 1698431365
transform 1 0 5488 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_101
timestamp 1698431365
transform 1 0 12656 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_107
timestamp 1698431365
transform 1 0 13328 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_171
timestamp 1698431365
transform 1 0 20496 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_177
timestamp 1698431365
transform 1 0 21168 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_183
timestamp 1698431365
transform 1 0 21840 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_243
timestamp 1698431365
transform 1 0 28560 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_247
timestamp 1698431365
transform 1 0 29008 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_251
timestamp 1698431365
transform 1 0 29456 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_311
timestamp 1698431365
transform 1 0 36176 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_325
timestamp 1698431365
transform 1 0 37744 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_329
timestamp 1698431365
transform 1 0 38192 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_375
timestamp 1698431365
transform 1 0 43344 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_416
timestamp 1698431365
transform 1 0 47936 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_448
timestamp 1698431365
transform 1 0 51520 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_452
timestamp 1698431365
transform 1 0 51968 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_454
timestamp 1698431365
transform 1 0 52192 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_457
timestamp 1698431365
transform 1 0 52528 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_489
timestamp 1698431365
transform 1 0 56112 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_505
timestamp 1698431365
transform 1 0 57904 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_2
timestamp 1698431365
transform 1 0 1568 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_66
timestamp 1698431365
transform 1 0 8736 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_72
timestamp 1698431365
transform 1 0 9408 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_136
timestamp 1698431365
transform 1 0 16576 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_9_142
timestamp 1698431365
transform 1 0 17248 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_158
timestamp 1698431365
transform 1 0 19040 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_166
timestamp 1698431365
transform 1 0 19936 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_170
timestamp 1698431365
transform 1 0 20384 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_172
timestamp 1698431365
transform 1 0 20608 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_9_212
timestamp 1698431365
transform 1 0 25088 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_265
timestamp 1698431365
transform 1 0 31024 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_267
timestamp 1698431365
transform 1 0 31248 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_336
timestamp 1698431365
transform 1 0 38976 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_340
timestamp 1698431365
transform 1 0 39424 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_344
timestamp 1698431365
transform 1 0 39872 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_348
timestamp 1698431365
transform 1 0 40320 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_352
timestamp 1698431365
transform 1 0 40768 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_356
timestamp 1698431365
transform 1 0 41216 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_360
timestamp 1698431365
transform 1 0 41664 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_418
timestamp 1698431365
transform 1 0 48160 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_422
timestamp 1698431365
transform 1 0 48608 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_486
timestamp 1698431365
transform 1 0 55776 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_9_492
timestamp 1698431365
transform 1 0 56448 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_508
timestamp 1698431365
transform 1 0 58240 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_2
timestamp 1698431365
transform 1 0 1568 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_34
timestamp 1698431365
transform 1 0 5152 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_37
timestamp 1698431365
transform 1 0 5488 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_101
timestamp 1698431365
transform 1 0 12656 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_107
timestamp 1698431365
transform 1 0 13328 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_139
timestamp 1698431365
transform 1 0 16912 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_147
timestamp 1698431365
transform 1 0 17808 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_177
timestamp 1698431365
transform 1 0 21168 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_181
timestamp 1698431365
transform 1 0 21616 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_191
timestamp 1698431365
transform 1 0 22736 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_247
timestamp 1698431365
transform 1 0 29008 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_351
timestamp 1698431365
transform 1 0 40656 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_379
timestamp 1698431365
transform 1 0 43792 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_387
timestamp 1698431365
transform 1 0 44688 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_395
timestamp 1698431365
transform 1 0 45584 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_397
timestamp 1698431365
transform 1 0 45808 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_431
timestamp 1698431365
transform 1 0 49616 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_447
timestamp 1698431365
transform 1 0 51408 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_457
timestamp 1698431365
transform 1 0 52528 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_489
timestamp 1698431365
transform 1 0 56112 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_505
timestamp 1698431365
transform 1 0 57904 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_2
timestamp 1698431365
transform 1 0 1568 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_66
timestamp 1698431365
transform 1 0 8736 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_72
timestamp 1698431365
transform 1 0 9408 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_136
timestamp 1698431365
transform 1 0 16576 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_142
timestamp 1698431365
transform 1 0 17248 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_158
timestamp 1698431365
transform 1 0 19040 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_162
timestamp 1698431365
transform 1 0 19488 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_164
timestamp 1698431365
transform 1 0 19712 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_167
timestamp 1698431365
transform 1 0 20048 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_204
timestamp 1698431365
transform 1 0 24192 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_219
timestamp 1698431365
transform 1 0 25872 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_223
timestamp 1698431365
transform 1 0 26320 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_227
timestamp 1698431365
transform 1 0 26768 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_229
timestamp 1698431365
transform 1 0 26992 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_270
timestamp 1698431365
transform 1 0 31584 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_274
timestamp 1698431365
transform 1 0 32032 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_278
timestamp 1698431365
transform 1 0 32480 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_282
timestamp 1698431365
transform 1 0 32928 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_294
timestamp 1698431365
transform 1 0 34272 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_296
timestamp 1698431365
transform 1 0 34496 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_345
timestamp 1698431365
transform 1 0 39984 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_349
timestamp 1698431365
transform 1 0 40432 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_352
timestamp 1698431365
transform 1 0 40768 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_356
timestamp 1698431365
transform 1 0 41216 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_360
timestamp 1698431365
transform 1 0 41664 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_364
timestamp 1698431365
transform 1 0 42112 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_366
timestamp 1698431365
transform 1 0 42336 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_377
timestamp 1698431365
transform 1 0 43568 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_379
timestamp 1698431365
transform 1 0 43792 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_419
timestamp 1698431365
transform 1 0 48272 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_422
timestamp 1698431365
transform 1 0 48608 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_426
timestamp 1698431365
transform 1 0 49056 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_492
timestamp 1698431365
transform 1 0 56448 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_508
timestamp 1698431365
transform 1 0 58240 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_2
timestamp 1698431365
transform 1 0 1568 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_34
timestamp 1698431365
transform 1 0 5152 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_37
timestamp 1698431365
transform 1 0 5488 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_101
timestamp 1698431365
transform 1 0 12656 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_107
timestamp 1698431365
transform 1 0 13328 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_171
timestamp 1698431365
transform 1 0 20496 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_177
timestamp 1698431365
transform 1 0 21168 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_227
timestamp 1698431365
transform 1 0 26768 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_231
timestamp 1698431365
transform 1 0 27216 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_235
timestamp 1698431365
transform 1 0 27664 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_241
timestamp 1698431365
transform 1 0 28336 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_247
timestamp 1698431365
transform 1 0 29008 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_251
timestamp 1698431365
transform 1 0 29456 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_255
timestamp 1698431365
transform 1 0 29904 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_257
timestamp 1698431365
transform 1 0 30128 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_280
timestamp 1698431365
transform 1 0 32704 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_282
timestamp 1698431365
transform 1 0 32928 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_291
timestamp 1698431365
transform 1 0 33936 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_295
timestamp 1698431365
transform 1 0 34384 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_300
timestamp 1698431365
transform 1 0 34944 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_304
timestamp 1698431365
transform 1 0 35392 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_306
timestamp 1698431365
transform 1 0 35616 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_317
timestamp 1698431365
transform 1 0 36848 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_387
timestamp 1698431365
transform 1 0 44688 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_389
timestamp 1698431365
transform 1 0 44912 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_427
timestamp 1698431365
transform 1 0 49168 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_431
timestamp 1698431365
transform 1 0 49616 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_447
timestamp 1698431365
transform 1 0 51408 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_457
timestamp 1698431365
transform 1 0 52528 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_489
timestamp 1698431365
transform 1 0 56112 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_505
timestamp 1698431365
transform 1 0 57904 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_2
timestamp 1698431365
transform 1 0 1568 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_66
timestamp 1698431365
transform 1 0 8736 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_72
timestamp 1698431365
transform 1 0 9408 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_136
timestamp 1698431365
transform 1 0 16576 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_142
timestamp 1698431365
transform 1 0 17248 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_150
timestamp 1698431365
transform 1 0 18144 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_225
timestamp 1698431365
transform 1 0 26544 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_245
timestamp 1698431365
transform 1 0 28784 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_279
timestamp 1698431365
transform 1 0 32592 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_282
timestamp 1698431365
transform 1 0 32928 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_284
timestamp 1698431365
transform 1 0 33152 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_304
timestamp 1698431365
transform 1 0 35392 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_310
timestamp 1698431365
transform 1 0 36064 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_314
timestamp 1698431365
transform 1 0 36512 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_318
timestamp 1698431365
transform 1 0 36960 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_341
timestamp 1698431365
transform 1 0 39536 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_369
timestamp 1698431365
transform 1 0 42672 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_373
timestamp 1698431365
transform 1 0 43120 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_377
timestamp 1698431365
transform 1 0 43568 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_387
timestamp 1698431365
transform 1 0 44688 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_418
timestamp 1698431365
transform 1 0 48160 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_430
timestamp 1698431365
transform 1 0 49504 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_13_434
timestamp 1698431365
transform 1 0 49952 0 -1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_466
timestamp 1698431365
transform 1 0 53536 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_482
timestamp 1698431365
transform 1 0 55328 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_492
timestamp 1698431365
transform 1 0 56448 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_508
timestamp 1698431365
transform 1 0 58240 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_2
timestamp 1698431365
transform 1 0 1568 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_34
timestamp 1698431365
transform 1 0 5152 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_37
timestamp 1698431365
transform 1 0 5488 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_69
timestamp 1698431365
transform 1 0 9072 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_71
timestamp 1698431365
transform 1 0 9296 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_99
timestamp 1698431365
transform 1 0 12432 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_103
timestamp 1698431365
transform 1 0 12880 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_107
timestamp 1698431365
transform 1 0 13328 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_139
timestamp 1698431365
transform 1 0 16912 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_174
timestamp 1698431365
transform 1 0 20832 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_197
timestamp 1698431365
transform 1 0 23408 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_199
timestamp 1698431365
transform 1 0 23632 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_227
timestamp 1698431365
transform 1 0 26768 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_231
timestamp 1698431365
transform 1 0 27216 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_237
timestamp 1698431365
transform 1 0 27888 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_241
timestamp 1698431365
transform 1 0 28336 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_247
timestamp 1698431365
transform 1 0 29008 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_307
timestamp 1698431365
transform 1 0 35728 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_309
timestamp 1698431365
transform 1 0 35952 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_374
timestamp 1698431365
transform 1 0 43232 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_378
timestamp 1698431365
transform 1 0 43680 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_382
timestamp 1698431365
transform 1 0 44128 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_384
timestamp 1698431365
transform 1 0 44352 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_392
timestamp 1698431365
transform 1 0 45248 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_396
timestamp 1698431365
transform 1 0 45696 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_443
timestamp 1698431365
transform 1 0 50960 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_451
timestamp 1698431365
transform 1 0 51856 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_457
timestamp 1698431365
transform 1 0 52528 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_489
timestamp 1698431365
transform 1 0 56112 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_505
timestamp 1698431365
transform 1 0 57904 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_2
timestamp 1698431365
transform 1 0 1568 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_66
timestamp 1698431365
transform 1 0 8736 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_72
timestamp 1698431365
transform 1 0 9408 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_88
timestamp 1698431365
transform 1 0 11200 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_119
timestamp 1698431365
transform 1 0 14672 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_127
timestamp 1698431365
transform 1 0 15568 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_131
timestamp 1698431365
transform 1 0 16016 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_133
timestamp 1698431365
transform 1 0 16240 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_142
timestamp 1698431365
transform 1 0 17248 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_173
timestamp 1698431365
transform 1 0 20720 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_181
timestamp 1698431365
transform 1 0 21616 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_185
timestamp 1698431365
transform 1 0 22064 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_217
timestamp 1698431365
transform 1 0 25648 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_245
timestamp 1698431365
transform 1 0 28784 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_249
timestamp 1698431365
transform 1 0 29232 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_273
timestamp 1698431365
transform 1 0 31920 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_279
timestamp 1698431365
transform 1 0 32592 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_314
timestamp 1698431365
transform 1 0 36512 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_318
timestamp 1698431365
transform 1 0 36960 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_340
timestamp 1698431365
transform 1 0 39424 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_367
timestamp 1698431365
transform 1 0 42448 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_415
timestamp 1698431365
transform 1 0 47824 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_419
timestamp 1698431365
transform 1 0 48272 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_430
timestamp 1698431365
transform 1 0 49504 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_434
timestamp 1698431365
transform 1 0 49952 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_492
timestamp 1698431365
transform 1 0 56448 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_508
timestamp 1698431365
transform 1 0 58240 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_2
timestamp 1698431365
transform 1 0 1568 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_6
timestamp 1698431365
transform 1 0 2016 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_22
timestamp 1698431365
transform 1 0 3808 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_30
timestamp 1698431365
transform 1 0 4704 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_34
timestamp 1698431365
transform 1 0 5152 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_37
timestamp 1698431365
transform 1 0 5488 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_53
timestamp 1698431365
transform 1 0 7280 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_90
timestamp 1698431365
transform 1 0 11424 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_98
timestamp 1698431365
transform 1 0 12320 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_104
timestamp 1698431365
transform 1 0 12992 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_107
timestamp 1698431365
transform 1 0 13328 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_144
timestamp 1698431365
transform 1 0 17472 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_177
timestamp 1698431365
transform 1 0 21168 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_185
timestamp 1698431365
transform 1 0 22064 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_189
timestamp 1698431365
transform 1 0 22512 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_191
timestamp 1698431365
transform 1 0 22736 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_194
timestamp 1698431365
transform 1 0 23072 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_196
timestamp 1698431365
transform 1 0 23296 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_212
timestamp 1698431365
transform 1 0 25088 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_252
timestamp 1698431365
transform 1 0 29568 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_308
timestamp 1698431365
transform 1 0 35840 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_312
timestamp 1698431365
transform 1 0 36288 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_314
timestamp 1698431365
transform 1 0 36512 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_317
timestamp 1698431365
transform 1 0 36848 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_321
timestamp 1698431365
transform 1 0 37296 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_323
timestamp 1698431365
transform 1 0 37520 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_329
timestamp 1698431365
transform 1 0 38192 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_333
timestamp 1698431365
transform 1 0 38640 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_408
timestamp 1698431365
transform 1 0 47040 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_432
timestamp 1698431365
transform 1 0 49728 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_436
timestamp 1698431365
transform 1 0 50176 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_440
timestamp 1698431365
transform 1 0 50624 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_448
timestamp 1698431365
transform 1 0 51520 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_452
timestamp 1698431365
transform 1 0 51968 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_454
timestamp 1698431365
transform 1 0 52192 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_457
timestamp 1698431365
transform 1 0 52528 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_489
timestamp 1698431365
transform 1 0 56112 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_505
timestamp 1698431365
transform 1 0 57904 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_8
timestamp 1698431365
transform 1 0 2240 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_12
timestamp 1698431365
transform 1 0 2688 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_44
timestamp 1698431365
transform 1 0 6272 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_60
timestamp 1698431365
transform 1 0 8064 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_64
timestamp 1698431365
transform 1 0 8512 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_72
timestamp 1698431365
transform 1 0 9408 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_103
timestamp 1698431365
transform 1 0 12880 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_105
timestamp 1698431365
transform 1 0 13104 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_110
timestamp 1698431365
transform 1 0 13664 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_192
timestamp 1698431365
transform 1 0 22848 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_196
timestamp 1698431365
transform 1 0 23296 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_208
timestamp 1698431365
transform 1 0 24640 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_217
timestamp 1698431365
transform 1 0 25648 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_248
timestamp 1698431365
transform 1 0 29120 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_256
timestamp 1698431365
transform 1 0 30016 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_266
timestamp 1698431365
transform 1 0 31136 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_270
timestamp 1698431365
transform 1 0 31584 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_277
timestamp 1698431365
transform 1 0 32368 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_279
timestamp 1698431365
transform 1 0 32592 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_282
timestamp 1698431365
transform 1 0 32928 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_286
timestamp 1698431365
transform 1 0 33376 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_305
timestamp 1698431365
transform 1 0 35504 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_309
timestamp 1698431365
transform 1 0 35952 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_311
timestamp 1698431365
transform 1 0 36176 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_340
timestamp 1698431365
transform 1 0 39424 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_344
timestamp 1698431365
transform 1 0 39872 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_348
timestamp 1698431365
transform 1 0 40320 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_359
timestamp 1698431365
transform 1 0 41552 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_368
timestamp 1698431365
transform 1 0 42560 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_372
timestamp 1698431365
transform 1 0 43008 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_405
timestamp 1698431365
transform 1 0 46704 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_409
timestamp 1698431365
transform 1 0 47152 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_413
timestamp 1698431365
transform 1 0 47600 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_417
timestamp 1698431365
transform 1 0 48048 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_419
timestamp 1698431365
transform 1 0 48272 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_430
timestamp 1698431365
transform 1 0 49504 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_434
timestamp 1698431365
transform 1 0 49952 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_466
timestamp 1698431365
transform 1 0 53536 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_482
timestamp 1698431365
transform 1 0 55328 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_492
timestamp 1698431365
transform 1 0 56448 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_508
timestamp 1698431365
transform 1 0 58240 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_14
timestamp 1698431365
transform 1 0 2912 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_18
timestamp 1698431365
transform 1 0 3360 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_34
timestamp 1698431365
transform 1 0 5152 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_37
timestamp 1698431365
transform 1 0 5488 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_45
timestamp 1698431365
transform 1 0 6384 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_49
timestamp 1698431365
transform 1 0 6832 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_79
timestamp 1698431365
transform 1 0 10192 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_83
timestamp 1698431365
transform 1 0 10640 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_89
timestamp 1698431365
transform 1 0 11312 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_93
timestamp 1698431365
transform 1 0 11760 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_165
timestamp 1698431365
transform 1 0 19824 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_169
timestamp 1698431365
transform 1 0 20272 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_173
timestamp 1698431365
transform 1 0 20720 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_212
timestamp 1698431365
transform 1 0 25088 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_216
timestamp 1698431365
transform 1 0 25536 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_232
timestamp 1698431365
transform 1 0 27328 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_242
timestamp 1698431365
transform 1 0 28448 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_244
timestamp 1698431365
transform 1 0 28672 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_247
timestamp 1698431365
transform 1 0 29008 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_251
timestamp 1698431365
transform 1 0 29456 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_286
timestamp 1698431365
transform 1 0 33376 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_295
timestamp 1698431365
transform 1 0 34384 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_305
timestamp 1698431365
transform 1 0 35504 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_346
timestamp 1698431365
transform 1 0 40096 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_363
timestamp 1698431365
transform 1 0 42000 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_367
timestamp 1698431365
transform 1 0 42448 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_370
timestamp 1698431365
transform 1 0 42784 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_374
timestamp 1698431365
transform 1 0 43232 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_378
timestamp 1698431365
transform 1 0 43680 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_382
timestamp 1698431365
transform 1 0 44128 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_384
timestamp 1698431365
transform 1 0 44352 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_399
timestamp 1698431365
transform 1 0 46032 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_403
timestamp 1698431365
transform 1 0 46480 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_407
timestamp 1698431365
transform 1 0 46928 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_430
timestamp 1698431365
transform 1 0 49504 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_434
timestamp 1698431365
transform 1 0 49952 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_438
timestamp 1698431365
transform 1 0 50400 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_454
timestamp 1698431365
transform 1 0 52192 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_457
timestamp 1698431365
transform 1 0 52528 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_489
timestamp 1698431365
transform 1 0 56112 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_505
timestamp 1698431365
transform 1 0 57904 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_8
timestamp 1698431365
transform 1 0 2240 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_12
timestamp 1698431365
transform 1 0 2688 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_28
timestamp 1698431365
transform 1 0 4480 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_36
timestamp 1698431365
transform 1 0 5376 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_40
timestamp 1698431365
transform 1 0 5824 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_42
timestamp 1698431365
transform 1 0 6048 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_84
timestamp 1698431365
transform 1 0 10752 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_86
timestamp 1698431365
transform 1 0 10976 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_139
timestamp 1698431365
transform 1 0 16912 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_142
timestamp 1698431365
transform 1 0 17248 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_183
timestamp 1698431365
transform 1 0 21840 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_212
timestamp 1698431365
transform 1 0 25088 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_216
timestamp 1698431365
transform 1 0 25536 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_220
timestamp 1698431365
transform 1 0 25984 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_236
timestamp 1698431365
transform 1 0 27776 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_240
timestamp 1698431365
transform 1 0 28224 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_242
timestamp 1698431365
transform 1 0 28448 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_274
timestamp 1698431365
transform 1 0 32032 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_278
timestamp 1698431365
transform 1 0 32480 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_282
timestamp 1698431365
transform 1 0 32928 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_284
timestamp 1698431365
transform 1 0 33152 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_326
timestamp 1698431365
transform 1 0 37856 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_360
timestamp 1698431365
transform 1 0 41664 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_362
timestamp 1698431365
transform 1 0 41888 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_392
timestamp 1698431365
transform 1 0 45248 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_408
timestamp 1698431365
transform 1 0 47040 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_418
timestamp 1698431365
transform 1 0 48160 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_451
timestamp 1698431365
transform 1 0 51856 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_483
timestamp 1698431365
transform 1 0 55440 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_487
timestamp 1698431365
transform 1 0 55888 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_489
timestamp 1698431365
transform 1 0 56112 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_492
timestamp 1698431365
transform 1 0 56448 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_508
timestamp 1698431365
transform 1 0 58240 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_2
timestamp 1698431365
transform 1 0 1568 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_34
timestamp 1698431365
transform 1 0 5152 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_37
timestamp 1698431365
transform 1 0 5488 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_45
timestamp 1698431365
transform 1 0 6384 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_107
timestamp 1698431365
transform 1 0 13328 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_163
timestamp 1698431365
transform 1 0 19600 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_167
timestamp 1698431365
transform 1 0 20048 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_171
timestamp 1698431365
transform 1 0 20496 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_205
timestamp 1698431365
transform 1 0 24304 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_243
timestamp 1698431365
transform 1 0 28560 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_247
timestamp 1698431365
transform 1 0 29008 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_265
timestamp 1698431365
transform 1 0 31024 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_271
timestamp 1698431365
transform 1 0 31696 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_312
timestamp 1698431365
transform 1 0 36288 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_314
timestamp 1698431365
transform 1 0 36512 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_322
timestamp 1698431365
transform 1 0 37408 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_326
timestamp 1698431365
transform 1 0 37856 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_330
timestamp 1698431365
transform 1 0 38304 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_334
timestamp 1698431365
transform 1 0 38752 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_383
timestamp 1698431365
transform 1 0 44240 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_392
timestamp 1698431365
transform 1 0 45248 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_396
timestamp 1698431365
transform 1 0 45696 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_437
timestamp 1698431365
transform 1 0 50288 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_453
timestamp 1698431365
transform 1 0 52080 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_457
timestamp 1698431365
transform 1 0 52528 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_489
timestamp 1698431365
transform 1 0 56112 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_505
timestamp 1698431365
transform 1 0 57904 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_8
timestamp 1698431365
transform 1 0 2240 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_12
timestamp 1698431365
transform 1 0 2688 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_28
timestamp 1698431365
transform 1 0 4480 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_36
timestamp 1698431365
transform 1 0 5376 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_40
timestamp 1698431365
transform 1 0 5824 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_138
timestamp 1698431365
transform 1 0 16800 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_146
timestamp 1698431365
transform 1 0 17696 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_150
timestamp 1698431365
transform 1 0 18144 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_212
timestamp 1698431365
transform 1 0 25088 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_271
timestamp 1698431365
transform 1 0 31696 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_275
timestamp 1698431365
transform 1 0 32144 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_279
timestamp 1698431365
transform 1 0 32592 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_288
timestamp 1698431365
transform 1 0 33600 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_300
timestamp 1698431365
transform 1 0 34944 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_331
timestamp 1698431365
transform 1 0 38416 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_335
timestamp 1698431365
transform 1 0 38864 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_347
timestamp 1698431365
transform 1 0 40208 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_349
timestamp 1698431365
transform 1 0 40432 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_352
timestamp 1698431365
transform 1 0 40768 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_354
timestamp 1698431365
transform 1 0 40992 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_365
timestamp 1698431365
transform 1 0 42224 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_369
timestamp 1698431365
transform 1 0 42672 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_397
timestamp 1698431365
transform 1 0 45808 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_401
timestamp 1698431365
transform 1 0 46256 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_417
timestamp 1698431365
transform 1 0 48048 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_419
timestamp 1698431365
transform 1 0 48272 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_422
timestamp 1698431365
transform 1 0 48608 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_426
timestamp 1698431365
transform 1 0 49056 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_492
timestamp 1698431365
transform 1 0 56448 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_508
timestamp 1698431365
transform 1 0 58240 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_8
timestamp 1698431365
transform 1 0 2240 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_12
timestamp 1698431365
transform 1 0 2688 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_28
timestamp 1698431365
transform 1 0 4480 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_32
timestamp 1698431365
transform 1 0 4928 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_34
timestamp 1698431365
transform 1 0 5152 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_37
timestamp 1698431365
transform 1 0 5488 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_107
timestamp 1698431365
transform 1 0 13328 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_109
timestamp 1698431365
transform 1 0 13552 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_172
timestamp 1698431365
transform 1 0 20608 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_174
timestamp 1698431365
transform 1 0 20832 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_233
timestamp 1698431365
transform 1 0 27440 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_247
timestamp 1698431365
transform 1 0 29008 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_276
timestamp 1698431365
transform 1 0 32256 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_292
timestamp 1698431365
transform 1 0 34048 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_302
timestamp 1698431365
transform 1 0 35168 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_312
timestamp 1698431365
transform 1 0 36288 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_314
timestamp 1698431365
transform 1 0 36512 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_317
timestamp 1698431365
transform 1 0 36848 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_321
timestamp 1698431365
transform 1 0 37296 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_349
timestamp 1698431365
transform 1 0 40432 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_353
timestamp 1698431365
transform 1 0 40880 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_355
timestamp 1698431365
transform 1 0 41104 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_362
timestamp 1698431365
transform 1 0 41888 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_364
timestamp 1698431365
transform 1 0 42112 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_373
timestamp 1698431365
transform 1 0 43120 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_379
timestamp 1698431365
transform 1 0 43792 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_383
timestamp 1698431365
transform 1 0 44240 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_387
timestamp 1698431365
transform 1 0 44688 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_391
timestamp 1698431365
transform 1 0 45136 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_394
timestamp 1698431365
transform 1 0 45472 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_396
timestamp 1698431365
transform 1 0 45696 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_399
timestamp 1698431365
transform 1 0 46032 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_403
timestamp 1698431365
transform 1 0 46480 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_405
timestamp 1698431365
transform 1 0 46704 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_408
timestamp 1698431365
transform 1 0 47040 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_417
timestamp 1698431365
transform 1 0 48048 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_421
timestamp 1698431365
transform 1 0 48496 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_453
timestamp 1698431365
transform 1 0 52080 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_457
timestamp 1698431365
transform 1 0 52528 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_489
timestamp 1698431365
transform 1 0 56112 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_505
timestamp 1698431365
transform 1 0 57904 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_8
timestamp 1698431365
transform 1 0 2240 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_12
timestamp 1698431365
transform 1 0 2688 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_16
timestamp 1698431365
transform 1 0 3136 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_32
timestamp 1698431365
transform 1 0 4928 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_40
timestamp 1698431365
transform 1 0 5824 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_42
timestamp 1698431365
transform 1 0 6048 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_76
timestamp 1698431365
transform 1 0 9856 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_142
timestamp 1698431365
transform 1 0 17248 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_189
timestamp 1698431365
transform 1 0 22512 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_217
timestamp 1698431365
transform 1 0 25648 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_267
timestamp 1698431365
transform 1 0 31248 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_271
timestamp 1698431365
transform 1 0 31696 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_298
timestamp 1698431365
transform 1 0 34720 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_300
timestamp 1698431365
transform 1 0 34944 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_315
timestamp 1698431365
transform 1 0 36624 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_317
timestamp 1698431365
transform 1 0 36848 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_349
timestamp 1698431365
transform 1 0 40432 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_352
timestamp 1698431365
transform 1 0 40768 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_356
timestamp 1698431365
transform 1 0 41216 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_360
timestamp 1698431365
transform 1 0 41664 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_372
timestamp 1698431365
transform 1 0 43008 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_413
timestamp 1698431365
transform 1 0 47600 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_417
timestamp 1698431365
transform 1 0 48048 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_419
timestamp 1698431365
transform 1 0 48272 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_422
timestamp 1698431365
transform 1 0 48608 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_486
timestamp 1698431365
transform 1 0 55776 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_492
timestamp 1698431365
transform 1 0 56448 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_508
timestamp 1698431365
transform 1 0 58240 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_14
timestamp 1698431365
transform 1 0 2912 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_18
timestamp 1698431365
transform 1 0 3360 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_34
timestamp 1698431365
transform 1 0 5152 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_37
timestamp 1698431365
transform 1 0 5488 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_45
timestamp 1698431365
transform 1 0 6384 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_53
timestamp 1698431365
transform 1 0 7280 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_55
timestamp 1698431365
transform 1 0 7504 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_99
timestamp 1698431365
transform 1 0 12432 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_103
timestamp 1698431365
transform 1 0 12880 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_233
timestamp 1698431365
transform 1 0 27440 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_237
timestamp 1698431365
transform 1 0 27888 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_241
timestamp 1698431365
transform 1 0 28336 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_247
timestamp 1698431365
transform 1 0 29008 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_255
timestamp 1698431365
transform 1 0 29904 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_284
timestamp 1698431365
transform 1 0 33152 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_317
timestamp 1698431365
transform 1 0 36848 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_321
timestamp 1698431365
transform 1 0 37296 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_379
timestamp 1698431365
transform 1 0 43792 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_384
timestamp 1698431365
transform 1 0 44352 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_402
timestamp 1698431365
transform 1 0 46368 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_406
timestamp 1698431365
transform 1 0 46816 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_436
timestamp 1698431365
transform 1 0 50176 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_452
timestamp 1698431365
transform 1 0 51968 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_454
timestamp 1698431365
transform 1 0 52192 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_457
timestamp 1698431365
transform 1 0 52528 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_489
timestamp 1698431365
transform 1 0 56112 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_497
timestamp 1698431365
transform 1 0 57008 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_8
timestamp 1698431365
transform 1 0 2240 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_12
timestamp 1698431365
transform 1 0 2688 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_28
timestamp 1698431365
transform 1 0 4480 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_32
timestamp 1698431365
transform 1 0 4928 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_63
timestamp 1698431365
transform 1 0 8400 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_67
timestamp 1698431365
transform 1 0 8848 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_69
timestamp 1698431365
transform 1 0 9072 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_113
timestamp 1698431365
transform 1 0 14000 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_121
timestamp 1698431365
transform 1 0 14896 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_125
timestamp 1698431365
transform 1 0 15344 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_133
timestamp 1698431365
transform 1 0 16240 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_135
timestamp 1698431365
transform 1 0 16464 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_177
timestamp 1698431365
transform 1 0 21168 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_181
timestamp 1698431365
transform 1 0 21616 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_185
timestamp 1698431365
transform 1 0 22064 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_188
timestamp 1698431365
transform 1 0 22400 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_192
timestamp 1698431365
transform 1 0 22848 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_196
timestamp 1698431365
transform 1 0 23296 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_200
timestamp 1698431365
transform 1 0 23744 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_212
timestamp 1698431365
transform 1 0 25088 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_238
timestamp 1698431365
transform 1 0 28000 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_242
timestamp 1698431365
transform 1 0 28448 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_244
timestamp 1698431365
transform 1 0 28672 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_274
timestamp 1698431365
transform 1 0 32032 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_278
timestamp 1698431365
transform 1 0 32480 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_282
timestamp 1698431365
transform 1 0 32928 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_336
timestamp 1698431365
transform 1 0 38976 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_345
timestamp 1698431365
transform 1 0 39984 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_349
timestamp 1698431365
transform 1 0 40432 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_419
timestamp 1698431365
transform 1 0 48272 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_439
timestamp 1698431365
transform 1 0 50512 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_471
timestamp 1698431365
transform 1 0 54096 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_487
timestamp 1698431365
transform 1 0 55888 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_489
timestamp 1698431365
transform 1 0 56112 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_492
timestamp 1698431365
transform 1 0 56448 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_508
timestamp 1698431365
transform 1 0 58240 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_8
timestamp 1698431365
transform 1 0 2240 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_12
timestamp 1698431365
transform 1 0 2688 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_28
timestamp 1698431365
transform 1 0 4480 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_32
timestamp 1698431365
transform 1 0 4928 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_34
timestamp 1698431365
transform 1 0 5152 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_37
timestamp 1698431365
transform 1 0 5488 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_45
timestamp 1698431365
transform 1 0 6384 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_64
timestamp 1698431365
transform 1 0 8512 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_72
timestamp 1698431365
transform 1 0 9408 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_163
timestamp 1698431365
transform 1 0 19600 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_167
timestamp 1698431365
transform 1 0 20048 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_171
timestamp 1698431365
transform 1 0 20496 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_177
timestamp 1698431365
transform 1 0 21168 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_181
timestamp 1698431365
transform 1 0 21616 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_201
timestamp 1698431365
transform 1 0 23856 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_203
timestamp 1698431365
transform 1 0 24080 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_237
timestamp 1698431365
transform 1 0 27888 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_241
timestamp 1698431365
transform 1 0 28336 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_257
timestamp 1698431365
transform 1 0 30128 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_265
timestamp 1698431365
transform 1 0 31024 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_269
timestamp 1698431365
transform 1 0 31472 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_271
timestamp 1698431365
transform 1 0 31696 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_309
timestamp 1698431365
transform 1 0 35952 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_313
timestamp 1698431365
transform 1 0 36400 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_325
timestamp 1698431365
transform 1 0 37744 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_329
timestamp 1698431365
transform 1 0 38192 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_333
timestamp 1698431365
transform 1 0 38640 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_365
timestamp 1698431365
transform 1 0 42224 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_383
timestamp 1698431365
transform 1 0 44240 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_443
timestamp 1698431365
transform 1 0 50960 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_451
timestamp 1698431365
transform 1 0 51856 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_457
timestamp 1698431365
transform 1 0 52528 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_489
timestamp 1698431365
transform 1 0 56112 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_497
timestamp 1698431365
transform 1 0 57008 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_8
timestamp 1698431365
transform 1 0 2240 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_12
timestamp 1698431365
transform 1 0 2688 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_28
timestamp 1698431365
transform 1 0 4480 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_69
timestamp 1698431365
transform 1 0 9072 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_72
timestamp 1698431365
transform 1 0 9408 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_81
timestamp 1698431365
transform 1 0 10416 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_85
timestamp 1698431365
transform 1 0 10864 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_123
timestamp 1698431365
transform 1 0 15120 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_127
timestamp 1698431365
transform 1 0 15568 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_135
timestamp 1698431365
transform 1 0 16464 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_139
timestamp 1698431365
transform 1 0 16912 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_142
timestamp 1698431365
transform 1 0 17248 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_152
timestamp 1698431365
transform 1 0 18368 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_156
timestamp 1698431365
transform 1 0 18816 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_160
timestamp 1698431365
transform 1 0 19264 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_164
timestamp 1698431365
transform 1 0 19712 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_260
timestamp 1698431365
transform 1 0 30464 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_282
timestamp 1698431365
transform 1 0 32928 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_288
timestamp 1698431365
transform 1 0 33600 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_294
timestamp 1698431365
transform 1 0 34272 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_296
timestamp 1698431365
transform 1 0 34496 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_299
timestamp 1698431365
transform 1 0 34832 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_408
timestamp 1698431365
transform 1 0 47040 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_412
timestamp 1698431365
transform 1 0 47488 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_414
timestamp 1698431365
transform 1 0 47712 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_443
timestamp 1698431365
transform 1 0 50960 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_475
timestamp 1698431365
transform 1 0 54544 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_483
timestamp 1698431365
transform 1 0 55440 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_487
timestamp 1698431365
transform 1 0 55888 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_489
timestamp 1698431365
transform 1 0 56112 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_492
timestamp 1698431365
transform 1 0 56448 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_500
timestamp 1698431365
transform 1 0 57344 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_8
timestamp 1698431365
transform 1 0 2240 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_12
timestamp 1698431365
transform 1 0 2688 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_28
timestamp 1698431365
transform 1 0 4480 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_32
timestamp 1698431365
transform 1 0 4928 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_34
timestamp 1698431365
transform 1 0 5152 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_37
timestamp 1698431365
transform 1 0 5488 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_41
timestamp 1698431365
transform 1 0 5936 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_43
timestamp 1698431365
transform 1 0 6160 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_73
timestamp 1698431365
transform 1 0 9520 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_77
timestamp 1698431365
transform 1 0 9968 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_154
timestamp 1698431365
transform 1 0 18592 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_156
timestamp 1698431365
transform 1 0 18816 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_167
timestamp 1698431365
transform 1 0 20048 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_169
timestamp 1698431365
transform 1 0 20272 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_227
timestamp 1698431365
transform 1 0 26768 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_235
timestamp 1698431365
transform 1 0 27664 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_243
timestamp 1698431365
transform 1 0 28560 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_247
timestamp 1698431365
transform 1 0 29008 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_263
timestamp 1698431365
transform 1 0 30800 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_305
timestamp 1698431365
transform 1 0 35504 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_309
timestamp 1698431365
transform 1 0 35952 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_313
timestamp 1698431365
transform 1 0 36400 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_351
timestamp 1698431365
transform 1 0 40656 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_384
timestamp 1698431365
transform 1 0 44352 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_416
timestamp 1698431365
transform 1 0 47936 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_448
timestamp 1698431365
transform 1 0 51520 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_452
timestamp 1698431365
transform 1 0 51968 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_454
timestamp 1698431365
transform 1 0 52192 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_457
timestamp 1698431365
transform 1 0 52528 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_489
timestamp 1698431365
transform 1 0 56112 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_497
timestamp 1698431365
transform 1 0 57008 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_8
timestamp 1698431365
transform 1 0 2240 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_12
timestamp 1698431365
transform 1 0 2688 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_16
timestamp 1698431365
transform 1 0 3136 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_48
timestamp 1698431365
transform 1 0 6720 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_56
timestamp 1698431365
transform 1 0 7616 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_64
timestamp 1698431365
transform 1 0 8512 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_68
timestamp 1698431365
transform 1 0 8960 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_72
timestamp 1698431365
transform 1 0 9408 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_80
timestamp 1698431365
transform 1 0 10304 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_84
timestamp 1698431365
transform 1 0 10752 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_129
timestamp 1698431365
transform 1 0 15792 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_131
timestamp 1698431365
transform 1 0 16016 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_209
timestamp 1698431365
transform 1 0 24752 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_225
timestamp 1698431365
transform 1 0 26544 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_229
timestamp 1698431365
transform 1 0 26992 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_233
timestamp 1698431365
transform 1 0 27440 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_237
timestamp 1698431365
transform 1 0 27888 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_241
timestamp 1698431365
transform 1 0 28336 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_248
timestamp 1698431365
transform 1 0 29120 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_282
timestamp 1698431365
transform 1 0 32928 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_286
timestamp 1698431365
transform 1 0 33376 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_319
timestamp 1698431365
transform 1 0 37072 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_324
timestamp 1698431365
transform 1 0 37632 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_328
timestamp 1698431365
transform 1 0 38080 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_340
timestamp 1698431365
transform 1 0 39424 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_348
timestamp 1698431365
transform 1 0 40320 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_352
timestamp 1698431365
transform 1 0 40768 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_368
timestamp 1698431365
transform 1 0 42560 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_397
timestamp 1698431365
transform 1 0 45808 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_401
timestamp 1698431365
transform 1 0 46256 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_411
timestamp 1698431365
transform 1 0 47376 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_438
timestamp 1698431365
transform 1 0 50400 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_470
timestamp 1698431365
transform 1 0 53984 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_486
timestamp 1698431365
transform 1 0 55776 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_492
timestamp 1698431365
transform 1 0 56448 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_508
timestamp 1698431365
transform 1 0 58240 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_14
timestamp 1698431365
transform 1 0 2912 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_18
timestamp 1698431365
transform 1 0 3360 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_34
timestamp 1698431365
transform 1 0 5152 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_37
timestamp 1698431365
transform 1 0 5488 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_53
timestamp 1698431365
transform 1 0 7280 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_90
timestamp 1698431365
transform 1 0 11424 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_98
timestamp 1698431365
transform 1 0 12320 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_102
timestamp 1698431365
transform 1 0 12768 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_104
timestamp 1698431365
transform 1 0 12992 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_134
timestamp 1698431365
transform 1 0 16352 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_169
timestamp 1698431365
transform 1 0 20272 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_177
timestamp 1698431365
transform 1 0 21168 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_217
timestamp 1698431365
transform 1 0 25648 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_221
timestamp 1698431365
transform 1 0 26096 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_225
timestamp 1698431365
transform 1 0 26544 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_229
timestamp 1698431365
transform 1 0 26992 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_240
timestamp 1698431365
transform 1 0 28224 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_244
timestamp 1698431365
transform 1 0 28672 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_276
timestamp 1698431365
transform 1 0 32256 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_280
timestamp 1698431365
transform 1 0 32704 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_309
timestamp 1698431365
transform 1 0 35952 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_313
timestamp 1698431365
transform 1 0 36400 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_317
timestamp 1698431365
transform 1 0 36848 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_319
timestamp 1698431365
transform 1 0 37072 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_337
timestamp 1698431365
transform 1 0 39088 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_351
timestamp 1698431365
transform 1 0 40656 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_378
timestamp 1698431365
transform 1 0 43680 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_382
timestamp 1698431365
transform 1 0 44128 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_384
timestamp 1698431365
transform 1 0 44352 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_391
timestamp 1698431365
transform 1 0 45136 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_449
timestamp 1698431365
transform 1 0 51632 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_453
timestamp 1698431365
transform 1 0 52080 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_457
timestamp 1698431365
transform 1 0 52528 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_489
timestamp 1698431365
transform 1 0 56112 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_505
timestamp 1698431365
transform 1 0 57904 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_8
timestamp 1698431365
transform 1 0 2240 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_31_12
timestamp 1698431365
transform 1 0 2688 0 -1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_44
timestamp 1698431365
transform 1 0 6272 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_60
timestamp 1698431365
transform 1 0 8064 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_68
timestamp 1698431365
transform 1 0 8960 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_72
timestamp 1698431365
transform 1 0 9408 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_74
timestamp 1698431365
transform 1 0 9632 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_79
timestamp 1698431365
transform 1 0 10192 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_83
timestamp 1698431365
transform 1 0 10640 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_114
timestamp 1698431365
transform 1 0 14112 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_118
timestamp 1698431365
transform 1 0 14560 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_126
timestamp 1698431365
transform 1 0 15456 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_142
timestamp 1698431365
transform 1 0 17248 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_146
timestamp 1698431365
transform 1 0 17696 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_150
timestamp 1698431365
transform 1 0 18144 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_153
timestamp 1698431365
transform 1 0 18480 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_200
timestamp 1698431365
transform 1 0 23744 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_206
timestamp 1698431365
transform 1 0 24416 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_225
timestamp 1698431365
transform 1 0 26544 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_229
timestamp 1698431365
transform 1 0 26992 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_239
timestamp 1698431365
transform 1 0 28112 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_241
timestamp 1698431365
transform 1 0 28336 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_244
timestamp 1698431365
transform 1 0 28672 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_248
timestamp 1698431365
transform 1 0 29120 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_263
timestamp 1698431365
transform 1 0 30800 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_311
timestamp 1698431365
transform 1 0 36176 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_319
timestamp 1698431365
transform 1 0 37072 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_364
timestamp 1698431365
transform 1 0 42112 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_394
timestamp 1698431365
transform 1 0 45472 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_398
timestamp 1698431365
transform 1 0 45920 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_402
timestamp 1698431365
transform 1 0 46368 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_405
timestamp 1698431365
transform 1 0 46704 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_413
timestamp 1698431365
transform 1 0 47600 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_419
timestamp 1698431365
transform 1 0 48272 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_31_440
timestamp 1698431365
transform 1 0 50624 0 -1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_472
timestamp 1698431365
transform 1 0 54208 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_488
timestamp 1698431365
transform 1 0 56000 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_492
timestamp 1698431365
transform 1 0 56448 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_508
timestamp 1698431365
transform 1 0 58240 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_8
timestamp 1698431365
transform 1 0 2240 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_12
timestamp 1698431365
transform 1 0 2688 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_28
timestamp 1698431365
transform 1 0 4480 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_32
timestamp 1698431365
transform 1 0 4928 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_34
timestamp 1698431365
transform 1 0 5152 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_37
timestamp 1698431365
transform 1 0 5488 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_53
timestamp 1698431365
transform 1 0 7280 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_104
timestamp 1698431365
transform 1 0 12992 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_111
timestamp 1698431365
transform 1 0 13776 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_113
timestamp 1698431365
transform 1 0 14000 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_172
timestamp 1698431365
transform 1 0 20608 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_174
timestamp 1698431365
transform 1 0 20832 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_177
timestamp 1698431365
transform 1 0 21168 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_199
timestamp 1698431365
transform 1 0 23632 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_252
timestamp 1698431365
transform 1 0 29568 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_284
timestamp 1698431365
transform 1 0 33152 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_286
timestamp 1698431365
transform 1 0 33376 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_325
timestamp 1698431365
transform 1 0 37744 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_331
timestamp 1698431365
transform 1 0 38416 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_335
timestamp 1698431365
transform 1 0 38864 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_339
timestamp 1698431365
transform 1 0 39312 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_345
timestamp 1698431365
transform 1 0 39984 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_347
timestamp 1698431365
transform 1 0 40208 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_373
timestamp 1698431365
transform 1 0 43120 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_403
timestamp 1698431365
transform 1 0 46480 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_405
timestamp 1698431365
transform 1 0 46704 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_413
timestamp 1698431365
transform 1 0 47600 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_417
timestamp 1698431365
transform 1 0 48048 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_449
timestamp 1698431365
transform 1 0 51632 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_453
timestamp 1698431365
transform 1 0 52080 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_457
timestamp 1698431365
transform 1 0 52528 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_473
timestamp 1698431365
transform 1 0 54320 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_8
timestamp 1698431365
transform 1 0 2240 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_33_12
timestamp 1698431365
transform 1 0 2688 0 -1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_33_44
timestamp 1698431365
transform 1 0 6272 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_60
timestamp 1698431365
transform 1 0 8064 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_64
timestamp 1698431365
transform 1 0 8512 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_72
timestamp 1698431365
transform 1 0 9408 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_139
timestamp 1698431365
transform 1 0 16912 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_192
timestamp 1698431365
transform 1 0 22848 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_194
timestamp 1698431365
transform 1 0 23072 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_212
timestamp 1698431365
transform 1 0 25088 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_222
timestamp 1698431365
transform 1 0 26208 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_265
timestamp 1698431365
transform 1 0 31024 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_279
timestamp 1698431365
transform 1 0 32592 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_282
timestamp 1698431365
transform 1 0 32928 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_286
timestamp 1698431365
transform 1 0 33376 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_290
timestamp 1698431365
transform 1 0 33824 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_317
timestamp 1698431365
transform 1 0 36848 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_325
timestamp 1698431365
transform 1 0 37744 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_336
timestamp 1698431365
transform 1 0 38976 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_342
timestamp 1698431365
transform 1 0 39648 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_344
timestamp 1698431365
transform 1 0 39872 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_417
timestamp 1698431365
transform 1 0 48048 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_419
timestamp 1698431365
transform 1 0 48272 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_422
timestamp 1698431365
transform 1 0 48608 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_426
timestamp 1698431365
transform 1 0 49056 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_33_492
timestamp 1698431365
transform 1 0 56448 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_508
timestamp 1698431365
transform 1 0 58240 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_8
timestamp 1698431365
transform 1 0 2240 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_12
timestamp 1698431365
transform 1 0 2688 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_34_16
timestamp 1698431365
transform 1 0 3136 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_32
timestamp 1698431365
transform 1 0 4928 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_34
timestamp 1698431365
transform 1 0 5152 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_34_37
timestamp 1698431365
transform 1 0 5488 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_53
timestamp 1698431365
transform 1 0 7280 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_86
timestamp 1698431365
transform 1 0 10976 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_96
timestamp 1698431365
transform 1 0 12096 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_100
timestamp 1698431365
transform 1 0 12544 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_104
timestamp 1698431365
transform 1 0 12992 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_136
timestamp 1698431365
transform 1 0 16576 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_144
timestamp 1698431365
transform 1 0 17472 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_148
timestamp 1698431365
transform 1 0 17920 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_154
timestamp 1698431365
transform 1 0 18592 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_158
timestamp 1698431365
transform 1 0 19040 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_160
timestamp 1698431365
transform 1 0 19264 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_171
timestamp 1698431365
transform 1 0 20496 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_193
timestamp 1698431365
transform 1 0 22960 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_228
timestamp 1698431365
transform 1 0 26880 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_247
timestamp 1698431365
transform 1 0 29008 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_290
timestamp 1698431365
transform 1 0 33824 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_294
timestamp 1698431365
transform 1 0 34272 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_304
timestamp 1698431365
transform 1 0 35392 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_306
timestamp 1698431365
transform 1 0 35616 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_309
timestamp 1698431365
transform 1 0 35952 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_313
timestamp 1698431365
transform 1 0 36400 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_322
timestamp 1698431365
transform 1 0 37408 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_344
timestamp 1698431365
transform 1 0 39872 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_346
timestamp 1698431365
transform 1 0 40096 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_377
timestamp 1698431365
transform 1 0 43568 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_381
timestamp 1698431365
transform 1 0 44016 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_408
timestamp 1698431365
transform 1 0 47040 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_443
timestamp 1698431365
transform 1 0 50960 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_451
timestamp 1698431365
transform 1 0 51856 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_457
timestamp 1698431365
transform 1 0 52528 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_461
timestamp 1698431365
transform 1 0 52976 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_34_490
timestamp 1698431365
transform 1 0 56224 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_506
timestamp 1698431365
transform 1 0 58016 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_508
timestamp 1698431365
transform 1 0 58240 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_14
timestamp 1698431365
transform 1 0 2912 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_35_18
timestamp 1698431365
transform 1 0 3360 0 -1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_35_50
timestamp 1698431365
transform 1 0 6944 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_66
timestamp 1698431365
transform 1 0 8736 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_72
timestamp 1698431365
transform 1 0 9408 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_138
timestamp 1698431365
transform 1 0 16800 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_35_147
timestamp 1698431365
transform 1 0 17808 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_163
timestamp 1698431365
transform 1 0 19600 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_165
timestamp 1698431365
transform 1 0 19824 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_208
timestamp 1698431365
transform 1 0 24640 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_267
timestamp 1698431365
transform 1 0 31248 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_316
timestamp 1698431365
transform 1 0 36736 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_320
timestamp 1698431365
transform 1 0 37184 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_324
timestamp 1698431365
transform 1 0 37632 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_326
timestamp 1698431365
transform 1 0 37856 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_343
timestamp 1698431365
transform 1 0 39760 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_347
timestamp 1698431365
transform 1 0 40208 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_349
timestamp 1698431365
transform 1 0 40432 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_352
timestamp 1698431365
transform 1 0 40768 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_35_375
timestamp 1698431365
transform 1 0 43344 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_407
timestamp 1698431365
transform 1 0 46928 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_419
timestamp 1698431365
transform 1 0 48272 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_35_472
timestamp 1698431365
transform 1 0 54208 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_488
timestamp 1698431365
transform 1 0 56000 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_35_492
timestamp 1698431365
transform 1 0 56448 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_508
timestamp 1698431365
transform 1 0 58240 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_28
timestamp 1698431365
transform 1 0 4480 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_32
timestamp 1698431365
transform 1 0 4928 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_34
timestamp 1698431365
transform 1 0 5152 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_36_37
timestamp 1698431365
transform 1 0 5488 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_53
timestamp 1698431365
transform 1 0 7280 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_86
timestamp 1698431365
transform 1 0 10976 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_103
timestamp 1698431365
transform 1 0 12880 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_107
timestamp 1698431365
transform 1 0 13328 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_134
timestamp 1698431365
transform 1 0 16352 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_165
timestamp 1698431365
transform 1 0 19824 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_173
timestamp 1698431365
transform 1 0 20720 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_177
timestamp 1698431365
transform 1 0 21168 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_179
timestamp 1698431365
transform 1 0 21392 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_192
timestamp 1698431365
transform 1 0 22848 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_196
timestamp 1698431365
transform 1 0 23296 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_200
timestamp 1698431365
transform 1 0 23744 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_204
timestamp 1698431365
transform 1 0 24192 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_208
timestamp 1698431365
transform 1 0 24640 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_225
timestamp 1698431365
transform 1 0 26544 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_237
timestamp 1698431365
transform 1 0 27888 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_241
timestamp 1698431365
transform 1 0 28336 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_247
timestamp 1698431365
transform 1 0 29008 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_249
timestamp 1698431365
transform 1 0 29232 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_310
timestamp 1698431365
transform 1 0 36064 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_314
timestamp 1698431365
transform 1 0 36512 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_325
timestamp 1698431365
transform 1 0 37744 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_333
timestamp 1698431365
transform 1 0 38640 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_347
timestamp 1698431365
transform 1 0 40208 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_351
timestamp 1698431365
transform 1 0 40656 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_353
timestamp 1698431365
transform 1 0 40880 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_383
timestamp 1698431365
transform 1 0 44240 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_387
timestamp 1698431365
transform 1 0 44688 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_389
timestamp 1698431365
transform 1 0 44912 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_441
timestamp 1698431365
transform 1 0 50736 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_449
timestamp 1698431365
transform 1 0 51632 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_453
timestamp 1698431365
transform 1 0 52080 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_8
timestamp 1698431365
transform 1 0 2240 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_37_12
timestamp 1698431365
transform 1 0 2688 0 -1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_37_44
timestamp 1698431365
transform 1 0 6272 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_60
timestamp 1698431365
transform 1 0 8064 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_64
timestamp 1698431365
transform 1 0 8512 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_72
timestamp 1698431365
transform 1 0 9408 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_74
timestamp 1698431365
transform 1 0 9632 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_79
timestamp 1698431365
transform 1 0 10192 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_87
timestamp 1698431365
transform 1 0 11088 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_116
timestamp 1698431365
transform 1 0 14336 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_125
timestamp 1698431365
transform 1 0 15344 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_129
timestamp 1698431365
transform 1 0 15792 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_139
timestamp 1698431365
transform 1 0 16912 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_142
timestamp 1698431365
transform 1 0 17248 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_195
timestamp 1698431365
transform 1 0 23184 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_199
timestamp 1698431365
transform 1 0 23632 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_217
timestamp 1698431365
transform 1 0 25648 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_256
timestamp 1698431365
transform 1 0 30016 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_260
timestamp 1698431365
transform 1 0 30464 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_277
timestamp 1698431365
transform 1 0 32368 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_279
timestamp 1698431365
transform 1 0 32592 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_290
timestamp 1698431365
transform 1 0 33824 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_316
timestamp 1698431365
transform 1 0 36736 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_320
timestamp 1698431365
transform 1 0 37184 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_37_352
timestamp 1698431365
transform 1 0 40768 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_368
timestamp 1698431365
transform 1 0 42560 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_370
timestamp 1698431365
transform 1 0 42784 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_410
timestamp 1698431365
transform 1 0 47264 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_418
timestamp 1698431365
transform 1 0 48160 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_422
timestamp 1698431365
transform 1 0 48608 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_426
timestamp 1698431365
transform 1 0 49056 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_37_429
timestamp 1698431365
transform 1 0 49392 0 -1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_461
timestamp 1698431365
transform 1 0 52976 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_463
timestamp 1698431365
transform 1 0 53200 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_37_492
timestamp 1698431365
transform 1 0 56448 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_508
timestamp 1698431365
transform 1 0 58240 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_8
timestamp 1698431365
transform 1 0 2240 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_38_12
timestamp 1698431365
transform 1 0 2688 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_28
timestamp 1698431365
transform 1 0 4480 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_32
timestamp 1698431365
transform 1 0 4928 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_34
timestamp 1698431365
transform 1 0 5152 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_38_37
timestamp 1698431365
transform 1 0 5488 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_53
timestamp 1698431365
transform 1 0 7280 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_57
timestamp 1698431365
transform 1 0 7728 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_59
timestamp 1698431365
transform 1 0 7952 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_38_89
timestamp 1698431365
transform 1 0 11312 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_107
timestamp 1698431365
transform 1 0 13328 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_115
timestamp 1698431365
transform 1 0 14224 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_117
timestamp 1698431365
transform 1 0 14448 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_125
timestamp 1698431365
transform 1 0 15344 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_133
timestamp 1698431365
transform 1 0 16240 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_137
timestamp 1698431365
transform 1 0 16688 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_141
timestamp 1698431365
transform 1 0 17136 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_151
timestamp 1698431365
transform 1 0 18256 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_161
timestamp 1698431365
transform 1 0 19376 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_165
timestamp 1698431365
transform 1 0 19824 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_173
timestamp 1698431365
transform 1 0 20720 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_177
timestamp 1698431365
transform 1 0 21168 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_181
timestamp 1698431365
transform 1 0 21616 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_183
timestamp 1698431365
transform 1 0 21840 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_186
timestamp 1698431365
transform 1 0 22176 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_190
timestamp 1698431365
transform 1 0 22624 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_192
timestamp 1698431365
transform 1 0 22848 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_222
timestamp 1698431365
transform 1 0 26208 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_224
timestamp 1698431365
transform 1 0 26432 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_227
timestamp 1698431365
transform 1 0 26768 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_260
timestamp 1698431365
transform 1 0 30464 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_262
timestamp 1698431365
transform 1 0 30688 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_277
timestamp 1698431365
transform 1 0 32368 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_281
timestamp 1698431365
transform 1 0 32816 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_289
timestamp 1698431365
transform 1 0 33712 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_322
timestamp 1698431365
transform 1 0 37408 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_326
timestamp 1698431365
transform 1 0 37856 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_330
timestamp 1698431365
transform 1 0 38304 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_338
timestamp 1698431365
transform 1 0 39200 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_340
timestamp 1698431365
transform 1 0 39424 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_343
timestamp 1698431365
transform 1 0 39760 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_347
timestamp 1698431365
transform 1 0 40208 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_349
timestamp 1698431365
transform 1 0 40432 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_38_357
timestamp 1698431365
transform 1 0 41328 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_373
timestamp 1698431365
transform 1 0 43120 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_377
timestamp 1698431365
transform 1 0 43568 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_387
timestamp 1698431365
transform 1 0 44688 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_395
timestamp 1698431365
transform 1 0 45584 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_404
timestamp 1698431365
transform 1 0 46592 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_412
timestamp 1698431365
transform 1 0 47488 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_420
timestamp 1698431365
transform 1 0 48384 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_442
timestamp 1698431365
transform 1 0 50848 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_450
timestamp 1698431365
transform 1 0 51744 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_454
timestamp 1698431365
transform 1 0 52192 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_38_457
timestamp 1698431365
transform 1 0 52528 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_473
timestamp 1698431365
transform 1 0 54320 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_28
timestamp 1698431365
transform 1 0 4480 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_39_32
timestamp 1698431365
transform 1 0 4928 0 -1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_64
timestamp 1698431365
transform 1 0 8512 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_68
timestamp 1698431365
transform 1 0 8960 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_72
timestamp 1698431365
transform 1 0 9408 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_80
timestamp 1698431365
transform 1 0 10304 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_116
timestamp 1698431365
transform 1 0 14336 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_120
timestamp 1698431365
transform 1 0 14784 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_135
timestamp 1698431365
transform 1 0 16464 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_139
timestamp 1698431365
transform 1 0 16912 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_39_142
timestamp 1698431365
transform 1 0 17248 0 -1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_39_174
timestamp 1698431365
transform 1 0 20832 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_190
timestamp 1698431365
transform 1 0 22624 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_194
timestamp 1698431365
transform 1 0 23072 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_231
timestamp 1698431365
transform 1 0 27216 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_233
timestamp 1698431365
transform 1 0 27440 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_236
timestamp 1698431365
transform 1 0 27776 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_260
timestamp 1698431365
transform 1 0 30464 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_262
timestamp 1698431365
transform 1 0 30688 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_269
timestamp 1698431365
transform 1 0 31472 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_273
timestamp 1698431365
transform 1 0 31920 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_279
timestamp 1698431365
transform 1 0 32592 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_282
timestamp 1698431365
transform 1 0 32928 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_286
timestamp 1698431365
transform 1 0 33376 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_288
timestamp 1698431365
transform 1 0 33600 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_291
timestamp 1698431365
transform 1 0 33936 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_332
timestamp 1698431365
transform 1 0 38528 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_336
timestamp 1698431365
transform 1 0 38976 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_348
timestamp 1698431365
transform 1 0 40320 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_386
timestamp 1698431365
transform 1 0 44576 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_390
timestamp 1698431365
transform 1 0 45024 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_394
timestamp 1698431365
transform 1 0 45472 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_408
timestamp 1698431365
transform 1 0 47040 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_410
timestamp 1698431365
transform 1 0 47264 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_416
timestamp 1698431365
transform 1 0 47936 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_451
timestamp 1698431365
transform 1 0 51856 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_459
timestamp 1698431365
transform 1 0 52752 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_463
timestamp 1698431365
transform 1 0 53200 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_39_492
timestamp 1698431365
transform 1 0 56448 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_508
timestamp 1698431365
transform 1 0 58240 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_8
timestamp 1698431365
transform 1 0 2240 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_12
timestamp 1698431365
transform 1 0 2688 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_40_16
timestamp 1698431365
transform 1 0 3136 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_32
timestamp 1698431365
transform 1 0 4928 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_34
timestamp 1698431365
transform 1 0 5152 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_40_37
timestamp 1698431365
transform 1 0 5488 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_53
timestamp 1698431365
transform 1 0 7280 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_90
timestamp 1698431365
transform 1 0 11424 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_94
timestamp 1698431365
transform 1 0 11872 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_144
timestamp 1698431365
transform 1 0 17472 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_156
timestamp 1698431365
transform 1 0 18816 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_160
timestamp 1698431365
transform 1 0 19264 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_168
timestamp 1698431365
transform 1 0 20160 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_177
timestamp 1698431365
transform 1 0 21168 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_179
timestamp 1698431365
transform 1 0 21392 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_188
timestamp 1698431365
transform 1 0 22400 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_224
timestamp 1698431365
transform 1 0 26432 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_244
timestamp 1698431365
transform 1 0 28672 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_247
timestamp 1698431365
transform 1 0 29008 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_251
timestamp 1698431365
transform 1 0 29456 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_259
timestamp 1698431365
transform 1 0 30352 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_263
timestamp 1698431365
transform 1 0 30800 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_265
timestamp 1698431365
transform 1 0 31024 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_288
timestamp 1698431365
transform 1 0 33600 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_292
timestamp 1698431365
transform 1 0 34048 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_311
timestamp 1698431365
transform 1 0 36176 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_317
timestamp 1698431365
transform 1 0 36848 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_322
timestamp 1698431365
transform 1 0 37408 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_326
timestamp 1698431365
transform 1 0 37856 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_330
timestamp 1698431365
transform 1 0 38304 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_336
timestamp 1698431365
transform 1 0 38976 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_344
timestamp 1698431365
transform 1 0 39872 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_351
timestamp 1698431365
transform 1 0 40656 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_353
timestamp 1698431365
transform 1 0 40880 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_382
timestamp 1698431365
transform 1 0 44128 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_384
timestamp 1698431365
transform 1 0 44352 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_392
timestamp 1698431365
transform 1 0 45248 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_40_429
timestamp 1698431365
transform 1 0 49392 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_445
timestamp 1698431365
transform 1 0 51184 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_453
timestamp 1698431365
transform 1 0 52080 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_40_457
timestamp 1698431365
transform 1 0 52528 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_473
timestamp 1698431365
transform 1 0 54320 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_481
timestamp 1698431365
transform 1 0 55216 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_14
timestamp 1698431365
transform 1 0 2912 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_41_18
timestamp 1698431365
transform 1 0 3360 0 -1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_41_50
timestamp 1698431365
transform 1 0 6944 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_66
timestamp 1698431365
transform 1 0 8736 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_72
timestamp 1698431365
transform 1 0 9408 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_76
timestamp 1698431365
transform 1 0 9856 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_137
timestamp 1698431365
transform 1 0 16688 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_139
timestamp 1698431365
transform 1 0 16912 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_166
timestamp 1698431365
transform 1 0 19936 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_168
timestamp 1698431365
transform 1 0 20160 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_195
timestamp 1698431365
transform 1 0 23184 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_199
timestamp 1698431365
transform 1 0 23632 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_203
timestamp 1698431365
transform 1 0 24080 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_207
timestamp 1698431365
transform 1 0 24528 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_209
timestamp 1698431365
transform 1 0 24752 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_212
timestamp 1698431365
transform 1 0 25088 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_222
timestamp 1698431365
transform 1 0 26208 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_226
timestamp 1698431365
transform 1 0 26656 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_230
timestamp 1698431365
transform 1 0 27104 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_41_234
timestamp 1698431365
transform 1 0 27552 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_250
timestamp 1698431365
transform 1 0 29344 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_282
timestamp 1698431365
transform 1 0 32928 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_292
timestamp 1698431365
transform 1 0 34048 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_298
timestamp 1698431365
transform 1 0 34720 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_300
timestamp 1698431365
transform 1 0 34944 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_336
timestamp 1698431365
transform 1 0 38976 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_338
timestamp 1698431365
transform 1 0 39200 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_348
timestamp 1698431365
transform 1 0 40320 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_385
timestamp 1698431365
transform 1 0 44464 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_389
timestamp 1698431365
transform 1 0 44912 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_408
timestamp 1698431365
transform 1 0 47040 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_410
timestamp 1698431365
transform 1 0 47264 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_451
timestamp 1698431365
transform 1 0 51856 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_459
timestamp 1698431365
transform 1 0 52752 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_461
timestamp 1698431365
transform 1 0 52976 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_41_492
timestamp 1698431365
transform 1 0 56448 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_508
timestamp 1698431365
transform 1 0 58240 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_28
timestamp 1698431365
transform 1 0 4480 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_32
timestamp 1698431365
transform 1 0 4928 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_34
timestamp 1698431365
transform 1 0 5152 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_37
timestamp 1698431365
transform 1 0 5488 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_53
timestamp 1698431365
transform 1 0 7280 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_61
timestamp 1698431365
transform 1 0 8176 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_91
timestamp 1698431365
transform 1 0 11536 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_99
timestamp 1698431365
transform 1 0 12432 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_141
timestamp 1698431365
transform 1 0 17136 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_172
timestamp 1698431365
transform 1 0 20608 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_174
timestamp 1698431365
transform 1 0 20832 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_193
timestamp 1698431365
transform 1 0 22960 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_197
timestamp 1698431365
transform 1 0 23408 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_201
timestamp 1698431365
transform 1 0 23856 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_205
timestamp 1698431365
transform 1 0 24304 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_208
timestamp 1698431365
transform 1 0 24640 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_235
timestamp 1698431365
transform 1 0 27664 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_266
timestamp 1698431365
transform 1 0 31136 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_303
timestamp 1698431365
transform 1 0 35280 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_314
timestamp 1698431365
transform 1 0 36512 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_373
timestamp 1698431365
transform 1 0 43120 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_378
timestamp 1698431365
transform 1 0 43680 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_380
timestamp 1698431365
transform 1 0 43904 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_445
timestamp 1698431365
transform 1 0 51184 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_8
timestamp 1698431365
transform 1 0 2240 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_43_12
timestamp 1698431365
transform 1 0 2688 0 -1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_44
timestamp 1698431365
transform 1 0 6272 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_60
timestamp 1698431365
transform 1 0 8064 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_68
timestamp 1698431365
transform 1 0 8960 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_72
timestamp 1698431365
transform 1 0 9408 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_76
timestamp 1698431365
transform 1 0 9856 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_82
timestamp 1698431365
transform 1 0 10528 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_142
timestamp 1698431365
transform 1 0 17248 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_164
timestamp 1698431365
transform 1 0 19712 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_179
timestamp 1698431365
transform 1 0 21392 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_188
timestamp 1698431365
transform 1 0 22400 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_194
timestamp 1698431365
transform 1 0 23072 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_196
timestamp 1698431365
transform 1 0 23296 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_225
timestamp 1698431365
transform 1 0 26544 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_227
timestamp 1698431365
transform 1 0 26768 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_266
timestamp 1698431365
transform 1 0 31136 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_272
timestamp 1698431365
transform 1 0 31808 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_282
timestamp 1698431365
transform 1 0 32928 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_286
timestamp 1698431365
transform 1 0 33376 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_289
timestamp 1698431365
transform 1 0 33712 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_291
timestamp 1698431365
transform 1 0 33936 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_352
timestamp 1698431365
transform 1 0 40768 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_356
timestamp 1698431365
transform 1 0 41216 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_418
timestamp 1698431365
transform 1 0 48160 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_43_431
timestamp 1698431365
transform 1 0 49616 0 -1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_463
timestamp 1698431365
transform 1 0 53200 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_492
timestamp 1698431365
transform 1 0 56448 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_508
timestamp 1698431365
transform 1 0 58240 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_8
timestamp 1698431365
transform 1 0 2240 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_44_12
timestamp 1698431365
transform 1 0 2688 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_28
timestamp 1698431365
transform 1 0 4480 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_32
timestamp 1698431365
transform 1 0 4928 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_34
timestamp 1698431365
transform 1 0 5152 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_44_37
timestamp 1698431365
transform 1 0 5488 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_53
timestamp 1698431365
transform 1 0 7280 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_61
timestamp 1698431365
transform 1 0 8176 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_65
timestamp 1698431365
transform 1 0 8624 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_96
timestamp 1698431365
transform 1 0 12096 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_104
timestamp 1698431365
transform 1 0 12992 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_140
timestamp 1698431365
transform 1 0 17024 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_157
timestamp 1698431365
transform 1 0 18928 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_177
timestamp 1698431365
transform 1 0 21168 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_188
timestamp 1698431365
transform 1 0 22400 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_232
timestamp 1698431365
transform 1 0 27328 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_244
timestamp 1698431365
transform 1 0 28672 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_293
timestamp 1698431365
transform 1 0 34160 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_301
timestamp 1698431365
transform 1 0 35056 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_305
timestamp 1698431365
transform 1 0 35504 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_313
timestamp 1698431365
transform 1 0 36400 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_317
timestamp 1698431365
transform 1 0 36848 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_350
timestamp 1698431365
transform 1 0 40544 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_358
timestamp 1698431365
transform 1 0 41440 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_362
timestamp 1698431365
transform 1 0 41888 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_372
timestamp 1698431365
transform 1 0 43008 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_376
timestamp 1698431365
transform 1 0 43456 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_381
timestamp 1698431365
transform 1 0 44016 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_44_387
timestamp 1698431365
transform 1 0 44688 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_403
timestamp 1698431365
transform 1 0 46480 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_417
timestamp 1698431365
transform 1 0 48048 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_423
timestamp 1698431365
transform 1 0 48720 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_44_457
timestamp 1698431365
transform 1 0 52528 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_473
timestamp 1698431365
transform 1 0 54320 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_45_28
timestamp 1698431365
transform 1 0 4480 0 -1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_60
timestamp 1698431365
transform 1 0 8064 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_68
timestamp 1698431365
transform 1 0 8960 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_72
timestamp 1698431365
transform 1 0 9408 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_80
timestamp 1698431365
transform 1 0 10304 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_115
timestamp 1698431365
transform 1 0 14224 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_117
timestamp 1698431365
transform 1 0 14448 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_138
timestamp 1698431365
transform 1 0 16800 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_142
timestamp 1698431365
transform 1 0 17248 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_146
timestamp 1698431365
transform 1 0 17696 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_148
timestamp 1698431365
transform 1 0 17920 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_151
timestamp 1698431365
transform 1 0 18256 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_155
timestamp 1698431365
transform 1 0 18704 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_163
timestamp 1698431365
transform 1 0 19600 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_212
timestamp 1698431365
transform 1 0 25088 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_216
timestamp 1698431365
transform 1 0 25536 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_224
timestamp 1698431365
transform 1 0 26432 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_228
timestamp 1698431365
transform 1 0 26880 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_261
timestamp 1698431365
transform 1 0 30576 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_332
timestamp 1698431365
transform 1 0 38528 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_336
timestamp 1698431365
transform 1 0 38976 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_342
timestamp 1698431365
transform 1 0 39648 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_356
timestamp 1698431365
transform 1 0 41216 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_422
timestamp 1698431365
transform 1 0 48608 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_45_433
timestamp 1698431365
transform 1 0 49840 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_449
timestamp 1698431365
transform 1 0 51632 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_457
timestamp 1698431365
transform 1 0 52528 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_461
timestamp 1698431365
transform 1 0 52976 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_45_492
timestamp 1698431365
transform 1 0 56448 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_508
timestamp 1698431365
transform 1 0 58240 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_8
timestamp 1698431365
transform 1 0 2240 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_46_12
timestamp 1698431365
transform 1 0 2688 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_28
timestamp 1698431365
transform 1 0 4480 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_32
timestamp 1698431365
transform 1 0 4928 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_34
timestamp 1698431365
transform 1 0 5152 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_46_37
timestamp 1698431365
transform 1 0 5488 0 1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_69
timestamp 1698431365
transform 1 0 9072 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_77
timestamp 1698431365
transform 1 0 9968 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_111
timestamp 1698431365
transform 1 0 13776 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_115
timestamp 1698431365
transform 1 0 14224 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_123
timestamp 1698431365
transform 1 0 15120 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_171
timestamp 1698431365
transform 1 0 20496 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_177
timestamp 1698431365
transform 1 0 21168 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_231
timestamp 1698431365
transform 1 0 27216 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_235
timestamp 1698431365
transform 1 0 27664 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_243
timestamp 1698431365
transform 1 0 28560 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_247
timestamp 1698431365
transform 1 0 29008 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_251
timestamp 1698431365
transform 1 0 29456 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_259
timestamp 1698431365
transform 1 0 30352 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_274
timestamp 1698431365
transform 1 0 32032 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_278
timestamp 1698431365
transform 1 0 32480 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_282
timestamp 1698431365
transform 1 0 32928 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_312
timestamp 1698431365
transform 1 0 36288 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_314
timestamp 1698431365
transform 1 0 36512 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_317
timestamp 1698431365
transform 1 0 36848 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_347
timestamp 1698431365
transform 1 0 40208 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_364
timestamp 1698431365
transform 1 0 42112 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_368
timestamp 1698431365
transform 1 0 42560 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_378
timestamp 1698431365
transform 1 0 43680 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_382
timestamp 1698431365
transform 1 0 44128 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_384
timestamp 1698431365
transform 1 0 44352 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_387
timestamp 1698431365
transform 1 0 44688 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_416
timestamp 1698431365
transform 1 0 47936 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_449
timestamp 1698431365
transform 1 0 51632 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_453
timestamp 1698431365
transform 1 0 52080 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_46_457
timestamp 1698431365
transform 1 0 52528 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_473
timestamp 1698431365
transform 1 0 54320 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_8
timestamp 1698431365
transform 1 0 2240 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_12
timestamp 1698431365
transform 1 0 2688 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_47_16
timestamp 1698431365
transform 1 0 3136 0 -1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_47_48
timestamp 1698431365
transform 1 0 6720 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_64
timestamp 1698431365
transform 1 0 8512 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_68
timestamp 1698431365
transform 1 0 8960 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_47_72
timestamp 1698431365
transform 1 0 9408 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_47_90
timestamp 1698431365
transform 1 0 11424 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_106
timestamp 1698431365
transform 1 0 13216 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_110
timestamp 1698431365
transform 1 0 13664 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_187
timestamp 1698431365
transform 1 0 22288 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_209
timestamp 1698431365
transform 1 0 24752 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_212
timestamp 1698431365
transform 1 0 25088 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_216
timestamp 1698431365
transform 1 0 25536 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_220
timestamp 1698431365
transform 1 0 25984 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_226
timestamp 1698431365
transform 1 0 26656 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_282
timestamp 1698431365
transform 1 0 32928 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_286
timestamp 1698431365
transform 1 0 33376 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_314
timestamp 1698431365
transform 1 0 36512 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_318
timestamp 1698431365
transform 1 0 36960 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_322
timestamp 1698431365
transform 1 0 37408 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_348
timestamp 1698431365
transform 1 0 40320 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_352
timestamp 1698431365
transform 1 0 40768 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_354
timestamp 1698431365
transform 1 0 40992 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_384
timestamp 1698431365
transform 1 0 44352 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_386
timestamp 1698431365
transform 1 0 44576 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_416
timestamp 1698431365
transform 1 0 47936 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_451
timestamp 1698431365
transform 1 0 51856 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_459
timestamp 1698431365
transform 1 0 52752 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_463
timestamp 1698431365
transform 1 0 53200 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_47_492
timestamp 1698431365
transform 1 0 56448 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_508
timestamp 1698431365
transform 1 0 58240 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_14
timestamp 1698431365
transform 1 0 2912 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_48_18
timestamp 1698431365
transform 1 0 3360 0 1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_34
timestamp 1698431365
transform 1 0 5152 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_48_37
timestamp 1698431365
transform 1 0 5488 0 1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_48_69
timestamp 1698431365
transform 1 0 9072 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_79
timestamp 1698431365
transform 1 0 10192 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_99
timestamp 1698431365
transform 1 0 12432 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_103
timestamp 1698431365
transform 1 0 12880 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_48_107
timestamp 1698431365
transform 1 0 13328 0 1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_123
timestamp 1698431365
transform 1 0 15120 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_48_139
timestamp 1698431365
transform 1 0 16912 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_147
timestamp 1698431365
transform 1 0 17808 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_151
timestamp 1698431365
transform 1 0 18256 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_168
timestamp 1698431365
transform 1 0 20160 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_172
timestamp 1698431365
transform 1 0 20608 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_174
timestamp 1698431365
transform 1 0 20832 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_177
timestamp 1698431365
transform 1 0 21168 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_181
timestamp 1698431365
transform 1 0 21616 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_186
timestamp 1698431365
transform 1 0 22176 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_188
timestamp 1698431365
transform 1 0 22400 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_195
timestamp 1698431365
transform 1 0 23184 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_205
timestamp 1698431365
transform 1 0 24304 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_207
timestamp 1698431365
transform 1 0 24528 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_236
timestamp 1698431365
transform 1 0 27776 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_240
timestamp 1698431365
transform 1 0 28224 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_242
timestamp 1698431365
transform 1 0 28448 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_48_280
timestamp 1698431365
transform 1 0 32704 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_288
timestamp 1698431365
transform 1 0 33600 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_292
timestamp 1698431365
transform 1 0 34048 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_296
timestamp 1698431365
transform 1 0 34496 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_300
timestamp 1698431365
transform 1 0 34944 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_48_304
timestamp 1698431365
transform 1 0 35392 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_312
timestamp 1698431365
transform 1 0 36288 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_314
timestamp 1698431365
transform 1 0 36512 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_48_317
timestamp 1698431365
transform 1 0 36848 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_325
timestamp 1698431365
transform 1 0 37744 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_327
timestamp 1698431365
transform 1 0 37968 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_48_330
timestamp 1698431365
transform 1 0 38304 0 1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_346
timestamp 1698431365
transform 1 0 40096 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_350
timestamp 1698431365
transform 1 0 40544 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_352
timestamp 1698431365
transform 1 0 40768 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_382
timestamp 1698431365
transform 1 0 44128 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_384
timestamp 1698431365
transform 1 0 44352 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_387
timestamp 1698431365
transform 1 0 44688 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_389
timestamp 1698431365
transform 1 0 44912 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_450
timestamp 1698431365
transform 1 0 51744 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_454
timestamp 1698431365
transform 1 0 52192 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_8
timestamp 1698431365
transform 1 0 2240 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_49_12
timestamp 1698431365
transform 1 0 2688 0 -1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_49_44
timestamp 1698431365
transform 1 0 6272 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_60
timestamp 1698431365
transform 1 0 8064 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_68
timestamp 1698431365
transform 1 0 8960 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_72
timestamp 1698431365
transform 1 0 9408 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_89
timestamp 1698431365
transform 1 0 11312 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_97
timestamp 1698431365
transform 1 0 12208 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_127
timestamp 1698431365
transform 1 0 15568 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_135
timestamp 1698431365
transform 1 0 16464 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_139
timestamp 1698431365
transform 1 0 16912 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_142
timestamp 1698431365
transform 1 0 17248 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_150
timestamp 1698431365
transform 1 0 18144 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_154
timestamp 1698431365
transform 1 0 18592 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_161
timestamp 1698431365
transform 1 0 19376 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_165
timestamp 1698431365
transform 1 0 19824 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_196
timestamp 1698431365
transform 1 0 23296 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_198
timestamp 1698431365
transform 1 0 23520 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_209
timestamp 1698431365
transform 1 0 24752 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_218
timestamp 1698431365
transform 1 0 25760 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_233
timestamp 1698431365
transform 1 0 27440 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_237
timestamp 1698431365
transform 1 0 27888 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_245
timestamp 1698431365
transform 1 0 28784 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_255
timestamp 1698431365
transform 1 0 29904 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_265
timestamp 1698431365
transform 1 0 31024 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_273
timestamp 1698431365
transform 1 0 31920 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_277
timestamp 1698431365
transform 1 0 32368 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_279
timestamp 1698431365
transform 1 0 32592 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_282
timestamp 1698431365
transform 1 0 32928 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_284
timestamp 1698431365
transform 1 0 33152 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_301
timestamp 1698431365
transform 1 0 35056 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_309
timestamp 1698431365
transform 1 0 35952 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_313
timestamp 1698431365
transform 1 0 36400 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_317
timestamp 1698431365
transform 1 0 36848 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_319
timestamp 1698431365
transform 1 0 37072 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_328
timestamp 1698431365
transform 1 0 38080 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_344
timestamp 1698431365
transform 1 0 39872 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_348
timestamp 1698431365
transform 1 0 40320 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_352
timestamp 1698431365
transform 1 0 40768 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_362
timestamp 1698431365
transform 1 0 41888 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_49_366
timestamp 1698431365
transform 1 0 42336 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_382
timestamp 1698431365
transform 1 0 44128 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_390
timestamp 1698431365
transform 1 0 45024 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_394
timestamp 1698431365
transform 1 0 45472 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_414
timestamp 1698431365
transform 1 0 47712 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_418
timestamp 1698431365
transform 1 0 48160 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_422
timestamp 1698431365
transform 1 0 48608 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_424
timestamp 1698431365
transform 1 0 48832 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_49_434
timestamp 1698431365
transform 1 0 49952 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_450
timestamp 1698431365
transform 1 0 51744 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_458
timestamp 1698431365
transform 1 0 52640 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_49_492
timestamp 1698431365
transform 1 0 56448 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_508
timestamp 1698431365
transform 1 0 58240 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_8
timestamp 1698431365
transform 1 0 2240 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_50_12
timestamp 1698431365
transform 1 0 2688 0 1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_28
timestamp 1698431365
transform 1 0 4480 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_32
timestamp 1698431365
transform 1 0 4928 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_34
timestamp 1698431365
transform 1 0 5152 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_50_37
timestamp 1698431365
transform 1 0 5488 0 1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_69
timestamp 1698431365
transform 1 0 9072 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_92
timestamp 1698431365
transform 1 0 11648 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_100
timestamp 1698431365
transform 1 0 12544 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_104
timestamp 1698431365
transform 1 0 12992 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_107
timestamp 1698431365
transform 1 0 13328 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_109
timestamp 1698431365
transform 1 0 13552 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_50_115
timestamp 1698431365
transform 1 0 14224 0 1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_131
timestamp 1698431365
transform 1 0 16016 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_139
timestamp 1698431365
transform 1 0 16912 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_143
timestamp 1698431365
transform 1 0 17360 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_155
timestamp 1698431365
transform 1 0 18704 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_157
timestamp 1698431365
transform 1 0 18928 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_168
timestamp 1698431365
transform 1 0 20160 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_172
timestamp 1698431365
transform 1 0 20608 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_177
timestamp 1698431365
transform 1 0 21168 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_215
timestamp 1698431365
transform 1 0 25424 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_240
timestamp 1698431365
transform 1 0 28224 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_244
timestamp 1698431365
transform 1 0 28672 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_247
timestamp 1698431365
transform 1 0 29008 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_249
timestamp 1698431365
transform 1 0 29232 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_258
timestamp 1698431365
transform 1 0 30240 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_260
timestamp 1698431365
transform 1 0 30464 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_275
timestamp 1698431365
transform 1 0 32144 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_277
timestamp 1698431365
transform 1 0 32368 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_304
timestamp 1698431365
transform 1 0 35392 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_306
timestamp 1698431365
transform 1 0 35616 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_323
timestamp 1698431365
transform 1 0 37520 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_372
timestamp 1698431365
transform 1 0 43008 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_380
timestamp 1698431365
transform 1 0 43904 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_384
timestamp 1698431365
transform 1 0 44352 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_434
timestamp 1698431365
transform 1 0 49952 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_442
timestamp 1698431365
transform 1 0 50848 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_450
timestamp 1698431365
transform 1 0 51744 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_454
timestamp 1698431365
transform 1 0 52192 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_50_457
timestamp 1698431365
transform 1 0 52528 0 1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_473
timestamp 1698431365
transform 1 0 54320 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_481
timestamp 1698431365
transform 1 0 55216 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_28
timestamp 1698431365
transform 1 0 4480 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_51_32
timestamp 1698431365
transform 1 0 4928 0 -1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_48
timestamp 1698431365
transform 1 0 6720 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_52
timestamp 1698431365
transform 1 0 7168 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_54
timestamp 1698431365
transform 1 0 7392 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_51_59
timestamp 1698431365
transform 1 0 7952 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_67
timestamp 1698431365
transform 1 0 8848 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_69
timestamp 1698431365
transform 1 0 9072 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_72
timestamp 1698431365
transform 1 0 9408 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_76
timestamp 1698431365
transform 1 0 9856 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_78
timestamp 1698431365
transform 1 0 10080 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_83
timestamp 1698431365
transform 1 0 10640 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_87
timestamp 1698431365
transform 1 0 11088 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_138
timestamp 1698431365
transform 1 0 16800 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_142
timestamp 1698431365
transform 1 0 17248 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_198
timestamp 1698431365
transform 1 0 23520 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_207
timestamp 1698431365
transform 1 0 24528 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_209
timestamp 1698431365
transform 1 0 24752 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_212
timestamp 1698431365
transform 1 0 25088 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_214
timestamp 1698431365
transform 1 0 25312 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_244
timestamp 1698431365
transform 1 0 28672 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_51_261
timestamp 1698431365
transform 1 0 30576 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_269
timestamp 1698431365
transform 1 0 31472 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_273
timestamp 1698431365
transform 1 0 31920 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_277
timestamp 1698431365
transform 1 0 32368 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_279
timestamp 1698431365
transform 1 0 32592 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_282
timestamp 1698431365
transform 1 0 32928 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_286
timestamp 1698431365
transform 1 0 33376 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_293
timestamp 1698431365
transform 1 0 34160 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_311
timestamp 1698431365
transform 1 0 36176 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_51_315
timestamp 1698431365
transform 1 0 36624 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_329
timestamp 1698431365
transform 1 0 38192 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_339
timestamp 1698431365
transform 1 0 39312 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_343
timestamp 1698431365
transform 1 0 39760 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_347
timestamp 1698431365
transform 1 0 40208 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_349
timestamp 1698431365
transform 1 0 40432 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_352
timestamp 1698431365
transform 1 0 40768 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_369
timestamp 1698431365
transform 1 0 42672 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_400
timestamp 1698431365
transform 1 0 46144 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_51_451
timestamp 1698431365
transform 1 0 51856 0 -1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_483
timestamp 1698431365
transform 1 0 55440 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_487
timestamp 1698431365
transform 1 0 55888 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_489
timestamp 1698431365
transform 1 0 56112 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_51_492
timestamp 1698431365
transform 1 0 56448 0 -1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_508
timestamp 1698431365
transform 1 0 58240 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_8
timestamp 1698431365
transform 1 0 2240 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_52_12
timestamp 1698431365
transform 1 0 2688 0 1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_28
timestamp 1698431365
transform 1 0 4480 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_32
timestamp 1698431365
transform 1 0 4928 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_34
timestamp 1698431365
transform 1 0 5152 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_37
timestamp 1698431365
transform 1 0 5488 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_52_71
timestamp 1698431365
transform 1 0 9296 0 1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_107
timestamp 1698431365
transform 1 0 13328 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_109
timestamp 1698431365
transform 1 0 13552 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_170
timestamp 1698431365
transform 1 0 20384 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_174
timestamp 1698431365
transform 1 0 20832 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_183
timestamp 1698431365
transform 1 0 21840 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_187
timestamp 1698431365
transform 1 0 22288 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_52_191
timestamp 1698431365
transform 1 0 22736 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_199
timestamp 1698431365
transform 1 0 23632 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_52_215
timestamp 1698431365
transform 1 0 25424 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_243
timestamp 1698431365
transform 1 0 28560 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_247
timestamp 1698431365
transform 1 0 29008 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_52_251
timestamp 1698431365
transform 1 0 29456 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_288
timestamp 1698431365
transform 1 0 33600 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_294
timestamp 1698431365
transform 1 0 34272 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_298
timestamp 1698431365
transform 1 0 34720 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_306
timestamp 1698431365
transform 1 0 35616 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_310
timestamp 1698431365
transform 1 0 36064 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_314
timestamp 1698431365
transform 1 0 36512 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_52_317
timestamp 1698431365
transform 1 0 36848 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_325
timestamp 1698431365
transform 1 0 37744 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_52_335
timestamp 1698431365
transform 1 0 38864 0 1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_52_351
timestamp 1698431365
transform 1 0 40656 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_52_361
timestamp 1698431365
transform 1 0 41776 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_369
timestamp 1698431365
transform 1 0 42672 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_373
timestamp 1698431365
transform 1 0 43120 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_52_377
timestamp 1698431365
transform 1 0 43568 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_387
timestamp 1698431365
transform 1 0 44688 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_391
timestamp 1698431365
transform 1 0 45136 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_52_395
timestamp 1698431365
transform 1 0 45584 0 1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_411
timestamp 1698431365
transform 1 0 47376 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_415
timestamp 1698431365
transform 1 0 47824 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_417
timestamp 1698431365
transform 1 0 48048 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_52_434
timestamp 1698431365
transform 1 0 49952 0 1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_450
timestamp 1698431365
transform 1 0 51744 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_454
timestamp 1698431365
transform 1 0 52192 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_52_457
timestamp 1698431365
transform 1 0 52528 0 1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_52_473
timestamp 1698431365
transform 1 0 54320 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_481
timestamp 1698431365
transform 1 0 55216 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_8
timestamp 1698431365
transform 1 0 2240 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_53_12
timestamp 1698431365
transform 1 0 2688 0 -1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_28
timestamp 1698431365
transform 1 0 4480 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_32
timestamp 1698431365
transform 1 0 4928 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_62
timestamp 1698431365
transform 1 0 8288 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_64
timestamp 1698431365
transform 1 0 8512 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_101
timestamp 1698431365
transform 1 0 12656 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_142
timestamp 1698431365
transform 1 0 17248 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_144
timestamp 1698431365
transform 1 0 17472 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_212
timestamp 1698431365
transform 1 0 25088 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_53_216
timestamp 1698431365
transform 1 0 25536 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_224
timestamp 1698431365
transform 1 0 26432 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_236
timestamp 1698431365
transform 1 0 27776 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_53_255
timestamp 1698431365
transform 1 0 29904 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_282
timestamp 1698431365
transform 1 0 32928 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_294
timestamp 1698431365
transform 1 0 34272 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_327
timestamp 1698431365
transform 1 0 37968 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_53_337
timestamp 1698431365
transform 1 0 39088 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_345
timestamp 1698431365
transform 1 0 39984 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_349
timestamp 1698431365
transform 1 0 40432 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_400
timestamp 1698431365
transform 1 0 46144 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_53_404
timestamp 1698431365
transform 1 0 46592 0 -1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_53_422
timestamp 1698431365
transform 1 0 48608 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_486
timestamp 1698431365
transform 1 0 55776 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_53_492
timestamp 1698431365
transform 1 0 56448 0 -1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_508
timestamp 1698431365
transform 1 0 58240 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_14
timestamp 1698431365
transform 1 0 2912 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_54_18
timestamp 1698431365
transform 1 0 3360 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_34
timestamp 1698431365
transform 1 0 5152 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_37
timestamp 1698431365
transform 1 0 5488 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_41
timestamp 1698431365
transform 1 0 5936 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_71
timestamp 1698431365
transform 1 0 9296 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_75
timestamp 1698431365
transform 1 0 9744 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_94
timestamp 1698431365
transform 1 0 11872 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_98
timestamp 1698431365
transform 1 0 12320 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_107
timestamp 1698431365
transform 1 0 13328 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_138
timestamp 1698431365
transform 1 0 16800 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_177
timestamp 1698431365
transform 1 0 21168 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_191
timestamp 1698431365
transform 1 0 22736 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_54_202
timestamp 1698431365
transform 1 0 23968 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_218
timestamp 1698431365
transform 1 0 25760 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_226
timestamp 1698431365
transform 1 0 26656 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_230
timestamp 1698431365
transform 1 0 27104 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_247
timestamp 1698431365
transform 1 0 29008 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_372
timestamp 1698431365
transform 1 0 43008 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_383
timestamp 1698431365
transform 1 0 44240 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_395
timestamp 1698431365
transform 1 0 45584 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_399
timestamp 1698431365
transform 1 0 46032 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_54_430
timestamp 1698431365
transform 1 0 49504 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_446
timestamp 1698431365
transform 1 0 51296 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_454
timestamp 1698431365
transform 1 0 52192 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_8
timestamp 1698431365
transform 1 0 2240 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_12
timestamp 1698431365
transform 1 0 2688 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_55_16
timestamp 1698431365
transform 1 0 3136 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_24
timestamp 1698431365
transform 1 0 4032 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_26
timestamp 1698431365
transform 1 0 4256 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_65
timestamp 1698431365
transform 1 0 8624 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_69
timestamp 1698431365
transform 1 0 9072 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_55_101
timestamp 1698431365
transform 1 0 12656 0 -1 47040
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_133
timestamp 1698431365
transform 1 0 16240 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_137
timestamp 1698431365
transform 1 0 16688 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_142
timestamp 1698431365
transform 1 0 17248 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_216
timestamp 1698431365
transform 1 0 25536 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_220
timestamp 1698431365
transform 1 0 25984 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_240
timestamp 1698431365
transform 1 0 28224 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_246
timestamp 1698431365
transform 1 0 28896 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_248
timestamp 1698431365
transform 1 0 29120 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_278
timestamp 1698431365
transform 1 0 32480 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_282
timestamp 1698431365
transform 1 0 32928 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_304
timestamp 1698431365
transform 1 0 35392 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_314
timestamp 1698431365
transform 1 0 36512 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_318
timestamp 1698431365
transform 1 0 36960 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_320
timestamp 1698431365
transform 1 0 37184 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_391
timestamp 1698431365
transform 1 0 45136 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_393
timestamp 1698431365
transform 1 0 45360 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_418
timestamp 1698431365
transform 1 0 48160 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_55_422
timestamp 1698431365
transform 1 0 48608 0 -1 47040
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_55_454
timestamp 1698431365
transform 1 0 52192 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_55_492
timestamp 1698431365
transform 1 0 56448 0 -1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_508
timestamp 1698431365
transform 1 0 58240 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_28
timestamp 1698431365
transform 1 0 4480 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_32
timestamp 1698431365
transform 1 0 4928 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_34
timestamp 1698431365
transform 1 0 5152 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_96
timestamp 1698431365
transform 1 0 12096 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_104
timestamp 1698431365
transform 1 0 12992 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_107
timestamp 1698431365
transform 1 0 13328 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_111
timestamp 1698431365
transform 1 0 13776 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_56_119
timestamp 1698431365
transform 1 0 14672 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_127
timestamp 1698431365
transform 1 0 15568 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_129
timestamp 1698431365
transform 1 0 15792 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_161
timestamp 1698431365
transform 1 0 19376 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_165
timestamp 1698431365
transform 1 0 19824 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_169
timestamp 1698431365
transform 1 0 20272 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_173
timestamp 1698431365
transform 1 0 20720 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_177
timestamp 1698431365
transform 1 0 21168 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_192
timestamp 1698431365
transform 1 0 22848 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_201
timestamp 1698431365
transform 1 0 23856 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_205
timestamp 1698431365
transform 1 0 24304 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_247
timestamp 1698431365
transform 1 0 29008 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_285
timestamp 1698431365
transform 1 0 33264 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_287
timestamp 1698431365
transform 1 0 33488 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_312
timestamp 1698431365
transform 1 0 36288 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_314
timestamp 1698431365
transform 1 0 36512 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_333
timestamp 1698431365
transform 1 0 38640 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_359
timestamp 1698431365
transform 1 0 41552 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_363
timestamp 1698431365
transform 1 0 42000 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_387
timestamp 1698431365
transform 1 0 44688 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_417
timestamp 1698431365
transform 1 0 48048 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_421
timestamp 1698431365
transform 1 0 48496 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_56_425
timestamp 1698431365
transform 1 0 48944 0 1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_56_441
timestamp 1698431365
transform 1 0 50736 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_449
timestamp 1698431365
transform 1 0 51632 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_453
timestamp 1698431365
transform 1 0 52080 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_56_457
timestamp 1698431365
transform 1 0 52528 0 1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_56_473
timestamp 1698431365
transform 1 0 54320 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_481
timestamp 1698431365
transform 1 0 55216 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_28
timestamp 1698431365
transform 1 0 4480 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_57_32
timestamp 1698431365
transform 1 0 4928 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_40
timestamp 1698431365
transform 1 0 5824 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_42
timestamp 1698431365
transform 1 0 6048 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_62
timestamp 1698431365
transform 1 0 8288 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_72
timestamp 1698431365
transform 1 0 9408 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_81
timestamp 1698431365
transform 1 0 10416 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_85
timestamp 1698431365
transform 1 0 10864 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_89
timestamp 1698431365
transform 1 0 11312 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_95
timestamp 1698431365
transform 1 0 11984 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_97
timestamp 1698431365
transform 1 0 12208 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_133
timestamp 1698431365
transform 1 0 16240 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_135
timestamp 1698431365
transform 1 0 16464 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_151
timestamp 1698431365
transform 1 0 18256 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_57_155
timestamp 1698431365
transform 1 0 18704 0 -1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_171
timestamp 1698431365
transform 1 0 20496 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_173
timestamp 1698431365
transform 1 0 20720 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_190
timestamp 1698431365
transform 1 0 22624 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_194
timestamp 1698431365
transform 1 0 23072 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_198
timestamp 1698431365
transform 1 0 23520 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_262
timestamp 1698431365
transform 1 0 30688 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_276
timestamp 1698431365
transform 1 0 32256 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_325
timestamp 1698431365
transform 1 0 37744 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_349
timestamp 1698431365
transform 1 0 40432 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_356
timestamp 1698431365
transform 1 0 41216 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_360
timestamp 1698431365
transform 1 0 41664 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_364
timestamp 1698431365
transform 1 0 42112 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_368
timestamp 1698431365
transform 1 0 42560 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_370
timestamp 1698431365
transform 1 0 42784 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_382
timestamp 1698431365
transform 1 0 44128 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_386
timestamp 1698431365
transform 1 0 44576 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_390
timestamp 1698431365
transform 1 0 45024 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_57_422
timestamp 1698431365
transform 1 0 48608 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_486
timestamp 1698431365
transform 1 0 55776 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_57_492
timestamp 1698431365
transform 1 0 56448 0 -1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_508
timestamp 1698431365
transform 1 0 58240 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_28
timestamp 1698431365
transform 1 0 4480 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_32
timestamp 1698431365
transform 1 0 4928 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_34
timestamp 1698431365
transform 1 0 5152 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_70
timestamp 1698431365
transform 1 0 9184 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_116
timestamp 1698431365
transform 1 0 14336 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_155
timestamp 1698431365
transform 1 0 18704 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_157
timestamp 1698431365
transform 1 0 18928 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_160
timestamp 1698431365
transform 1 0 19264 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_177
timestamp 1698431365
transform 1 0 21168 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_58_181
timestamp 1698431365
transform 1 0 21616 0 1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_226
timestamp 1698431365
transform 1 0 26656 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_242
timestamp 1698431365
transform 1 0 28448 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_244
timestamp 1698431365
transform 1 0 28672 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_281
timestamp 1698431365
transform 1 0 32816 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_291
timestamp 1698431365
transform 1 0 33936 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_293
timestamp 1698431365
transform 1 0 34160 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_302
timestamp 1698431365
transform 1 0 35168 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_304
timestamp 1698431365
transform 1 0 35392 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_330
timestamp 1698431365
transform 1 0 38304 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_332
timestamp 1698431365
transform 1 0 38528 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_345
timestamp 1698431365
transform 1 0 39984 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_349
timestamp 1698431365
transform 1 0 40432 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_353
timestamp 1698431365
transform 1 0 40880 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_375
timestamp 1698431365
transform 1 0 43344 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_384
timestamp 1698431365
transform 1 0 44352 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_387
timestamp 1698431365
transform 1 0 44688 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_58_440
timestamp 1698431365
transform 1 0 50624 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_448
timestamp 1698431365
transform 1 0 51520 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_452
timestamp 1698431365
transform 1 0 51968 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_454
timestamp 1698431365
transform 1 0 52192 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_58_457
timestamp 1698431365
transform 1 0 52528 0 1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_58_489
timestamp 1698431365
transform 1 0 56112 0 1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_505
timestamp 1698431365
transform 1 0 57904 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_8
timestamp 1698431365
transform 1 0 2240 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_59_12
timestamp 1698431365
transform 1 0 2688 0 -1 50176
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_44
timestamp 1698431365
transform 1 0 6272 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_48
timestamp 1698431365
transform 1 0 6720 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_66
timestamp 1698431365
transform 1 0 8736 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_139
timestamp 1698431365
transform 1 0 16912 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_142
timestamp 1698431365
transform 1 0 17248 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_59_188
timestamp 1698431365
transform 1 0 22400 0 -1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_204
timestamp 1698431365
transform 1 0 24192 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_208
timestamp 1698431365
transform 1 0 24640 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_216
timestamp 1698431365
transform 1 0 25536 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_220
timestamp 1698431365
transform 1 0 25984 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_242
timestamp 1698431365
transform 1 0 28448 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_246
timestamp 1698431365
transform 1 0 28896 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_250
timestamp 1698431365
transform 1 0 29344 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_254
timestamp 1698431365
transform 1 0 29792 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_263
timestamp 1698431365
transform 1 0 30800 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_273
timestamp 1698431365
transform 1 0 31920 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_277
timestamp 1698431365
transform 1 0 32368 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_279
timestamp 1698431365
transform 1 0 32592 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_59_282
timestamp 1698431365
transform 1 0 32928 0 -1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_305
timestamp 1698431365
transform 1 0 35504 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_309
timestamp 1698431365
transform 1 0 35952 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_331
timestamp 1698431365
transform 1 0 38416 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_335
timestamp 1698431365
transform 1 0 38864 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_349
timestamp 1698431365
transform 1 0 40432 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_59_352
timestamp 1698431365
transform 1 0 40768 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_360
timestamp 1698431365
transform 1 0 41664 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_362
timestamp 1698431365
transform 1 0 41888 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_368
timestamp 1698431365
transform 1 0 42560 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_388
timestamp 1698431365
transform 1 0 44800 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_392
timestamp 1698431365
transform 1 0 45248 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_395
timestamp 1698431365
transform 1 0 45584 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_59_399
timestamp 1698431365
transform 1 0 46032 0 -1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_415
timestamp 1698431365
transform 1 0 47824 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_419
timestamp 1698431365
transform 1 0 48272 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_422
timestamp 1698431365
transform 1 0 48608 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_426
timestamp 1698431365
transform 1 0 49056 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_59_480
timestamp 1698431365
transform 1 0 55104 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_488
timestamp 1698431365
transform 1 0 56000 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_59_492
timestamp 1698431365
transform 1 0 56448 0 -1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_508
timestamp 1698431365
transform 1 0 58240 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_14
timestamp 1698431365
transform 1 0 2912 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_60_18
timestamp 1698431365
transform 1 0 3360 0 1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_34
timestamp 1698431365
transform 1 0 5152 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_60_37
timestamp 1698431365
transform 1 0 5488 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_45
timestamp 1698431365
transform 1 0 6384 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_60_54
timestamp 1698431365
transform 1 0 7392 0 1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_70
timestamp 1698431365
transform 1 0 9184 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_92
timestamp 1698431365
transform 1 0 11648 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_94
timestamp 1698431365
transform 1 0 11872 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_113
timestamp 1698431365
transform 1 0 14000 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_115
timestamp 1698431365
transform 1 0 14224 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_193
timestamp 1698431365
transform 1 0 22960 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_197
timestamp 1698431365
transform 1 0 23408 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_60_201
timestamp 1698431365
transform 1 0 23856 0 1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_217
timestamp 1698431365
transform 1 0 25648 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_221
timestamp 1698431365
transform 1 0 26096 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_60_230
timestamp 1698431365
transform 1 0 27104 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_238
timestamp 1698431365
transform 1 0 28000 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_242
timestamp 1698431365
transform 1 0 28448 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_244
timestamp 1698431365
transform 1 0 28672 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_247
timestamp 1698431365
transform 1 0 29008 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_251
timestamp 1698431365
transform 1 0 29456 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_253
timestamp 1698431365
transform 1 0 29680 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_258
timestamp 1698431365
transform 1 0 30240 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_262
timestamp 1698431365
transform 1 0 30688 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_60_269
timestamp 1698431365
transform 1 0 31472 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_277
timestamp 1698431365
transform 1 0 32368 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_281
timestamp 1698431365
transform 1 0 32816 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_283
timestamp 1698431365
transform 1 0 33040 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_60_292
timestamp 1698431365
transform 1 0 34048 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_300
timestamp 1698431365
transform 1 0 34944 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_304
timestamp 1698431365
transform 1 0 35392 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_364
timestamp 1698431365
transform 1 0 42112 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_368
timestamp 1698431365
transform 1 0 42560 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_372
timestamp 1698431365
transform 1 0 43008 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_383
timestamp 1698431365
transform 1 0 44240 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_60_387
timestamp 1698431365
transform 1 0 44688 0 1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_403
timestamp 1698431365
transform 1 0 46480 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_60_436
timestamp 1698431365
transform 1 0 50176 0 1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_452
timestamp 1698431365
transform 1 0 51968 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_454
timestamp 1698431365
transform 1 0 52192 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_60_457
timestamp 1698431365
transform 1 0 52528 0 1 50176
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_60_489
timestamp 1698431365
transform 1 0 56112 0 1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_505
timestamp 1698431365
transform 1 0 57904 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_8
timestamp 1698431365
transform 1 0 2240 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_12
timestamp 1698431365
transform 1 0 2688 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_61_16
timestamp 1698431365
transform 1 0 3136 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_24
timestamp 1698431365
transform 1 0 4032 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_26
timestamp 1698431365
transform 1 0 4256 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_61_56
timestamp 1698431365
transform 1 0 7616 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_64
timestamp 1698431365
transform 1 0 8512 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_68
timestamp 1698431365
transform 1 0 8960 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_72
timestamp 1698431365
transform 1 0 9408 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_74
timestamp 1698431365
transform 1 0 9632 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_142
timestamp 1698431365
transform 1 0 17248 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_154
timestamp 1698431365
transform 1 0 18592 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_158
timestamp 1698431365
transform 1 0 19040 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_202
timestamp 1698431365
transform 1 0 23968 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_206
timestamp 1698431365
transform 1 0 24416 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_274
timestamp 1698431365
transform 1 0 32032 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_278
timestamp 1698431365
transform 1 0 32480 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_282
timestamp 1698431365
transform 1 0 32928 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_318
timestamp 1698431365
transform 1 0 36960 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_322
timestamp 1698431365
transform 1 0 37408 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_324
timestamp 1698431365
transform 1 0 37632 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_348
timestamp 1698431365
transform 1 0 40320 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_352
timestamp 1698431365
transform 1 0 40768 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_354
timestamp 1698431365
transform 1 0 40992 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_384
timestamp 1698431365
transform 1 0 44352 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_386
timestamp 1698431365
transform 1 0 44576 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_395
timestamp 1698431365
transform 1 0 45584 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_430
timestamp 1698431365
transform 1 0 49504 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_61_434
timestamp 1698431365
transform 1 0 49952 0 -1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_61_466
timestamp 1698431365
transform 1 0 53536 0 -1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_61_482
timestamp 1698431365
transform 1 0 55328 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_61_492
timestamp 1698431365
transform 1 0 56448 0 -1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_508
timestamp 1698431365
transform 1 0 58240 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_8
timestamp 1698431365
transform 1 0 2240 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_62_12
timestamp 1698431365
transform 1 0 2688 0 1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_28
timestamp 1698431365
transform 1 0 4480 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_32
timestamp 1698431365
transform 1 0 4928 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_34
timestamp 1698431365
transform 1 0 5152 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_62_37
timestamp 1698431365
transform 1 0 5488 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_62_63
timestamp 1698431365
transform 1 0 8400 0 1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_79
timestamp 1698431365
transform 1 0 10192 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_83
timestamp 1698431365
transform 1 0 10640 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_85
timestamp 1698431365
transform 1 0 10864 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_97
timestamp 1698431365
transform 1 0 12208 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_101
timestamp 1698431365
transform 1 0 12656 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_107
timestamp 1698431365
transform 1 0 13328 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_109
timestamp 1698431365
transform 1 0 13552 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_145
timestamp 1698431365
transform 1 0 17584 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_147
timestamp 1698431365
transform 1 0 17808 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_174
timestamp 1698431365
transform 1 0 20832 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_177
timestamp 1698431365
transform 1 0 21168 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_181
timestamp 1698431365
transform 1 0 21616 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_196
timestamp 1698431365
transform 1 0 23296 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_200
timestamp 1698431365
transform 1 0 23744 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_207
timestamp 1698431365
transform 1 0 24528 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_211
timestamp 1698431365
transform 1 0 24976 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_62_267
timestamp 1698431365
transform 1 0 31248 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_275
timestamp 1698431365
transform 1 0 32144 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_282
timestamp 1698431365
transform 1 0 32928 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_292
timestamp 1698431365
transform 1 0 34048 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_296
timestamp 1698431365
transform 1 0 34496 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_62_301
timestamp 1698431365
transform 1 0 35056 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_309
timestamp 1698431365
transform 1 0 35952 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_313
timestamp 1698431365
transform 1 0 36400 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_62_317
timestamp 1698431365
transform 1 0 36848 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_325
timestamp 1698431365
transform 1 0 37744 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_327
timestamp 1698431365
transform 1 0 37968 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_62_348
timestamp 1698431365
transform 1 0 40320 0 1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_380
timestamp 1698431365
transform 1 0 43904 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_382
timestamp 1698431365
transform 1 0 44128 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_62_437
timestamp 1698431365
transform 1 0 50288 0 1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_453
timestamp 1698431365
transform 1 0 52080 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_62_457
timestamp 1698431365
transform 1 0 52528 0 1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_62_489
timestamp 1698431365
transform 1 0 56112 0 1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_505
timestamp 1698431365
transform 1 0 57904 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_8
timestamp 1698431365
transform 1 0 2240 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_63_12
timestamp 1698431365
transform 1 0 2688 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_20
timestamp 1698431365
transform 1 0 3584 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_24
timestamp 1698431365
transform 1 0 4032 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_26
timestamp 1698431365
transform 1 0 4256 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_68
timestamp 1698431365
transform 1 0 8960 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_72
timestamp 1698431365
transform 1 0 9408 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_63_79
timestamp 1698431365
transform 1 0 10192 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_87
timestamp 1698431365
transform 1 0 11088 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_63_97
timestamp 1698431365
transform 1 0 12208 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_105
timestamp 1698431365
transform 1 0 13104 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_107
timestamp 1698431365
transform 1 0 13328 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_132
timestamp 1698431365
transform 1 0 16128 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_185
timestamp 1698431365
transform 1 0 22064 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_189
timestamp 1698431365
transform 1 0 22512 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_197
timestamp 1698431365
transform 1 0 23408 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_199
timestamp 1698431365
transform 1 0 23632 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_212
timestamp 1698431365
transform 1 0 25088 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_228
timestamp 1698431365
transform 1 0 26880 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_238
timestamp 1698431365
transform 1 0 28000 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_252
timestamp 1698431365
transform 1 0 29568 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_254
timestamp 1698431365
transform 1 0 29792 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_269
timestamp 1698431365
transform 1 0 31472 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_278
timestamp 1698431365
transform 1 0 32480 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_288
timestamp 1698431365
transform 1 0 33600 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_292
timestamp 1698431365
transform 1 0 34048 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_306
timestamp 1698431365
transform 1 0 35616 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_310
timestamp 1698431365
transform 1 0 36064 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_312
timestamp 1698431365
transform 1 0 36288 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_63_325
timestamp 1698431365
transform 1 0 37744 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_333
timestamp 1698431365
transform 1 0 38640 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_335
timestamp 1698431365
transform 1 0 38864 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_344
timestamp 1698431365
transform 1 0 39872 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_348
timestamp 1698431365
transform 1 0 40320 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_63_352
timestamp 1698431365
transform 1 0 40768 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_360
timestamp 1698431365
transform 1 0 41664 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_364
timestamp 1698431365
transform 1 0 42112 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_63_376
timestamp 1698431365
transform 1 0 43456 0 -1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_392
timestamp 1698431365
transform 1 0 45248 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_422
timestamp 1698431365
transform 1 0 48608 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_424
timestamp 1698431365
transform 1 0 48832 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_63_431
timestamp 1698431365
transform 1 0 49616 0 -1 53312
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_63_463
timestamp 1698431365
transform 1 0 53200 0 -1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_63_479
timestamp 1698431365
transform 1 0 54992 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_487
timestamp 1698431365
transform 1 0 55888 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_489
timestamp 1698431365
transform 1 0 56112 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_63_492
timestamp 1698431365
transform 1 0 56448 0 -1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_508
timestamp 1698431365
transform 1 0 58240 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_8
timestamp 1698431365
transform 1 0 2240 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_64_12
timestamp 1698431365
transform 1 0 2688 0 1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_28
timestamp 1698431365
transform 1 0 4480 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_32
timestamp 1698431365
transform 1 0 4928 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_34
timestamp 1698431365
transform 1 0 5152 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_64_37
timestamp 1698431365
transform 1 0 5488 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_64_63
timestamp 1698431365
transform 1 0 8400 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_64_90
timestamp 1698431365
transform 1 0 11424 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_98
timestamp 1698431365
transform 1 0 12320 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_102
timestamp 1698431365
transform 1 0 12768 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_104
timestamp 1698431365
transform 1 0 12992 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_64_107
timestamp 1698431365
transform 1 0 13328 0 1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_64_123
timestamp 1698431365
transform 1 0 15120 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_131
timestamp 1698431365
transform 1 0 16016 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_137
timestamp 1698431365
transform 1 0 16688 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_141
timestamp 1698431365
transform 1 0 17136 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_143
timestamp 1698431365
transform 1 0 17360 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_234
timestamp 1698431365
transform 1 0 27552 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_242
timestamp 1698431365
transform 1 0 28448 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_244
timestamp 1698431365
transform 1 0 28672 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_247
timestamp 1698431365
transform 1 0 29008 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_251
timestamp 1698431365
transform 1 0 29456 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_64_261
timestamp 1698431365
transform 1 0 30576 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_314
timestamp 1698431365
transform 1 0 36512 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_64_330
timestamp 1698431365
transform 1 0 38304 0 1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_64_391
timestamp 1698431365
transform 1 0 45136 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_399
timestamp 1698431365
transform 1 0 46032 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_401
timestamp 1698431365
transform 1 0 46256 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_410
timestamp 1698431365
transform 1 0 47264 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_440
timestamp 1698431365
transform 1 0 50624 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_64_444
timestamp 1698431365
transform 1 0 51072 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_452
timestamp 1698431365
transform 1 0 51968 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_454
timestamp 1698431365
transform 1 0 52192 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_64_457
timestamp 1698431365
transform 1 0 52528 0 1 53312
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_64_489
timestamp 1698431365
transform 1 0 56112 0 1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_505
timestamp 1698431365
transform 1 0 57904 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_8
timestamp 1698431365
transform 1 0 2240 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_65_12
timestamp 1698431365
transform 1 0 2688 0 -1 54880
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_44
timestamp 1698431365
transform 1 0 6272 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_59
timestamp 1698431365
transform 1 0 7952 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_63
timestamp 1698431365
transform 1 0 8400 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_65_101
timestamp 1698431365
transform 1 0 12656 0 -1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_117
timestamp 1698431365
transform 1 0 14448 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_130
timestamp 1698431365
transform 1 0 15904 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_137
timestamp 1698431365
transform 1 0 16688 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_139
timestamp 1698431365
transform 1 0 16912 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_142
timestamp 1698431365
transform 1 0 17248 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_146
timestamp 1698431365
transform 1 0 17696 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_150
timestamp 1698431365
transform 1 0 18144 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_204
timestamp 1698431365
transform 1 0 24192 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_231
timestamp 1698431365
transform 1 0 27216 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_235
timestamp 1698431365
transform 1 0 27664 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_239
timestamp 1698431365
transform 1 0 28112 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_243
timestamp 1698431365
transform 1 0 28560 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_247
timestamp 1698431365
transform 1 0 29008 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_268
timestamp 1698431365
transform 1 0 31360 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_270
timestamp 1698431365
transform 1 0 31584 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_277
timestamp 1698431365
transform 1 0 32368 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_279
timestamp 1698431365
transform 1 0 32592 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_282
timestamp 1698431365
transform 1 0 32928 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_288
timestamp 1698431365
transform 1 0 33600 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_344
timestamp 1698431365
transform 1 0 39872 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_348
timestamp 1698431365
transform 1 0 40320 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_410
timestamp 1698431365
transform 1 0 47264 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_65_451
timestamp 1698431365
transform 1 0 51856 0 -1 54880
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_483
timestamp 1698431365
transform 1 0 55440 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_487
timestamp 1698431365
transform 1 0 55888 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_489
timestamp 1698431365
transform 1 0 56112 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_65_492
timestamp 1698431365
transform 1 0 56448 0 -1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_508
timestamp 1698431365
transform 1 0 58240 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_66_2
timestamp 1698431365
transform 1 0 1568 0 1 54880
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_34
timestamp 1698431365
transform 1 0 5152 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_66
timestamp 1698431365
transform 1 0 8736 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_99
timestamp 1698431365
transform 1 0 12432 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_103
timestamp 1698431365
transform 1 0 12880 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_136
timestamp 1698431365
transform 1 0 16576 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_140
timestamp 1698431365
transform 1 0 17024 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_150
timestamp 1698431365
transform 1 0 18144 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_66_154
timestamp 1698431365
transform 1 0 18592 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_162
timestamp 1698431365
transform 1 0 19488 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_168
timestamp 1698431365
transform 1 0 20160 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_174
timestamp 1698431365
transform 1 0 20832 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_233
timestamp 1698431365
transform 1 0 27440 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_251
timestamp 1698431365
transform 1 0 29456 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_253
timestamp 1698431365
transform 1 0 29680 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_260
timestamp 1698431365
transform 1 0 30464 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_264
timestamp 1698431365
transform 1 0 30912 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_66_279
timestamp 1698431365
transform 1 0 32592 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_287
timestamp 1698431365
transform 1 0 33488 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_289
timestamp 1698431365
transform 1 0 33712 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_298
timestamp 1698431365
transform 1 0 34720 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_346
timestamp 1698431365
transform 1 0 40096 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_350
timestamp 1698431365
transform 1 0 40544 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_352
timestamp 1698431365
transform 1 0 40768 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_387
timestamp 1698431365
transform 1 0 44688 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_389
timestamp 1698431365
transform 1 0 44912 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_66_440
timestamp 1698431365
transform 1 0 50624 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_448
timestamp 1698431365
transform 1 0 51520 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_452
timestamp 1698431365
transform 1 0 51968 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_454
timestamp 1698431365
transform 1 0 52192 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_66_457
timestamp 1698431365
transform 1 0 52528 0 1 54880
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_66_489
timestamp 1698431365
transform 1 0 56112 0 1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_505
timestamp 1698431365
transform 1 0 57904 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_67_2
timestamp 1698431365
transform 1 0 1568 0 -1 56448
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_34
timestamp 1698431365
transform 1 0 5152 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_42
timestamp 1698431365
transform 1 0 6048 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_46
timestamp 1698431365
transform 1 0 6496 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_72
timestamp 1698431365
transform 1 0 9408 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_74
timestamp 1698431365
transform 1 0 9632 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_84
timestamp 1698431365
transform 1 0 10752 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_86
timestamp 1698431365
transform 1 0 10976 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_93
timestamp 1698431365
transform 1 0 11760 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_95
timestamp 1698431365
transform 1 0 11984 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_139
timestamp 1698431365
transform 1 0 16912 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_146
timestamp 1698431365
transform 1 0 17696 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_67_150
timestamp 1698431365
transform 1 0 18144 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_166
timestamp 1698431365
transform 1 0 19936 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_172
timestamp 1698431365
transform 1 0 20608 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_182
timestamp 1698431365
transform 1 0 21728 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_192
timestamp 1698431365
transform 1 0 22848 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_209
timestamp 1698431365
transform 1 0 24752 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_220
timestamp 1698431365
transform 1 0 25984 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_253
timestamp 1698431365
transform 1 0 29680 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_257
timestamp 1698431365
transform 1 0 30128 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_261
timestamp 1698431365
transform 1 0 30576 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_269
timestamp 1698431365
transform 1 0 31472 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_273
timestamp 1698431365
transform 1 0 31920 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_277
timestamp 1698431365
transform 1 0 32368 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_346
timestamp 1698431365
transform 1 0 40096 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_352
timestamp 1698431365
transform 1 0 40768 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_356
timestamp 1698431365
transform 1 0 41216 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_364
timestamp 1698431365
transform 1 0 42112 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_375
timestamp 1698431365
transform 1 0 43344 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_400
timestamp 1698431365
transform 1 0 46144 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_404
timestamp 1698431365
transform 1 0 46592 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_408
timestamp 1698431365
transform 1 0 47040 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_419
timestamp 1698431365
transform 1 0 48272 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_67_432
timestamp 1698431365
transform 1 0 49728 0 -1 56448
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_67_464
timestamp 1698431365
transform 1 0 53312 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_480
timestamp 1698431365
transform 1 0 55104 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_488
timestamp 1698431365
transform 1 0 56000 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_67_492
timestamp 1698431365
transform 1 0 56448 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_508
timestamp 1698431365
transform 1 0 58240 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_68_2
timestamp 1698431365
transform 1 0 1568 0 1 56448
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_68_34
timestamp 1698431365
transform 1 0 5152 0 1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_75
timestamp 1698431365
transform 1 0 9744 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_68_95
timestamp 1698431365
transform 1 0 11984 0 1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_103
timestamp 1698431365
transform 1 0 12880 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_107
timestamp 1698431365
transform 1 0 13328 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_68_119
timestamp 1698431365
transform 1 0 14672 0 1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_68_163
timestamp 1698431365
transform 1 0 19600 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_68_167
timestamp 1698431365
transform 1 0 20048 0 1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_172
timestamp 1698431365
transform 1 0 20608 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_68_174
timestamp 1698431365
transform 1 0 20832 0 1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_182
timestamp 1698431365
transform 1 0 21728 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_68_184
timestamp 1698431365
transform 1 0 21952 0 1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_212
timestamp 1698431365
transform 1 0 25088 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_253
timestamp 1698431365
transform 1 0 29680 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_68_255
timestamp 1698431365
transform 1 0 29904 0 1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_262
timestamp 1698431365
transform 1 0 30688 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_266
timestamp 1698431365
transform 1 0 31136 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_68_268
timestamp 1698431365
transform 1 0 31360 0 1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_68_289
timestamp 1698431365
transform 1 0 33712 0 1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_68_304
timestamp 1698431365
transform 1 0 35392 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_308
timestamp 1698431365
transform 1 0 35840 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_68_310
timestamp 1698431365
transform 1 0 36064 0 1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_68_325
timestamp 1698431365
transform 1 0 37744 0 1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_68_367
timestamp 1698431365
transform 1 0 42448 0 1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_375
timestamp 1698431365
transform 1 0 43344 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_68_377
timestamp 1698431365
transform 1 0 43568 0 1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_383
timestamp 1698431365
transform 1 0 44240 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_68_387
timestamp 1698431365
transform 1 0 44688 0 1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_395
timestamp 1698431365
transform 1 0 45584 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_68_399
timestamp 1698431365
transform 1 0 46032 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_403
timestamp 1698431365
transform 1 0 46480 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_407
timestamp 1698431365
transform 1 0 46928 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_68_414
timestamp 1698431365
transform 1 0 47712 0 1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_421
timestamp 1698431365
transform 1 0 48496 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_68_425
timestamp 1698431365
transform 1 0 48944 0 1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_68_441
timestamp 1698431365
transform 1 0 50736 0 1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_68_449
timestamp 1698431365
transform 1 0 51632 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_68_453
timestamp 1698431365
transform 1 0 52080 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_68_457
timestamp 1698431365
transform 1 0 52528 0 1 56448
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_68_489
timestamp 1698431365
transform 1 0 56112 0 1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_68_505
timestamp 1698431365
transform 1 0 57904 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_69_2
timestamp 1698431365
transform 1 0 1568 0 -1 58016
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_69_34
timestamp 1698431365
transform 1 0 5152 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_69_38
timestamp 1698431365
transform 1 0 5600 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_69_40
timestamp 1698431365
transform 1 0 5824 0 -1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_69_77
timestamp 1698431365
transform 1 0 9968 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_69_138
timestamp 1698431365
transform 1 0 16800 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_69_142
timestamp 1698431365
transform 1 0 17248 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_69_186
timestamp 1698431365
transform 1 0 22176 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_69_188
timestamp 1698431365
transform 1 0 22400 0 -1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_69_266
timestamp 1698431365
transform 1 0 31136 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_69_270
timestamp 1698431365
transform 1 0 31584 0 -1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_69_290
timestamp 1698431365
transform 1 0 33824 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_69_294
timestamp 1698431365
transform 1 0 34272 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_69_346
timestamp 1698431365
transform 1 0 40096 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_69_368
timestamp 1698431365
transform 1 0 42560 0 -1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_69_381
timestamp 1698431365
transform 1 0 44016 0 -1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_69_422
timestamp 1698431365
transform 1 0 48608 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_69_426
timestamp 1698431365
transform 1 0 49056 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_69_430
timestamp 1698431365
transform 1 0 49504 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_69_434
timestamp 1698431365
transform 1 0 49952 0 -1 58016
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_69_466
timestamp 1698431365
transform 1 0 53536 0 -1 58016
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_69_482
timestamp 1698431365
transform 1 0 55328 0 -1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_69_492
timestamp 1698431365
transform 1 0 56448 0 -1 58016
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_69_508
timestamp 1698431365
transform 1 0 58240 0 -1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_70_2
timestamp 1698431365
transform 1 0 1568 0 1 58016
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_70_34
timestamp 1698431365
transform 1 0 5152 0 1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_70_37
timestamp 1698431365
transform 1 0 5488 0 1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_70_45
timestamp 1698431365
transform 1 0 6384 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_99
timestamp 1698431365
transform 1 0 12432 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_103
timestamp 1698431365
transform 1 0 12880 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_70_107
timestamp 1698431365
transform 1 0 13328 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_70_111
timestamp 1698431365
transform 1 0 13776 0 1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_70_118
timestamp 1698431365
transform 1 0 14560 0 1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_137
timestamp 1698431365
transform 1 0 16688 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_70_139
timestamp 1698431365
transform 1 0 16912 0 1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_150
timestamp 1698431365
transform 1 0 18144 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_70_152
timestamp 1698431365
transform 1 0 18368 0 1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_159
timestamp 1698431365
transform 1 0 19152 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_70_161
timestamp 1698431365
transform 1 0 19376 0 1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_177
timestamp 1698431365
transform 1 0 21168 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_231
timestamp 1698431365
transform 1 0 27216 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_70_233
timestamp 1698431365
transform 1 0 27440 0 1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_70_244
timestamp 1698431365
transform 1 0 28672 0 1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_247
timestamp 1698431365
transform 1 0 29008 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_70_249
timestamp 1698431365
transform 1 0 29232 0 1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_260
timestamp 1698431365
transform 1 0 30464 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_70_262
timestamp 1698431365
transform 1 0 30688 0 1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_271
timestamp 1698431365
transform 1 0 31696 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_70_275
timestamp 1698431365
transform 1 0 32144 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_289
timestamp 1698431365
transform 1 0 33712 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_70_291
timestamp 1698431365
transform 1 0 33936 0 1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_70_297
timestamp 1698431365
transform 1 0 34608 0 1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_304
timestamp 1698431365
transform 1 0 35392 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_308
timestamp 1698431365
transform 1 0 35840 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_312
timestamp 1698431365
transform 1 0 36288 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_70_314
timestamp 1698431365
transform 1 0 36512 0 1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_317
timestamp 1698431365
transform 1 0 36848 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_332
timestamp 1698431365
transform 1 0 38528 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_364
timestamp 1698431365
transform 1 0 42112 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_70_366
timestamp 1698431365
transform 1 0 42336 0 1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_373
timestamp 1698431365
transform 1 0 43120 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_70_375
timestamp 1698431365
transform 1 0 43344 0 1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_381
timestamp 1698431365
transform 1 0 44016 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_70_437
timestamp 1698431365
transform 1 0 50288 0 1 58016
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_453
timestamp 1698431365
transform 1 0 52080 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_70_457
timestamp 1698431365
transform 1 0 52528 0 1 58016
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_70_489
timestamp 1698431365
transform 1 0 56112 0 1 58016
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_70_505
timestamp 1698431365
transform 1 0 57904 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_71_2
timestamp 1698431365
transform 1 0 1568 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_71_101
timestamp 1698431365
transform 1 0 12656 0 -1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_109
timestamp 1698431365
transform 1 0 13552 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_142
timestamp 1698431365
transform 1 0 17248 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_71_146
timestamp 1698431365
transform 1 0 17696 0 -1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_71_154
timestamp 1698431365
transform 1 0 18592 0 -1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_185
timestamp 1698431365
transform 1 0 22064 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_189
timestamp 1698431365
transform 1 0 22512 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_71_193
timestamp 1698431365
transform 1 0 22960 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_197
timestamp 1698431365
transform 1 0 23408 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_201
timestamp 1698431365
transform 1 0 23856 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_225
timestamp 1698431365
transform 1 0 26544 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_235
timestamp 1698431365
transform 1 0 27664 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_71_239
timestamp 1698431365
transform 1 0 28112 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_71_243
timestamp 1698431365
transform 1 0 28560 0 -1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_71_279
timestamp 1698431365
transform 1 0 32592 0 -1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_71_336
timestamp 1698431365
transform 1 0 38976 0 -1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_347
timestamp 1698431365
transform 1 0 40208 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_71_349
timestamp 1698431365
transform 1 0 40432 0 -1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_71_365
timestamp 1698431365
transform 1 0 42224 0 -1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_371
timestamp 1698431365
transform 1 0 42896 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_71_398
timestamp 1698431365
transform 1 0 45920 0 -1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_417
timestamp 1698431365
transform 1 0 48048 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_71_419
timestamp 1698431365
transform 1 0 48272 0 -1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_427
timestamp 1698431365
transform 1 0 49168 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_431
timestamp 1698431365
transform 1 0 49616 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_435
timestamp 1698431365
transform 1 0 50064 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_71_439
timestamp 1698431365
transform 1 0 50512 0 -1 59584
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_71_471
timestamp 1698431365
transform 1 0 54096 0 -1 59584
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_487
timestamp 1698431365
transform 1 0 55888 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_71_489
timestamp 1698431365
transform 1 0 56112 0 -1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_71_492
timestamp 1698431365
transform 1 0 56448 0 -1 59584
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_71_508
timestamp 1698431365
transform 1 0 58240 0 -1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_72_2
timestamp 1698431365
transform 1 0 1568 0 1 59584
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_72_34
timestamp 1698431365
transform 1 0 5152 0 1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_72_37
timestamp 1698431365
transform 1 0 5488 0 1 59584
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_72_69
timestamp 1698431365
transform 1 0 9072 0 1 59584
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_72_85
timestamp 1698431365
transform 1 0 10864 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_72_89
timestamp 1698431365
transform 1 0 11312 0 1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_72_99
timestamp 1698431365
transform 1 0 12432 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_72_103
timestamp 1698431365
transform 1 0 12880 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_72_107
timestamp 1698431365
transform 1 0 13328 0 1 59584
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_72_123
timestamp 1698431365
transform 1 0 15120 0 1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_72_137
timestamp 1698431365
transform 1 0 16688 0 1 59584
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_72_153
timestamp 1698431365
transform 1 0 18480 0 1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_72_161
timestamp 1698431365
transform 1 0 19376 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_72_165
timestamp 1698431365
transform 1 0 19824 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_72_177
timestamp 1698431365
transform 1 0 21168 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_72_179
timestamp 1698431365
transform 1 0 21392 0 1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_72_188
timestamp 1698431365
transform 1 0 22400 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_72_192
timestamp 1698431365
transform 1 0 22848 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_72_196
timestamp 1698431365
transform 1 0 23296 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_72_208
timestamp 1698431365
transform 1 0 24640 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_72_212
timestamp 1698431365
transform 1 0 25088 0 1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_72_215
timestamp 1698431365
transform 1 0 25424 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_72_243
timestamp 1698431365
transform 1 0 28560 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_72_247
timestamp 1698431365
transform 1 0 29008 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_72_251
timestamp 1698431365
transform 1 0 29456 0 1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_72_254
timestamp 1698431365
transform 1 0 29792 0 1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_72_262
timestamp 1698431365
transform 1 0 30688 0 1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_72_269
timestamp 1698431365
transform 1 0 31472 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_72_302
timestamp 1698431365
transform 1 0 35168 0 1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_72_313
timestamp 1698431365
transform 1 0 36400 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_72_352
timestamp 1698431365
transform 1 0 40768 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_72_356
timestamp 1698431365
transform 1 0 41216 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_72_360
timestamp 1698431365
transform 1 0 41664 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_72_383
timestamp 1698431365
transform 1 0 44240 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_72_397
timestamp 1698431365
transform 1 0 45808 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_72_401
timestamp 1698431365
transform 1 0 46256 0 1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_72_419
timestamp 1698431365
transform 1 0 48272 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_72_421
timestamp 1698431365
transform 1 0 48496 0 1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_72_430
timestamp 1698431365
transform 1 0 49504 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_72_434
timestamp 1698431365
transform 1 0 49952 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_72_438
timestamp 1698431365
transform 1 0 50400 0 1 59584
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_72_454
timestamp 1698431365
transform 1 0 52192 0 1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_72_457
timestamp 1698431365
transform 1 0 52528 0 1 59584
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_72_489
timestamp 1698431365
transform 1 0 56112 0 1 59584
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_72_505
timestamp 1698431365
transform 1 0 57904 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_73_2
timestamp 1698431365
transform 1 0 1568 0 -1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_73_66
timestamp 1698431365
transform 1 0 8736 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_73_107
timestamp 1698431365
transform 1 0 13328 0 -1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_73_115
timestamp 1698431365
transform 1 0 14224 0 -1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_73_122
timestamp 1698431365
transform 1 0 15008 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_73_126
timestamp 1698431365
transform 1 0 15456 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_73_128
timestamp 1698431365
transform 1 0 15680 0 -1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_73_146
timestamp 1698431365
transform 1 0 17696 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_73_150
timestamp 1698431365
transform 1 0 18144 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_73_154
timestamp 1698431365
transform 1 0 18592 0 -1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_73_159
timestamp 1698431365
transform 1 0 19152 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_73_176
timestamp 1698431365
transform 1 0 21056 0 -1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_73_197
timestamp 1698431365
transform 1 0 23408 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_73_201
timestamp 1698431365
transform 1 0 23856 0 -1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_73_249
timestamp 1698431365
transform 1 0 29232 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_73_263
timestamp 1698431365
transform 1 0 30800 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_73_267
timestamp 1698431365
transform 1 0 31248 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_73_271
timestamp 1698431365
transform 1 0 31696 0 -1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_73_342
timestamp 1698431365
transform 1 0 39648 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_73_346
timestamp 1698431365
transform 1 0 40096 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_73_352
timestamp 1698431365
transform 1 0 40768 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_73_356
timestamp 1698431365
transform 1 0 41216 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_73_362
timestamp 1698431365
transform 1 0 41888 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_73_368
timestamp 1698431365
transform 1 0 42560 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_73_370
timestamp 1698431365
transform 1 0 42784 0 -1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_73_402
timestamp 1698431365
transform 1 0 46368 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_73_404
timestamp 1698431365
transform 1 0 46592 0 -1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_73_435
timestamp 1698431365
transform 1 0 50064 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_73_439
timestamp 1698431365
transform 1 0 50512 0 -1 61152
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_73_471
timestamp 1698431365
transform 1 0 54096 0 -1 61152
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_73_487
timestamp 1698431365
transform 1 0 55888 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_73_489
timestamp 1698431365
transform 1 0 56112 0 -1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_73_492
timestamp 1698431365
transform 1 0 56448 0 -1 61152
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_73_508
timestamp 1698431365
transform 1 0 58240 0 -1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_74_2
timestamp 1698431365
transform 1 0 1568 0 1 61152
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_74_34
timestamp 1698431365
transform 1 0 5152 0 1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_74_37
timestamp 1698431365
transform 1 0 5488 0 1 61152
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_74_69
timestamp 1698431365
transform 1 0 9072 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_74_73
timestamp 1698431365
transform 1 0 9520 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_74_75
timestamp 1698431365
transform 1 0 9744 0 1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_74_98
timestamp 1698431365
transform 1 0 12320 0 1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_74_107
timestamp 1698431365
transform 1 0 13328 0 1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_74_172
timestamp 1698431365
transform 1 0 20608 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_74_174
timestamp 1698431365
transform 1 0 20832 0 1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_74_219
timestamp 1698431365
transform 1 0 25872 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_74_242
timestamp 1698431365
transform 1 0 28448 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_74_244
timestamp 1698431365
transform 1 0 28672 0 1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_74_283
timestamp 1698431365
transform 1 0 33040 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_74_285
timestamp 1698431365
transform 1 0 33264 0 1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_74_305
timestamp 1698431365
transform 1 0 35504 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_74_309
timestamp 1698431365
transform 1 0 35952 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_74_313
timestamp 1698431365
transform 1 0 36400 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_74_317
timestamp 1698431365
transform 1 0 36848 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_74_319
timestamp 1698431365
transform 1 0 37072 0 1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_74_341
timestamp 1698431365
transform 1 0 39536 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_74_343
timestamp 1698431365
transform 1 0 39760 0 1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_74_367
timestamp 1698431365
transform 1 0 42448 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_74_371
timestamp 1698431365
transform 1 0 42896 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_74_375
timestamp 1698431365
transform 1 0 43344 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_74_379
timestamp 1698431365
transform 1 0 43792 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_74_405
timestamp 1698431365
transform 1 0 46704 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_74_444
timestamp 1698431365
transform 1 0 51072 0 1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_74_452
timestamp 1698431365
transform 1 0 51968 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_74_454
timestamp 1698431365
transform 1 0 52192 0 1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_74_457
timestamp 1698431365
transform 1 0 52528 0 1 61152
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_74_489
timestamp 1698431365
transform 1 0 56112 0 1 61152
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_74_505
timestamp 1698431365
transform 1 0 57904 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_75_2
timestamp 1698431365
transform 1 0 1568 0 -1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_75_66
timestamp 1698431365
transform 1 0 8736 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_75_106
timestamp 1698431365
transform 1 0 13216 0 -1 62720
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_75_122
timestamp 1698431365
transform 1 0 15008 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_75_142
timestamp 1698431365
transform 1 0 17248 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_75_146
timestamp 1698431365
transform 1 0 17696 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_75_206
timestamp 1698431365
transform 1 0 24416 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_75_212
timestamp 1698431365
transform 1 0 25088 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_75_216
timestamp 1698431365
transform 1 0 25536 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_75_218
timestamp 1698431365
transform 1 0 25760 0 -1 62720
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_75_221
timestamp 1698431365
transform 1 0 26096 0 -1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_75_229
timestamp 1698431365
transform 1 0 26992 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_75_231
timestamp 1698431365
transform 1 0 27216 0 -1 62720
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_75_234
timestamp 1698431365
transform 1 0 27552 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_75_274
timestamp 1698431365
transform 1 0 32032 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_75_278
timestamp 1698431365
transform 1 0 32480 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_75_296
timestamp 1698431365
transform 1 0 34496 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_75_300
timestamp 1698431365
transform 1 0 34944 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_75_304
timestamp 1698431365
transform 1 0 35392 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_75_308
timestamp 1698431365
transform 1 0 35840 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_75_312
timestamp 1698431365
transform 1 0 36288 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_75_316
timestamp 1698431365
transform 1 0 36736 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_75_322
timestamp 1698431365
transform 1 0 37408 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_75_326
timestamp 1698431365
transform 1 0 37856 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_75_330
timestamp 1698431365
transform 1 0 38304 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_75_334
timestamp 1698431365
transform 1 0 38752 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_75_338
timestamp 1698431365
transform 1 0 39200 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_75_384
timestamp 1698431365
transform 1 0 44352 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_75_388
timestamp 1698431365
transform 1 0 44800 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_75_390
timestamp 1698431365
transform 1 0 45024 0 -1 62720
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_75_472
timestamp 1698431365
transform 1 0 54208 0 -1 62720
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_75_488
timestamp 1698431365
transform 1 0 56000 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_75_492
timestamp 1698431365
transform 1 0 56448 0 -1 62720
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_75_508
timestamp 1698431365
transform 1 0 58240 0 -1 62720
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_76_2
timestamp 1698431365
transform 1 0 1568 0 1 62720
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_76_34
timestamp 1698431365
transform 1 0 5152 0 1 62720
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_76_37
timestamp 1698431365
transform 1 0 5488 0 1 62720
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_76_69
timestamp 1698431365
transform 1 0 9072 0 1 62720
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_76_85
timestamp 1698431365
transform 1 0 10864 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_76_89
timestamp 1698431365
transform 1 0 11312 0 1 62720
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_76_95
timestamp 1698431365
transform 1 0 11984 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_76_103
timestamp 1698431365
transform 1 0 12880 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_76_157
timestamp 1698431365
transform 1 0 18928 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_76_161
timestamp 1698431365
transform 1 0 19376 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_76_171
timestamp 1698431365
transform 1 0 20496 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_76_177
timestamp 1698431365
transform 1 0 21168 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_76_179
timestamp 1698431365
transform 1 0 21392 0 1 62720
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_76_218
timestamp 1698431365
transform 1 0 25760 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_76_222
timestamp 1698431365
transform 1 0 26208 0 1 62720
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_76_238
timestamp 1698431365
transform 1 0 28000 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_76_244
timestamp 1698431365
transform 1 0 28672 0 1 62720
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_76_247
timestamp 1698431365
transform 1 0 29008 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_76_249
timestamp 1698431365
transform 1 0 29232 0 1 62720
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_76_300
timestamp 1698431365
transform 1 0 34944 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_76_312
timestamp 1698431365
transform 1 0 36288 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_76_314
timestamp 1698431365
transform 1 0 36512 0 1 62720
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_76_322
timestamp 1698431365
transform 1 0 37408 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_76_324
timestamp 1698431365
transform 1 0 37632 0 1 62720
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_76_333
timestamp 1698431365
transform 1 0 38640 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_76_337
timestamp 1698431365
transform 1 0 39088 0 1 62720
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_76_375
timestamp 1698431365
transform 1 0 43344 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_76_377
timestamp 1698431365
transform 1 0 43568 0 1 62720
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_76_437
timestamp 1698431365
transform 1 0 50288 0 1 62720
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_76_453
timestamp 1698431365
transform 1 0 52080 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_76_457
timestamp 1698431365
transform 1 0 52528 0 1 62720
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_76_489
timestamp 1698431365
transform 1 0 56112 0 1 62720
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_76_505
timestamp 1698431365
transform 1 0 57904 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_77_2
timestamp 1698431365
transform 1 0 1568 0 -1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_77_66
timestamp 1698431365
transform 1 0 8736 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_77_72
timestamp 1698431365
transform 1 0 9408 0 -1 64288
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_77_115
timestamp 1698431365
transform 1 0 14224 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_77_117
timestamp 1698431365
transform 1 0 14448 0 -1 64288
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_77_138
timestamp 1698431365
transform 1 0 16800 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_77_146
timestamp 1698431365
transform 1 0 17696 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_77_150
timestamp 1698431365
transform 1 0 18144 0 -1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_77_158
timestamp 1698431365
transform 1 0 19040 0 -1 64288
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_77_163
timestamp 1698431365
transform 1 0 19600 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_77_172
timestamp 1698431365
transform 1 0 20608 0 -1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_77_180
timestamp 1698431365
transform 1 0 21504 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_77_184
timestamp 1698431365
transform 1 0 21952 0 -1 64288
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_77_208
timestamp 1698431365
transform 1 0 24640 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_77_212
timestamp 1698431365
transform 1 0 25088 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_77_214
timestamp 1698431365
transform 1 0 25312 0 -1 64288
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_77_228
timestamp 1698431365
transform 1 0 26880 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_77_232
timestamp 1698431365
transform 1 0 27328 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_77_234
timestamp 1698431365
transform 1 0 27552 0 -1 64288
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_77_248
timestamp 1698431365
transform 1 0 29120 0 -1 64288
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_77_267
timestamp 1698431365
transform 1 0 31248 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_77_348
timestamp 1698431365
transform 1 0 40320 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_77_370
timestamp 1698431365
transform 1 0 42784 0 -1 64288
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_77_400
timestamp 1698431365
transform 1 0 46144 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_77_404
timestamp 1698431365
transform 1 0 46592 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_77_406
timestamp 1698431365
transform 1 0 46816 0 -1 64288
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_77_422
timestamp 1698431365
transform 1 0 48608 0 -1 64288
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_77_427
timestamp 1698431365
transform 1 0 49168 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_77_431
timestamp 1698431365
transform 1 0 49616 0 -1 64288
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_77_463
timestamp 1698431365
transform 1 0 53200 0 -1 64288
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_77_479
timestamp 1698431365
transform 1 0 54992 0 -1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_77_487
timestamp 1698431365
transform 1 0 55888 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_77_489
timestamp 1698431365
transform 1 0 56112 0 -1 64288
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_77_492
timestamp 1698431365
transform 1 0 56448 0 -1 64288
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_77_508
timestamp 1698431365
transform 1 0 58240 0 -1 64288
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_78_2
timestamp 1698431365
transform 1 0 1568 0 1 64288
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_78_34
timestamp 1698431365
transform 1 0 5152 0 1 64288
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_78_37
timestamp 1698431365
transform 1 0 5488 0 1 64288
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_78_69
timestamp 1698431365
transform 1 0 9072 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_78_73
timestamp 1698431365
transform 1 0 9520 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_78_75
timestamp 1698431365
transform 1 0 9744 0 1 64288
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_78_107
timestamp 1698431365
transform 1 0 13328 0 1 64288
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_78_182
timestamp 1698431365
transform 1 0 21728 0 1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_78_255
timestamp 1698431365
transform 1 0 29904 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_78_259
timestamp 1698431365
transform 1 0 30352 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_78_263
timestamp 1698431365
transform 1 0 30800 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_78_302
timestamp 1698431365
transform 1 0 35168 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_78_304
timestamp 1698431365
transform 1 0 35392 0 1 64288
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_78_317
timestamp 1698431365
transform 1 0 36848 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_78_370
timestamp 1698431365
transform 1 0 42784 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_78_374
timestamp 1698431365
transform 1 0 43232 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_78_376
timestamp 1698431365
transform 1 0 43456 0 1 64288
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_78_383
timestamp 1698431365
transform 1 0 44240 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_78_395
timestamp 1698431365
transform 1 0 45584 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_78_399
timestamp 1698431365
transform 1 0 46032 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_78_403
timestamp 1698431365
transform 1 0 46480 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_78_407
timestamp 1698431365
transform 1 0 46928 0 1 64288
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_78_439
timestamp 1698431365
transform 1 0 50512 0 1 64288
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_78_457
timestamp 1698431365
transform 1 0 52528 0 1 64288
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_78_489
timestamp 1698431365
transform 1 0 56112 0 1 64288
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_78_505
timestamp 1698431365
transform 1 0 57904 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_79_2
timestamp 1698431365
transform 1 0 1568 0 -1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_79_66
timestamp 1698431365
transform 1 0 8736 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_79_72
timestamp 1698431365
transform 1 0 9408 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_79_137
timestamp 1698431365
transform 1 0 16688 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_79_139
timestamp 1698431365
transform 1 0 16912 0 -1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_79_155
timestamp 1698431365
transform 1 0 18704 0 -1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_79_163
timestamp 1698431365
transform 1 0 19600 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_79_200
timestamp 1698431365
transform 1 0 23744 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_79_202
timestamp 1698431365
transform 1 0 23968 0 -1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_79_209
timestamp 1698431365
transform 1 0 24752 0 -1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_79_263
timestamp 1698431365
transform 1 0 30800 0 -1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_79_271
timestamp 1698431365
transform 1 0 31696 0 -1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_79_298
timestamp 1698431365
transform 1 0 34720 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_79_358
timestamp 1698431365
transform 1 0 41440 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_79_362
timestamp 1698431365
transform 1 0 41888 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_79_366
timestamp 1698431365
transform 1 0 42336 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_79_370
timestamp 1698431365
transform 1 0 42784 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_79_374
timestamp 1698431365
transform 1 0 43232 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_79_376
timestamp 1698431365
transform 1 0 43456 0 -1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_79_387
timestamp 1698431365
transform 1 0 44688 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_79_395
timestamp 1698431365
transform 1 0 45584 0 -1 65856
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_79_417
timestamp 1698431365
transform 1 0 48048 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_79_419
timestamp 1698431365
transform 1 0 48272 0 -1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_79_422
timestamp 1698431365
transform 1 0 48608 0 -1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_79_486
timestamp 1698431365
transform 1 0 55776 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_79_492
timestamp 1698431365
transform 1 0 56448 0 -1 65856
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_79_508
timestamp 1698431365
transform 1 0 58240 0 -1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_80_2
timestamp 1698431365
transform 1 0 1568 0 1 65856
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_80_34
timestamp 1698431365
transform 1 0 5152 0 1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_80_37
timestamp 1698431365
transform 1 0 5488 0 1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_80_101
timestamp 1698431365
transform 1 0 12656 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_80_107
timestamp 1698431365
transform 1 0 13328 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_80_145
timestamp 1698431365
transform 1 0 17584 0 1 65856
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_80_161
timestamp 1698431365
transform 1 0 19376 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_80_163
timestamp 1698431365
transform 1 0 19600 0 1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_80_170
timestamp 1698431365
transform 1 0 20384 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_80_174
timestamp 1698431365
transform 1 0 20832 0 1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_80_188
timestamp 1698431365
transform 1 0 22400 0 1 65856
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_80_204
timestamp 1698431365
transform 1 0 24192 0 1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_80_224
timestamp 1698431365
transform 1 0 26432 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_80_226
timestamp 1698431365
transform 1 0 26656 0 1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_80_243
timestamp 1698431365
transform 1 0 28560 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_80_247
timestamp 1698431365
transform 1 0 29008 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_80_251
timestamp 1698431365
transform 1 0 29456 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_80_268
timestamp 1698431365
transform 1 0 31360 0 1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_80_276
timestamp 1698431365
transform 1 0 32256 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_80_282
timestamp 1698431365
transform 1 0 32928 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_80_284
timestamp 1698431365
transform 1 0 33152 0 1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_80_294
timestamp 1698431365
transform 1 0 34272 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_80_298
timestamp 1698431365
transform 1 0 34720 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_80_300
timestamp 1698431365
transform 1 0 34944 0 1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_80_325
timestamp 1698431365
transform 1 0 37744 0 1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_80_346
timestamp 1698431365
transform 1 0 40096 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_80_350
timestamp 1698431365
transform 1 0 40544 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_80_352
timestamp 1698431365
transform 1 0 40768 0 1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_80_383
timestamp 1698431365
transform 1 0 44240 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_80_387
timestamp 1698431365
transform 1 0 44688 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_80_389
timestamp 1698431365
transform 1 0 44912 0 1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_80_419
timestamp 1698431365
transform 1 0 48272 0 1 65856
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_80_451
timestamp 1698431365
transform 1 0 51856 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_80_457
timestamp 1698431365
transform 1 0 52528 0 1 65856
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_80_489
timestamp 1698431365
transform 1 0 56112 0 1 65856
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_80_505
timestamp 1698431365
transform 1 0 57904 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_81_2
timestamp 1698431365
transform 1 0 1568 0 -1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_81_66
timestamp 1698431365
transform 1 0 8736 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_81_72
timestamp 1698431365
transform 1 0 9408 0 -1 67424
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_81_104
timestamp 1698431365
transform 1 0 12992 0 -1 67424
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_81_120
timestamp 1698431365
transform 1 0 14784 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_81_122
timestamp 1698431365
transform 1 0 15008 0 -1 67424
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_81_127
timestamp 1698431365
transform 1 0 15568 0 -1 67424
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_81_135
timestamp 1698431365
transform 1 0 16464 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_81_139
timestamp 1698431365
transform 1 0 16912 0 -1 67424
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_81_142
timestamp 1698431365
transform 1 0 17248 0 -1 67424
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_81_158
timestamp 1698431365
transform 1 0 19040 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_81_162
timestamp 1698431365
transform 1 0 19488 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_81_164
timestamp 1698431365
transform 1 0 19712 0 -1 67424
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_81_173
timestamp 1698431365
transform 1 0 20720 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_81_175
timestamp 1698431365
transform 1 0 20944 0 -1 67424
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_81_196
timestamp 1698431365
transform 1 0 23296 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_81_200
timestamp 1698431365
transform 1 0 23744 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_81_207
timestamp 1698431365
transform 1 0 24528 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_81_209
timestamp 1698431365
transform 1 0 24752 0 -1 67424
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_81_212
timestamp 1698431365
transform 1 0 25088 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_81_218
timestamp 1698431365
transform 1 0 25760 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_81_222
timestamp 1698431365
transform 1 0 26208 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_81_226
timestamp 1698431365
transform 1 0 26656 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_81_230
timestamp 1698431365
transform 1 0 27104 0 -1 67424
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_81_238
timestamp 1698431365
transform 1 0 28000 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_81_242
timestamp 1698431365
transform 1 0 28448 0 -1 67424
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_81_245
timestamp 1698431365
transform 1 0 28784 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_81_272
timestamp 1698431365
transform 1 0 31808 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_81_276
timestamp 1698431365
transform 1 0 32256 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_81_282
timestamp 1698431365
transform 1 0 32928 0 -1 67424
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_81_290
timestamp 1698431365
transform 1 0 33824 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_81_296
timestamp 1698431365
transform 1 0 34496 0 -1 67424
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_81_312
timestamp 1698431365
transform 1 0 36288 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_81_314
timestamp 1698431365
transform 1 0 36512 0 -1 67424
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_81_317
timestamp 1698431365
transform 1 0 36848 0 -1 67424
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_81_333
timestamp 1698431365
transform 1 0 38640 0 -1 67424
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_81_341
timestamp 1698431365
transform 1 0 39536 0 -1 67424
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_81_344
timestamp 1698431365
transform 1 0 39872 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_81_348
timestamp 1698431365
transform 1 0 40320 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_81_352
timestamp 1698431365
transform 1 0 40768 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_81_397
timestamp 1698431365
transform 1 0 45808 0 -1 67424
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_81_413
timestamp 1698431365
transform 1 0 47600 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_81_417
timestamp 1698431365
transform 1 0 48048 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_81_419
timestamp 1698431365
transform 1 0 48272 0 -1 67424
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_81_422
timestamp 1698431365
transform 1 0 48608 0 -1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_81_486
timestamp 1698431365
transform 1 0 55776 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_81_492
timestamp 1698431365
transform 1 0 56448 0 -1 67424
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_81_508
timestamp 1698431365
transform 1 0 58240 0 -1 67424
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_82_2
timestamp 1698431365
transform 1 0 1568 0 1 67424
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_82_34
timestamp 1698431365
transform 1 0 5152 0 1 67424
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_82_37
timestamp 1698431365
transform 1 0 5488 0 1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_82_101
timestamp 1698431365
transform 1 0 12656 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_82_107
timestamp 1698431365
transform 1 0 13328 0 1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_82_171
timestamp 1698431365
transform 1 0 20496 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_82_181
timestamp 1698431365
transform 1 0 21616 0 1 67424
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_82_202
timestamp 1698431365
transform 1 0 23968 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_82_204
timestamp 1698431365
transform 1 0 24192 0 1 67424
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_82_225
timestamp 1698431365
transform 1 0 26544 0 1 67424
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_82_233
timestamp 1698431365
transform 1 0 27440 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_82_280
timestamp 1698431365
transform 1 0 32704 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_82_288
timestamp 1698431365
transform 1 0 33600 0 1 67424
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_82_304
timestamp 1698431365
transform 1 0 35392 0 1 67424
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_82_313
timestamp 1698431365
transform 1 0 36400 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_82_317
timestamp 1698431365
transform 1 0 36848 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_82_319
timestamp 1698431365
transform 1 0 37072 0 1 67424
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_82_325
timestamp 1698431365
transform 1 0 37744 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_82_327
timestamp 1698431365
transform 1 0 37968 0 1 67424
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_82_336
timestamp 1698431365
transform 1 0 38976 0 1 67424
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_82_344
timestamp 1698431365
transform 1 0 39872 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_82_346
timestamp 1698431365
transform 1 0 40096 0 1 67424
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_82_416
timestamp 1698431365
transform 1 0 47936 0 1 67424
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_82_448
timestamp 1698431365
transform 1 0 51520 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_82_452
timestamp 1698431365
transform 1 0 51968 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_82_454
timestamp 1698431365
transform 1 0 52192 0 1 67424
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_82_457
timestamp 1698431365
transform 1 0 52528 0 1 67424
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_82_489
timestamp 1698431365
transform 1 0 56112 0 1 67424
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_82_505
timestamp 1698431365
transform 1 0 57904 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_83_2
timestamp 1698431365
transform 1 0 1568 0 -1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_83_66
timestamp 1698431365
transform 1 0 8736 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_83_72
timestamp 1698431365
transform 1 0 9408 0 -1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_83_136
timestamp 1698431365
transform 1 0 16576 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_83_142
timestamp 1698431365
transform 1 0 17248 0 -1 68992
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_83_158
timestamp 1698431365
transform 1 0 19040 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_83_162
timestamp 1698431365
transform 1 0 19488 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_83_193
timestamp 1698431365
transform 1 0 22960 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_83_262
timestamp 1698431365
transform 1 0 30688 0 -1 68992
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_83_278
timestamp 1698431365
transform 1 0 32480 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_83_289
timestamp 1698431365
transform 1 0 33712 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_83_293
timestamp 1698431365
transform 1 0 34160 0 -1 68992
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_83_300
timestamp 1698431365
transform 1 0 34944 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_83_302
timestamp 1698431365
transform 1 0 35168 0 -1 68992
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_83_341
timestamp 1698431365
transform 1 0 39536 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_83_360
timestamp 1698431365
transform 1 0 41664 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_83_412
timestamp 1698431365
transform 1 0 47488 0 -1 68992
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_83_422
timestamp 1698431365
transform 1 0 48608 0 -1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_83_486
timestamp 1698431365
transform 1 0 55776 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_83_492
timestamp 1698431365
transform 1 0 56448 0 -1 68992
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_83_508
timestamp 1698431365
transform 1 0 58240 0 -1 68992
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_84_2
timestamp 1698431365
transform 1 0 1568 0 1 68992
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_84_34
timestamp 1698431365
transform 1 0 5152 0 1 68992
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_84_37
timestamp 1698431365
transform 1 0 5488 0 1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_84_101
timestamp 1698431365
transform 1 0 12656 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_84_107
timestamp 1698431365
transform 1 0 13328 0 1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_84_171
timestamp 1698431365
transform 1 0 20496 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_84_177
timestamp 1698431365
transform 1 0 21168 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_84_181
timestamp 1698431365
transform 1 0 21616 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_84_183
timestamp 1698431365
transform 1 0 21840 0 1 68992
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_84_242
timestamp 1698431365
transform 1 0 28448 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_84_244
timestamp 1698431365
transform 1 0 28672 0 1 68992
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_84_274
timestamp 1698431365
transform 1 0 32032 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_84_278
timestamp 1698431365
transform 1 0 32480 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_84_288
timestamp 1698431365
transform 1 0 33600 0 1 68992
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_84_309
timestamp 1698431365
transform 1 0 35952 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_84_317
timestamp 1698431365
transform 1 0 36848 0 1 68992
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_84_334
timestamp 1698431365
transform 1 0 38752 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_84_336
timestamp 1698431365
transform 1 0 38976 0 1 68992
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_84_380
timestamp 1698431365
transform 1 0 43904 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_84_384
timestamp 1698431365
transform 1 0 44352 0 1 68992
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_84_387
timestamp 1698431365
transform 1 0 44688 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_84_395
timestamp 1698431365
transform 1 0 45584 0 1 68992
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_84_427
timestamp 1698431365
transform 1 0 49168 0 1 68992
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_84_443
timestamp 1698431365
transform 1 0 50960 0 1 68992
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_84_451
timestamp 1698431365
transform 1 0 51856 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_84_457
timestamp 1698431365
transform 1 0 52528 0 1 68992
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_84_489
timestamp 1698431365
transform 1 0 56112 0 1 68992
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_84_505
timestamp 1698431365
transform 1 0 57904 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_85_2
timestamp 1698431365
transform 1 0 1568 0 -1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_85_66
timestamp 1698431365
transform 1 0 8736 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_85_72
timestamp 1698431365
transform 1 0 9408 0 -1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_85_136
timestamp 1698431365
transform 1 0 16576 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_85_142
timestamp 1698431365
transform 1 0 17248 0 -1 70560
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_85_174
timestamp 1698431365
transform 1 0 20832 0 -1 70560
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_85_190
timestamp 1698431365
transform 1 0 22624 0 -1 70560
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_85_198
timestamp 1698431365
transform 1 0 23520 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_85_204
timestamp 1698431365
transform 1 0 24192 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_85_208
timestamp 1698431365
transform 1 0 24640 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_85_212
timestamp 1698431365
transform 1 0 25088 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_85_216
timestamp 1698431365
transform 1 0 25536 0 -1 70560
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_85_221
timestamp 1698431365
transform 1 0 26096 0 -1 70560
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_85_229
timestamp 1698431365
transform 1 0 26992 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_85_233
timestamp 1698431365
transform 1 0 27440 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_85_268
timestamp 1698431365
transform 1 0 31360 0 -1 70560
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_85_282
timestamp 1698431365
transform 1 0 32928 0 -1 70560
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_85_341
timestamp 1698431365
transform 1 0 39536 0 -1 70560
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_85_381
timestamp 1698431365
transform 1 0 44016 0 -1 70560
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_85_413
timestamp 1698431365
transform 1 0 47600 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_85_417
timestamp 1698431365
transform 1 0 48048 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_85_419
timestamp 1698431365
transform 1 0 48272 0 -1 70560
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_85_422
timestamp 1698431365
transform 1 0 48608 0 -1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_85_486
timestamp 1698431365
transform 1 0 55776 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_85_492
timestamp 1698431365
transform 1 0 56448 0 -1 70560
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_85_508
timestamp 1698431365
transform 1 0 58240 0 -1 70560
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_86_2
timestamp 1698431365
transform 1 0 1568 0 1 70560
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_86_34
timestamp 1698431365
transform 1 0 5152 0 1 70560
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_86_37
timestamp 1698431365
transform 1 0 5488 0 1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_86_101
timestamp 1698431365
transform 1 0 12656 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_86_107
timestamp 1698431365
transform 1 0 13328 0 1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_86_171
timestamp 1698431365
transform 1 0 20496 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_86_177
timestamp 1698431365
transform 1 0 21168 0 1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_86_241
timestamp 1698431365
transform 1 0 28336 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_86_247
timestamp 1698431365
transform 1 0 29008 0 1 70560
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_86_263
timestamp 1698431365
transform 1 0 30800 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_86_267
timestamp 1698431365
transform 1 0 31248 0 1 70560
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_86_301
timestamp 1698431365
transform 1 0 35056 0 1 70560
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_86_309
timestamp 1698431365
transform 1 0 35952 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_86_313
timestamp 1698431365
transform 1 0 36400 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_86_367
timestamp 1698431365
transform 1 0 42448 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_86_371
timestamp 1698431365
transform 1 0 42896 0 1 70560
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_86_379
timestamp 1698431365
transform 1 0 43792 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_86_383
timestamp 1698431365
transform 1 0 44240 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_86_387
timestamp 1698431365
transform 1 0 44688 0 1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_86_451
timestamp 1698431365
transform 1 0 51856 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_86_457
timestamp 1698431365
transform 1 0 52528 0 1 70560
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_86_489
timestamp 1698431365
transform 1 0 56112 0 1 70560
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_86_505
timestamp 1698431365
transform 1 0 57904 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_87_2
timestamp 1698431365
transform 1 0 1568 0 -1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_87_66
timestamp 1698431365
transform 1 0 8736 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_87_72
timestamp 1698431365
transform 1 0 9408 0 -1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_87_136
timestamp 1698431365
transform 1 0 16576 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_87_142
timestamp 1698431365
transform 1 0 17248 0 -1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_87_206
timestamp 1698431365
transform 1 0 24416 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_87_212
timestamp 1698431365
transform 1 0 25088 0 -1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_87_276
timestamp 1698431365
transform 1 0 32256 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_87_282
timestamp 1698431365
transform 1 0 32928 0 -1 72128
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_87_314
timestamp 1698431365
transform 1 0 36512 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_87_316
timestamp 1698431365
transform 1 0 36736 0 -1 72128
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_87_356
timestamp 1698431365
transform 1 0 41216 0 -1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_87_422
timestamp 1698431365
transform 1 0 48608 0 -1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_87_486
timestamp 1698431365
transform 1 0 55776 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_87_492
timestamp 1698431365
transform 1 0 56448 0 -1 72128
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_87_508
timestamp 1698431365
transform 1 0 58240 0 -1 72128
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_88_2
timestamp 1698431365
transform 1 0 1568 0 1 72128
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_88_34
timestamp 1698431365
transform 1 0 5152 0 1 72128
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_88_37
timestamp 1698431365
transform 1 0 5488 0 1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_88_101
timestamp 1698431365
transform 1 0 12656 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_88_107
timestamp 1698431365
transform 1 0 13328 0 1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_88_171
timestamp 1698431365
transform 1 0 20496 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_88_177
timestamp 1698431365
transform 1 0 21168 0 1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_88_241
timestamp 1698431365
transform 1 0 28336 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_88_247
timestamp 1698431365
transform 1 0 29008 0 1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_88_311
timestamp 1698431365
transform 1 0 36176 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_88_317
timestamp 1698431365
transform 1 0 36848 0 1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_88_381
timestamp 1698431365
transform 1 0 44016 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_88_387
timestamp 1698431365
transform 1 0 44688 0 1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_88_451
timestamp 1698431365
transform 1 0 51856 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_88_457
timestamp 1698431365
transform 1 0 52528 0 1 72128
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_88_489
timestamp 1698431365
transform 1 0 56112 0 1 72128
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_88_505
timestamp 1698431365
transform 1 0 57904 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_89_2
timestamp 1698431365
transform 1 0 1568 0 -1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_89_66
timestamp 1698431365
transform 1 0 8736 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_89_72
timestamp 1698431365
transform 1 0 9408 0 -1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_89_136
timestamp 1698431365
transform 1 0 16576 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_89_142
timestamp 1698431365
transform 1 0 17248 0 -1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_89_206
timestamp 1698431365
transform 1 0 24416 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_89_212
timestamp 1698431365
transform 1 0 25088 0 -1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_89_276
timestamp 1698431365
transform 1 0 32256 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_89_282
timestamp 1698431365
transform 1 0 32928 0 -1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_89_346
timestamp 1698431365
transform 1 0 40096 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_89_352
timestamp 1698431365
transform 1 0 40768 0 -1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_89_416
timestamp 1698431365
transform 1 0 47936 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_89_422
timestamp 1698431365
transform 1 0 48608 0 -1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_89_486
timestamp 1698431365
transform 1 0 55776 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_89_492
timestamp 1698431365
transform 1 0 56448 0 -1 73696
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_89_508
timestamp 1698431365
transform 1 0 58240 0 -1 73696
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_90_2
timestamp 1698431365
transform 1 0 1568 0 1 73696
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_90_34
timestamp 1698431365
transform 1 0 5152 0 1 73696
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_90_37
timestamp 1698431365
transform 1 0 5488 0 1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_90_101
timestamp 1698431365
transform 1 0 12656 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_90_107
timestamp 1698431365
transform 1 0 13328 0 1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_90_171
timestamp 1698431365
transform 1 0 20496 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_90_177
timestamp 1698431365
transform 1 0 21168 0 1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_90_241
timestamp 1698431365
transform 1 0 28336 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_90_247
timestamp 1698431365
transform 1 0 29008 0 1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_90_311
timestamp 1698431365
transform 1 0 36176 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_90_317
timestamp 1698431365
transform 1 0 36848 0 1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_90_381
timestamp 1698431365
transform 1 0 44016 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_90_387
timestamp 1698431365
transform 1 0 44688 0 1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_90_451
timestamp 1698431365
transform 1 0 51856 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_90_457
timestamp 1698431365
transform 1 0 52528 0 1 73696
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_90_489
timestamp 1698431365
transform 1 0 56112 0 1 73696
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_90_505
timestamp 1698431365
transform 1 0 57904 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_91_2
timestamp 1698431365
transform 1 0 1568 0 -1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_91_66
timestamp 1698431365
transform 1 0 8736 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_91_72
timestamp 1698431365
transform 1 0 9408 0 -1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_91_136
timestamp 1698431365
transform 1 0 16576 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_91_142
timestamp 1698431365
transform 1 0 17248 0 -1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_91_206
timestamp 1698431365
transform 1 0 24416 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_91_212
timestamp 1698431365
transform 1 0 25088 0 -1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_91_276
timestamp 1698431365
transform 1 0 32256 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_91_282
timestamp 1698431365
transform 1 0 32928 0 -1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_91_346
timestamp 1698431365
transform 1 0 40096 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_91_352
timestamp 1698431365
transform 1 0 40768 0 -1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_91_416
timestamp 1698431365
transform 1 0 47936 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_91_422
timestamp 1698431365
transform 1 0 48608 0 -1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_91_486
timestamp 1698431365
transform 1 0 55776 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_91_492
timestamp 1698431365
transform 1 0 56448 0 -1 75264
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_91_508
timestamp 1698431365
transform 1 0 58240 0 -1 75264
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_92_2
timestamp 1698431365
transform 1 0 1568 0 1 75264
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_92_34
timestamp 1698431365
transform 1 0 5152 0 1 75264
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_92_37
timestamp 1698431365
transform 1 0 5488 0 1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_92_101
timestamp 1698431365
transform 1 0 12656 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_92_107
timestamp 1698431365
transform 1 0 13328 0 1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_92_171
timestamp 1698431365
transform 1 0 20496 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_92_177
timestamp 1698431365
transform 1 0 21168 0 1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_92_241
timestamp 1698431365
transform 1 0 28336 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_92_247
timestamp 1698431365
transform 1 0 29008 0 1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_92_311
timestamp 1698431365
transform 1 0 36176 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_92_317
timestamp 1698431365
transform 1 0 36848 0 1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_92_381
timestamp 1698431365
transform 1 0 44016 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_92_387
timestamp 1698431365
transform 1 0 44688 0 1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_92_451
timestamp 1698431365
transform 1 0 51856 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_92_457
timestamp 1698431365
transform 1 0 52528 0 1 75264
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_92_489
timestamp 1698431365
transform 1 0 56112 0 1 75264
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_92_505
timestamp 1698431365
transform 1 0 57904 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_93_2
timestamp 1698431365
transform 1 0 1568 0 -1 76832
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_93_36
timestamp 1698431365
transform 1 0 5376 0 -1 76832
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_93_70
timestamp 1698431365
transform 1 0 9184 0 -1 76832
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_93_104
timestamp 1698431365
transform 1 0 12992 0 -1 76832
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_93_138
timestamp 1698431365
transform 1 0 16800 0 -1 76832
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_93_172
timestamp 1698431365
transform 1 0 20608 0 -1 76832
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_93_206
timestamp 1698431365
transform 1 0 24416 0 -1 76832
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_93_240
timestamp 1698431365
transform 1 0 28224 0 -1 76832
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_93_274
timestamp 1698431365
transform 1 0 32032 0 -1 76832
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_93_308
timestamp 1698431365
transform 1 0 35840 0 -1 76832
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_93_342
timestamp 1698431365
transform 1 0 39648 0 -1 76832
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_93_376
timestamp 1698431365
transform 1 0 43456 0 -1 76832
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_93_410
timestamp 1698431365
transform 1 0 47264 0 -1 76832
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_93_444
timestamp 1698431365
transform 1 0 51072 0 -1 76832
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_93_478
timestamp 1698431365
transform 1 0 54880 0 -1 76832
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_93_494
timestamp 1698431365
transform 1 0 56672 0 -1 76832
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_93_502
timestamp 1698431365
transform 1 0 57568 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_93_506
timestamp 1698431365
transform 1 0 58016 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_93_508
timestamp 1698431365
transform 1 0 58240 0 -1 76832
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input1
timestamp 1698431365
transform 1 0 1568 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input2
timestamp 1698431365
transform 1 0 1568 0 -1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input3
timestamp 1698431365
transform 1 0 1568 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input4
timestamp 1698431365
transform 1 0 2240 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input5
timestamp 1698431365
transform 1 0 1568 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input6
timestamp 1698431365
transform 1 0 1568 0 1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input7
timestamp 1698431365
transform 1 0 2240 0 1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input8
timestamp 1698431365
transform 1 0 1568 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input9
timestamp 1698431365
transform 1 0 1568 0 1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input10
timestamp 1698431365
transform 1 0 1568 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input11
timestamp 1698431365
transform 1 0 1568 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input12
timestamp 1698431365
transform 1 0 1568 0 1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input13
timestamp 1698431365
transform 1 0 1568 0 -1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input14
timestamp 1698431365
transform 1 0 1568 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input15
timestamp 1698431365
transform 1 0 1568 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input16
timestamp 1698431365
transform 1 0 2240 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input17
timestamp 1698431365
transform 1 0 1568 0 -1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input18
timestamp 1698431365
transform 1 0 1568 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input19
timestamp 1698431365
transform 1 0 24416 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input20
timestamp 1698431365
transform 1 0 12992 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input21
timestamp 1698431365
transform 1 0 1568 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input22
timestamp 1698431365
transform 1 0 2240 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input23
timestamp 1698431365
transform 1 0 1568 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input24
timestamp 1698431365
transform 1 0 1568 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input25
timestamp 1698431365
transform 1 0 1568 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input26
timestamp 1698431365
transform 1 0 1568 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input27
timestamp 1698431365
transform 1 0 1568 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input28
timestamp 1698431365
transform 1 0 1568 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input29
timestamp 1698431365
transform 1 0 1568 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input30
timestamp 1698431365
transform -1 0 20384 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input31
timestamp 1698431365
transform 1 0 1568 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input32
timestamp 1698431365
transform 1 0 2240 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input33
timestamp 1698431365
transform 1 0 1568 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input34
timestamp 1698431365
transform 1 0 1568 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input35
timestamp 1698431365
transform 1 0 2240 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input36
timestamp 1698431365
transform 1 0 1568 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input37
timestamp 1698431365
transform 1 0 1568 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input38
timestamp 1698431365
transform 1 0 1568 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input39
timestamp 1698431365
transform 1 0 1568 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input40
timestamp 1698431365
transform 1 0 1568 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input41
timestamp 1698431365
transform -1 0 19712 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input42
timestamp 1698431365
transform 1 0 2240 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input43
timestamp 1698431365
transform 1 0 1568 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input44
timestamp 1698431365
transform 1 0 18368 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input45
timestamp 1698431365
transform 1 0 17696 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input46
timestamp 1698431365
transform -1 0 17584 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input47
timestamp 1698431365
transform -1 0 16576 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input48
timestamp 1698431365
transform 1 0 1568 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input49
timestamp 1698431365
transform 1 0 2240 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input50
timestamp 1698431365
transform 1 0 1568 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input51
timestamp 1698431365
transform 1 0 1568 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input52
timestamp 1698431365
transform -1 0 31808 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input53
timestamp 1698431365
transform 1 0 33040 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input54
timestamp 1698431365
transform 1 0 34384 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input55
timestamp 1698431365
transform 1 0 36512 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input56
timestamp 1698431365
transform 1 0 38528 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input57
timestamp 1698431365
transform 1 0 39760 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input58
timestamp 1698431365
transform 1 0 41104 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input59
timestamp 1698431365
transform 1 0 42448 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input60
timestamp 1698431365
transform -1 0 44128 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input61
timestamp 1698431365
transform 1 0 44128 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input62
timestamp 1698431365
transform 1 0 1568 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input63
timestamp 1698431365
transform -1 0 58352 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input64
timestamp 1698431365
transform -1 0 58352 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input65
timestamp 1698431365
transform -1 0 58352 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input66
timestamp 1698431365
transform -1 0 58352 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input67
timestamp 1698431365
transform 1 0 40432 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input68
timestamp 1698431365
transform -1 0 38528 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input69
timestamp 1698431365
transform 1 0 37184 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input70
timestamp 1698431365
transform 1 0 35840 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input71
timestamp 1698431365
transform 1 0 33712 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input72
timestamp 1698431365
transform 1 0 30352 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input73
timestamp 1698431365
transform 1 0 1568 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input74
timestamp 1698431365
transform 1 0 29008 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input75
timestamp 1698431365
transform 1 0 1568 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input76
timestamp 1698431365
transform 1 0 1568 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input77
timestamp 1698431365
transform 1 0 20944 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input78
timestamp 1698431365
transform -1 0 23520 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input79
timestamp 1698431365
transform -1 0 24192 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input80
timestamp 1698431365
transform -1 0 26320 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input81
timestamp 1698431365
transform 1 0 27328 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input82
timestamp 1698431365
transform -1 0 30352 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input83
timestamp 1698431365
transform 1 0 1568 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output84 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 4480 0 1 48608
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output85
timestamp 1698431365
transform 1 0 53312 0 -1 47040
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output86
timestamp 1698431365
transform 1 0 53312 0 1 29792
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output87
timestamp 1698431365
transform 1 0 55440 0 1 28224
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output88
timestamp 1698431365
transform 1 0 53312 0 -1 32928
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output89
timestamp 1698431365
transform 1 0 55440 0 1 36064
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output90
timestamp 1698431365
transform 1 0 55440 0 1 34496
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output91
timestamp 1698431365
transform 1 0 52528 0 1 31360
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output92
timestamp 1698431365
transform 1 0 55440 0 1 31360
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output93
timestamp 1698431365
transform 1 0 53312 0 -1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output94
timestamp 1698431365
transform 1 0 53312 0 -1 34496
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output95
timestamp 1698431365
transform -1 0 4480 0 -1 48608
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output96
timestamp 1698431365
transform 1 0 52528 0 1 45472
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output97
timestamp 1698431365
transform 1 0 55440 0 1 45472
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output98
timestamp 1698431365
transform 1 0 55440 0 1 43904
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output99
timestamp 1698431365
transform 1 0 55440 0 1 47040
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output100
timestamp 1698431365
transform 1 0 53312 0 -1 40768
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output101
timestamp 1698431365
transform 1 0 55440 0 1 42336
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output102
timestamp 1698431365
transform 1 0 55440 0 1 39200
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output103
timestamp 1698431365
transform 1 0 52528 0 1 40768
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output104
timestamp 1698431365
transform 1 0 53312 0 -1 39200
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output105
timestamp 1698431365
transform 1 0 55440 0 1 40768
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output106
timestamp 1698431365
transform -1 0 4480 0 1 47040
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output107
timestamp 1698431365
transform 1 0 53312 0 -1 42336
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output108
timestamp 1698431365
transform -1 0 4480 0 1 36064
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output109
timestamp 1698431365
transform -1 0 4480 0 -1 43904
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output110
timestamp 1698431365
transform -1 0 4480 0 1 31360
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output111
timestamp 1698431365
transform -1 0 4480 0 -1 34496
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output112
timestamp 1698431365
transform 1 0 28224 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output113
timestamp 1698431365
transform 1 0 26992 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output114
timestamp 1698431365
transform 1 0 55440 0 1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output115
timestamp 1698431365
transform 1 0 52528 0 1 36064
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output116
timestamp 1698431365
transform 1 0 53312 0 -1 36064
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output117
timestamp 1698431365
transform -1 0 4480 0 -1 39200
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output118
timestamp 1698431365
transform 1 0 55440 0 1 32928
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_94 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698431365
transform -1 0 58576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_95
timestamp 1698431365
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698431365
transform -1 0 58576 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_96
timestamp 1698431365
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698431365
transform -1 0 58576 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_97
timestamp 1698431365
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698431365
transform -1 0 58576 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_98
timestamp 1698431365
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698431365
transform -1 0 58576 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_99
timestamp 1698431365
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698431365
transform -1 0 58576 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_100
timestamp 1698431365
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698431365
transform -1 0 58576 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_101
timestamp 1698431365
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698431365
transform -1 0 58576 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_102
timestamp 1698431365
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698431365
transform -1 0 58576 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_103
timestamp 1698431365
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698431365
transform -1 0 58576 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_104
timestamp 1698431365
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698431365
transform -1 0 58576 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_105
timestamp 1698431365
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698431365
transform -1 0 58576 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_106
timestamp 1698431365
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698431365
transform -1 0 58576 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_107
timestamp 1698431365
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698431365
transform -1 0 58576 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_108
timestamp 1698431365
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698431365
transform -1 0 58576 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_109
timestamp 1698431365
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698431365
transform -1 0 58576 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_110
timestamp 1698431365
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698431365
transform -1 0 58576 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_111
timestamp 1698431365
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698431365
transform -1 0 58576 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_112
timestamp 1698431365
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698431365
transform -1 0 58576 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_113
timestamp 1698431365
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698431365
transform -1 0 58576 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_114
timestamp 1698431365
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698431365
transform -1 0 58576 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_115
timestamp 1698431365
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698431365
transform -1 0 58576 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_116
timestamp 1698431365
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1698431365
transform -1 0 58576 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_117
timestamp 1698431365
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1698431365
transform -1 0 58576 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_118
timestamp 1698431365
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1698431365
transform -1 0 58576 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_119
timestamp 1698431365
transform 1 0 1344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1698431365
transform -1 0 58576 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_120
timestamp 1698431365
transform 1 0 1344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1698431365
transform -1 0 58576 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_121
timestamp 1698431365
transform 1 0 1344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1698431365
transform -1 0 58576 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_122
timestamp 1698431365
transform 1 0 1344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1698431365
transform -1 0 58576 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_123
timestamp 1698431365
transform 1 0 1344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1698431365
transform -1 0 58576 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Left_124
timestamp 1698431365
transform 1 0 1344 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1698431365
transform -1 0 58576 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Left_125
timestamp 1698431365
transform 1 0 1344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1698431365
transform -1 0 58576 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Left_126
timestamp 1698431365
transform 1 0 1344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1698431365
transform -1 0 58576 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Left_127
timestamp 1698431365
transform 1 0 1344 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1698431365
transform -1 0 58576 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Left_128
timestamp 1698431365
transform 1 0 1344 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1698431365
transform -1 0 58576 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Left_129
timestamp 1698431365
transform 1 0 1344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Right_35
timestamp 1698431365
transform -1 0 58576 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Left_130
timestamp 1698431365
transform 1 0 1344 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Right_36
timestamp 1698431365
transform -1 0 58576 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Left_131
timestamp 1698431365
transform 1 0 1344 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Right_37
timestamp 1698431365
transform -1 0 58576 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Left_132
timestamp 1698431365
transform 1 0 1344 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Right_38
timestamp 1698431365
transform -1 0 58576 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Left_133
timestamp 1698431365
transform 1 0 1344 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Right_39
timestamp 1698431365
transform -1 0 58576 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Left_134
timestamp 1698431365
transform 1 0 1344 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Right_40
timestamp 1698431365
transform -1 0 58576 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Left_135
timestamp 1698431365
transform 1 0 1344 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Right_41
timestamp 1698431365
transform -1 0 58576 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Left_136
timestamp 1698431365
transform 1 0 1344 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Right_42
timestamp 1698431365
transform -1 0 58576 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Left_137
timestamp 1698431365
transform 1 0 1344 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Right_43
timestamp 1698431365
transform -1 0 58576 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Left_138
timestamp 1698431365
transform 1 0 1344 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Right_44
timestamp 1698431365
transform -1 0 58576 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_45_Left_139
timestamp 1698431365
transform 1 0 1344 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_45_Right_45
timestamp 1698431365
transform -1 0 58576 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_46_Left_140
timestamp 1698431365
transform 1 0 1344 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_46_Right_46
timestamp 1698431365
transform -1 0 58576 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_47_Left_141
timestamp 1698431365
transform 1 0 1344 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_47_Right_47
timestamp 1698431365
transform -1 0 58576 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_48_Left_142
timestamp 1698431365
transform 1 0 1344 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_48_Right_48
timestamp 1698431365
transform -1 0 58576 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_49_Left_143
timestamp 1698431365
transform 1 0 1344 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_49_Right_49
timestamp 1698431365
transform -1 0 58576 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_50_Left_144
timestamp 1698431365
transform 1 0 1344 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_50_Right_50
timestamp 1698431365
transform -1 0 58576 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_51_Left_145
timestamp 1698431365
transform 1 0 1344 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_51_Right_51
timestamp 1698431365
transform -1 0 58576 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_52_Left_146
timestamp 1698431365
transform 1 0 1344 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_52_Right_52
timestamp 1698431365
transform -1 0 58576 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_53_Left_147
timestamp 1698431365
transform 1 0 1344 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_53_Right_53
timestamp 1698431365
transform -1 0 58576 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_54_Left_148
timestamp 1698431365
transform 1 0 1344 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_54_Right_54
timestamp 1698431365
transform -1 0 58576 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_55_Left_149
timestamp 1698431365
transform 1 0 1344 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_55_Right_55
timestamp 1698431365
transform -1 0 58576 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_56_Left_150
timestamp 1698431365
transform 1 0 1344 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_56_Right_56
timestamp 1698431365
transform -1 0 58576 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_57_Left_151
timestamp 1698431365
transform 1 0 1344 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_57_Right_57
timestamp 1698431365
transform -1 0 58576 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_58_Left_152
timestamp 1698431365
transform 1 0 1344 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_58_Right_58
timestamp 1698431365
transform -1 0 58576 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_59_Left_153
timestamp 1698431365
transform 1 0 1344 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_59_Right_59
timestamp 1698431365
transform -1 0 58576 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_60_Left_154
timestamp 1698431365
transform 1 0 1344 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_60_Right_60
timestamp 1698431365
transform -1 0 58576 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_61_Left_155
timestamp 1698431365
transform 1 0 1344 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_61_Right_61
timestamp 1698431365
transform -1 0 58576 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_62_Left_156
timestamp 1698431365
transform 1 0 1344 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_62_Right_62
timestamp 1698431365
transform -1 0 58576 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_63_Left_157
timestamp 1698431365
transform 1 0 1344 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_63_Right_63
timestamp 1698431365
transform -1 0 58576 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_64_Left_158
timestamp 1698431365
transform 1 0 1344 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_64_Right_64
timestamp 1698431365
transform -1 0 58576 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_65_Left_159
timestamp 1698431365
transform 1 0 1344 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_65_Right_65
timestamp 1698431365
transform -1 0 58576 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_66_Left_160
timestamp 1698431365
transform 1 0 1344 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_66_Right_66
timestamp 1698431365
transform -1 0 58576 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_67_Left_161
timestamp 1698431365
transform 1 0 1344 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_67_Right_67
timestamp 1698431365
transform -1 0 58576 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_68_Left_162
timestamp 1698431365
transform 1 0 1344 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_68_Right_68
timestamp 1698431365
transform -1 0 58576 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_69_Left_163
timestamp 1698431365
transform 1 0 1344 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_69_Right_69
timestamp 1698431365
transform -1 0 58576 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_70_Left_164
timestamp 1698431365
transform 1 0 1344 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_70_Right_70
timestamp 1698431365
transform -1 0 58576 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_71_Left_165
timestamp 1698431365
transform 1 0 1344 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_71_Right_71
timestamp 1698431365
transform -1 0 58576 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_72_Left_166
timestamp 1698431365
transform 1 0 1344 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_72_Right_72
timestamp 1698431365
transform -1 0 58576 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_73_Left_167
timestamp 1698431365
transform 1 0 1344 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_73_Right_73
timestamp 1698431365
transform -1 0 58576 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_74_Left_168
timestamp 1698431365
transform 1 0 1344 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_74_Right_74
timestamp 1698431365
transform -1 0 58576 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_75_Left_169
timestamp 1698431365
transform 1 0 1344 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_75_Right_75
timestamp 1698431365
transform -1 0 58576 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_76_Left_170
timestamp 1698431365
transform 1 0 1344 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_76_Right_76
timestamp 1698431365
transform -1 0 58576 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_77_Left_171
timestamp 1698431365
transform 1 0 1344 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_77_Right_77
timestamp 1698431365
transform -1 0 58576 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_78_Left_172
timestamp 1698431365
transform 1 0 1344 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_78_Right_78
timestamp 1698431365
transform -1 0 58576 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_79_Left_173
timestamp 1698431365
transform 1 0 1344 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_79_Right_79
timestamp 1698431365
transform -1 0 58576 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_80_Left_174
timestamp 1698431365
transform 1 0 1344 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_80_Right_80
timestamp 1698431365
transform -1 0 58576 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_81_Left_175
timestamp 1698431365
transform 1 0 1344 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_81_Right_81
timestamp 1698431365
transform -1 0 58576 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_82_Left_176
timestamp 1698431365
transform 1 0 1344 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_82_Right_82
timestamp 1698431365
transform -1 0 58576 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_83_Left_177
timestamp 1698431365
transform 1 0 1344 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_83_Right_83
timestamp 1698431365
transform -1 0 58576 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_84_Left_178
timestamp 1698431365
transform 1 0 1344 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_84_Right_84
timestamp 1698431365
transform -1 0 58576 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_85_Left_179
timestamp 1698431365
transform 1 0 1344 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_85_Right_85
timestamp 1698431365
transform -1 0 58576 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_86_Left_180
timestamp 1698431365
transform 1 0 1344 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_86_Right_86
timestamp 1698431365
transform -1 0 58576 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_87_Left_181
timestamp 1698431365
transform 1 0 1344 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_87_Right_87
timestamp 1698431365
transform -1 0 58576 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_88_Left_182
timestamp 1698431365
transform 1 0 1344 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_88_Right_88
timestamp 1698431365
transform -1 0 58576 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_89_Left_183
timestamp 1698431365
transform 1 0 1344 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_89_Right_89
timestamp 1698431365
transform -1 0 58576 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_90_Left_184
timestamp 1698431365
transform 1 0 1344 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_90_Right_90
timestamp 1698431365
transform -1 0 58576 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_91_Left_185
timestamp 1698431365
transform 1 0 1344 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_91_Right_91
timestamp 1698431365
transform -1 0 58576 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_92_Left_186
timestamp 1698431365
transform 1 0 1344 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_92_Right_92
timestamp 1698431365
transform -1 0 58576 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_93_Left_187
timestamp 1698431365
transform 1 0 1344 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_93_Right_93
timestamp 1698431365
transform -1 0 58576 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_188 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5152 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_189
timestamp 1698431365
transform 1 0 8960 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_190
timestamp 1698431365
transform 1 0 12768 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_191
timestamp 1698431365
transform 1 0 16576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_192
timestamp 1698431365
transform 1 0 20384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_193
timestamp 1698431365
transform 1 0 24192 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_194
timestamp 1698431365
transform 1 0 28000 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_195
timestamp 1698431365
transform 1 0 31808 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_196
timestamp 1698431365
transform 1 0 35616 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_197
timestamp 1698431365
transform 1 0 39424 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_198
timestamp 1698431365
transform 1 0 43232 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_199
timestamp 1698431365
transform 1 0 47040 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_200
timestamp 1698431365
transform 1 0 50848 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_201
timestamp 1698431365
transform 1 0 54656 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_202
timestamp 1698431365
transform 1 0 9184 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_203
timestamp 1698431365
transform 1 0 17024 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_204
timestamp 1698431365
transform 1 0 24864 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_205
timestamp 1698431365
transform 1 0 32704 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_206
timestamp 1698431365
transform 1 0 40544 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_207
timestamp 1698431365
transform 1 0 48384 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_208
timestamp 1698431365
transform 1 0 56224 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_209
timestamp 1698431365
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_210
timestamp 1698431365
transform 1 0 13104 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_211
timestamp 1698431365
transform 1 0 20944 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_212
timestamp 1698431365
transform 1 0 28784 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_213
timestamp 1698431365
transform 1 0 36624 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_214
timestamp 1698431365
transform 1 0 44464 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_215
timestamp 1698431365
transform 1 0 52304 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_216
timestamp 1698431365
transform 1 0 9184 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_217
timestamp 1698431365
transform 1 0 17024 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_218
timestamp 1698431365
transform 1 0 24864 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_219
timestamp 1698431365
transform 1 0 32704 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_220
timestamp 1698431365
transform 1 0 40544 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_221
timestamp 1698431365
transform 1 0 48384 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_222
timestamp 1698431365
transform 1 0 56224 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_223
timestamp 1698431365
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_224
timestamp 1698431365
transform 1 0 13104 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_225
timestamp 1698431365
transform 1 0 20944 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_226
timestamp 1698431365
transform 1 0 28784 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_227
timestamp 1698431365
transform 1 0 36624 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_228
timestamp 1698431365
transform 1 0 44464 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_229
timestamp 1698431365
transform 1 0 52304 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_230
timestamp 1698431365
transform 1 0 9184 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_231
timestamp 1698431365
transform 1 0 17024 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_232
timestamp 1698431365
transform 1 0 24864 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_233
timestamp 1698431365
transform 1 0 32704 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_234
timestamp 1698431365
transform 1 0 40544 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_235
timestamp 1698431365
transform 1 0 48384 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_236
timestamp 1698431365
transform 1 0 56224 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_237
timestamp 1698431365
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_238
timestamp 1698431365
transform 1 0 13104 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_239
timestamp 1698431365
transform 1 0 20944 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_240
timestamp 1698431365
transform 1 0 28784 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_241
timestamp 1698431365
transform 1 0 36624 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_242
timestamp 1698431365
transform 1 0 44464 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_243
timestamp 1698431365
transform 1 0 52304 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_244
timestamp 1698431365
transform 1 0 9184 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_245
timestamp 1698431365
transform 1 0 17024 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_246
timestamp 1698431365
transform 1 0 24864 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_247
timestamp 1698431365
transform 1 0 32704 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_248
timestamp 1698431365
transform 1 0 40544 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_249
timestamp 1698431365
transform 1 0 48384 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_250
timestamp 1698431365
transform 1 0 56224 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_251
timestamp 1698431365
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_252
timestamp 1698431365
transform 1 0 13104 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_253
timestamp 1698431365
transform 1 0 20944 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_254
timestamp 1698431365
transform 1 0 28784 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_255
timestamp 1698431365
transform 1 0 36624 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_256
timestamp 1698431365
transform 1 0 44464 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_257
timestamp 1698431365
transform 1 0 52304 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_258
timestamp 1698431365
transform 1 0 9184 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_259
timestamp 1698431365
transform 1 0 17024 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_260
timestamp 1698431365
transform 1 0 24864 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_261
timestamp 1698431365
transform 1 0 32704 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_262
timestamp 1698431365
transform 1 0 40544 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_263
timestamp 1698431365
transform 1 0 48384 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_264
timestamp 1698431365
transform 1 0 56224 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_265
timestamp 1698431365
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_266
timestamp 1698431365
transform 1 0 13104 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_267
timestamp 1698431365
transform 1 0 20944 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_268
timestamp 1698431365
transform 1 0 28784 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_269
timestamp 1698431365
transform 1 0 36624 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_270
timestamp 1698431365
transform 1 0 44464 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_271
timestamp 1698431365
transform 1 0 52304 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_272
timestamp 1698431365
transform 1 0 9184 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_273
timestamp 1698431365
transform 1 0 17024 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_274
timestamp 1698431365
transform 1 0 24864 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_275
timestamp 1698431365
transform 1 0 32704 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_276
timestamp 1698431365
transform 1 0 40544 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_277
timestamp 1698431365
transform 1 0 48384 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_278
timestamp 1698431365
transform 1 0 56224 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_279
timestamp 1698431365
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_280
timestamp 1698431365
transform 1 0 13104 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_281
timestamp 1698431365
transform 1 0 20944 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_282
timestamp 1698431365
transform 1 0 28784 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_283
timestamp 1698431365
transform 1 0 36624 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_284
timestamp 1698431365
transform 1 0 44464 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_285
timestamp 1698431365
transform 1 0 52304 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_286
timestamp 1698431365
transform 1 0 9184 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_287
timestamp 1698431365
transform 1 0 17024 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_288
timestamp 1698431365
transform 1 0 24864 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_289
timestamp 1698431365
transform 1 0 32704 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_290
timestamp 1698431365
transform 1 0 40544 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_291
timestamp 1698431365
transform 1 0 48384 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_292
timestamp 1698431365
transform 1 0 56224 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_293
timestamp 1698431365
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_294
timestamp 1698431365
transform 1 0 13104 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_295
timestamp 1698431365
transform 1 0 20944 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_296
timestamp 1698431365
transform 1 0 28784 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_297
timestamp 1698431365
transform 1 0 36624 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_298
timestamp 1698431365
transform 1 0 44464 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_299
timestamp 1698431365
transform 1 0 52304 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_300
timestamp 1698431365
transform 1 0 9184 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_301
timestamp 1698431365
transform 1 0 17024 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_302
timestamp 1698431365
transform 1 0 24864 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_303
timestamp 1698431365
transform 1 0 32704 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_304
timestamp 1698431365
transform 1 0 40544 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_305
timestamp 1698431365
transform 1 0 48384 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_306
timestamp 1698431365
transform 1 0 56224 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_307
timestamp 1698431365
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_308
timestamp 1698431365
transform 1 0 13104 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_309
timestamp 1698431365
transform 1 0 20944 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_310
timestamp 1698431365
transform 1 0 28784 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_311
timestamp 1698431365
transform 1 0 36624 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_312
timestamp 1698431365
transform 1 0 44464 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_313
timestamp 1698431365
transform 1 0 52304 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_314
timestamp 1698431365
transform 1 0 9184 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_315
timestamp 1698431365
transform 1 0 17024 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_316
timestamp 1698431365
transform 1 0 24864 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_317
timestamp 1698431365
transform 1 0 32704 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_318
timestamp 1698431365
transform 1 0 40544 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_319
timestamp 1698431365
transform 1 0 48384 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_320
timestamp 1698431365
transform 1 0 56224 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_321
timestamp 1698431365
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_322
timestamp 1698431365
transform 1 0 13104 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_323
timestamp 1698431365
transform 1 0 20944 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_324
timestamp 1698431365
transform 1 0 28784 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_325
timestamp 1698431365
transform 1 0 36624 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_326
timestamp 1698431365
transform 1 0 44464 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_327
timestamp 1698431365
transform 1 0 52304 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_328
timestamp 1698431365
transform 1 0 9184 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_329
timestamp 1698431365
transform 1 0 17024 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_330
timestamp 1698431365
transform 1 0 24864 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_331
timestamp 1698431365
transform 1 0 32704 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_332
timestamp 1698431365
transform 1 0 40544 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_333
timestamp 1698431365
transform 1 0 48384 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_334
timestamp 1698431365
transform 1 0 56224 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_335
timestamp 1698431365
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_336
timestamp 1698431365
transform 1 0 13104 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_337
timestamp 1698431365
transform 1 0 20944 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_338
timestamp 1698431365
transform 1 0 28784 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_339
timestamp 1698431365
transform 1 0 36624 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_340
timestamp 1698431365
transform 1 0 44464 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_341
timestamp 1698431365
transform 1 0 52304 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_342
timestamp 1698431365
transform 1 0 9184 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_343
timestamp 1698431365
transform 1 0 17024 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_344
timestamp 1698431365
transform 1 0 24864 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_345
timestamp 1698431365
transform 1 0 32704 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_346
timestamp 1698431365
transform 1 0 40544 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_347
timestamp 1698431365
transform 1 0 48384 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_348
timestamp 1698431365
transform 1 0 56224 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_349
timestamp 1698431365
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_350
timestamp 1698431365
transform 1 0 13104 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_351
timestamp 1698431365
transform 1 0 20944 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_352
timestamp 1698431365
transform 1 0 28784 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_353
timestamp 1698431365
transform 1 0 36624 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_354
timestamp 1698431365
transform 1 0 44464 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_355
timestamp 1698431365
transform 1 0 52304 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_356
timestamp 1698431365
transform 1 0 9184 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_357
timestamp 1698431365
transform 1 0 17024 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_358
timestamp 1698431365
transform 1 0 24864 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_359
timestamp 1698431365
transform 1 0 32704 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_360
timestamp 1698431365
transform 1 0 40544 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_361
timestamp 1698431365
transform 1 0 48384 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_362
timestamp 1698431365
transform 1 0 56224 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_363
timestamp 1698431365
transform 1 0 5264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_364
timestamp 1698431365
transform 1 0 13104 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_365
timestamp 1698431365
transform 1 0 20944 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_366
timestamp 1698431365
transform 1 0 28784 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_367
timestamp 1698431365
transform 1 0 36624 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_368
timestamp 1698431365
transform 1 0 44464 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_369
timestamp 1698431365
transform 1 0 52304 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_370
timestamp 1698431365
transform 1 0 9184 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_371
timestamp 1698431365
transform 1 0 17024 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_372
timestamp 1698431365
transform 1 0 24864 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_373
timestamp 1698431365
transform 1 0 32704 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_374
timestamp 1698431365
transform 1 0 40544 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_375
timestamp 1698431365
transform 1 0 48384 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_376
timestamp 1698431365
transform 1 0 56224 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_377
timestamp 1698431365
transform 1 0 5264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_378
timestamp 1698431365
transform 1 0 13104 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_379
timestamp 1698431365
transform 1 0 20944 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_380
timestamp 1698431365
transform 1 0 28784 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_381
timestamp 1698431365
transform 1 0 36624 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_382
timestamp 1698431365
transform 1 0 44464 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_383
timestamp 1698431365
transform 1 0 52304 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_384
timestamp 1698431365
transform 1 0 9184 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_385
timestamp 1698431365
transform 1 0 17024 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_386
timestamp 1698431365
transform 1 0 24864 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_387
timestamp 1698431365
transform 1 0 32704 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_388
timestamp 1698431365
transform 1 0 40544 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_389
timestamp 1698431365
transform 1 0 48384 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_390
timestamp 1698431365
transform 1 0 56224 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_391
timestamp 1698431365
transform 1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_392
timestamp 1698431365
transform 1 0 13104 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_393
timestamp 1698431365
transform 1 0 20944 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_394
timestamp 1698431365
transform 1 0 28784 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_395
timestamp 1698431365
transform 1 0 36624 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_396
timestamp 1698431365
transform 1 0 44464 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_397
timestamp 1698431365
transform 1 0 52304 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_398
timestamp 1698431365
transform 1 0 9184 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_399
timestamp 1698431365
transform 1 0 17024 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_400
timestamp 1698431365
transform 1 0 24864 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_401
timestamp 1698431365
transform 1 0 32704 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_402
timestamp 1698431365
transform 1 0 40544 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_403
timestamp 1698431365
transform 1 0 48384 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_404
timestamp 1698431365
transform 1 0 56224 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_405
timestamp 1698431365
transform 1 0 5264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_406
timestamp 1698431365
transform 1 0 13104 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_407
timestamp 1698431365
transform 1 0 20944 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_408
timestamp 1698431365
transform 1 0 28784 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_409
timestamp 1698431365
transform 1 0 36624 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_410
timestamp 1698431365
transform 1 0 44464 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_411
timestamp 1698431365
transform 1 0 52304 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_412
timestamp 1698431365
transform 1 0 9184 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_413
timestamp 1698431365
transform 1 0 17024 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_414
timestamp 1698431365
transform 1 0 24864 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_415
timestamp 1698431365
transform 1 0 32704 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_416
timestamp 1698431365
transform 1 0 40544 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_417
timestamp 1698431365
transform 1 0 48384 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_418
timestamp 1698431365
transform 1 0 56224 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_419
timestamp 1698431365
transform 1 0 5264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_420
timestamp 1698431365
transform 1 0 13104 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_421
timestamp 1698431365
transform 1 0 20944 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_422
timestamp 1698431365
transform 1 0 28784 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_423
timestamp 1698431365
transform 1 0 36624 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_424
timestamp 1698431365
transform 1 0 44464 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_425
timestamp 1698431365
transform 1 0 52304 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_426
timestamp 1698431365
transform 1 0 9184 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_427
timestamp 1698431365
transform 1 0 17024 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_428
timestamp 1698431365
transform 1 0 24864 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_429
timestamp 1698431365
transform 1 0 32704 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_430
timestamp 1698431365
transform 1 0 40544 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_431
timestamp 1698431365
transform 1 0 48384 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_432
timestamp 1698431365
transform 1 0 56224 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_433
timestamp 1698431365
transform 1 0 5264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_434
timestamp 1698431365
transform 1 0 13104 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_435
timestamp 1698431365
transform 1 0 20944 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_436
timestamp 1698431365
transform 1 0 28784 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_437
timestamp 1698431365
transform 1 0 36624 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_438
timestamp 1698431365
transform 1 0 44464 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_439
timestamp 1698431365
transform 1 0 52304 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_440
timestamp 1698431365
transform 1 0 9184 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_441
timestamp 1698431365
transform 1 0 17024 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_442
timestamp 1698431365
transform 1 0 24864 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_443
timestamp 1698431365
transform 1 0 32704 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_444
timestamp 1698431365
transform 1 0 40544 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_445
timestamp 1698431365
transform 1 0 48384 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_446
timestamp 1698431365
transform 1 0 56224 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_447
timestamp 1698431365
transform 1 0 5264 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_448
timestamp 1698431365
transform 1 0 13104 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_449
timestamp 1698431365
transform 1 0 20944 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_450
timestamp 1698431365
transform 1 0 28784 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_451
timestamp 1698431365
transform 1 0 36624 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_452
timestamp 1698431365
transform 1 0 44464 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_453
timestamp 1698431365
transform 1 0 52304 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_454
timestamp 1698431365
transform 1 0 9184 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_455
timestamp 1698431365
transform 1 0 17024 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_456
timestamp 1698431365
transform 1 0 24864 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_457
timestamp 1698431365
transform 1 0 32704 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_458
timestamp 1698431365
transform 1 0 40544 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_459
timestamp 1698431365
transform 1 0 48384 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_460
timestamp 1698431365
transform 1 0 56224 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_461
timestamp 1698431365
transform 1 0 5264 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_462
timestamp 1698431365
transform 1 0 13104 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_463
timestamp 1698431365
transform 1 0 20944 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_464
timestamp 1698431365
transform 1 0 28784 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_465
timestamp 1698431365
transform 1 0 36624 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_466
timestamp 1698431365
transform 1 0 44464 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_467
timestamp 1698431365
transform 1 0 52304 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_468
timestamp 1698431365
transform 1 0 9184 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_469
timestamp 1698431365
transform 1 0 17024 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_470
timestamp 1698431365
transform 1 0 24864 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_471
timestamp 1698431365
transform 1 0 32704 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_472
timestamp 1698431365
transform 1 0 40544 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_473
timestamp 1698431365
transform 1 0 48384 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_474
timestamp 1698431365
transform 1 0 56224 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_475
timestamp 1698431365
transform 1 0 5264 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_476
timestamp 1698431365
transform 1 0 13104 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_477
timestamp 1698431365
transform 1 0 20944 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_478
timestamp 1698431365
transform 1 0 28784 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_479
timestamp 1698431365
transform 1 0 36624 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_480
timestamp 1698431365
transform 1 0 44464 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_481
timestamp 1698431365
transform 1 0 52304 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_482
timestamp 1698431365
transform 1 0 9184 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_483
timestamp 1698431365
transform 1 0 17024 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_484
timestamp 1698431365
transform 1 0 24864 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_485
timestamp 1698431365
transform 1 0 32704 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_486
timestamp 1698431365
transform 1 0 40544 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_487
timestamp 1698431365
transform 1 0 48384 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_488
timestamp 1698431365
transform 1 0 56224 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_489
timestamp 1698431365
transform 1 0 5264 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_490
timestamp 1698431365
transform 1 0 13104 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_491
timestamp 1698431365
transform 1 0 20944 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_492
timestamp 1698431365
transform 1 0 28784 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_493
timestamp 1698431365
transform 1 0 36624 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_494
timestamp 1698431365
transform 1 0 44464 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_495
timestamp 1698431365
transform 1 0 52304 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_496
timestamp 1698431365
transform 1 0 9184 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_497
timestamp 1698431365
transform 1 0 17024 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_498
timestamp 1698431365
transform 1 0 24864 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_499
timestamp 1698431365
transform 1 0 32704 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_500
timestamp 1698431365
transform 1 0 40544 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_501
timestamp 1698431365
transform 1 0 48384 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_502
timestamp 1698431365
transform 1 0 56224 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_503
timestamp 1698431365
transform 1 0 5264 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_504
timestamp 1698431365
transform 1 0 13104 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_505
timestamp 1698431365
transform 1 0 20944 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_506
timestamp 1698431365
transform 1 0 28784 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_507
timestamp 1698431365
transform 1 0 36624 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_508
timestamp 1698431365
transform 1 0 44464 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_509
timestamp 1698431365
transform 1 0 52304 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_510
timestamp 1698431365
transform 1 0 9184 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_511
timestamp 1698431365
transform 1 0 17024 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_512
timestamp 1698431365
transform 1 0 24864 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_513
timestamp 1698431365
transform 1 0 32704 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_514
timestamp 1698431365
transform 1 0 40544 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_515
timestamp 1698431365
transform 1 0 48384 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_516
timestamp 1698431365
transform 1 0 56224 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_517
timestamp 1698431365
transform 1 0 5264 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_518
timestamp 1698431365
transform 1 0 13104 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_519
timestamp 1698431365
transform 1 0 20944 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_520
timestamp 1698431365
transform 1 0 28784 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_521
timestamp 1698431365
transform 1 0 36624 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_522
timestamp 1698431365
transform 1 0 44464 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_523
timestamp 1698431365
transform 1 0 52304 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_524
timestamp 1698431365
transform 1 0 9184 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_525
timestamp 1698431365
transform 1 0 17024 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_526
timestamp 1698431365
transform 1 0 24864 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_527
timestamp 1698431365
transform 1 0 32704 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_528
timestamp 1698431365
transform 1 0 40544 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_529
timestamp 1698431365
transform 1 0 48384 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_530
timestamp 1698431365
transform 1 0 56224 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_531
timestamp 1698431365
transform 1 0 5264 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_532
timestamp 1698431365
transform 1 0 13104 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_533
timestamp 1698431365
transform 1 0 20944 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_534
timestamp 1698431365
transform 1 0 28784 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_535
timestamp 1698431365
transform 1 0 36624 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_536
timestamp 1698431365
transform 1 0 44464 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_537
timestamp 1698431365
transform 1 0 52304 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_538
timestamp 1698431365
transform 1 0 9184 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_539
timestamp 1698431365
transform 1 0 17024 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_540
timestamp 1698431365
transform 1 0 24864 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_541
timestamp 1698431365
transform 1 0 32704 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_542
timestamp 1698431365
transform 1 0 40544 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_543
timestamp 1698431365
transform 1 0 48384 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_544
timestamp 1698431365
transform 1 0 56224 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_545
timestamp 1698431365
transform 1 0 5264 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_546
timestamp 1698431365
transform 1 0 13104 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_547
timestamp 1698431365
transform 1 0 20944 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_548
timestamp 1698431365
transform 1 0 28784 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_549
timestamp 1698431365
transform 1 0 36624 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_550
timestamp 1698431365
transform 1 0 44464 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_551
timestamp 1698431365
transform 1 0 52304 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_552
timestamp 1698431365
transform 1 0 9184 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_553
timestamp 1698431365
transform 1 0 17024 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_554
timestamp 1698431365
transform 1 0 24864 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_555
timestamp 1698431365
transform 1 0 32704 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_556
timestamp 1698431365
transform 1 0 40544 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_557
timestamp 1698431365
transform 1 0 48384 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_558
timestamp 1698431365
transform 1 0 56224 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_559
timestamp 1698431365
transform 1 0 5264 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_560
timestamp 1698431365
transform 1 0 13104 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_561
timestamp 1698431365
transform 1 0 20944 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_562
timestamp 1698431365
transform 1 0 28784 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_563
timestamp 1698431365
transform 1 0 36624 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_564
timestamp 1698431365
transform 1 0 44464 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_565
timestamp 1698431365
transform 1 0 52304 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_566
timestamp 1698431365
transform 1 0 9184 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_567
timestamp 1698431365
transform 1 0 17024 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_568
timestamp 1698431365
transform 1 0 24864 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_569
timestamp 1698431365
transform 1 0 32704 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_570
timestamp 1698431365
transform 1 0 40544 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_571
timestamp 1698431365
transform 1 0 48384 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_572
timestamp 1698431365
transform 1 0 56224 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_573
timestamp 1698431365
transform 1 0 5264 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_574
timestamp 1698431365
transform 1 0 13104 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_575
timestamp 1698431365
transform 1 0 20944 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_576
timestamp 1698431365
transform 1 0 28784 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_577
timestamp 1698431365
transform 1 0 36624 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_578
timestamp 1698431365
transform 1 0 44464 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_579
timestamp 1698431365
transform 1 0 52304 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_580
timestamp 1698431365
transform 1 0 9184 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_581
timestamp 1698431365
transform 1 0 17024 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_582
timestamp 1698431365
transform 1 0 24864 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_583
timestamp 1698431365
transform 1 0 32704 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_584
timestamp 1698431365
transform 1 0 40544 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_585
timestamp 1698431365
transform 1 0 48384 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_586
timestamp 1698431365
transform 1 0 56224 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_587
timestamp 1698431365
transform 1 0 5264 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_588
timestamp 1698431365
transform 1 0 13104 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_589
timestamp 1698431365
transform 1 0 20944 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_590
timestamp 1698431365
transform 1 0 28784 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_591
timestamp 1698431365
transform 1 0 36624 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_592
timestamp 1698431365
transform 1 0 44464 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_593
timestamp 1698431365
transform 1 0 52304 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_594
timestamp 1698431365
transform 1 0 9184 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_595
timestamp 1698431365
transform 1 0 17024 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_596
timestamp 1698431365
transform 1 0 24864 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_597
timestamp 1698431365
transform 1 0 32704 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_598
timestamp 1698431365
transform 1 0 40544 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_599
timestamp 1698431365
transform 1 0 48384 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_600
timestamp 1698431365
transform 1 0 56224 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_601
timestamp 1698431365
transform 1 0 5264 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_602
timestamp 1698431365
transform 1 0 13104 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_603
timestamp 1698431365
transform 1 0 20944 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_604
timestamp 1698431365
transform 1 0 28784 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_605
timestamp 1698431365
transform 1 0 36624 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_606
timestamp 1698431365
transform 1 0 44464 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_607
timestamp 1698431365
transform 1 0 52304 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_608
timestamp 1698431365
transform 1 0 9184 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_609
timestamp 1698431365
transform 1 0 17024 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_610
timestamp 1698431365
transform 1 0 24864 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_611
timestamp 1698431365
transform 1 0 32704 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_612
timestamp 1698431365
transform 1 0 40544 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_613
timestamp 1698431365
transform 1 0 48384 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_614
timestamp 1698431365
transform 1 0 56224 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_615
timestamp 1698431365
transform 1 0 5264 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_616
timestamp 1698431365
transform 1 0 13104 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_617
timestamp 1698431365
transform 1 0 20944 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_618
timestamp 1698431365
transform 1 0 28784 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_619
timestamp 1698431365
transform 1 0 36624 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_620
timestamp 1698431365
transform 1 0 44464 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_621
timestamp 1698431365
transform 1 0 52304 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_622
timestamp 1698431365
transform 1 0 9184 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_623
timestamp 1698431365
transform 1 0 17024 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_624
timestamp 1698431365
transform 1 0 24864 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_625
timestamp 1698431365
transform 1 0 32704 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_626
timestamp 1698431365
transform 1 0 40544 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_627
timestamp 1698431365
transform 1 0 48384 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_628
timestamp 1698431365
transform 1 0 56224 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_629
timestamp 1698431365
transform 1 0 5264 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_630
timestamp 1698431365
transform 1 0 13104 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_631
timestamp 1698431365
transform 1 0 20944 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_632
timestamp 1698431365
transform 1 0 28784 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_633
timestamp 1698431365
transform 1 0 36624 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_634
timestamp 1698431365
transform 1 0 44464 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_635
timestamp 1698431365
transform 1 0 52304 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_636
timestamp 1698431365
transform 1 0 9184 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_637
timestamp 1698431365
transform 1 0 17024 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_638
timestamp 1698431365
transform 1 0 24864 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_639
timestamp 1698431365
transform 1 0 32704 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_640
timestamp 1698431365
transform 1 0 40544 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_641
timestamp 1698431365
transform 1 0 48384 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_642
timestamp 1698431365
transform 1 0 56224 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_643
timestamp 1698431365
transform 1 0 5264 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_644
timestamp 1698431365
transform 1 0 13104 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_645
timestamp 1698431365
transform 1 0 20944 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_646
timestamp 1698431365
transform 1 0 28784 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_647
timestamp 1698431365
transform 1 0 36624 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_648
timestamp 1698431365
transform 1 0 44464 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_649
timestamp 1698431365
transform 1 0 52304 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_650
timestamp 1698431365
transform 1 0 9184 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_651
timestamp 1698431365
transform 1 0 17024 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_652
timestamp 1698431365
transform 1 0 24864 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_653
timestamp 1698431365
transform 1 0 32704 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_654
timestamp 1698431365
transform 1 0 40544 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_655
timestamp 1698431365
transform 1 0 48384 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_656
timestamp 1698431365
transform 1 0 56224 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_657
timestamp 1698431365
transform 1 0 5264 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_658
timestamp 1698431365
transform 1 0 13104 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_659
timestamp 1698431365
transform 1 0 20944 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_660
timestamp 1698431365
transform 1 0 28784 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_661
timestamp 1698431365
transform 1 0 36624 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_662
timestamp 1698431365
transform 1 0 44464 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_663
timestamp 1698431365
transform 1 0 52304 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_664
timestamp 1698431365
transform 1 0 9184 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_665
timestamp 1698431365
transform 1 0 17024 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_666
timestamp 1698431365
transform 1 0 24864 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_667
timestamp 1698431365
transform 1 0 32704 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_668
timestamp 1698431365
transform 1 0 40544 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_669
timestamp 1698431365
transform 1 0 48384 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_670
timestamp 1698431365
transform 1 0 56224 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_68_671
timestamp 1698431365
transform 1 0 5264 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_68_672
timestamp 1698431365
transform 1 0 13104 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_68_673
timestamp 1698431365
transform 1 0 20944 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_68_674
timestamp 1698431365
transform 1 0 28784 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_68_675
timestamp 1698431365
transform 1 0 36624 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_68_676
timestamp 1698431365
transform 1 0 44464 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_68_677
timestamp 1698431365
transform 1 0 52304 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_69_678
timestamp 1698431365
transform 1 0 9184 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_69_679
timestamp 1698431365
transform 1 0 17024 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_69_680
timestamp 1698431365
transform 1 0 24864 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_69_681
timestamp 1698431365
transform 1 0 32704 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_69_682
timestamp 1698431365
transform 1 0 40544 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_69_683
timestamp 1698431365
transform 1 0 48384 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_69_684
timestamp 1698431365
transform 1 0 56224 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_685
timestamp 1698431365
transform 1 0 5264 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_686
timestamp 1698431365
transform 1 0 13104 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_687
timestamp 1698431365
transform 1 0 20944 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_688
timestamp 1698431365
transform 1 0 28784 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_689
timestamp 1698431365
transform 1 0 36624 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_690
timestamp 1698431365
transform 1 0 44464 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_691
timestamp 1698431365
transform 1 0 52304 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_71_692
timestamp 1698431365
transform 1 0 9184 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_71_693
timestamp 1698431365
transform 1 0 17024 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_71_694
timestamp 1698431365
transform 1 0 24864 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_71_695
timestamp 1698431365
transform 1 0 32704 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_71_696
timestamp 1698431365
transform 1 0 40544 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_71_697
timestamp 1698431365
transform 1 0 48384 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_71_698
timestamp 1698431365
transform 1 0 56224 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_72_699
timestamp 1698431365
transform 1 0 5264 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_72_700
timestamp 1698431365
transform 1 0 13104 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_72_701
timestamp 1698431365
transform 1 0 20944 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_72_702
timestamp 1698431365
transform 1 0 28784 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_72_703
timestamp 1698431365
transform 1 0 36624 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_72_704
timestamp 1698431365
transform 1 0 44464 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_72_705
timestamp 1698431365
transform 1 0 52304 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_73_706
timestamp 1698431365
transform 1 0 9184 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_73_707
timestamp 1698431365
transform 1 0 17024 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_73_708
timestamp 1698431365
transform 1 0 24864 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_73_709
timestamp 1698431365
transform 1 0 32704 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_73_710
timestamp 1698431365
transform 1 0 40544 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_73_711
timestamp 1698431365
transform 1 0 48384 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_73_712
timestamp 1698431365
transform 1 0 56224 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_74_713
timestamp 1698431365
transform 1 0 5264 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_74_714
timestamp 1698431365
transform 1 0 13104 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_74_715
timestamp 1698431365
transform 1 0 20944 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_74_716
timestamp 1698431365
transform 1 0 28784 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_74_717
timestamp 1698431365
transform 1 0 36624 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_74_718
timestamp 1698431365
transform 1 0 44464 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_74_719
timestamp 1698431365
transform 1 0 52304 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_75_720
timestamp 1698431365
transform 1 0 9184 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_75_721
timestamp 1698431365
transform 1 0 17024 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_75_722
timestamp 1698431365
transform 1 0 24864 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_75_723
timestamp 1698431365
transform 1 0 32704 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_75_724
timestamp 1698431365
transform 1 0 40544 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_75_725
timestamp 1698431365
transform 1 0 48384 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_75_726
timestamp 1698431365
transform 1 0 56224 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_76_727
timestamp 1698431365
transform 1 0 5264 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_76_728
timestamp 1698431365
transform 1 0 13104 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_76_729
timestamp 1698431365
transform 1 0 20944 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_76_730
timestamp 1698431365
transform 1 0 28784 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_76_731
timestamp 1698431365
transform 1 0 36624 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_76_732
timestamp 1698431365
transform 1 0 44464 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_76_733
timestamp 1698431365
transform 1 0 52304 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_77_734
timestamp 1698431365
transform 1 0 9184 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_77_735
timestamp 1698431365
transform 1 0 17024 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_77_736
timestamp 1698431365
transform 1 0 24864 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_77_737
timestamp 1698431365
transform 1 0 32704 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_77_738
timestamp 1698431365
transform 1 0 40544 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_77_739
timestamp 1698431365
transform 1 0 48384 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_77_740
timestamp 1698431365
transform 1 0 56224 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_78_741
timestamp 1698431365
transform 1 0 5264 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_78_742
timestamp 1698431365
transform 1 0 13104 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_78_743
timestamp 1698431365
transform 1 0 20944 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_78_744
timestamp 1698431365
transform 1 0 28784 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_78_745
timestamp 1698431365
transform 1 0 36624 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_78_746
timestamp 1698431365
transform 1 0 44464 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_78_747
timestamp 1698431365
transform 1 0 52304 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_79_748
timestamp 1698431365
transform 1 0 9184 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_79_749
timestamp 1698431365
transform 1 0 17024 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_79_750
timestamp 1698431365
transform 1 0 24864 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_79_751
timestamp 1698431365
transform 1 0 32704 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_79_752
timestamp 1698431365
transform 1 0 40544 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_79_753
timestamp 1698431365
transform 1 0 48384 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_79_754
timestamp 1698431365
transform 1 0 56224 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_80_755
timestamp 1698431365
transform 1 0 5264 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_80_756
timestamp 1698431365
transform 1 0 13104 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_80_757
timestamp 1698431365
transform 1 0 20944 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_80_758
timestamp 1698431365
transform 1 0 28784 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_80_759
timestamp 1698431365
transform 1 0 36624 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_80_760
timestamp 1698431365
transform 1 0 44464 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_80_761
timestamp 1698431365
transform 1 0 52304 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_81_762
timestamp 1698431365
transform 1 0 9184 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_81_763
timestamp 1698431365
transform 1 0 17024 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_81_764
timestamp 1698431365
transform 1 0 24864 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_81_765
timestamp 1698431365
transform 1 0 32704 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_81_766
timestamp 1698431365
transform 1 0 40544 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_81_767
timestamp 1698431365
transform 1 0 48384 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_81_768
timestamp 1698431365
transform 1 0 56224 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_82_769
timestamp 1698431365
transform 1 0 5264 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_82_770
timestamp 1698431365
transform 1 0 13104 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_82_771
timestamp 1698431365
transform 1 0 20944 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_82_772
timestamp 1698431365
transform 1 0 28784 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_82_773
timestamp 1698431365
transform 1 0 36624 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_82_774
timestamp 1698431365
transform 1 0 44464 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_82_775
timestamp 1698431365
transform 1 0 52304 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_83_776
timestamp 1698431365
transform 1 0 9184 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_83_777
timestamp 1698431365
transform 1 0 17024 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_83_778
timestamp 1698431365
transform 1 0 24864 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_83_779
timestamp 1698431365
transform 1 0 32704 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_83_780
timestamp 1698431365
transform 1 0 40544 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_83_781
timestamp 1698431365
transform 1 0 48384 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_83_782
timestamp 1698431365
transform 1 0 56224 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_84_783
timestamp 1698431365
transform 1 0 5264 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_84_784
timestamp 1698431365
transform 1 0 13104 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_84_785
timestamp 1698431365
transform 1 0 20944 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_84_786
timestamp 1698431365
transform 1 0 28784 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_84_787
timestamp 1698431365
transform 1 0 36624 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_84_788
timestamp 1698431365
transform 1 0 44464 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_84_789
timestamp 1698431365
transform 1 0 52304 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_85_790
timestamp 1698431365
transform 1 0 9184 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_85_791
timestamp 1698431365
transform 1 0 17024 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_85_792
timestamp 1698431365
transform 1 0 24864 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_85_793
timestamp 1698431365
transform 1 0 32704 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_85_794
timestamp 1698431365
transform 1 0 40544 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_85_795
timestamp 1698431365
transform 1 0 48384 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_85_796
timestamp 1698431365
transform 1 0 56224 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_86_797
timestamp 1698431365
transform 1 0 5264 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_86_798
timestamp 1698431365
transform 1 0 13104 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_86_799
timestamp 1698431365
transform 1 0 20944 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_86_800
timestamp 1698431365
transform 1 0 28784 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_86_801
timestamp 1698431365
transform 1 0 36624 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_86_802
timestamp 1698431365
transform 1 0 44464 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_86_803
timestamp 1698431365
transform 1 0 52304 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_87_804
timestamp 1698431365
transform 1 0 9184 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_87_805
timestamp 1698431365
transform 1 0 17024 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_87_806
timestamp 1698431365
transform 1 0 24864 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_87_807
timestamp 1698431365
transform 1 0 32704 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_87_808
timestamp 1698431365
transform 1 0 40544 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_87_809
timestamp 1698431365
transform 1 0 48384 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_87_810
timestamp 1698431365
transform 1 0 56224 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_88_811
timestamp 1698431365
transform 1 0 5264 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_88_812
timestamp 1698431365
transform 1 0 13104 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_88_813
timestamp 1698431365
transform 1 0 20944 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_88_814
timestamp 1698431365
transform 1 0 28784 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_88_815
timestamp 1698431365
transform 1 0 36624 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_88_816
timestamp 1698431365
transform 1 0 44464 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_88_817
timestamp 1698431365
transform 1 0 52304 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_89_818
timestamp 1698431365
transform 1 0 9184 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_89_819
timestamp 1698431365
transform 1 0 17024 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_89_820
timestamp 1698431365
transform 1 0 24864 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_89_821
timestamp 1698431365
transform 1 0 32704 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_89_822
timestamp 1698431365
transform 1 0 40544 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_89_823
timestamp 1698431365
transform 1 0 48384 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_89_824
timestamp 1698431365
transform 1 0 56224 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_90_825
timestamp 1698431365
transform 1 0 5264 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_90_826
timestamp 1698431365
transform 1 0 13104 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_90_827
timestamp 1698431365
transform 1 0 20944 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_90_828
timestamp 1698431365
transform 1 0 28784 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_90_829
timestamp 1698431365
transform 1 0 36624 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_90_830
timestamp 1698431365
transform 1 0 44464 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_90_831
timestamp 1698431365
transform 1 0 52304 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_91_832
timestamp 1698431365
transform 1 0 9184 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_91_833
timestamp 1698431365
transform 1 0 17024 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_91_834
timestamp 1698431365
transform 1 0 24864 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_91_835
timestamp 1698431365
transform 1 0 32704 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_91_836
timestamp 1698431365
transform 1 0 40544 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_91_837
timestamp 1698431365
transform 1 0 48384 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_91_838
timestamp 1698431365
transform 1 0 56224 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_92_839
timestamp 1698431365
transform 1 0 5264 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_92_840
timestamp 1698431365
transform 1 0 13104 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_92_841
timestamp 1698431365
transform 1 0 20944 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_92_842
timestamp 1698431365
transform 1 0 28784 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_92_843
timestamp 1698431365
transform 1 0 36624 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_92_844
timestamp 1698431365
transform 1 0 44464 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_92_845
timestamp 1698431365
transform 1 0 52304 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_93_846
timestamp 1698431365
transform 1 0 5152 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_93_847
timestamp 1698431365
transform 1 0 8960 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_93_848
timestamp 1698431365
transform 1 0 12768 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_93_849
timestamp 1698431365
transform 1 0 16576 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_93_850
timestamp 1698431365
transform 1 0 20384 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_93_851
timestamp 1698431365
transform 1 0 24192 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_93_852
timestamp 1698431365
transform 1 0 28000 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_93_853
timestamp 1698431365
transform 1 0 31808 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_93_854
timestamp 1698431365
transform 1 0 35616 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_93_855
timestamp 1698431365
transform 1 0 39424 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_93_856
timestamp 1698431365
transform 1 0 43232 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_93_857
timestamp 1698431365
transform 1 0 47040 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_93_858
timestamp 1698431365
transform 1 0 50848 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_93_859
timestamp 1698431365
transform 1 0 54656 0 -1 76832
box -86 -86 310 870
<< labels >>
flabel metal3 s 0 70560 800 70672 0 FreeSans 448 0 0 0 clk
port 0 nsew signal input
flabel metal3 s 0 30912 800 31024 0 FreeSans 448 0 0 0 pcpi_insn[0]
port 1 nsew signal input
flabel metal2 s 0 0 112 800 0 FreeSans 448 90 0 0 pcpi_insn[10]
port 2 nsew signal input
flabel metal2 s 672 0 784 800 0 FreeSans 448 90 0 0 pcpi_insn[11]
port 3 nsew signal input
flabel metal3 s 0 53760 800 53872 0 FreeSans 448 0 0 0 pcpi_insn[12]
port 4 nsew signal input
flabel metal3 s 0 46368 800 46480 0 FreeSans 448 0 0 0 pcpi_insn[13]
port 5 nsew signal input
flabel metal3 s 0 45696 800 45808 0 FreeSans 448 0 0 0 pcpi_insn[14]
port 6 nsew signal input
flabel metal2 s 1344 0 1456 800 0 FreeSans 448 90 0 0 pcpi_insn[15]
port 7 nsew signal input
flabel metal2 s 2016 0 2128 800 0 FreeSans 448 90 0 0 pcpi_insn[16]
port 8 nsew signal input
flabel metal2 s 2688 0 2800 800 0 FreeSans 448 90 0 0 pcpi_insn[17]
port 9 nsew signal input
flabel metal2 s 3360 0 3472 800 0 FreeSans 448 90 0 0 pcpi_insn[18]
port 10 nsew signal input
flabel metal2 s 4032 0 4144 800 0 FreeSans 448 90 0 0 pcpi_insn[19]
port 11 nsew signal input
flabel metal3 s 0 40992 800 41104 0 FreeSans 448 0 0 0 pcpi_insn[1]
port 12 nsew signal input
flabel metal2 s 4704 0 4816 800 0 FreeSans 448 90 0 0 pcpi_insn[20]
port 13 nsew signal input
flabel metal2 s 5376 0 5488 800 0 FreeSans 448 90 0 0 pcpi_insn[21]
port 14 nsew signal input
flabel metal2 s 6048 0 6160 800 0 FreeSans 448 90 0 0 pcpi_insn[22]
port 15 nsew signal input
flabel metal2 s 6720 0 6832 800 0 FreeSans 448 90 0 0 pcpi_insn[23]
port 16 nsew signal input
flabel metal2 s 7392 0 7504 800 0 FreeSans 448 90 0 0 pcpi_insn[24]
port 17 nsew signal input
flabel metal3 s 0 51744 800 51856 0 FreeSans 448 0 0 0 pcpi_insn[25]
port 18 nsew signal input
flabel metal3 s 0 50400 800 50512 0 FreeSans 448 0 0 0 pcpi_insn[26]
port 19 nsew signal input
flabel metal3 s 0 49056 800 49168 0 FreeSans 448 0 0 0 pcpi_insn[27]
port 20 nsew signal input
flabel metal3 s 0 53088 800 53200 0 FreeSans 448 0 0 0 pcpi_insn[28]
port 21 nsew signal input
flabel metal3 s 0 43680 800 43792 0 FreeSans 448 0 0 0 pcpi_insn[29]
port 22 nsew signal input
flabel metal3 s 0 42336 800 42448 0 FreeSans 448 0 0 0 pcpi_insn[2]
port 23 nsew signal input
flabel metal3 s 0 49728 800 49840 0 FreeSans 448 0 0 0 pcpi_insn[30]
port 24 nsew signal input
flabel metal3 s 0 52416 800 52528 0 FreeSans 448 0 0 0 pcpi_insn[31]
port 25 nsew signal input
flabel metal3 s 0 38976 800 39088 0 FreeSans 448 0 0 0 pcpi_insn[3]
port 26 nsew signal input
flabel metal3 s 0 41664 800 41776 0 FreeSans 448 0 0 0 pcpi_insn[4]
port 27 nsew signal input
flabel metal3 s 0 40320 800 40432 0 FreeSans 448 0 0 0 pcpi_insn[5]
port 28 nsew signal input
flabel metal3 s 0 51072 800 51184 0 FreeSans 448 0 0 0 pcpi_insn[6]
port 29 nsew signal input
flabel metal2 s 8064 0 8176 800 0 FreeSans 448 90 0 0 pcpi_insn[7]
port 30 nsew signal input
flabel metal2 s 8736 0 8848 800 0 FreeSans 448 90 0 0 pcpi_insn[8]
port 31 nsew signal input
flabel metal2 s 9408 0 9520 800 0 FreeSans 448 90 0 0 pcpi_insn[9]
port 32 nsew signal input
flabel metal3 s 0 48384 800 48496 0 FreeSans 448 0 0 0 pcpi_mul_rd[0]
port 33 nsew signal tristate
flabel metal3 s 59200 46368 60000 46480 0 FreeSans 448 0 0 0 pcpi_mul_rd[10]
port 34 nsew signal tristate
flabel metal3 s 59200 30240 60000 30352 0 FreeSans 448 0 0 0 pcpi_mul_rd[11]
port 35 nsew signal tristate
flabel metal3 s 59200 31584 60000 31696 0 FreeSans 448 0 0 0 pcpi_mul_rd[12]
port 36 nsew signal tristate
flabel metal3 s 59200 32256 60000 32368 0 FreeSans 448 0 0 0 pcpi_mul_rd[13]
port 37 nsew signal tristate
flabel metal3 s 59200 37632 60000 37744 0 FreeSans 448 0 0 0 pcpi_mul_rd[14]
port 38 nsew signal tristate
flabel metal3 s 59200 36288 60000 36400 0 FreeSans 448 0 0 0 pcpi_mul_rd[15]
port 39 nsew signal tristate
flabel metal3 s 59200 30912 60000 31024 0 FreeSans 448 0 0 0 pcpi_mul_rd[16]
port 40 nsew signal tristate
flabel metal3 s 59200 32928 60000 33040 0 FreeSans 448 0 0 0 pcpi_mul_rd[17]
port 41 nsew signal tristate
flabel metal3 s 59200 36960 60000 37072 0 FreeSans 448 0 0 0 pcpi_mul_rd[18]
port 42 nsew signal tristate
flabel metal3 s 59200 33600 60000 33712 0 FreeSans 448 0 0 0 pcpi_mul_rd[19]
port 43 nsew signal tristate
flabel metal3 s 0 47712 800 47824 0 FreeSans 448 0 0 0 pcpi_mul_rd[1]
port 44 nsew signal tristate
flabel metal3 s 59200 45696 60000 45808 0 FreeSans 448 0 0 0 pcpi_mul_rd[20]
port 45 nsew signal tristate
flabel metal3 s 59200 44352 60000 44464 0 FreeSans 448 0 0 0 pcpi_mul_rd[21]
port 46 nsew signal tristate
flabel metal3 s 59200 43680 60000 43792 0 FreeSans 448 0 0 0 pcpi_mul_rd[22]
port 47 nsew signal tristate
flabel metal3 s 59200 45024 60000 45136 0 FreeSans 448 0 0 0 pcpi_mul_rd[23]
port 48 nsew signal tristate
flabel metal3 s 59200 39648 60000 39760 0 FreeSans 448 0 0 0 pcpi_mul_rd[24]
port 49 nsew signal tristate
flabel metal3 s 59200 43008 60000 43120 0 FreeSans 448 0 0 0 pcpi_mul_rd[25]
port 50 nsew signal tristate
flabel metal3 s 59200 40992 60000 41104 0 FreeSans 448 0 0 0 pcpi_mul_rd[26]
port 51 nsew signal tristate
flabel metal3 s 59200 40320 60000 40432 0 FreeSans 448 0 0 0 pcpi_mul_rd[27]
port 52 nsew signal tristate
flabel metal3 s 59200 38304 60000 38416 0 FreeSans 448 0 0 0 pcpi_mul_rd[28]
port 53 nsew signal tristate
flabel metal3 s 59200 42336 60000 42448 0 FreeSans 448 0 0 0 pcpi_mul_rd[29]
port 54 nsew signal tristate
flabel metal3 s 0 47040 800 47152 0 FreeSans 448 0 0 0 pcpi_mul_rd[2]
port 55 nsew signal tristate
flabel metal3 s 59200 41664 60000 41776 0 FreeSans 448 0 0 0 pcpi_mul_rd[30]
port 56 nsew signal tristate
flabel metal3 s 0 36288 800 36400 0 FreeSans 448 0 0 0 pcpi_mul_rd[31]
port 57 nsew signal tristate
flabel metal3 s 0 43008 800 43120 0 FreeSans 448 0 0 0 pcpi_mul_rd[3]
port 58 nsew signal tristate
flabel metal3 s 0 31584 800 31696 0 FreeSans 448 0 0 0 pcpi_mul_rd[4]
port 59 nsew signal tristate
flabel metal3 s 0 33600 800 33712 0 FreeSans 448 0 0 0 pcpi_mul_rd[5]
port 60 nsew signal tristate
flabel metal2 s 26208 0 26320 800 0 FreeSans 448 90 0 0 pcpi_mul_rd[6]
port 61 nsew signal tristate
flabel metal2 s 26880 0 26992 800 0 FreeSans 448 90 0 0 pcpi_mul_rd[7]
port 62 nsew signal tristate
flabel metal3 s 59200 38976 60000 39088 0 FreeSans 448 0 0 0 pcpi_mul_rd[8]
port 63 nsew signal tristate
flabel metal3 s 59200 35616 60000 35728 0 FreeSans 448 0 0 0 pcpi_mul_rd[9]
port 64 nsew signal tristate
flabel metal3 s 59200 34944 60000 35056 0 FreeSans 448 0 0 0 pcpi_mul_ready
port 65 nsew signal tristate
flabel metal3 s 0 34272 800 34384 0 FreeSans 448 0 0 0 pcpi_mul_valid
port 66 nsew signal input
flabel metal3 s 0 38304 800 38416 0 FreeSans 448 0 0 0 pcpi_mul_wait
port 67 nsew signal tristate
flabel metal3 s 59200 34272 60000 34384 0 FreeSans 448 0 0 0 pcpi_mul_wr
port 68 nsew signal tristate
flabel metal2 s 24192 0 24304 800 0 FreeSans 448 90 0 0 pcpi_rs1[0]
port 69 nsew signal input
flabel metal2 s 12768 0 12880 800 0 FreeSans 448 90 0 0 pcpi_rs1[10]
port 70 nsew signal input
flabel metal3 s 0 16128 800 16240 0 FreeSans 448 0 0 0 pcpi_rs1[11]
port 71 nsew signal input
flabel metal3 s 0 16800 800 16912 0 FreeSans 448 0 0 0 pcpi_rs1[12]
port 72 nsew signal input
flabel metal3 s 0 17472 800 17584 0 FreeSans 448 0 0 0 pcpi_rs1[13]
port 73 nsew signal input
flabel metal3 s 0 18144 800 18256 0 FreeSans 448 0 0 0 pcpi_rs1[14]
port 74 nsew signal input
flabel metal3 s 0 19488 800 19600 0 FreeSans 448 0 0 0 pcpi_rs1[15]
port 75 nsew signal input
flabel metal3 s 0 22176 800 22288 0 FreeSans 448 0 0 0 pcpi_rs1[16]
port 76 nsew signal input
flabel metal3 s 0 22848 800 22960 0 FreeSans 448 0 0 0 pcpi_rs1[17]
port 77 nsew signal input
flabel metal3 s 0 23520 800 23632 0 FreeSans 448 0 0 0 pcpi_rs1[18]
port 78 nsew signal input
flabel metal3 s 0 24192 800 24304 0 FreeSans 448 0 0 0 pcpi_rs1[19]
port 79 nsew signal input
flabel metal2 s 20160 0 20272 800 0 FreeSans 448 90 0 0 pcpi_rs1[1]
port 80 nsew signal input
flabel metal3 s 0 24864 800 24976 0 FreeSans 448 0 0 0 pcpi_rs1[20]
port 81 nsew signal input
flabel metal3 s 0 26208 800 26320 0 FreeSans 448 0 0 0 pcpi_rs1[21]
port 82 nsew signal input
flabel metal3 s 0 27552 800 27664 0 FreeSans 448 0 0 0 pcpi_rs1[22]
port 83 nsew signal input
flabel metal3 s 0 29568 800 29680 0 FreeSans 448 0 0 0 pcpi_rs1[23]
port 84 nsew signal input
flabel metal3 s 0 30240 800 30352 0 FreeSans 448 0 0 0 pcpi_rs1[24]
port 85 nsew signal input
flabel metal3 s 0 32256 800 32368 0 FreeSans 448 0 0 0 pcpi_rs1[25]
port 86 nsew signal input
flabel metal3 s 0 32928 800 33040 0 FreeSans 448 0 0 0 pcpi_rs1[26]
port 87 nsew signal input
flabel metal3 s 0 35616 800 35728 0 FreeSans 448 0 0 0 pcpi_rs1[27]
port 88 nsew signal input
flabel metal3 s 0 36960 800 37072 0 FreeSans 448 0 0 0 pcpi_rs1[28]
port 89 nsew signal input
flabel metal3 s 0 37632 800 37744 0 FreeSans 448 0 0 0 pcpi_rs1[29]
port 90 nsew signal input
flabel metal2 s 19488 0 19600 800 0 FreeSans 448 90 0 0 pcpi_rs1[2]
port 91 nsew signal input
flabel metal3 s 0 34944 800 35056 0 FreeSans 448 0 0 0 pcpi_rs1[30]
port 92 nsew signal input
flabel metal3 s 0 45024 800 45136 0 FreeSans 448 0 0 0 pcpi_rs1[31]
port 93 nsew signal input
flabel metal2 s 18816 0 18928 800 0 FreeSans 448 90 0 0 pcpi_rs1[3]
port 94 nsew signal input
flabel metal2 s 18144 0 18256 800 0 FreeSans 448 90 0 0 pcpi_rs1[4]
port 95 nsew signal input
flabel metal2 s 16800 0 16912 800 0 FreeSans 448 90 0 0 pcpi_rs1[5]
port 96 nsew signal input
flabel metal2 s 16128 0 16240 800 0 FreeSans 448 90 0 0 pcpi_rs1[6]
port 97 nsew signal input
flabel metal3 s 0 20832 800 20944 0 FreeSans 448 0 0 0 pcpi_rs1[7]
port 98 nsew signal input
flabel metal3 s 0 21504 800 21616 0 FreeSans 448 0 0 0 pcpi_rs1[8]
port 99 nsew signal input
flabel metal3 s 0 20160 800 20272 0 FreeSans 448 0 0 0 pcpi_rs1[9]
port 100 nsew signal input
flabel metal3 s 0 28896 800 29008 0 FreeSans 448 0 0 0 pcpi_rs2[0]
port 101 nsew signal input
flabel metal2 s 30912 0 31024 800 0 FreeSans 448 90 0 0 pcpi_rs2[10]
port 102 nsew signal input
flabel metal2 s 32928 0 33040 800 0 FreeSans 448 90 0 0 pcpi_rs2[11]
port 103 nsew signal input
flabel metal2 s 34272 0 34384 800 0 FreeSans 448 90 0 0 pcpi_rs2[12]
port 104 nsew signal input
flabel metal2 s 36288 0 36400 800 0 FreeSans 448 90 0 0 pcpi_rs2[13]
port 105 nsew signal input
flabel metal2 s 38304 0 38416 800 0 FreeSans 448 90 0 0 pcpi_rs2[14]
port 106 nsew signal input
flabel metal2 s 39648 0 39760 800 0 FreeSans 448 90 0 0 pcpi_rs2[15]
port 107 nsew signal input
flabel metal2 s 40992 0 41104 800 0 FreeSans 448 90 0 0 pcpi_rs2[16]
port 108 nsew signal input
flabel metal2 s 42336 0 42448 800 0 FreeSans 448 90 0 0 pcpi_rs2[17]
port 109 nsew signal input
flabel metal2 s 43008 0 43120 800 0 FreeSans 448 90 0 0 pcpi_rs2[18]
port 110 nsew signal input
flabel metal2 s 43680 0 43792 800 0 FreeSans 448 90 0 0 pcpi_rs2[19]
port 111 nsew signal input
flabel metal3 s 0 28224 800 28336 0 FreeSans 448 0 0 0 pcpi_rs2[1]
port 112 nsew signal input
flabel metal3 s 59200 21504 60000 21616 0 FreeSans 448 0 0 0 pcpi_rs2[20]
port 113 nsew signal input
flabel metal3 s 59200 23520 60000 23632 0 FreeSans 448 0 0 0 pcpi_rs2[21]
port 114 nsew signal input
flabel metal3 s 59200 24192 60000 24304 0 FreeSans 448 0 0 0 pcpi_rs2[22]
port 115 nsew signal input
flabel metal3 s 59200 24864 60000 24976 0 FreeSans 448 0 0 0 pcpi_rs2[23]
port 116 nsew signal input
flabel metal2 s 40320 0 40432 800 0 FreeSans 448 90 0 0 pcpi_rs2[24]
port 117 nsew signal input
flabel metal2 s 37632 0 37744 800 0 FreeSans 448 90 0 0 pcpi_rs2[25]
port 118 nsew signal input
flabel metal2 s 36960 0 37072 800 0 FreeSans 448 90 0 0 pcpi_rs2[26]
port 119 nsew signal input
flabel metal2 s 35616 0 35728 800 0 FreeSans 448 90 0 0 pcpi_rs2[27]
port 120 nsew signal input
flabel metal2 s 33600 0 33712 800 0 FreeSans 448 90 0 0 pcpi_rs2[28]
port 121 nsew signal input
flabel metal2 s 30240 0 30352 800 0 FreeSans 448 90 0 0 pcpi_rs2[29]
port 122 nsew signal input
flabel metal3 s 0 26880 800 26992 0 FreeSans 448 0 0 0 pcpi_rs2[2]
port 123 nsew signal input
flabel metal2 s 28896 0 29008 800 0 FreeSans 448 90 0 0 pcpi_rs2[30]
port 124 nsew signal input
flabel metal3 s 0 44352 800 44464 0 FreeSans 448 0 0 0 pcpi_rs2[31]
port 125 nsew signal input
flabel metal3 s 0 25536 800 25648 0 FreeSans 448 0 0 0 pcpi_rs2[3]
port 126 nsew signal input
flabel metal2 s 20832 0 20944 800 0 FreeSans 448 90 0 0 pcpi_rs2[4]
port 127 nsew signal input
flabel metal2 s 22848 0 22960 800 0 FreeSans 448 90 0 0 pcpi_rs2[5]
port 128 nsew signal input
flabel metal2 s 23520 0 23632 800 0 FreeSans 448 90 0 0 pcpi_rs2[6]
port 129 nsew signal input
flabel metal2 s 25536 0 25648 800 0 FreeSans 448 90 0 0 pcpi_rs2[7]
port 130 nsew signal input
flabel metal2 s 27552 0 27664 800 0 FreeSans 448 90 0 0 pcpi_rs2[8]
port 131 nsew signal input
flabel metal2 s 29568 0 29680 800 0 FreeSans 448 90 0 0 pcpi_rs2[9]
port 132 nsew signal input
flabel metal3 s 0 39648 800 39760 0 FreeSans 448 0 0 0 resetn
port 133 nsew signal input
flabel metal4 s 4448 3076 4768 76892 0 FreeSans 1280 90 0 0 vdd
port 134 nsew power bidirectional
flabel metal4 s 35168 3076 35488 76892 0 FreeSans 1280 90 0 0 vdd
port 134 nsew power bidirectional
flabel metal4 s 19808 3076 20128 76892 0 FreeSans 1280 90 0 0 vss
port 135 nsew ground bidirectional
flabel metal4 s 50528 3076 50848 76892 0 FreeSans 1280 90 0 0 vss
port 135 nsew ground bidirectional
rlabel metal1 29960 76048 29960 76048 0 vdd
rlabel metal1 29960 76832 29960 76832 0 vss
rlabel metal3 30352 36456 30352 36456 0 _0000_
rlabel metal2 14448 43624 14448 43624 0 _0001_
rlabel metal2 13328 42056 13328 42056 0 _0002_
rlabel metal2 19656 36792 19656 36792 0 _0003_
rlabel metal2 22120 39704 22120 39704 0 _0004_
rlabel metal2 12936 44744 12936 44744 0 _0005_
rlabel metal2 18872 31920 18872 31920 0 _0006_
rlabel metal3 15540 29288 15540 29288 0 _0007_
rlabel metal2 14896 31080 14896 31080 0 _0008_
rlabel metal2 14616 34160 14616 34160 0 _0009_
rlabel metal2 15400 38416 15400 38416 0 _0010_
rlabel metal2 14616 44968 14616 44968 0 _0011_
rlabel metal2 18312 29344 18312 29344 0 _0012_
rlabel metal3 16632 26936 16632 26936 0 _0013_
rlabel metal2 18200 23856 18200 23856 0 _0014_
rlabel metal2 19320 14056 19320 14056 0 _0015_
rlabel metal2 22904 9856 22904 9856 0 _0016_
rlabel metal2 24472 9464 24472 9464 0 _0017_
rlabel metal2 26488 9072 26488 9072 0 _0018_
rlabel metal2 28056 9408 28056 9408 0 _0019_
rlabel metal2 30856 9632 30856 9632 0 _0020_
rlabel metal2 31528 9352 31528 9352 0 _0021_
rlabel metal2 33936 8456 33936 8456 0 _0022_
rlabel metal2 34328 12096 34328 12096 0 _0023_
rlabel metal3 37128 8120 37128 8120 0 _0024_
rlabel metal2 39592 8176 39592 8176 0 _0025_
rlabel metal2 40208 9240 40208 9240 0 _0026_
rlabel metal2 42280 11816 42280 11816 0 _0027_
rlabel metal2 42280 7728 42280 7728 0 _0028_
rlabel metal2 45752 8372 45752 8372 0 _0029_
rlabel metal2 45640 9464 45640 9464 0 _0030_
rlabel metal2 44072 21896 44072 21896 0 _0031_
rlabel metal2 43624 22960 43624 22960 0 _0032_
rlabel metal3 45304 26824 45304 26824 0 _0033_
rlabel metal2 43512 24752 43512 24752 0 _0034_
rlabel metal3 42616 23800 42616 23800 0 _0035_
rlabel metal2 38360 22008 38360 22008 0 _0036_
rlabel metal2 37800 25816 37800 25816 0 _0037_
rlabel metal3 36232 22456 36232 22456 0 _0038_
rlabel metal3 33040 24024 33040 24024 0 _0039_
rlabel metal2 31080 22400 31080 22400 0 _0040_
rlabel metal2 29288 24360 29288 24360 0 _0041_
rlabel metal2 21448 44856 21448 44856 0 _0042_
rlabel metal2 20328 55552 20328 55552 0 _0043_
rlabel metal2 20552 52584 20552 52584 0 _0044_
rlabel metal2 18872 61152 18872 61152 0 _0045_
rlabel metal2 19320 64344 19320 64344 0 _0046_
rlabel metal2 20776 65800 20776 65800 0 _0047_
rlabel metal2 21448 68264 21448 68264 0 _0048_
rlabel metal2 22904 69720 22904 69720 0 _0049_
rlabel metal2 26152 69720 26152 69720 0 _0050_
rlabel metal2 30352 67928 30352 67928 0 _0051_
rlabel metal2 29008 67928 29008 67928 0 _0052_
rlabel metal2 32368 70392 32368 70392 0 _0053_
rlabel metal2 33992 70504 33992 70504 0 _0054_
rlabel metal3 36848 69608 36848 69608 0 _0055_
rlabel metal2 39144 71904 39144 71904 0 _0056_
rlabel metal2 41720 70896 41720 70896 0 _0057_
rlabel metal3 39928 69272 39928 69272 0 _0058_
rlabel metal2 45416 65912 45416 65912 0 _0059_
rlabel metal2 46984 68544 46984 68544 0 _0060_
rlabel metal2 43568 67928 43568 67928 0 _0061_
rlabel metal2 43848 64232 43848 64232 0 _0062_
rlabel metal2 45976 55608 45976 55608 0 _0063_
rlabel metal2 44968 54152 44968 54152 0 _0064_
rlabel metal2 41720 54656 41720 54656 0 _0065_
rlabel metal2 43344 51464 43344 51464 0 _0066_
rlabel metal2 33992 51632 33992 51632 0 _0067_
rlabel metal2 37576 55608 37576 55608 0 _0068_
rlabel metal2 37800 56000 37800 56000 0 _0069_
rlabel metal2 33656 53704 33656 53704 0 _0070_
rlabel metal2 29960 51016 29960 51016 0 _0071_
rlabel metal2 28504 51800 28504 51800 0 _0072_
rlabel metal2 26040 51912 26040 51912 0 _0073_
rlabel metal2 24360 49336 24360 49336 0 _0074_
rlabel metal2 14392 47824 14392 47824 0 _0075_
rlabel metal2 15848 28280 15848 28280 0 _0076_
rlabel metal2 20888 31528 20888 31528 0 _0077_
rlabel metal2 19880 32704 19880 32704 0 _0078_
rlabel metal3 21168 27720 21168 27720 0 _0079_
rlabel metal3 23184 26824 23184 26824 0 _0080_
rlabel metal2 22120 18368 22120 18368 0 _0081_
rlabel metal2 22568 14056 22568 14056 0 _0082_
rlabel metal2 26376 15736 26376 15736 0 _0083_
rlabel metal2 25648 19208 25648 19208 0 _0084_
rlabel metal2 29736 18480 29736 18480 0 _0085_
rlabel metal3 32368 15176 32368 15176 0 _0086_
rlabel metal2 34104 15148 34104 15148 0 _0087_
rlabel metal3 33320 18424 33320 18424 0 _0088_
rlabel metal2 37800 17920 37800 17920 0 _0089_
rlabel metal2 37968 13048 37968 13048 0 _0090_
rlabel metal3 41440 15960 41440 15960 0 _0091_
rlabel metal3 40544 18312 40544 18312 0 _0092_
rlabel metal2 43848 15344 43848 15344 0 _0093_
rlabel metal2 48664 11760 48664 11760 0 _0094_
rlabel metal2 48608 13048 48608 13048 0 _0095_
rlabel metal2 50904 17640 50904 17640 0 _0096_
rlabel metal2 47880 22512 47880 22512 0 _0097_
rlabel metal2 49784 26712 49784 26712 0 _0098_
rlabel metal2 48888 30968 48888 30968 0 _0099_
rlabel metal2 45528 31920 45528 31920 0 _0100_
rlabel metal2 38472 26908 38472 26908 0 _0101_
rlabel metal2 42168 31416 42168 31416 0 _0102_
rlabel metal2 38248 32144 38248 32144 0 _0103_
rlabel metal2 36008 33712 36008 33712 0 _0104_
rlabel metal2 33936 27160 33936 27160 0 _0105_
rlabel metal2 30016 27160 30016 27160 0 _0106_
rlabel metal2 27720 29288 27720 29288 0 _0107_
rlabel metal2 29176 32648 29176 32648 0 _0108_
rlabel metal3 24416 53816 24416 53816 0 _0109_
rlabel metal2 20440 49336 20440 49336 0 _0110_
rlabel metal2 18424 57960 18424 57960 0 _0111_
rlabel metal3 28000 60648 28000 60648 0 _0112_
rlabel metal2 22792 58072 22792 58072 0 _0113_
rlabel metal2 22176 61656 22176 61656 0 _0114_
rlabel metal2 24024 64792 24024 64792 0 _0115_
rlabel metal2 27384 65800 27384 65800 0 _0116_
rlabel metal2 32872 60368 32872 60368 0 _0117_
rlabel metal3 29008 62328 29008 62328 0 _0118_
rlabel metal2 32088 64792 32088 64792 0 _0119_
rlabel metal2 36008 63504 36008 63504 0 _0120_
rlabel metal3 37744 60648 37744 60648 0 _0121_
rlabel metal2 41496 57568 41496 57568 0 _0122_
rlabel metal2 42616 62776 42616 62776 0 _0123_
rlabel metal2 38248 64176 38248 64176 0 _0124_
rlabel metal2 47768 62972 47768 62972 0 _0125_
rlabel metal2 47656 56784 47656 56784 0 _0126_
rlabel metal2 45192 60256 45192 60256 0 _0127_
rlabel metal2 48552 46256 48552 46256 0 _0128_
rlabel metal2 50904 54824 50904 54824 0 _0129_
rlabel metal2 49224 50904 49224 50904 0 _0130_
rlabel metal2 46088 48552 46088 48552 0 _0131_
rlabel metal2 44296 44324 44296 44324 0 _0132_
rlabel metal2 35280 47208 35280 47208 0 _0133_
rlabel metal2 39256 50848 39256 50848 0 _0134_
rlabel metal2 38528 45304 38528 45304 0 _0135_
rlabel metal2 35672 45864 35672 45864 0 _0136_
rlabel metal2 32648 48216 32648 48216 0 _0137_
rlabel metal2 26824 43064 26824 43064 0 _0138_
rlabel metal2 25592 46928 25592 46928 0 _0139_
rlabel metal2 26264 37688 26264 37688 0 _0140_
rlabel metal2 22568 20384 22568 20384 0 _0141_
rlabel metal2 28168 21168 28168 21168 0 _0142_
rlabel metal2 36120 20216 36120 20216 0 _0143_
rlabel metal2 42952 18480 42952 18480 0 _0144_
rlabel metal2 47992 19740 47992 19740 0 _0145_
rlabel metal2 44352 27944 44352 27944 0 _0146_
rlabel metal3 34664 31080 34664 31080 0 _0147_
rlabel metal2 28056 55664 28056 55664 0 _0148_
rlabel metal2 26488 57568 26488 57568 0 _0149_
rlabel metal2 30072 58800 30072 58800 0 _0150_
rlabel metal2 35616 59304 35616 59304 0 _0151_
rlabel metal2 46088 62188 46088 62188 0 _0152_
rlabel metal3 47208 48888 47208 48888 0 _0153_
rlabel metal2 41720 45864 41720 45864 0 _0154_
rlabel metal2 31360 44408 31360 44408 0 _0155_
rlabel metal2 18648 40712 18648 40712 0 _0156_
rlabel metal3 25032 23800 25032 23800 0 _0157_
rlabel metal2 20272 21000 20272 21000 0 _0158_
rlabel metal2 17864 20832 17864 20832 0 _0159_
rlabel metal3 19096 16184 19096 16184 0 _0160_
rlabel metal2 18424 16688 18424 16688 0 _0161_
rlabel metal2 16744 15736 16744 15736 0 _0162_
rlabel metal2 14728 17584 14728 17584 0 _0163_
rlabel metal2 16968 22680 16968 22680 0 _0164_
rlabel metal2 14280 21896 14280 21896 0 _0165_
rlabel metal2 11032 21896 11032 21896 0 _0166_
rlabel metal2 13384 17696 13384 17696 0 _0167_
rlabel metal2 13720 15624 13720 15624 0 _0168_
rlabel metal2 10584 17192 10584 17192 0 _0169_
rlabel metal2 9072 16184 9072 16184 0 _0170_
rlabel metal2 7896 17976 7896 17976 0 _0171_
rlabel metal2 6888 19656 6888 19656 0 _0172_
rlabel metal2 6888 21112 6888 21112 0 _0173_
rlabel metal2 7000 22792 7000 22792 0 _0174_
rlabel metal3 7560 24584 7560 24584 0 _0175_
rlabel metal2 7224 25816 7224 25816 0 _0176_
rlabel metal3 11704 24024 11704 24024 0 _0177_
rlabel metal3 13160 25704 13160 25704 0 _0178_
rlabel metal2 11816 28280 11816 28280 0 _0179_
rlabel metal2 9128 27384 9128 27384 0 _0180_
rlabel metal2 8904 29848 8904 29848 0 _0181_
rlabel metal2 8680 32088 8680 32088 0 _0182_
rlabel metal2 9800 32760 9800 32760 0 _0183_
rlabel metal2 9128 35224 9128 35224 0 _0184_
rlabel metal2 9240 36792 9240 36792 0 _0185_
rlabel metal3 10248 38696 10248 38696 0 _0186_
rlabel metal2 11928 39144 11928 39144 0 _0187_
rlabel metal2 18424 47600 18424 47600 0 _0188_
rlabel metal2 15400 49168 15400 49168 0 _0189_
rlabel metal2 15288 52696 15288 52696 0 _0190_
rlabel metal2 13720 52696 13720 52696 0 _0191_
rlabel metal2 15624 55412 15624 55412 0 _0192_
rlabel metal2 13048 57344 13048 57344 0 _0193_
rlabel metal2 15736 57736 15736 57736 0 _0194_
rlabel metal2 14728 59528 14728 59528 0 _0195_
rlabel metal3 15512 62216 15512 62216 0 _0196_
rlabel metal3 15848 64120 15848 64120 0 _0197_
rlabel metal3 16520 65464 16520 65464 0 _0198_
rlabel metal2 13888 64792 13888 64792 0 _0199_
rlabel metal3 11536 63784 11536 63784 0 _0200_
rlabel metal2 11704 64344 11704 64344 0 _0201_
rlabel metal2 10472 62216 10472 62216 0 _0202_
rlabel metal2 10360 61096 10360 61096 0 _0203_
rlabel metal2 10696 58464 10696 58464 0 _0204_
rlabel metal2 10416 53816 10416 53816 0 _0205_
rlabel metal3 11088 55160 11088 55160 0 _0206_
rlabel metal3 7952 56952 7952 56952 0 _0207_
rlabel metal2 7224 56224 7224 56224 0 _0208_
rlabel metal2 6608 54376 6608 54376 0 _0209_
rlabel metal2 5320 53424 5320 53424 0 _0210_
rlabel metal2 5320 51856 5320 51856 0 _0211_
rlabel metal3 6776 48440 6776 48440 0 _0212_
rlabel metal3 6720 46536 6720 46536 0 _0213_
rlabel metal2 5992 45584 5992 45584 0 _0214_
rlabel metal2 6608 44408 6608 44408 0 _0215_
rlabel metal2 11704 45248 11704 45248 0 _0216_
rlabel metal2 11648 46760 11648 46760 0 _0217_
rlabel metal2 13608 49392 13608 49392 0 _0218_
rlabel metal2 10584 50680 10584 50680 0 _0219_
rlabel metal2 23688 46256 23688 46256 0 _0220_
rlabel metal2 22456 46256 22456 46256 0 _0221_
rlabel metal2 21616 43624 21616 43624 0 _0222_
rlabel metal2 22344 42448 22344 42448 0 _0223_
rlabel metal2 25424 33432 25424 33432 0 _0224_
rlabel metal2 24360 34552 24360 34552 0 _0225_
rlabel metal2 25928 31024 25928 31024 0 _0226_
rlabel metal2 24696 29008 24696 29008 0 _0227_
rlabel metal2 34048 39704 34048 39704 0 _0228_
rlabel metal2 33544 36120 33544 36120 0 _0229_
rlabel metal2 35056 37352 35056 37352 0 _0230_
rlabel metal2 36008 36008 36008 36008 0 _0231_
rlabel metal2 38248 36512 38248 36512 0 _0232_
rlabel metal2 42280 34272 42280 34272 0 _0233_
rlabel metal2 42560 37352 42560 37352 0 _0234_
rlabel metal2 42504 34552 42504 34552 0 _0235_
rlabel metal2 46536 36512 46536 36512 0 _0236_
rlabel metal2 49560 35840 49560 35840 0 _0237_
rlabel metal2 47208 35000 47208 35000 0 _0238_
rlabel metal3 48776 34216 48776 34216 0 _0239_
rlabel metal2 49336 39256 49336 39256 0 _0240_
rlabel metal2 49504 40488 49504 40488 0 _0241_
rlabel metal2 49560 43120 49560 43120 0 _0242_
rlabel metal2 46200 39592 46200 39592 0 _0243_
rlabel metal2 39816 39648 39816 39648 0 _0244_
rlabel metal2 41608 40040 41608 40040 0 _0245_
rlabel metal2 41832 41384 41832 41384 0 _0246_
rlabel metal2 37912 39984 37912 39984 0 _0247_
rlabel metal2 31472 38136 31472 38136 0 _0248_
rlabel metal2 31304 40376 31304 40376 0 _0249_
rlabel metal3 29512 38920 29512 38920 0 _0250_
rlabel metal2 29232 37352 29232 37352 0 _0251_
rlabel metal2 14280 37576 14280 37576 0 _0252_
rlabel metal3 24416 24024 24416 24024 0 _0253_
rlabel metal3 23912 27048 23912 27048 0 _0254_
rlabel metal2 23968 26152 23968 26152 0 _0255_
rlabel metal2 24696 25984 24696 25984 0 _0256_
rlabel metal2 24360 25256 24360 25256 0 _0257_
rlabel metal2 20720 25704 20720 25704 0 _0258_
rlabel metal2 24696 18648 24696 18648 0 _0259_
rlabel metal3 23464 18312 23464 18312 0 _0260_
rlabel metal2 22456 18704 22456 18704 0 _0261_
rlabel metal2 26376 22064 26376 22064 0 _0262_
rlabel metal3 24640 17752 24640 17752 0 _0263_
rlabel metal3 23016 19096 23016 19096 0 _0264_
rlabel metal2 22344 19488 22344 19488 0 _0265_
rlabel metal2 25368 21840 25368 21840 0 _0266_
rlabel metal3 23856 18424 23856 18424 0 _0267_
rlabel metal2 23912 16352 23912 16352 0 _0268_
rlabel metal3 23352 15512 23352 15512 0 _0269_
rlabel metal2 24584 16352 24584 16352 0 _0270_
rlabel metal3 24808 14392 24808 14392 0 _0271_
rlabel metal2 26600 12992 26600 12992 0 _0272_
rlabel metal2 26264 13104 26264 13104 0 _0273_
rlabel metal2 25256 14168 25256 14168 0 _0274_
rlabel metal2 24360 14784 24360 14784 0 _0275_
rlabel metal2 24192 14504 24192 14504 0 _0276_
rlabel metal3 25088 16632 25088 16632 0 _0277_
rlabel metal2 25816 12096 25816 12096 0 _0278_
rlabel metal2 25648 12040 25648 12040 0 _0279_
rlabel metal2 26320 14504 26320 14504 0 _0280_
rlabel metal2 26488 16464 26488 16464 0 _0281_
rlabel metal3 35112 21560 35112 21560 0 _0282_
rlabel metal2 27720 15568 27720 15568 0 _0283_
rlabel metal2 26824 16128 26824 16128 0 _0284_
rlabel metal2 26264 15624 26264 15624 0 _0285_
rlabel metal2 46760 26488 46760 26488 0 _0286_
rlabel metal3 32536 15848 32536 15848 0 _0287_
rlabel metal2 26544 15512 26544 15512 0 _0288_
rlabel metal2 25704 15288 25704 15288 0 _0289_
rlabel metal2 34216 17696 34216 17696 0 _0290_
rlabel metal2 27496 16968 27496 16968 0 _0291_
rlabel metal2 26264 18760 26264 18760 0 _0292_
rlabel metal2 26824 20888 26824 20888 0 _0293_
rlabel metal2 26936 22792 26936 22792 0 _0294_
rlabel metal2 27160 19432 27160 19432 0 _0295_
rlabel metal3 26208 19096 26208 19096 0 _0296_
rlabel metal3 25928 18984 25928 18984 0 _0297_
rlabel metal2 25144 20384 25144 20384 0 _0298_
rlabel metal2 31528 19264 31528 19264 0 _0299_
rlabel metal3 30408 17752 30408 17752 0 _0300_
rlabel metal3 30072 18984 30072 18984 0 _0301_
rlabel metal2 47992 21784 47992 21784 0 _0302_
rlabel metal2 31640 18872 31640 18872 0 _0303_
rlabel metal2 30296 19600 30296 19600 0 _0304_
rlabel metal2 47208 30632 47208 30632 0 _0305_
rlabel metal2 32872 17584 32872 17584 0 _0306_
rlabel metal2 31080 19208 31080 19208 0 _0307_
rlabel metal2 30968 15960 30968 15960 0 _0308_
rlabel metal2 30352 15288 30352 15288 0 _0309_
rlabel metal2 31864 15960 31864 15960 0 _0310_
rlabel metal2 31304 14728 31304 14728 0 _0311_
rlabel metal2 31080 12712 31080 12712 0 _0312_
rlabel metal3 31024 14392 31024 14392 0 _0313_
rlabel metal3 31360 15512 31360 15512 0 _0314_
rlabel metal3 31976 15400 31976 15400 0 _0315_
rlabel metal2 33544 15344 33544 15344 0 _0316_
rlabel metal2 32424 13328 32424 13328 0 _0317_
rlabel metal2 32256 13496 32256 13496 0 _0318_
rlabel metal2 33376 15288 33376 15288 0 _0319_
rlabel metal2 45976 14056 45976 14056 0 _0320_
rlabel metal2 34720 13720 34720 13720 0 _0321_
rlabel metal2 33600 13608 33600 13608 0 _0322_
rlabel metal2 33768 13552 33768 13552 0 _0323_
rlabel metal3 34664 15288 34664 15288 0 _0324_
rlabel metal2 34664 15568 34664 15568 0 _0325_
rlabel metal2 36680 14728 36680 14728 0 _0326_
rlabel metal2 35784 17920 35784 17920 0 _0327_
rlabel metal3 45472 28056 45472 28056 0 _0328_
rlabel metal3 35056 19432 35056 19432 0 _0329_
rlabel metal2 35000 48104 35000 48104 0 _0330_
rlabel metal2 47432 17192 47432 17192 0 _0331_
rlabel metal2 34832 17752 34832 17752 0 _0332_
rlabel metal2 34216 20160 34216 20160 0 _0333_
rlabel metal2 34496 18424 34496 18424 0 _0334_
rlabel metal2 39648 13720 39648 13720 0 _0335_
rlabel metal2 33656 18872 33656 18872 0 _0336_
rlabel metal2 34104 18200 34104 18200 0 _0337_
rlabel metal2 45360 20888 45360 20888 0 _0338_
rlabel metal2 39592 32536 39592 32536 0 _0339_
rlabel metal2 36456 17472 36456 17472 0 _0340_
rlabel metal2 36008 17808 36008 17808 0 _0341_
rlabel metal2 36400 16968 36400 16968 0 _0342_
rlabel metal2 36568 16744 36568 16744 0 _0343_
rlabel metal3 42056 15064 42056 15064 0 _0344_
rlabel metal2 38920 17528 38920 17528 0 _0345_
rlabel metal2 38696 16464 38696 16464 0 _0346_
rlabel metal3 37128 15288 37128 15288 0 _0347_
rlabel metal2 37688 15568 37688 15568 0 _0348_
rlabel metal2 38136 14784 38136 14784 0 _0349_
rlabel metal2 37464 12824 37464 12824 0 _0350_
rlabel metal2 38696 12880 38696 12880 0 _0351_
rlabel metal3 38752 13720 38752 13720 0 _0352_
rlabel metal2 38248 14112 38248 14112 0 _0353_
rlabel metal2 39256 14504 39256 14504 0 _0354_
rlabel metal2 40488 12152 40488 12152 0 _0355_
rlabel metal2 40376 13272 40376 13272 0 _0356_
rlabel metal2 40152 14336 40152 14336 0 _0357_
rlabel metal2 41160 13272 41160 13272 0 _0358_
rlabel metal2 40432 13944 40432 13944 0 _0359_
rlabel metal2 40376 16184 40376 16184 0 _0360_
rlabel metal2 40264 14112 40264 14112 0 _0361_
rlabel metal2 42280 16856 42280 16856 0 _0362_
rlabel metal2 40824 17192 40824 17192 0 _0363_
rlabel metal2 41048 15568 41048 15568 0 _0364_
rlabel metal2 40152 18704 40152 18704 0 _0365_
rlabel metal3 41944 20664 41944 20664 0 _0366_
rlabel metal3 42168 19320 42168 19320 0 _0367_
rlabel metal3 42280 20776 42280 20776 0 _0368_
rlabel metal2 41216 17864 41216 17864 0 _0369_
rlabel metal2 40264 18480 40264 18480 0 _0370_
rlabel metal2 41496 18032 41496 18032 0 _0371_
rlabel metal2 47824 16744 47824 16744 0 _0372_
rlabel metal2 44296 17304 44296 17304 0 _0373_
rlabel metal3 44296 16072 44296 16072 0 _0374_
rlabel metal2 45080 17360 45080 17360 0 _0375_
rlabel metal2 46312 17192 46312 17192 0 _0376_
rlabel metal2 44856 16464 44856 16464 0 _0377_
rlabel metal2 48104 14280 48104 14280 0 _0378_
rlabel metal2 45528 16744 45528 16744 0 _0379_
rlabel metal2 46648 15456 46648 15456 0 _0380_
rlabel metal2 44856 14560 44856 14560 0 _0381_
rlabel metal3 45864 15176 45864 15176 0 _0382_
rlabel metal2 47264 15288 47264 15288 0 _0383_
rlabel metal2 46760 14448 46760 14448 0 _0384_
rlabel metal2 44632 12712 44632 12712 0 _0385_
rlabel metal2 47096 13664 47096 13664 0 _0386_
rlabel metal3 47488 12824 47488 12824 0 _0387_
rlabel metal3 48552 13944 48552 13944 0 _0388_
rlabel metal2 47544 13272 47544 13272 0 _0389_
rlabel metal2 48216 12656 48216 12656 0 _0390_
rlabel metal3 45808 11256 45808 11256 0 _0391_
rlabel metal2 46200 12600 46200 12600 0 _0392_
rlabel metal3 47880 13720 47880 13720 0 _0393_
rlabel metal2 46480 14504 46480 14504 0 _0394_
rlabel metal3 48328 15512 48328 15512 0 _0395_
rlabel metal2 48496 12712 48496 12712 0 _0396_
rlabel metal2 48440 13272 48440 13272 0 _0397_
rlabel metal2 49112 13608 49112 13608 0 _0398_
rlabel metal2 49336 15792 49336 15792 0 _0399_
rlabel metal2 48776 17248 48776 17248 0 _0400_
rlabel metal2 46928 18984 46928 18984 0 _0401_
rlabel metal2 46760 18480 46760 18480 0 _0402_
rlabel metal2 48104 18536 48104 18536 0 _0403_
rlabel metal2 49112 17248 49112 17248 0 _0404_
rlabel metal3 48832 17080 48832 17080 0 _0405_
rlabel metal2 48888 17248 48888 17248 0 _0406_
rlabel metal2 49896 24360 49896 24360 0 _0407_
rlabel metal2 46200 22680 46200 22680 0 _0408_
rlabel metal2 45864 22624 45864 22624 0 _0409_
rlabel metal2 45304 22848 45304 22848 0 _0410_
rlabel metal2 47544 23016 47544 23016 0 _0411_
rlabel metal2 50344 26936 50344 26936 0 _0412_
rlabel metal2 46872 23464 46872 23464 0 _0413_
rlabel metal3 50008 24696 50008 24696 0 _0414_
rlabel metal2 47544 22064 47544 22064 0 _0415_
rlabel metal2 50008 24024 50008 24024 0 _0416_
rlabel metal2 48776 25480 48776 25480 0 _0417_
rlabel metal2 47432 27104 47432 27104 0 _0418_
rlabel metal2 49000 26572 49000 26572 0 _0419_
rlabel metal2 49560 26040 49560 26040 0 _0420_
rlabel metal3 48888 26488 48888 26488 0 _0421_
rlabel metal2 50120 27160 50120 27160 0 _0422_
rlabel metal2 46872 27496 46872 27496 0 _0423_
rlabel metal3 48440 27832 48440 27832 0 _0424_
rlabel metal2 49672 28952 49672 28952 0 _0425_
rlabel metal2 47656 28616 47656 28616 0 _0426_
rlabel metal2 48440 29848 48440 29848 0 _0427_
rlabel metal3 49616 29960 49616 29960 0 _0428_
rlabel metal2 43176 30800 43176 30800 0 _0429_
rlabel metal3 48384 30184 48384 30184 0 _0430_
rlabel metal3 49952 30184 49952 30184 0 _0431_
rlabel metal2 47208 29288 47208 29288 0 _0432_
rlabel metal2 45976 30352 45976 30352 0 _0433_
rlabel metal2 46312 29344 46312 29344 0 _0434_
rlabel metal2 45976 29400 45976 29400 0 _0435_
rlabel metal2 45584 30184 45584 30184 0 _0436_
rlabel metal2 46200 31472 46200 31472 0 _0437_
rlabel metal2 45752 31248 45752 31248 0 _0438_
rlabel metal2 46816 30408 46816 30408 0 _0439_
rlabel metal2 39480 29288 39480 29288 0 _0440_
rlabel metal2 39312 27048 39312 27048 0 _0441_
rlabel metal2 38808 26544 38808 26544 0 _0442_
rlabel metal2 25816 59528 25816 59528 0 _0443_
rlabel metal2 38024 27832 38024 27832 0 _0444_
rlabel metal2 38360 27720 38360 27720 0 _0445_
rlabel metal3 31528 50344 31528 50344 0 _0446_
rlabel metal2 34776 32480 34776 32480 0 _0447_
rlabel metal2 39032 28224 39032 28224 0 _0448_
rlabel metal2 41384 28168 41384 28168 0 _0449_
rlabel metal2 40600 26180 40600 26180 0 _0450_
rlabel metal2 41832 27832 41832 27832 0 _0451_
rlabel metal2 41384 29960 41384 29960 0 _0452_
rlabel metal2 40600 29624 40600 29624 0 _0453_
rlabel metal2 42728 29624 42728 29624 0 _0454_
rlabel metal2 42392 29904 42392 29904 0 _0455_
rlabel metal2 42504 31192 42504 31192 0 _0456_
rlabel metal2 41384 30744 41384 30744 0 _0457_
rlabel metal2 43232 27272 43232 27272 0 _0458_
rlabel metal3 41944 30184 41944 30184 0 _0459_
rlabel metal3 39928 29960 39928 29960 0 _0460_
rlabel metal2 37632 30184 37632 30184 0 _0461_
rlabel metal3 38752 30968 38752 30968 0 _0462_
rlabel metal2 39088 31192 39088 31192 0 _0463_
rlabel metal3 39088 30184 39088 30184 0 _0464_
rlabel metal2 39592 31752 39592 31752 0 _0465_
rlabel metal2 38696 30128 38696 30128 0 _0466_
rlabel metal2 37576 31472 37576 31472 0 _0467_
rlabel metal3 34104 41944 34104 41944 0 _0468_
rlabel metal3 34888 33096 34888 33096 0 _0469_
rlabel metal2 27328 44072 27328 44072 0 _0470_
rlabel metal2 34440 33600 34440 33600 0 _0471_
rlabel metal3 35000 32536 35000 32536 0 _0472_
rlabel metal2 37016 32088 37016 32088 0 _0473_
rlabel metal2 33208 46480 33208 46480 0 _0474_
rlabel metal2 31192 32984 31192 32984 0 _0475_
rlabel metal2 35560 32816 35560 32816 0 _0476_
rlabel metal2 36736 33320 36736 33320 0 _0477_
rlabel metal2 32760 29120 32760 29120 0 _0478_
rlabel metal2 34888 27608 34888 27608 0 _0479_
rlabel metal2 33880 26908 33880 26908 0 _0480_
rlabel metal2 33880 28224 33880 28224 0 _0481_
rlabel metal2 34104 27944 34104 27944 0 _0482_
rlabel metal3 32592 29624 32592 29624 0 _0483_
rlabel metal2 33432 27720 33432 27720 0 _0484_
rlabel metal2 35672 29064 35672 29064 0 _0485_
rlabel metal2 34216 25312 34216 25312 0 _0486_
rlabel metal2 36120 28672 36120 28672 0 _0487_
rlabel metal3 32984 29512 32984 29512 0 _0488_
rlabel metal2 29904 27608 29904 27608 0 _0489_
rlabel metal2 31304 29904 31304 29904 0 _0490_
rlabel metal2 31192 28224 31192 28224 0 _0491_
rlabel metal2 29960 28896 29960 28896 0 _0492_
rlabel metal3 31472 28616 31472 28616 0 _0493_
rlabel metal2 32424 28112 32424 28112 0 _0494_
rlabel metal2 32256 28392 32256 28392 0 _0495_
rlabel metal3 30744 30184 30744 30184 0 _0496_
rlabel metal2 29288 29120 29288 29120 0 _0497_
rlabel metal2 29848 29904 29848 29904 0 _0498_
rlabel metal2 28168 28840 28168 28840 0 _0499_
rlabel metal2 27832 30184 27832 30184 0 _0500_
rlabel metal2 28728 30576 28728 30576 0 _0501_
rlabel metal2 29176 30856 29176 30856 0 _0502_
rlabel metal2 28392 32480 28392 32480 0 _0503_
rlabel metal2 28952 34216 28952 34216 0 _0504_
rlabel metal3 28448 34664 28448 34664 0 _0505_
rlabel metal2 28392 34160 28392 34160 0 _0506_
rlabel metal3 28280 33208 28280 33208 0 _0507_
rlabel metal3 28840 33096 28840 33096 0 _0508_
rlabel metal3 30016 33096 30016 33096 0 _0509_
rlabel metal3 25928 55104 25928 55104 0 _0510_
rlabel metal2 23240 52416 23240 52416 0 _0511_
rlabel metal3 25088 54264 25088 54264 0 _0512_
rlabel metal3 32984 56056 32984 56056 0 _0513_
rlabel metal2 24024 56280 24024 56280 0 _0514_
rlabel metal2 25368 54040 25368 54040 0 _0515_
rlabel metal3 26208 53480 26208 53480 0 _0516_
rlabel metal2 26824 54768 26824 54768 0 _0517_
rlabel metal2 26824 53984 26824 53984 0 _0518_
rlabel metal2 24640 54712 24640 54712 0 _0519_
rlabel metal2 26152 53816 26152 53816 0 _0520_
rlabel metal2 20496 50344 20496 50344 0 _0521_
rlabel metal2 23352 53424 23352 53424 0 _0522_
rlabel metal3 24136 52024 24136 52024 0 _0523_
rlabel metal2 38696 56056 38696 56056 0 _0524_
rlabel metal2 23352 50736 23352 50736 0 _0525_
rlabel metal2 22568 51072 22568 51072 0 _0526_
rlabel metal3 23576 51352 23576 51352 0 _0527_
rlabel metal3 21336 51576 21336 51576 0 _0528_
rlabel metal3 22064 51464 22064 51464 0 _0529_
rlabel metal3 22624 51352 22624 51352 0 _0530_
rlabel metal2 20776 49168 20776 49168 0 _0531_
rlabel metal2 17864 55412 17864 55412 0 _0532_
rlabel metal2 19712 58184 19712 58184 0 _0533_
rlabel metal3 18928 56728 18928 56728 0 _0534_
rlabel metal2 21672 57344 21672 57344 0 _0535_
rlabel metal3 23800 59416 23800 59416 0 _0536_
rlabel metal3 21280 59192 21280 59192 0 _0537_
rlabel metal2 20720 57848 20720 57848 0 _0538_
rlabel metal2 19544 57512 19544 57512 0 _0539_
rlabel metal2 21448 58464 21448 58464 0 _0540_
rlabel metal2 22008 58072 22008 58072 0 _0541_
rlabel metal2 21560 58072 21560 58072 0 _0542_
rlabel metal2 19208 57624 19208 57624 0 _0543_
rlabel metal2 18872 57736 18872 57736 0 _0544_
rlabel metal2 26040 59920 26040 59920 0 _0545_
rlabel metal2 27664 59752 27664 59752 0 _0546_
rlabel metal2 28392 60592 28392 60592 0 _0547_
rlabel metal3 26544 60200 26544 60200 0 _0548_
rlabel metal2 26600 60480 26600 60480 0 _0549_
rlabel metal2 38696 65912 38696 65912 0 _0550_
rlabel metal2 28504 60984 28504 60984 0 _0551_
rlabel metal2 26600 61152 26600 61152 0 _0552_
rlabel metal2 25704 58184 25704 58184 0 _0553_
rlabel metal2 24024 53256 24024 53256 0 _0554_
rlabel metal2 24920 57176 24920 57176 0 _0555_
rlabel metal2 25816 58744 25816 58744 0 _0556_
rlabel metal2 22904 58352 22904 58352 0 _0557_
rlabel metal2 23688 57176 23688 57176 0 _0558_
rlabel metal2 22848 57624 22848 57624 0 _0559_
rlabel metal2 23352 58296 23352 58296 0 _0560_
rlabel metal2 22512 60984 22512 60984 0 _0561_
rlabel metal2 23016 57232 23016 57232 0 _0562_
rlabel metal2 25704 61264 25704 61264 0 _0563_
rlabel metal2 24472 61544 24472 61544 0 _0564_
rlabel metal3 23296 62888 23296 62888 0 _0565_
rlabel metal2 25368 61208 25368 61208 0 _0566_
rlabel metal3 23464 60984 23464 60984 0 _0567_
rlabel metal2 22680 63840 22680 63840 0 _0568_
rlabel metal2 24752 60984 24752 60984 0 _0569_
rlabel metal2 26544 64904 26544 64904 0 _0570_
rlabel metal2 23576 64232 23576 64232 0 _0571_
rlabel metal2 25144 61908 25144 61908 0 _0572_
rlabel via2 25592 66024 25592 66024 0 _0573_
rlabel metal2 42616 64120 42616 64120 0 _0574_
rlabel metal2 26712 65240 26712 65240 0 _0575_
rlabel metal2 26600 63784 26600 63784 0 _0576_
rlabel metal3 25424 65688 25424 65688 0 _0577_
rlabel metal2 25648 63112 25648 63112 0 _0578_
rlabel metal2 25144 63448 25144 63448 0 _0579_
rlabel metal3 23744 64120 23744 64120 0 _0580_
rlabel metal2 27496 64288 27496 64288 0 _0581_
rlabel metal2 28896 64568 28896 64568 0 _0582_
rlabel metal2 27944 63672 27944 63672 0 _0583_
rlabel metal2 29960 64680 29960 64680 0 _0584_
rlabel metal2 26936 65464 26936 65464 0 _0585_
rlabel metal3 28840 65464 28840 65464 0 _0586_
rlabel metal3 27832 64120 27832 64120 0 _0587_
rlabel metal2 32424 58688 32424 58688 0 _0588_
rlabel metal2 34664 48328 34664 48328 0 _0589_
rlabel metal2 47656 59808 47656 59808 0 _0590_
rlabel metal2 33152 58632 33152 58632 0 _0591_
rlabel metal2 49112 61040 49112 61040 0 _0592_
rlabel metal2 32536 60144 32536 60144 0 _0593_
rlabel metal2 33544 58744 33544 58744 0 _0594_
rlabel metal3 46368 64120 46368 64120 0 _0595_
rlabel metal2 34216 59556 34216 59556 0 _0596_
rlabel metal2 34552 60088 34552 60088 0 _0597_
rlabel metal2 39816 64736 39816 64736 0 _0598_
rlabel metal2 34328 58800 34328 58800 0 _0599_
rlabel metal2 29064 61656 29064 61656 0 _0600_
rlabel metal2 40040 60088 40040 60088 0 _0601_
rlabel metal2 32984 61432 32984 61432 0 _0602_
rlabel metal3 30576 61432 30576 61432 0 _0603_
rlabel metal2 30856 61656 30856 61656 0 _0604_
rlabel metal2 30408 62384 30408 62384 0 _0605_
rlabel metal2 30408 64064 30408 64064 0 _0606_
rlabel metal3 31248 63000 31248 63000 0 _0607_
rlabel metal2 28168 63112 28168 63112 0 _0608_
rlabel metal2 33544 65800 33544 65800 0 _0609_
rlabel metal2 32424 64120 32424 64120 0 _0610_
rlabel metal3 32592 63896 32592 63896 0 _0611_
rlabel metal2 31752 64176 31752 64176 0 _0612_
rlabel metal2 33880 65128 33880 65128 0 _0613_
rlabel metal2 31640 65016 31640 65016 0 _0614_
rlabel metal3 32816 64008 32816 64008 0 _0615_
rlabel metal2 33208 64232 33208 64232 0 _0616_
rlabel metal3 34104 64120 34104 64120 0 _0617_
rlabel metal2 35000 65184 35000 65184 0 _0618_
rlabel metal2 37408 66248 37408 66248 0 _0619_
rlabel metal2 44800 49112 44800 49112 0 _0620_
rlabel metal3 36624 66136 36624 66136 0 _0621_
rlabel metal2 44408 48048 44408 48048 0 _0622_
rlabel metal2 38416 63224 38416 63224 0 _0623_
rlabel metal2 37688 65184 37688 65184 0 _0624_
rlabel metal2 35896 63616 35896 63616 0 _0625_
rlabel metal2 36120 63224 36120 63224 0 _0626_
rlabel metal3 36288 62888 36288 62888 0 _0627_
rlabel metal2 37128 58632 37128 58632 0 _0628_
rlabel metal2 38864 44968 38864 44968 0 _0629_
rlabel metal2 38024 59472 38024 59472 0 _0630_
rlabel metal2 38136 60872 38136 60872 0 _0631_
rlabel metal2 37464 60256 37464 60256 0 _0632_
rlabel metal2 38136 58128 38136 58128 0 _0633_
rlabel metal2 38808 59864 38808 59864 0 _0634_
rlabel metal2 39704 60088 39704 60088 0 _0635_
rlabel metal2 39144 47880 39144 47880 0 _0636_
rlabel metal3 40040 59416 40040 59416 0 _0637_
rlabel metal2 39368 60032 39368 60032 0 _0638_
rlabel metal2 41608 59584 41608 59584 0 _0639_
rlabel metal2 46424 57624 46424 57624 0 _0640_
rlabel metal2 40992 58632 40992 58632 0 _0641_
rlabel metal2 44968 56448 44968 56448 0 _0642_
rlabel metal3 40544 58520 40544 58520 0 _0643_
rlabel metal2 41832 58912 41832 58912 0 _0644_
rlabel metal2 40992 55944 40992 55944 0 _0645_
rlabel metal2 42280 57680 42280 57680 0 _0646_
rlabel metal3 41272 57848 41272 57848 0 _0647_
rlabel metal2 41888 63112 41888 63112 0 _0648_
rlabel metal2 41496 61712 41496 61712 0 _0649_
rlabel metal2 40040 62440 40040 62440 0 _0650_
rlabel metal2 38696 49392 38696 49392 0 _0651_
rlabel metal3 40936 62664 40936 62664 0 _0652_
rlabel metal2 42168 63896 42168 63896 0 _0653_
rlabel metal2 40320 62888 40320 62888 0 _0654_
rlabel metal2 39648 62328 39648 62328 0 _0655_
rlabel metal2 40376 62608 40376 62608 0 _0656_
rlabel metal3 40376 62216 40376 62216 0 _0657_
rlabel metal3 42056 62328 42056 62328 0 _0658_
rlabel via2 40152 64568 40152 64568 0 _0659_
rlabel metal3 41496 64904 41496 64904 0 _0660_
rlabel metal2 40992 64120 40992 64120 0 _0661_
rlabel metal3 40208 65352 40208 65352 0 _0662_
rlabel metal2 39480 64120 39480 64120 0 _0663_
rlabel metal2 38696 64624 38696 64624 0 _0664_
rlabel metal2 39536 63896 39536 63896 0 _0665_
rlabel metal2 49000 63672 49000 63672 0 _0666_
rlabel metal3 48944 42840 48944 42840 0 _0667_
rlabel metal2 48104 60312 48104 60312 0 _0668_
rlabel metal2 47432 60984 47432 60984 0 _0669_
rlabel metal3 48440 63000 48440 63000 0 _0670_
rlabel metal3 46200 64008 46200 64008 0 _0671_
rlabel metal2 47208 63784 47208 63784 0 _0672_
rlabel metal2 45024 45080 45024 45080 0 _0673_
rlabel metal3 49280 47544 49280 47544 0 _0674_
rlabel metal2 48328 63028 48328 63028 0 _0675_
rlabel metal2 47432 56840 47432 56840 0 _0676_
rlabel metal2 46984 60424 46984 60424 0 _0677_
rlabel metal2 47432 59416 47432 59416 0 _0678_
rlabel metal2 45976 58128 45976 58128 0 _0679_
rlabel metal2 45136 57848 45136 57848 0 _0680_
rlabel metal3 47152 59192 47152 59192 0 _0681_
rlabel metal2 47712 59304 47712 59304 0 _0682_
rlabel metal3 47376 58072 47376 58072 0 _0683_
rlabel metal2 43736 58268 43736 58268 0 _0684_
rlabel metal2 43512 59808 43512 59808 0 _0685_
rlabel metal3 45528 58184 45528 58184 0 _0686_
rlabel metal3 43792 59192 43792 59192 0 _0687_
rlabel metal2 42952 59192 42952 59192 0 _0688_
rlabel metal2 43904 57736 43904 57736 0 _0689_
rlabel metal2 43512 59136 43512 59136 0 _0690_
rlabel metal2 45304 58576 45304 58576 0 _0691_
rlabel metal2 43736 59696 43736 59696 0 _0692_
rlabel metal2 44856 59808 44856 59808 0 _0693_
rlabel metal2 46424 47880 46424 47880 0 _0694_
rlabel metal3 46200 47432 46200 47432 0 _0695_
rlabel metal3 45472 47208 45472 47208 0 _0696_
rlabel metal2 46760 46844 46760 46844 0 _0697_
rlabel metal3 47376 46760 47376 46760 0 _0698_
rlabel metal2 45416 46088 45416 46088 0 _0699_
rlabel metal3 46760 46648 46760 46648 0 _0700_
rlabel metal2 47992 46928 47992 46928 0 _0701_
rlabel metal3 48496 48776 48496 48776 0 _0702_
rlabel metal2 49168 45640 49168 45640 0 _0703_
rlabel metal2 49560 54880 49560 54880 0 _0704_
rlabel metal2 48664 54600 48664 54600 0 _0705_
rlabel metal2 49896 54096 49896 54096 0 _0706_
rlabel metal2 47992 53256 47992 53256 0 _0707_
rlabel metal2 48384 53144 48384 53144 0 _0708_
rlabel metal2 50512 53704 50512 53704 0 _0709_
rlabel metal2 47936 51576 47936 51576 0 _0710_
rlabel metal2 47768 54768 47768 54768 0 _0711_
rlabel metal3 47320 53816 47320 53816 0 _0712_
rlabel metal2 46536 52528 46536 52528 0 _0713_
rlabel metal2 45080 52192 45080 52192 0 _0714_
rlabel metal3 46760 53144 46760 53144 0 _0715_
rlabel metal3 47992 51576 47992 51576 0 _0716_
rlabel metal2 47824 51352 47824 51352 0 _0717_
rlabel metal2 42392 48664 42392 48664 0 _0718_
rlabel metal3 42952 48888 42952 48888 0 _0719_
rlabel metal3 43848 49896 43848 49896 0 _0720_
rlabel metal2 43176 49448 43176 49448 0 _0721_
rlabel metal2 41832 49392 41832 49392 0 _0722_
rlabel metal3 42896 48328 42896 48328 0 _0723_
rlabel metal2 43736 49224 43736 49224 0 _0724_
rlabel metal2 44464 49784 44464 49784 0 _0725_
rlabel metal2 43848 49280 43848 49280 0 _0726_
rlabel metal2 45304 48832 45304 48832 0 _0727_
rlabel metal2 43512 47936 43512 47936 0 _0728_
rlabel metal2 43064 46760 43064 46760 0 _0729_
rlabel metal2 44520 47096 44520 47096 0 _0730_
rlabel metal2 42840 47124 42840 47124 0 _0731_
rlabel metal2 44408 45864 44408 45864 0 _0732_
rlabel metal3 44576 45304 44576 45304 0 _0733_
rlabel metal3 45248 45080 45248 45080 0 _0734_
rlabel metal2 41608 47040 41608 47040 0 _0735_
rlabel metal3 39032 49000 39032 49000 0 _0736_
rlabel metal2 37240 48216 37240 48216 0 _0737_
rlabel metal2 37072 48776 37072 48776 0 _0738_
rlabel metal3 36512 47208 36512 47208 0 _0739_
rlabel metal2 37128 49448 37128 49448 0 _0740_
rlabel metal2 35168 47432 35168 47432 0 _0741_
rlabel metal2 37128 45472 37128 45472 0 _0742_
rlabel metal2 34776 47656 34776 47656 0 _0743_
rlabel metal2 41832 51128 41832 51128 0 _0744_
rlabel metal2 36792 50288 36792 50288 0 _0745_
rlabel metal2 38752 51352 38752 51352 0 _0746_
rlabel metal3 39984 51352 39984 51352 0 _0747_
rlabel metal2 39256 52416 39256 52416 0 _0748_
rlabel metal2 39480 50456 39480 50456 0 _0749_
rlabel metal3 38808 52248 38808 52248 0 _0750_
rlabel metal3 38416 51352 38416 51352 0 _0751_
rlabel metal2 41048 48608 41048 48608 0 _0752_
rlabel metal3 40488 47320 40488 47320 0 _0753_
rlabel metal2 40096 48440 40096 48440 0 _0754_
rlabel metal2 41048 47152 41048 47152 0 _0755_
rlabel metal2 39256 49000 39256 49000 0 _0756_
rlabel metal2 41160 46872 41160 46872 0 _0757_
rlabel metal3 39816 48216 39816 48216 0 _0758_
rlabel metal2 40152 47768 40152 47768 0 _0759_
rlabel metal3 40096 47544 40096 47544 0 _0760_
rlabel metal2 39088 45192 39088 45192 0 _0761_
rlabel metal2 35784 47768 35784 47768 0 _0762_
rlabel metal2 33432 45864 33432 45864 0 _0763_
rlabel metal2 33656 45248 33656 45248 0 _0764_
rlabel metal2 35560 45640 35560 45640 0 _0765_
rlabel metal2 35952 46088 35952 46088 0 _0766_
rlabel metal2 35728 46872 35728 46872 0 _0767_
rlabel metal2 36904 46032 36904 46032 0 _0768_
rlabel metal3 32648 45192 32648 45192 0 _0769_
rlabel metal3 31696 45080 31696 45080 0 _0770_
rlabel metal3 31192 47432 31192 47432 0 _0771_
rlabel metal2 31640 47768 31640 47768 0 _0772_
rlabel metal2 32368 47432 32368 47432 0 _0773_
rlabel metal2 29736 47152 29736 47152 0 _0774_
rlabel metal3 30800 47208 30800 47208 0 _0775_
rlabel metal2 32704 45304 32704 45304 0 _0776_
rlabel metal2 26992 42168 26992 42168 0 _0777_
rlabel metal2 30408 48104 30408 48104 0 _0778_
rlabel metal3 29456 45752 29456 45752 0 _0779_
rlabel metal2 28000 45304 28000 45304 0 _0780_
rlabel metal2 28392 44632 28392 44632 0 _0781_
rlabel metal2 27608 45696 27608 45696 0 _0782_
rlabel metal2 17752 18088 17752 18088 0 _0783_
rlabel metal2 27160 44800 27160 44800 0 _0784_
rlabel metal2 27160 43456 27160 43456 0 _0785_
rlabel metal2 26600 48216 26600 48216 0 _0786_
rlabel metal2 28168 49336 28168 49336 0 _0787_
rlabel metal2 26824 47040 26824 47040 0 _0788_
rlabel metal3 27440 46872 27440 46872 0 _0789_
rlabel metal2 27552 46872 27552 46872 0 _0790_
rlabel metal2 28280 46648 28280 46648 0 _0791_
rlabel metal2 27048 49672 27048 49672 0 _0792_
rlabel metal2 26096 41720 26096 41720 0 _0793_
rlabel metal2 27272 36400 27272 36400 0 _0794_
rlabel metal2 26376 36904 26376 36904 0 _0795_
rlabel metal2 25368 20160 25368 20160 0 _0796_
rlabel metal2 25368 37072 25368 37072 0 _0797_
rlabel metal2 23576 24416 23576 24416 0 _0798_
rlabel metal2 22904 22400 22904 22400 0 _0799_
rlabel metal3 23968 21560 23968 21560 0 _0800_
rlabel metal2 28056 19768 28056 19768 0 _0801_
rlabel metal2 28728 21056 28728 21056 0 _0802_
rlabel metal2 43736 19432 43736 19432 0 _0803_
rlabel metal2 35560 19488 35560 19488 0 _0804_
rlabel metal3 36680 19432 36680 19432 0 _0805_
rlabel metal2 43512 18928 43512 18928 0 _0806_
rlabel metal3 44520 19096 44520 19096 0 _0807_
rlabel metal3 44352 18984 44352 18984 0 _0808_
rlabel metal2 47880 19320 47880 19320 0 _0809_
rlabel metal2 47488 20216 47488 20216 0 _0810_
rlabel metal2 44296 28840 44296 28840 0 _0811_
rlabel metal2 43624 27832 43624 27832 0 _0812_
rlabel metal3 34664 31528 34664 31528 0 _0813_
rlabel metal2 35336 31864 35336 31864 0 _0814_
rlabel metal2 36344 30744 36344 30744 0 _0815_
rlabel metal2 30128 58184 30128 58184 0 _0816_
rlabel metal2 28616 54600 28616 54600 0 _0817_
rlabel metal2 27720 59024 27720 59024 0 _0818_
rlabel metal2 29680 64120 29680 64120 0 _0819_
rlabel metal2 46032 63000 46032 63000 0 _0820_
rlabel metal2 37072 65688 37072 65688 0 _0821_
rlabel metal2 45416 49112 45416 49112 0 _0822_
rlabel metal3 44240 63336 44240 63336 0 _0823_
rlabel metal2 46312 48216 46312 48216 0 _0824_
rlabel metal2 42280 46480 42280 46480 0 _0825_
rlabel metal2 20664 23800 20664 23800 0 _0826_
rlabel metal2 31976 45360 31976 45360 0 _0827_
rlabel metal3 18536 39592 18536 39592 0 _0828_
rlabel metal3 19376 39704 19376 39704 0 _0829_
rlabel metal2 21336 21560 21336 21560 0 _0830_
rlabel metal2 24360 23128 24360 23128 0 _0831_
rlabel metal2 18984 18144 18984 18144 0 _0832_
rlabel metal2 20496 20888 20496 20888 0 _0833_
rlabel metal2 16744 20832 16744 20832 0 _0834_
rlabel metal3 18704 17640 18704 17640 0 _0835_
rlabel metal2 19656 17976 19656 17976 0 _0836_
rlabel metal2 20104 14504 20104 14504 0 _0837_
rlabel metal2 18704 18312 18704 18312 0 _0838_
rlabel metal2 15176 21112 15176 21112 0 _0839_
rlabel metal3 16072 18200 16072 18200 0 _0840_
rlabel metal2 16912 15400 16912 15400 0 _0841_
rlabel metal2 16800 18200 16800 18200 0 _0842_
rlabel metal2 16632 19768 16632 19768 0 _0843_
rlabel metal2 16688 23016 16688 23016 0 _0844_
rlabel metal2 12376 20496 12376 20496 0 _0845_
rlabel metal2 16576 19096 16576 19096 0 _0846_
rlabel metal2 14728 21224 14728 21224 0 _0847_
rlabel metal3 17192 19880 17192 19880 0 _0848_
rlabel metal2 14056 18928 14056 18928 0 _0849_
rlabel metal2 13552 16968 13552 16968 0 _0850_
rlabel metal2 12376 17584 12376 17584 0 _0851_
rlabel metal2 12768 16184 12768 16184 0 _0852_
rlabel metal2 11368 17752 11368 17752 0 _0853_
rlabel metal3 10472 17752 10472 17752 0 _0854_
rlabel metal2 7000 18256 7000 18256 0 _0855_
rlabel metal3 9520 16744 9520 16744 0 _0856_
rlabel metal2 8232 18256 8232 18256 0 _0857_
rlabel metal3 12432 24920 12432 24920 0 _0858_
rlabel via2 9240 21560 9240 21560 0 _0859_
rlabel metal2 6776 20160 6776 20160 0 _0860_
rlabel metal2 11872 22456 11872 22456 0 _0861_
rlabel metal2 9016 21392 9016 21392 0 _0862_
rlabel metal2 10360 24248 10360 24248 0 _0863_
rlabel metal3 7448 22456 7448 22456 0 _0864_
rlabel metal2 8904 24360 8904 24360 0 _0865_
rlabel metal2 11704 26320 11704 26320 0 _0866_
rlabel metal2 8344 25480 8344 25480 0 _0867_
rlabel metal2 15512 28168 15512 28168 0 _0868_
rlabel metal2 11144 25256 11144 25256 0 _0869_
rlabel metal2 12208 24696 12208 24696 0 _0870_
rlabel metal2 14056 27160 14056 27160 0 _0871_
rlabel metal2 13440 27048 13440 27048 0 _0872_
rlabel metal2 11256 29512 11256 29512 0 _0873_
rlabel metal2 10024 28392 10024 28392 0 _0874_
rlabel metal2 12488 30184 12488 30184 0 _0875_
rlabel metal2 9016 29232 9016 29232 0 _0876_
rlabel metal2 12152 31360 12152 31360 0 _0877_
rlabel metal2 9016 31584 9016 31584 0 _0878_
rlabel metal2 10024 32368 10024 32368 0 _0879_
rlabel metal3 13160 38136 13160 38136 0 _0880_
rlabel metal2 10248 34720 10248 34720 0 _0881_
rlabel metal2 10360 36288 10360 36288 0 _0882_
rlabel metal3 12152 38248 12152 38248 0 _0883_
rlabel metal3 13272 39704 13272 39704 0 _0884_
rlabel metal2 14504 61152 14504 61152 0 _0885_
rlabel metal2 16520 49392 16520 49392 0 _0886_
rlabel metal2 18200 48216 18200 48216 0 _0887_
rlabel metal3 17640 50568 17640 50568 0 _0888_
rlabel metal2 17752 48664 17752 48664 0 _0889_
rlabel metal2 17864 47880 17864 47880 0 _0890_
rlabel metal2 16744 49112 16744 49112 0 _0891_
rlabel metal2 16408 52528 16408 52528 0 _0892_
rlabel metal2 16072 50624 16072 50624 0 _0893_
rlabel metal2 16744 52080 16744 52080 0 _0894_
rlabel metal2 15960 53256 15960 53256 0 _0895_
rlabel metal2 14448 50792 14448 50792 0 _0896_
rlabel metal2 14952 53760 14952 53760 0 _0897_
rlabel metal2 16072 58576 16072 58576 0 _0898_
rlabel metal2 15568 54712 15568 54712 0 _0899_
rlabel metal2 16296 58128 16296 58128 0 _0900_
rlabel metal2 16296 56056 16296 56056 0 _0901_
rlabel metal2 13832 57736 13832 57736 0 _0902_
rlabel metal3 17584 58184 17584 58184 0 _0903_
rlabel metal3 16576 58408 16576 58408 0 _0904_
rlabel metal3 16688 56280 16688 56280 0 _0905_
rlabel metal3 17024 58296 17024 58296 0 _0906_
rlabel metal2 15736 59976 15736 59976 0 _0907_
rlabel metal2 16072 60256 16072 60256 0 _0908_
rlabel metal2 16408 64512 16408 64512 0 _0909_
rlabel metal3 16576 60536 16576 60536 0 _0910_
rlabel metal2 13832 64344 13832 64344 0 _0911_
rlabel metal2 16408 62328 16408 62328 0 _0912_
rlabel metal3 17024 63896 17024 63896 0 _0913_
rlabel metal2 14840 64904 14840 64904 0 _0914_
rlabel metal2 16072 64680 16072 64680 0 _0915_
rlabel metal2 18256 65464 18256 65464 0 _0916_
rlabel metal2 14840 63728 14840 63728 0 _0917_
rlabel metal2 14280 65744 14280 65744 0 _0918_
rlabel metal2 13720 65576 13720 65576 0 _0919_
rlabel metal3 12096 63896 12096 63896 0 _0920_
rlabel metal3 13216 64008 13216 64008 0 _0921_
rlabel metal2 11816 64176 11816 64176 0 _0922_
rlabel metal3 13384 63896 13384 63896 0 _0923_
rlabel metal3 12040 63336 12040 63336 0 _0924_
rlabel metal2 8680 49784 8680 49784 0 _0925_
rlabel metal2 11704 62720 11704 62720 0 _0926_
rlabel metal2 12600 62552 12600 62552 0 _0927_
rlabel metal2 10304 61544 10304 61544 0 _0928_
rlabel metal2 11312 62888 11312 62888 0 _0929_
rlabel metal2 12152 60872 12152 60872 0 _0930_
rlabel metal2 11480 60704 11480 60704 0 _0931_
rlabel metal3 8064 50344 8064 50344 0 _0932_
rlabel metal2 10360 56112 10360 56112 0 _0933_
rlabel metal2 11704 57344 11704 57344 0 _0934_
rlabel metal3 8680 50456 8680 50456 0 _0935_
rlabel metal3 10528 56056 10528 56056 0 _0936_
rlabel metal2 11032 57232 11032 57232 0 _0937_
rlabel metal2 10976 53704 10976 53704 0 _0938_
rlabel metal3 8176 54712 8176 54712 0 _0939_
rlabel metal2 10248 54992 10248 54992 0 _0940_
rlabel metal2 10584 56336 10584 56336 0 _0941_
rlabel metal2 9912 56896 9912 56896 0 _0942_
rlabel metal2 8904 57904 8904 57904 0 _0943_
rlabel metal2 9184 56280 9184 56280 0 _0944_
rlabel metal2 6776 54824 6776 54824 0 _0945_
rlabel metal2 8232 56056 8232 56056 0 _0946_
rlabel metal2 7168 54712 7168 54712 0 _0947_
rlabel metal2 7448 55384 7448 55384 0 _0948_
rlabel metal2 6664 55272 6664 55272 0 _0949_
rlabel metal2 8120 50008 8120 50008 0 _0950_
rlabel metal2 7448 54096 7448 54096 0 _0951_
rlabel metal3 7392 53480 7392 53480 0 _0952_
rlabel metal2 7392 52136 7392 52136 0 _0953_
rlabel metal2 6552 52248 6552 52248 0 _0954_
rlabel metal2 7112 51464 7112 51464 0 _0955_
rlabel metal3 7056 45752 7056 45752 0 _0956_
rlabel metal2 7448 48496 7448 48496 0 _0957_
rlabel metal2 7000 48832 7000 48832 0 _0958_
rlabel metal2 6888 49000 6888 49000 0 _0959_
rlabel metal2 7784 46760 7784 46760 0 _0960_
rlabel metal3 9408 48328 9408 48328 0 _0961_
rlabel metal2 9016 46368 9016 46368 0 _0962_
rlabel metal2 7672 43680 7672 43680 0 _0963_
rlabel metal2 7000 45920 7000 45920 0 _0964_
rlabel metal3 8232 44184 8232 44184 0 _0965_
rlabel metal3 8344 45304 8344 45304 0 _0966_
rlabel metal3 11144 47208 11144 47208 0 _0967_
rlabel metal3 10976 45864 10976 45864 0 _0968_
rlabel metal2 11480 47096 11480 47096 0 _0969_
rlabel metal2 10080 45864 10080 45864 0 _0970_
rlabel metal2 11704 46312 11704 46312 0 _0971_
rlabel metal2 11368 47824 11368 47824 0 _0972_
rlabel metal2 12824 47824 12824 47824 0 _0973_
rlabel metal3 12936 51464 12936 51464 0 _0974_
rlabel metal3 11872 50456 11872 50456 0 _0975_
rlabel metal2 12600 49112 12600 49112 0 _0976_
rlabel metal2 23576 46144 23576 46144 0 _0977_
rlabel metal2 46760 41664 46760 41664 0 _0978_
rlabel metal2 25144 43960 25144 43960 0 _0979_
rlabel metal2 22568 46368 22568 46368 0 _0980_
rlabel metal2 38864 34328 38864 34328 0 _0981_
rlabel metal2 26600 34776 26600 34776 0 _0982_
rlabel metal3 23688 37240 23688 37240 0 _0983_
rlabel metal2 23072 37464 23072 37464 0 _0984_
rlabel metal2 25480 41832 25480 41832 0 _0985_
rlabel metal3 24248 43960 24248 43960 0 _0986_
rlabel metal2 23240 46536 23240 46536 0 _0987_
rlabel metal2 22344 46536 22344 46536 0 _0988_
rlabel metal2 21896 37800 21896 37800 0 _0989_
rlabel metal2 22120 45864 22120 45864 0 _0990_
rlabel metal2 21560 46564 21560 46564 0 _0991_
rlabel metal2 21056 42952 21056 42952 0 _0992_
rlabel metal2 21560 47488 21560 47488 0 _0993_
rlabel metal2 22120 43008 22120 43008 0 _0994_
rlabel metal2 24304 37464 24304 37464 0 _0995_
rlabel metal2 23800 43120 23800 43120 0 _0996_
rlabel metal3 23632 43512 23632 43512 0 _0997_
rlabel metal3 26320 34104 26320 34104 0 _0998_
rlabel metal2 26264 35392 26264 35392 0 _0999_
rlabel metal2 25816 31416 25816 31416 0 _1000_
rlabel metal2 24472 29288 24472 29288 0 _1001_
rlabel metal2 24808 33432 24808 33432 0 _1002_
rlabel metal3 25648 42616 25648 42616 0 _1003_
rlabel metal2 24808 41720 24808 41720 0 _1004_
rlabel metal3 24080 34104 24080 34104 0 _1005_
rlabel metal3 24696 32760 24696 32760 0 _1006_
rlabel metal2 23968 41384 23968 41384 0 _1007_
rlabel metal3 25984 31528 25984 31528 0 _1008_
rlabel metal2 22512 28840 22512 28840 0 _1009_
rlabel metal2 24808 42336 24808 42336 0 _1010_
rlabel metal2 25592 30016 25592 30016 0 _1011_
rlabel metal3 25312 29400 25312 29400 0 _1012_
rlabel metal2 26712 42672 26712 42672 0 _1013_
rlabel metal3 26152 42504 26152 42504 0 _1014_
rlabel metal3 35000 40488 35000 40488 0 _1015_
rlabel metal3 34608 40376 34608 40376 0 _1016_
rlabel metal3 35616 34776 35616 34776 0 _1017_
rlabel metal3 33040 40376 33040 40376 0 _1018_
rlabel metal2 34216 42672 34216 42672 0 _1019_
rlabel metal2 33880 41440 33880 41440 0 _1020_
rlabel metal2 34440 35952 34440 35952 0 _1021_
rlabel metal2 33320 35392 33320 35392 0 _1022_
rlabel metal2 32984 40572 32984 40572 0 _1023_
rlabel metal3 35728 40376 35728 40376 0 _1024_
rlabel metal2 35000 34888 35000 34888 0 _1025_
rlabel metal2 34888 40880 34888 40880 0 _1026_
rlabel metal3 36512 35112 36512 35112 0 _1027_
rlabel metal2 36120 35560 36120 35560 0 _1028_
rlabel metal2 46200 41048 46200 41048 0 _1029_
rlabel metal2 38808 43120 38808 43120 0 _1030_
rlabel metal2 36400 42056 36400 42056 0 _1031_
rlabel metal3 40432 35672 40432 35672 0 _1032_
rlabel metal2 42672 36344 42672 36344 0 _1033_
rlabel metal2 45752 34608 45752 34608 0 _1034_
rlabel metal3 44408 34776 44408 34776 0 _1035_
rlabel metal2 39816 35000 39816 35000 0 _1036_
rlabel metal2 38696 42952 38696 42952 0 _1037_
rlabel metal2 39536 38696 39536 38696 0 _1038_
rlabel metal2 41608 35560 41608 35560 0 _1039_
rlabel metal2 41328 33320 41328 33320 0 _1040_
rlabel metal2 41216 39032 41216 39032 0 _1041_
rlabel metal3 43176 37800 43176 37800 0 _1042_
rlabel metal2 44968 36008 44968 36008 0 _1043_
rlabel metal2 42336 38024 42336 38024 0 _1044_
rlabel metal2 42616 35168 42616 35168 0 _1045_
rlabel metal3 43008 34664 43008 34664 0 _1046_
rlabel metal2 46424 42952 46424 42952 0 _1047_
rlabel metal2 42112 40600 42112 40600 0 _1048_
rlabel metal2 46424 36848 46424 36848 0 _1049_
rlabel metal2 47768 37632 47768 37632 0 _1050_
rlabel metal2 46872 34440 46872 34440 0 _1051_
rlabel metal2 46592 34328 46592 34328 0 _1052_
rlabel metal2 48216 43120 48216 43120 0 _1053_
rlabel metal2 46704 39592 46704 39592 0 _1054_
rlabel metal2 49224 36960 49224 36960 0 _1055_
rlabel metal2 48160 33544 48160 33544 0 _1056_
rlabel metal3 48720 40488 48720 40488 0 _1057_
rlabel metal3 48048 37800 48048 37800 0 _1058_
rlabel metal2 47432 36064 47432 36064 0 _1059_
rlabel metal2 46928 40376 46928 40376 0 _1060_
rlabel metal2 47992 36064 47992 36064 0 _1061_
rlabel metal2 48888 34216 48888 34216 0 _1062_
rlabel metal3 48216 44184 48216 44184 0 _1063_
rlabel metal2 47824 40488 47824 40488 0 _1064_
rlabel metal2 49224 39984 49224 39984 0 _1065_
rlabel metal2 49784 42336 49784 42336 0 _1066_
rlabel metal2 50680 33376 50680 33376 0 _1067_
rlabel metal2 49504 38808 49504 38808 0 _1068_
rlabel metal3 49056 44296 49056 44296 0 _1069_
rlabel metal2 49336 43876 49336 43876 0 _1070_
rlabel metal3 50288 41384 50288 41384 0 _1071_
rlabel metal2 50512 33544 50512 33544 0 _1072_
rlabel metal3 48272 41944 48272 41944 0 _1073_
rlabel metal3 50064 42504 50064 42504 0 _1074_
rlabel metal2 49168 42504 49168 42504 0 _1075_
rlabel metal2 48776 43876 48776 43876 0 _1076_
rlabel metal3 47040 39368 47040 39368 0 _1077_
rlabel metal2 46200 39004 46200 39004 0 _1078_
rlabel metal2 45416 42672 45416 42672 0 _1079_
rlabel metal2 45976 41048 45976 41048 0 _1080_
rlabel metal3 40432 38808 40432 38808 0 _1081_
rlabel metal2 40936 40656 40936 40656 0 _1082_
rlabel metal2 40936 34496 40936 34496 0 _1083_
rlabel metal2 39928 39508 39928 39508 0 _1084_
rlabel metal3 40992 42728 40992 42728 0 _1085_
rlabel metal2 40040 41440 40040 41440 0 _1086_
rlabel metal2 41496 39648 41496 39648 0 _1087_
rlabel metal2 43288 36064 43288 36064 0 _1088_
rlabel metal2 41944 40600 41944 40600 0 _1089_
rlabel metal2 42952 40880 42952 40880 0 _1090_
rlabel metal2 41440 39144 41440 39144 0 _1091_
rlabel metal2 40992 42056 40992 42056 0 _1092_
rlabel metal2 39368 39256 39368 39256 0 _1093_
rlabel metal2 38640 40376 38640 40376 0 _1094_
rlabel metal2 37352 42672 37352 42672 0 _1095_
rlabel metal2 38472 40992 38472 40992 0 _1096_
rlabel metal3 32760 38248 32760 38248 0 _1097_
rlabel metal3 30520 39592 30520 39592 0 _1098_
rlabel metal3 30968 37352 30968 37352 0 _1099_
rlabel metal2 31416 38724 31416 38724 0 _1100_
rlabel metal2 31136 38920 31136 38920 0 _1101_
rlabel metal2 31472 39368 31472 39368 0 _1102_
rlabel metal2 30968 39004 30968 39004 0 _1103_
rlabel metal2 30744 39760 30744 39760 0 _1104_
rlabel metal3 29400 41160 29400 41160 0 _1105_
rlabel metal2 30240 37240 30240 37240 0 _1106_
rlabel metal2 29176 42280 29176 42280 0 _1107_
rlabel metal2 29400 38080 29400 38080 0 _1108_
rlabel metal2 29288 36792 29288 36792 0 _1109_
rlabel metal2 29792 37800 29792 37800 0 _1110_
rlabel metal2 18536 36232 18536 36232 0 _1111_
rlabel metal3 17024 38248 17024 38248 0 _1112_
rlabel metal2 22456 42504 22456 42504 0 _1113_
rlabel metal2 26488 41552 26488 41552 0 _1114_
rlabel metal3 19208 41048 19208 41048 0 _1115_
rlabel metal2 16632 41216 16632 41216 0 _1116_
rlabel metal2 19712 41160 19712 41160 0 _1117_
rlabel via3 29848 40712 29848 40712 0 _1118_
rlabel metal2 45416 39424 45416 39424 0 _1119_
rlabel metal3 12992 42616 12992 42616 0 _1120_
rlabel metal2 13496 43960 13496 43960 0 _1121_
rlabel metal2 11816 43680 11816 43680 0 _1122_
rlabel metal2 10976 41384 10976 41384 0 _1123_
rlabel metal2 16184 24752 16184 24752 0 _1124_
rlabel metal2 11592 41384 11592 41384 0 _1125_
rlabel metal2 10696 41832 10696 41832 0 _1126_
rlabel metal2 10920 42392 10920 42392 0 _1127_
rlabel metal2 10136 43120 10136 43120 0 _1128_
rlabel metal2 11032 42560 11032 42560 0 _1129_
rlabel metal2 11704 43232 11704 43232 0 _1130_
rlabel metal2 12992 43512 12992 43512 0 _1131_
rlabel metal2 19096 42112 19096 42112 0 _1132_
rlabel metal2 18088 34664 18088 34664 0 _1133_
rlabel metal3 17920 35112 17920 35112 0 _1134_
rlabel metal2 18088 36568 18088 36568 0 _1135_
rlabel metal2 19768 48776 19768 48776 0 _1136_
rlabel metal2 17976 36400 17976 36400 0 _1137_
rlabel metal3 24584 52136 24584 52136 0 _1138_
rlabel metal2 25592 41104 25592 41104 0 _1139_
rlabel metal2 25816 41664 25816 41664 0 _1140_
rlabel metal2 21448 39872 21448 39872 0 _1141_
rlabel metal2 18648 37184 18648 37184 0 _1142_
rlabel metal2 19208 37128 19208 37128 0 _1143_
rlabel metal3 24136 38696 24136 38696 0 _1144_
rlabel metal2 23240 35616 23240 35616 0 _1145_
rlabel metal3 39928 49112 39928 49112 0 _1146_
rlabel metal3 23352 24920 23352 24920 0 _1147_
rlabel metal3 21336 39144 21336 39144 0 _1148_
rlabel metal2 12488 44688 12488 44688 0 _1149_
rlabel metal2 21448 24248 21448 24248 0 _1150_
rlabel metal2 19544 38136 19544 38136 0 _1151_
rlabel metal2 17528 43008 17528 43008 0 _1152_
rlabel metal2 17976 32592 17976 32592 0 _1153_
rlabel metal2 16408 31248 16408 31248 0 _1154_
rlabel metal2 16296 30184 16296 30184 0 _1155_
rlabel metal2 16072 31416 16072 31416 0 _1156_
rlabel metal2 16072 39368 16072 39368 0 _1157_
rlabel metal2 15288 39312 15288 39312 0 _1158_
rlabel metal2 15288 32648 15288 32648 0 _1159_
rlabel metal2 24920 32256 24920 32256 0 _1160_
rlabel metal2 16296 33432 16296 33432 0 _1161_
rlabel metal2 14112 31976 14112 31976 0 _1162_
rlabel metal2 14952 33600 14952 33600 0 _1163_
rlabel metal2 15176 34832 15176 34832 0 _1164_
rlabel metal2 17304 36456 17304 36456 0 _1165_
rlabel metal2 23800 59976 23800 59976 0 _1166_
rlabel metal2 24696 47992 24696 47992 0 _1167_
rlabel metal2 18704 59192 18704 59192 0 _1168_
rlabel metal3 16464 37912 16464 37912 0 _1169_
rlabel metal2 15792 39480 15792 39480 0 _1170_
rlabel metal2 20160 26488 20160 26488 0 _1171_
rlabel metal2 21392 36232 21392 36232 0 _1172_
rlabel metal2 15176 25592 15176 25592 0 _1173_
rlabel metal2 22344 13552 22344 13552 0 _1174_
rlabel metal2 21952 14616 21952 14616 0 _1175_
rlabel metal3 19264 26264 19264 26264 0 _1176_
rlabel metal2 18424 28672 18424 28672 0 _1177_
rlabel metal3 17528 26040 17528 26040 0 _1178_
rlabel metal2 24024 12600 24024 12600 0 _1179_
rlabel metal2 18088 25424 18088 25424 0 _1180_
rlabel metal2 23800 12208 23800 12208 0 _1181_
rlabel metal2 20832 12152 20832 12152 0 _1182_
rlabel metal2 21448 10080 21448 10080 0 _1183_
rlabel metal2 24136 12376 24136 12376 0 _1184_
rlabel metal2 21504 14392 21504 14392 0 _1185_
rlabel metal2 25032 12600 25032 12600 0 _1186_
rlabel metal2 19656 10360 19656 10360 0 _1187_
rlabel metal2 24584 10080 24584 10080 0 _1188_
rlabel metal2 42840 11872 42840 11872 0 _1189_
rlabel metal2 29288 11032 29288 11032 0 _1190_
rlabel metal2 26600 8568 26600 8568 0 _1191_
rlabel metal3 30744 17528 30744 17528 0 _1192_
rlabel metal3 28728 11368 28728 11368 0 _1193_
rlabel metal2 28168 9184 28168 9184 0 _1194_
rlabel metal2 34776 10528 34776 10528 0 _1195_
rlabel metal2 32536 11536 32536 11536 0 _1196_
rlabel metal2 31640 10248 31640 10248 0 _1197_
rlabel metal2 36792 10920 36792 10920 0 _1198_
rlabel metal2 34104 9352 34104 9352 0 _1199_
rlabel metal2 36680 11172 36680 11172 0 _1200_
rlabel metal3 40320 11256 40320 11256 0 _1201_
rlabel metal2 34832 12824 34832 12824 0 _1202_
rlabel metal2 42672 11368 42672 11368 0 _1203_
rlabel metal2 36344 8512 36344 8512 0 _1204_
rlabel metal2 38696 11536 38696 11536 0 _1205_
rlabel metal3 45416 7336 45416 7336 0 _1206_
rlabel metal2 40376 10360 40376 10360 0 _1207_
rlabel metal2 43904 13608 43904 13608 0 _1208_
rlabel metal2 44184 10864 44184 10864 0 _1209_
rlabel metal2 42448 10472 42448 10472 0 _1210_
rlabel metal2 42560 23688 42560 23688 0 _1211_
rlabel metal2 45696 7672 45696 7672 0 _1212_
rlabel metal2 42168 7280 42168 7280 0 _1213_
rlabel metal2 45080 6328 45080 6328 0 _1214_
rlabel metal2 44352 11144 44352 11144 0 _1215_
rlabel metal2 45528 10024 45528 10024 0 _1216_
rlabel metal2 45248 22120 45248 22120 0 _1217_
rlabel metal2 18536 20888 18536 20888 0 _1218_
rlabel metal2 43624 25032 43624 25032 0 _1219_
rlabel metal2 44184 21280 44184 21280 0 _1220_
rlabel metal3 43792 23128 43792 23128 0 _1221_
rlabel metal2 43512 22680 43512 22680 0 _1222_
rlabel metal2 44856 26488 44856 26488 0 _1223_
rlabel metal2 19096 23856 19096 23856 0 _1224_
rlabel metal2 41608 23968 41608 23968 0 _1225_
rlabel metal3 43344 24472 43344 24472 0 _1226_
rlabel metal2 39032 26600 39032 26600 0 _1227_
rlabel metal2 40936 23016 40936 23016 0 _1228_
rlabel metal2 42840 23296 42840 23296 0 _1229_
rlabel metal2 34776 26208 34776 26208 0 _1230_
rlabel metal2 40264 21224 40264 21224 0 _1231_
rlabel metal2 38696 22568 38696 22568 0 _1232_
rlabel metal2 32312 21616 32312 21616 0 _1233_
rlabel metal2 35896 26096 35896 26096 0 _1234_
rlabel metal2 33992 25256 33992 25256 0 _1235_
rlabel metal2 24024 21000 24024 21000 0 _1236_
rlabel metal2 33488 24808 33488 24808 0 _1237_
rlabel metal2 23240 21784 23240 21784 0 _1238_
rlabel metal2 30968 22120 30968 22120 0 _1239_
rlabel metal2 29176 22904 29176 22904 0 _1240_
rlabel metal2 24024 52248 24024 52248 0 _1241_
rlabel metal2 21000 52864 21000 52864 0 _1242_
rlabel metal2 21392 50456 21392 50456 0 _1243_
rlabel metal2 19656 44800 19656 44800 0 _1244_
rlabel metal3 20832 44072 20832 44072 0 _1245_
rlabel metal2 21336 44800 21336 44800 0 _1246_
rlabel metal2 21672 52528 21672 52528 0 _1247_
rlabel metal2 20664 54096 20664 54096 0 _1248_
rlabel metal3 32704 53144 32704 53144 0 _1249_
rlabel metal2 20328 51968 20328 51968 0 _1250_
rlabel metal2 19264 51464 19264 51464 0 _1251_
rlabel metal3 21112 59976 21112 59976 0 _1252_
rlabel metal2 20664 60312 20664 60312 0 _1253_
rlabel metal2 19432 51632 19432 51632 0 _1254_
rlabel metal2 19656 51688 19656 51688 0 _1255_
rlabel metal2 20216 53480 20216 53480 0 _1256_
rlabel metal2 19432 53592 19432 53592 0 _1257_
rlabel metal2 19208 52640 19208 52640 0 _1258_
rlabel metal2 20664 52304 20664 52304 0 _1259_
rlabel metal2 22120 58688 22120 58688 0 _1260_
rlabel metal2 21784 61544 21784 61544 0 _1261_
rlabel metal3 20244 60760 20244 60760 0 _1262_
rlabel metal2 20216 60648 20216 60648 0 _1263_
rlabel metal2 18984 60928 18984 60928 0 _1264_
rlabel metal2 21336 67032 21336 67032 0 _1265_
rlabel metal2 20888 63896 20888 63896 0 _1266_
rlabel metal2 21392 62888 21392 62888 0 _1267_
rlabel metal2 19880 63504 19880 63504 0 _1268_
rlabel metal2 22120 67424 22120 67424 0 _1269_
rlabel metal3 23520 56728 23520 56728 0 _1270_
rlabel metal2 22904 67312 22904 67312 0 _1271_
rlabel metal2 21672 65464 21672 65464 0 _1272_
rlabel metal2 22344 66752 22344 66752 0 _1273_
rlabel metal3 21672 66360 21672 66360 0 _1274_
rlabel metal3 22120 67032 22120 67032 0 _1275_
rlabel metal2 22568 67536 22568 67536 0 _1276_
rlabel metal3 21672 67704 21672 67704 0 _1277_
rlabel metal2 41160 66976 41160 66976 0 _1278_
rlabel metal2 24472 67536 24472 67536 0 _1279_
rlabel metal3 23688 67144 23688 67144 0 _1280_
rlabel metal2 23912 68544 23912 68544 0 _1281_
rlabel metal2 24584 69440 24584 69440 0 _1282_
rlabel metal2 26264 67424 26264 67424 0 _1283_
rlabel metal2 26432 67592 26432 67592 0 _1284_
rlabel metal2 25144 67872 25144 67872 0 _1285_
rlabel metal2 25760 67928 25760 67928 0 _1286_
rlabel metal2 33096 69104 33096 69104 0 _1287_
rlabel metal2 30408 67256 30408 67256 0 _1288_
rlabel metal2 33320 69048 33320 69048 0 _1289_
rlabel metal2 29512 67200 29512 67200 0 _1290_
rlabel metal2 30968 68264 30968 68264 0 _1291_
rlabel metal2 30520 68320 30520 68320 0 _1292_
rlabel metal3 30464 69272 30464 69272 0 _1293_
rlabel metal2 30408 69496 30408 69496 0 _1294_
rlabel metal2 29456 67928 29456 67928 0 _1295_
rlabel metal3 37744 68824 37744 68824 0 _1296_
rlabel metal2 31080 67536 31080 67536 0 _1297_
rlabel metal2 33432 68936 33432 68936 0 _1298_
rlabel metal2 32984 69776 32984 69776 0 _1299_
rlabel metal2 26712 53200 26712 53200 0 _1300_
rlabel metal3 39256 68656 39256 68656 0 _1301_
rlabel metal2 35504 69608 35504 69608 0 _1302_
rlabel metal3 34328 69160 34328 69160 0 _1303_
rlabel metal2 34328 69720 34328 69720 0 _1304_
rlabel metal2 42392 56448 42392 56448 0 _1305_
rlabel metal2 40152 69552 40152 69552 0 _1306_
rlabel metal2 38808 68264 38808 68264 0 _1307_
rlabel metal2 40152 68544 40152 68544 0 _1308_
rlabel metal2 36736 68712 36736 68712 0 _1309_
rlabel metal2 37240 68824 37240 68824 0 _1310_
rlabel metal3 36960 69272 36960 69272 0 _1311_
rlabel metal2 37464 68320 37464 68320 0 _1312_
rlabel metal2 38248 68992 38248 68992 0 _1313_
rlabel metal2 40376 71120 40376 71120 0 _1314_
rlabel metal2 42504 66976 42504 66976 0 _1315_
rlabel metal2 39648 68600 39648 68600 0 _1316_
rlabel metal2 39816 69720 39816 69720 0 _1317_
rlabel metal2 40264 71008 40264 71008 0 _1318_
rlabel metal3 44128 65688 44128 65688 0 _1319_
rlabel metal2 41104 66472 41104 66472 0 _1320_
rlabel metal2 40936 68320 40936 68320 0 _1321_
rlabel metal3 40264 68824 40264 68824 0 _1322_
rlabel metal2 43512 67256 43512 67256 0 _1323_
rlabel metal2 43960 65520 43960 65520 0 _1324_
rlabel metal3 42112 55272 42112 55272 0 _1325_
rlabel metal3 43512 62888 43512 62888 0 _1326_
rlabel metal2 42728 66192 42728 66192 0 _1327_
rlabel metal3 43736 66472 43736 66472 0 _1328_
rlabel metal2 45304 65800 45304 65800 0 _1329_
rlabel metal2 43624 65744 43624 65744 0 _1330_
rlabel metal2 42840 66976 42840 66976 0 _1331_
rlabel metal2 45528 67172 45528 67172 0 _1332_
rlabel metal2 44184 57344 44184 57344 0 _1333_
rlabel metal2 44184 65968 44184 65968 0 _1334_
rlabel metal2 43960 66752 43960 66752 0 _1335_
rlabel metal2 43512 66920 43512 66920 0 _1336_
rlabel metal2 43904 56616 43904 56616 0 _1337_
rlabel metal2 43848 62776 43848 62776 0 _1338_
rlabel metal2 44408 64008 44408 64008 0 _1339_
rlabel metal3 44688 64456 44688 64456 0 _1340_
rlabel metal2 43960 54376 43960 54376 0 _1341_
rlabel metal2 44072 56280 44072 56280 0 _1342_
rlabel metal4 41832 54040 41832 54040 0 _1343_
rlabel metal2 45136 56168 45136 56168 0 _1344_
rlabel metal2 44408 55552 44408 55552 0 _1345_
rlabel metal2 43848 55440 43848 55440 0 _1346_
rlabel metal2 43736 56392 43736 56392 0 _1347_
rlabel metal2 44296 54768 44296 54768 0 _1348_
rlabel metal3 44352 53592 44352 53592 0 _1349_
rlabel metal2 42840 52948 42840 52948 0 _1350_
rlabel metal2 43064 54208 43064 54208 0 _1351_
rlabel metal2 42728 55608 42728 55608 0 _1352_
rlabel metal3 41664 55160 41664 55160 0 _1353_
rlabel metal2 40488 53312 40488 53312 0 _1354_
rlabel metal2 42224 52920 42224 52920 0 _1355_
rlabel metal2 42504 53144 42504 53144 0 _1356_
rlabel metal2 43176 53088 43176 53088 0 _1357_
rlabel metal2 35112 53984 35112 53984 0 _1358_
rlabel metal2 35784 53816 35784 53816 0 _1359_
rlabel metal3 36008 53144 36008 53144 0 _1360_
rlabel metal2 41048 53256 41048 53256 0 _1361_
rlabel metal2 36456 53424 36456 53424 0 _1362_
rlabel metal2 34944 52248 34944 52248 0 _1363_
rlabel metal3 37408 53704 37408 53704 0 _1364_
rlabel metal2 37128 54320 37128 54320 0 _1365_
rlabel metal2 37464 55272 37464 55272 0 _1366_
rlabel metal2 35448 53200 35448 53200 0 _1367_
rlabel metal3 36456 52920 36456 52920 0 _1368_
rlabel metal3 35616 54264 35616 54264 0 _1369_
rlabel metal2 36344 55104 36344 55104 0 _1370_
rlabel metal3 26460 53032 26460 53032 0 _1371_
rlabel metal2 34888 52808 34888 52808 0 _1372_
rlabel metal2 35560 53424 35560 53424 0 _1373_
rlabel metal2 35000 54096 35000 54096 0 _1374_
rlabel metal3 23408 50680 23408 50680 0 _1375_
rlabel metal3 30800 49896 30800 49896 0 _1376_
rlabel metal2 29512 54152 29512 54152 0 _1377_
rlabel metal2 32424 52528 32424 52528 0 _1378_
rlabel metal2 30408 52360 30408 52360 0 _1379_
rlabel metal2 30072 51296 30072 51296 0 _1380_
rlabel metal2 30688 52136 30688 52136 0 _1381_
rlabel metal2 29512 52864 29512 52864 0 _1382_
rlabel metal2 28616 51744 28616 51744 0 _1383_
rlabel metal2 28280 53032 28280 53032 0 _1384_
rlabel metal2 29064 52416 29064 52416 0 _1385_
rlabel metal2 29288 52640 29288 52640 0 _1386_
rlabel metal2 25256 52528 25256 52528 0 _1387_
rlabel metal2 17528 54264 17528 54264 0 _1388_
rlabel metal2 27608 53704 27608 53704 0 _1389_
rlabel metal2 27048 52192 27048 52192 0 _1390_
rlabel metal2 26376 50344 26376 50344 0 _1391_
rlabel metal2 18200 44968 18200 44968 0 _1392_
rlabel metal2 17528 50400 17528 50400 0 _1393_
rlabel metal3 13160 53032 13160 53032 0 _1394_
rlabel metal2 15680 52920 15680 52920 0 _1395_
rlabel metal2 15848 47880 15848 47880 0 _1396_
rlabel metal2 15960 28336 15960 28336 0 _1397_
rlabel metal3 26516 40936 26516 40936 0 _1398_
rlabel metal2 20664 24640 20664 24640 0 _1399_
rlabel metal2 16520 27888 16520 27888 0 _1400_
rlabel metal2 29736 45752 29736 45752 0 _1401_
rlabel metal2 29960 45920 29960 45920 0 _1402_
rlabel metal3 34048 49000 34048 49000 0 _1403_
rlabel metal3 22568 57736 22568 57736 0 _1404_
rlabel metal2 25368 52752 25368 52752 0 _1405_
rlabel metal2 25816 19152 25816 19152 0 _1406_
rlabel metal3 22064 30184 22064 30184 0 _1407_
rlabel metal2 32088 24528 32088 24528 0 _1408_
rlabel metal2 24696 15400 24696 15400 0 _1409_
rlabel metal2 45584 27048 45584 27048 0 _1410_
rlabel metal2 22792 52584 22792 52584 0 _1411_
rlabel metal3 22400 30856 22400 30856 0 _1412_
rlabel metal2 22064 31976 22064 31976 0 _1413_
rlabel metal2 21560 59640 21560 59640 0 _1414_
rlabel metal3 22120 35672 22120 35672 0 _1415_
rlabel metal2 20664 35504 20664 35504 0 _1416_
rlabel metal2 21672 35896 21672 35896 0 _1417_
rlabel metal2 22120 35448 22120 35448 0 _1418_
rlabel metal3 24024 51352 24024 51352 0 _1419_
rlabel metal2 22344 35000 22344 35000 0 _1420_
rlabel metal3 21280 34776 21280 34776 0 _1421_
rlabel metal2 28392 17528 28392 17528 0 _1422_
rlabel metal3 34888 23688 34888 23688 0 _1423_
rlabel metal2 22680 15512 22680 15512 0 _1424_
rlabel metal2 21672 28952 21672 28952 0 _1425_
rlabel metal2 25144 27160 25144 27160 0 _1426_
rlabel metal2 25480 27048 25480 27048 0 _1427_
rlabel metal2 22904 29344 22904 29344 0 _1428_
rlabel metal2 21560 27608 21560 27608 0 _1429_
rlabel metal3 23408 27160 23408 27160 0 _1430_
rlabel metal2 22568 27440 22568 27440 0 _1431_
rlabel metal3 22960 28056 22960 28056 0 _1432_
rlabel metal2 24024 26488 24024 26488 0 _1433_
rlabel metal3 23296 26264 23296 26264 0 _1434_
rlabel metal3 24304 27832 24304 27832 0 _1435_
rlabel metal3 40656 48888 40656 48888 0 _1436_
rlabel metal2 26376 23240 26376 23240 0 _1437_
rlabel metal2 24808 26656 24808 26656 0 _1438_
rlabel metal2 26600 24864 26600 24864 0 _1439_
rlabel metal3 2478 70616 2478 70616 0 clk
rlabel metal2 26376 55608 26376 55608 0 clknet_0_clk
rlabel metal2 22792 11480 22792 11480 0 clknet_2_0__leaf_clk
rlabel metal2 50736 15512 50736 15512 0 clknet_2_1__leaf_clk
rlabel metal2 23800 50456 23800 50456 0 clknet_2_2__leaf_clk
rlabel metal2 49504 49784 49504 49784 0 clknet_2_3__leaf_clk
rlabel metal2 6048 20776 6048 20776 0 clknet_leaf_0_clk
rlabel metal3 12320 49784 12320 49784 0 clknet_leaf_10_clk
rlabel metal2 9576 59976 9576 59976 0 clknet_leaf_11_clk
rlabel metal2 6216 58072 6216 58072 0 clknet_leaf_12_clk
rlabel metal2 14616 64736 14616 64736 0 clknet_leaf_13_clk
rlabel metal2 17696 61544 17696 61544 0 clknet_leaf_14_clk
rlabel metal2 23016 65072 23016 65072 0 clknet_leaf_15_clk
rlabel metal2 25704 57008 25704 57008 0 clknet_leaf_16_clk
rlabel metal2 21336 54040 21336 54040 0 clknet_leaf_17_clk
rlabel metal2 25200 51352 25200 51352 0 clknet_leaf_18_clk
rlabel metal2 30408 44296 30408 44296 0 clknet_leaf_19_clk
rlabel metal2 13496 20832 13496 20832 0 clknet_leaf_1_clk
rlabel metal2 34440 53648 34440 53648 0 clknet_leaf_20_clk
rlabel metal2 31192 64792 31192 64792 0 clknet_leaf_21_clk
rlabel metal2 39592 69944 39592 69944 0 clknet_leaf_22_clk
rlabel metal2 37464 65016 37464 65016 0 clknet_leaf_23_clk
rlabel metal2 45416 62664 45416 62664 0 clknet_leaf_25_clk
rlabel metal2 40936 70224 40936 70224 0 clknet_leaf_26_clk
rlabel metal2 47544 67816 47544 67816 0 clknet_leaf_27_clk
rlabel metal2 45472 48216 45472 48216 0 clknet_leaf_28_clk
rlabel metal2 51688 52192 51688 52192 0 clknet_leaf_29_clk
rlabel metal2 5656 25088 5656 25088 0 clknet_leaf_2_clk
rlabel metal2 48664 41328 48664 41328 0 clknet_leaf_30_clk
rlabel metal2 40936 45528 40936 45528 0 clknet_leaf_31_clk
rlabel metal2 33320 39144 33320 39144 0 clknet_leaf_32_clk
rlabel metal2 35560 33824 35560 33824 0 clknet_leaf_33_clk
rlabel metal2 41160 30632 41160 30632 0 clknet_leaf_34_clk
rlabel metal2 48776 36008 48776 36008 0 clknet_leaf_35_clk
rlabel metal2 51352 29064 51352 29064 0 clknet_leaf_36_clk
rlabel metal2 47096 20776 47096 20776 0 clknet_leaf_37_clk
rlabel metal2 51688 16744 51688 16744 0 clknet_leaf_38_clk
rlabel metal2 44968 8316 44968 8316 0 clknet_leaf_39_clk
rlabel metal2 8456 35672 8456 35672 0 clknet_leaf_3_clk
rlabel metal2 39368 10752 39368 10752 0 clknet_leaf_40_clk
rlabel metal3 36680 8904 36680 8904 0 clknet_leaf_41_clk
rlabel metal3 29848 16184 29848 16184 0 clknet_leaf_42_clk
rlabel metal2 31976 24304 31976 24304 0 clknet_leaf_43_clk
rlabel metal2 26712 30688 26712 30688 0 clknet_leaf_44_clk
rlabel metal2 26600 29400 26600 29400 0 clknet_leaf_45_clk
rlabel metal2 23352 23576 23352 23576 0 clknet_leaf_46_clk
rlabel metal2 24920 22904 24920 22904 0 clknet_leaf_47_clk
rlabel metal2 21896 11172 21896 11172 0 clknet_leaf_48_clk
rlabel metal2 17640 16912 17640 16912 0 clknet_leaf_49_clk
rlabel metal2 15512 26180 15512 26180 0 clknet_leaf_4_clk
rlabel metal2 23240 40824 23240 40824 0 clknet_leaf_5_clk
rlabel metal2 17864 40544 17864 40544 0 clknet_leaf_6_clk
rlabel metal2 16632 51408 16632 51408 0 clknet_leaf_7_clk
rlabel metal2 15960 41664 15960 41664 0 clknet_leaf_8_clk
rlabel metal2 5656 49056 5656 49056 0 clknet_leaf_9_clk
rlabel metal2 11256 40152 11256 40152 0 net1
rlabel metal3 8624 41832 8624 41832 0 net10
rlabel metal2 45304 39816 45304 39816 0 net100
rlabel metal3 53816 40096 53816 40096 0 net101
rlabel metal2 43960 40432 43960 40432 0 net102
rlabel metal2 52696 40040 52696 40040 0 net103
rlabel metal2 53256 38416 53256 38416 0 net104
rlabel metal2 55496 40320 55496 40320 0 net105
rlabel metal2 19376 43400 19376 43400 0 net106
rlabel metal2 53256 41664 53256 41664 0 net107
rlabel metal2 4872 36736 4872 36736 0 net108
rlabel metal2 4872 43176 4872 43176 0 net109
rlabel metal3 2072 42168 2072 42168 0 net11
rlabel metal2 23128 33264 23128 33264 0 net110
rlabel metal2 23408 33992 23408 33992 0 net111
rlabel metal2 23800 30128 23800 30128 0 net112
rlabel metal2 27160 4536 27160 4536 0 net113
rlabel metal2 55496 38024 55496 38024 0 net114
rlabel metal2 52136 36008 52136 36008 0 net115
rlabel metal2 53256 35504 53256 35504 0 net116
rlabel metal2 17416 39984 17416 39984 0 net117
rlabel metal3 55440 33264 55440 33264 0 net118
rlabel metal2 2072 50568 2072 50568 0 net12
rlabel metal3 1848 53032 1848 53032 0 net13
rlabel metal2 10584 40320 10584 40320 0 net14
rlabel metal2 2072 42000 2072 42000 0 net15
rlabel metal2 9800 41496 9800 41496 0 net16
rlabel metal2 1960 45472 1960 45472 0 net17
rlabel metal3 2716 34664 2716 34664 0 net18
rlabel metal2 24920 9268 24920 9268 0 net19
rlabel metal2 3304 50848 3304 50848 0 net2
rlabel metal3 14952 3416 14952 3416 0 net20
rlabel metal2 2072 16856 2072 16856 0 net21
rlabel metal2 7448 18368 7448 18368 0 net22
rlabel metal3 7504 14504 7504 14504 0 net23
rlabel metal2 2072 18424 2072 18424 0 net24
rlabel metal2 9576 20440 9576 20440 0 net25
rlabel metal2 2128 22120 2128 22120 0 net26
rlabel metal2 2072 22792 2072 22792 0 net27
rlabel metal3 4536 23800 4536 23800 0 net28
rlabel metal2 2184 23968 2184 23968 0 net29
rlabel metal2 12600 44184 12600 44184 0 net3
rlabel metal3 19768 3416 19768 3416 0 net30
rlabel metal2 2072 25424 2072 25424 0 net31
rlabel metal2 2744 27272 2744 27272 0 net32
rlabel metal3 10416 24696 10416 24696 0 net33
rlabel metal2 2072 30296 2072 30296 0 net34
rlabel metal3 2744 30352 2744 30352 0 net35
rlabel metal2 2072 32088 2072 32088 0 net36
rlabel metal2 11816 32816 11816 32816 0 net37
rlabel metal2 11032 34944 11032 34944 0 net38
rlabel metal2 2184 36456 2184 36456 0 net39
rlabel metal2 2744 45024 2744 45024 0 net4
rlabel metal3 15428 38024 15428 38024 0 net40
rlabel metal3 18480 3416 18480 3416 0 net41
rlabel metal2 2744 36792 2744 36792 0 net42
rlabel metal3 2072 45528 2072 45528 0 net43
rlabel metal2 19040 14728 19040 14728 0 net44
rlabel metal2 18200 8960 18200 8960 0 net45
rlabel metal2 17024 3416 17024 3416 0 net46
rlabel metal2 16072 5908 16072 5908 0 net47
rlabel metal3 14280 21560 14280 21560 0 net48
rlabel metal2 2744 20944 2744 20944 0 net49
rlabel metal3 11592 40992 11592 40992 0 net5
rlabel metal2 2128 20552 2128 20552 0 net50
rlabel metal3 9408 29512 9408 29512 0 net51
rlabel metal2 30576 9800 30576 9800 0 net52
rlabel metal2 33432 10136 33432 10136 0 net53
rlabel metal2 34888 4200 34888 4200 0 net54
rlabel metal2 37128 3416 37128 3416 0 net55
rlabel metal2 39088 3416 39088 3416 0 net56
rlabel metal3 40824 9016 40824 9016 0 net57
rlabel metal2 41664 3416 41664 3416 0 net58
rlabel metal2 42952 5432 42952 5432 0 net59
rlabel metal2 2128 51912 2128 51912 0 net6
rlabel metal2 43456 5880 43456 5880 0 net60
rlabel metal2 44520 3416 44520 3416 0 net61
rlabel metal2 2072 28504 2072 28504 0 net62
rlabel metal2 53816 21000 53816 21000 0 net63
rlabel metal3 55440 23520 55440 23520 0 net64
rlabel metal3 57456 24920 57456 24920 0 net65
rlabel metal3 55440 25088 55440 25088 0 net66
rlabel metal2 40992 3416 40992 3416 0 net67
rlabel metal2 38024 19712 38024 19712 0 net68
rlabel metal2 37632 3416 37632 3416 0 net69
rlabel metal3 2128 50568 2128 50568 0 net7
rlabel metal3 36232 26264 36232 26264 0 net70
rlabel metal3 34440 24584 34440 24584 0 net71
rlabel metal2 30744 21280 30744 21280 0 net72
rlabel metal3 1960 26712 1960 26712 0 net73
rlabel metal2 29568 20776 29568 20776 0 net74
rlabel metal2 19208 43008 19208 43008 0 net75
rlabel metal2 2128 26488 2128 26488 0 net76
rlabel metal2 21392 3416 21392 3416 0 net77
rlabel metal2 20552 10136 20552 10136 0 net78
rlabel metal2 23688 8176 23688 8176 0 net79
rlabel metal2 2072 49560 2072 49560 0 net8
rlabel metal2 25816 6216 25816 6216 0 net80
rlabel metal2 27720 7784 27720 7784 0 net81
rlabel metal2 29848 8176 29848 8176 0 net82
rlabel metal2 2072 40376 2072 40376 0 net83
rlabel metal2 21784 46592 21784 46592 0 net84
rlabel metal2 53480 46592 53480 46592 0 net85
rlabel metal2 53368 30184 53368 30184 0 net86
rlabel metal2 55272 31696 55272 31696 0 net87
rlabel metal2 53480 33096 53480 33096 0 net88
rlabel metal3 53816 36960 53816 36960 0 net89
rlabel metal2 2576 48552 2576 48552 0 net9
rlabel metal3 53928 35112 53928 35112 0 net90
rlabel metal2 52696 34440 52696 34440 0 net91
rlabel metal2 50512 36344 50512 36344 0 net92
rlabel metal2 48552 37576 48552 37576 0 net93
rlabel metal3 51352 33992 51352 33992 0 net94
rlabel metal2 18536 46984 18536 46984 0 net95
rlabel metal2 51632 41160 51632 41160 0 net96
rlabel metal2 51688 40488 51688 40488 0 net97
rlabel metal3 51184 43736 51184 43736 0 net98
rlabel metal3 49952 40264 49952 40264 0 net99
rlabel metal3 1246 30968 1246 30968 0 pcpi_insn[0]
rlabel metal2 1736 54152 1736 54152 0 pcpi_insn[12]
rlabel metal2 1736 46536 1736 46536 0 pcpi_insn[13]
rlabel metal3 1582 45752 1582 45752 0 pcpi_insn[14]
rlabel metal3 1246 41048 1246 41048 0 pcpi_insn[1]
rlabel metal2 1736 51968 1736 51968 0 pcpi_insn[25]
rlabel metal3 1582 50456 1582 50456 0 pcpi_insn[26]
rlabel metal2 1736 49448 1736 49448 0 pcpi_insn[27]
rlabel metal2 1736 53368 1736 53368 0 pcpi_insn[28]
rlabel metal2 1736 43960 1736 43960 0 pcpi_insn[29]
rlabel metal2 1736 42504 1736 42504 0 pcpi_insn[2]
rlabel metal2 1848 50176 1848 50176 0 pcpi_insn[30]
rlabel metal2 1736 52696 1736 52696 0 pcpi_insn[31]
rlabel metal2 1736 39256 1736 39256 0 pcpi_insn[3]
rlabel metal2 1736 41832 1736 41832 0 pcpi_insn[4]
rlabel metal2 2408 40712 2408 40712 0 pcpi_insn[5]
rlabel metal2 1736 51240 1736 51240 0 pcpi_insn[6]
rlabel metal3 1358 48440 1358 48440 0 pcpi_mul_rd[0]
rlabel metal3 57330 46424 57330 46424 0 pcpi_mul_rd[10]
rlabel metal3 57330 30296 57330 30296 0 pcpi_mul_rd[11]
rlabel metal2 57960 30240 57960 30240 0 pcpi_mul_rd[12]
rlabel metal3 57330 32312 57330 32312 0 pcpi_mul_rd[13]
rlabel metal2 57960 37184 57960 37184 0 pcpi_mul_rd[14]
rlabel metal2 55272 35728 55272 35728 0 pcpi_mul_rd[15]
rlabel metal2 55048 31416 55048 31416 0 pcpi_mul_rd[16]
rlabel metal3 58618 32984 58618 32984 0 pcpi_mul_rd[17]
rlabel metal3 57330 37016 57330 37016 0 pcpi_mul_rd[18]
rlabel metal3 55412 33880 55412 33880 0 pcpi_mul_rd[19]
rlabel metal3 1358 47768 1358 47768 0 pcpi_mul_rd[1]
rlabel metal2 55048 45864 55048 45864 0 pcpi_mul_rd[20]
rlabel metal2 57848 45192 57848 45192 0 pcpi_mul_rd[21]
rlabel metal2 57960 44072 57960 44072 0 pcpi_mul_rd[22]
rlabel metal2 57960 46312 57960 46312 0 pcpi_mul_rd[23]
rlabel metal2 55384 39928 55384 39928 0 pcpi_mul_rd[24]
rlabel metal2 57960 43008 57960 43008 0 pcpi_mul_rd[25]
rlabel metal2 57960 40432 57960 40432 0 pcpi_mul_rd[26]
rlabel metal2 55048 40824 55048 40824 0 pcpi_mul_rd[27]
rlabel metal3 55412 38584 55412 38584 0 pcpi_mul_rd[28]
rlabel metal2 57960 41888 57960 41888 0 pcpi_mul_rd[29]
rlabel metal3 1358 47096 1358 47096 0 pcpi_mul_rd[2]
rlabel metal3 57330 41720 57330 41720 0 pcpi_mul_rd[30]
rlabel metal3 1358 36344 1358 36344 0 pcpi_mul_rd[31]
rlabel metal3 1358 43064 1358 43064 0 pcpi_mul_rd[3]
rlabel metal3 1358 31640 1358 31640 0 pcpi_mul_rd[4]
rlabel metal3 1358 33656 1358 33656 0 pcpi_mul_rd[5]
rlabel metal2 26264 2198 26264 2198 0 pcpi_mul_rd[6]
rlabel metal2 26936 2058 26936 2058 0 pcpi_mul_rd[7]
rlabel metal2 57960 38640 57960 38640 0 pcpi_mul_rd[8]
rlabel metal2 55048 36120 55048 36120 0 pcpi_mul_rd[9]
rlabel metal2 55384 35224 55384 35224 0 pcpi_mul_ready
rlabel metal2 1736 34552 1736 34552 0 pcpi_mul_valid
rlabel metal3 1358 38360 1358 38360 0 pcpi_mul_wait
rlabel metal2 57960 33936 57960 33936 0 pcpi_mul_wr
rlabel metal2 24584 2968 24584 2968 0 pcpi_rs1[0]
rlabel metal2 12768 3416 12768 3416 0 pcpi_rs1[10]
rlabel metal3 1302 16184 1302 16184 0 pcpi_rs1[11]
rlabel metal2 2408 17192 2408 17192 0 pcpi_rs1[12]
rlabel metal3 1246 17528 1246 17528 0 pcpi_rs1[13]
rlabel metal2 1736 18312 1736 18312 0 pcpi_rs1[14]
rlabel metal2 1736 19768 1736 19768 0 pcpi_rs1[15]
rlabel metal3 1246 22232 1246 22232 0 pcpi_rs1[16]
rlabel metal2 1736 23016 1736 23016 0 pcpi_rs1[17]
rlabel metal2 1736 23688 1736 23688 0 pcpi_rs1[18]
rlabel metal2 1736 24472 1736 24472 0 pcpi_rs1[19]
rlabel metal2 20216 2086 20216 2086 0 pcpi_rs1[1]
rlabel metal2 1736 25144 1736 25144 0 pcpi_rs1[20]
rlabel metal2 2408 26600 2408 26600 0 pcpi_rs1[21]
rlabel metal2 1736 27720 1736 27720 0 pcpi_rs1[22]
rlabel metal2 1736 29848 1736 29848 0 pcpi_rs1[23]
rlabel metal2 2408 30632 2408 30632 0 pcpi_rs1[24]
rlabel metal2 1736 32424 1736 32424 0 pcpi_rs1[25]
rlabel metal2 1736 33096 1736 33096 0 pcpi_rs1[26]
rlabel metal3 1246 35672 1246 35672 0 pcpi_rs1[27]
rlabel metal2 1736 37128 1736 37128 0 pcpi_rs1[28]
rlabel metal2 1736 37800 1736 37800 0 pcpi_rs1[29]
rlabel metal2 19544 2086 19544 2086 0 pcpi_rs1[2]
rlabel metal2 2408 35336 2408 35336 0 pcpi_rs1[30]
rlabel metal2 1848 45472 1848 45472 0 pcpi_rs1[31]
rlabel metal2 18648 3024 18648 3024 0 pcpi_rs1[3]
rlabel metal2 17976 3024 17976 3024 0 pcpi_rs1[4]
rlabel metal2 17304 3024 17304 3024 0 pcpi_rs1[5]
rlabel metal2 16240 3528 16240 3528 0 pcpi_rs1[6]
rlabel metal2 1736 21224 1736 21224 0 pcpi_rs1[7]
rlabel metal2 2408 22008 2408 22008 0 pcpi_rs1[8]
rlabel metal2 1736 20440 1736 20440 0 pcpi_rs1[9]
rlabel metal2 1736 29176 1736 29176 0 pcpi_rs2[0]
rlabel metal2 31248 2520 31248 2520 0 pcpi_rs2[10]
rlabel metal2 33096 3416 33096 3416 0 pcpi_rs2[11]
rlabel metal2 34440 3528 34440 3528 0 pcpi_rs2[12]
rlabel metal2 36512 2520 36512 2520 0 pcpi_rs2[13]
rlabel metal2 38472 2744 38472 2744 0 pcpi_rs2[14]
rlabel metal2 39816 3416 39816 3416 0 pcpi_rs2[15]
rlabel metal2 41272 2968 41272 2968 0 pcpi_rs2[16]
rlabel metal2 42392 2086 42392 2086 0 pcpi_rs2[17]
rlabel metal2 43064 2086 43064 2086 0 pcpi_rs2[18]
rlabel metal2 44296 2968 44296 2968 0 pcpi_rs2[19]
rlabel metal2 1736 28448 1736 28448 0 pcpi_rs2[1]
rlabel metal2 58184 21896 58184 21896 0 pcpi_rs2[20]
rlabel metal2 58184 23688 58184 23688 0 pcpi_rs2[21]
rlabel metal2 58184 24472 58184 24472 0 pcpi_rs2[22]
rlabel metal2 58184 25144 58184 25144 0 pcpi_rs2[23]
rlabel metal2 40488 3416 40488 3416 0 pcpi_rs2[24]
rlabel metal2 37968 2520 37968 2520 0 pcpi_rs2[25]
rlabel metal2 37184 2520 37184 2520 0 pcpi_rs2[26]
rlabel metal2 35840 3416 35840 3416 0 pcpi_rs2[27]
rlabel metal2 33768 3528 33768 3528 0 pcpi_rs2[28]
rlabel metal2 30520 4256 30520 4256 0 pcpi_rs2[29]
rlabel metal3 1246 26936 1246 26936 0 pcpi_rs2[2]
rlabel metal2 28952 2058 28952 2058 0 pcpi_rs2[30]
rlabel metal2 1736 44744 1736 44744 0 pcpi_rs2[31]
rlabel metal2 1736 25928 1736 25928 0 pcpi_rs2[3]
rlabel metal2 21000 3416 21000 3416 0 pcpi_rs2[4]
rlabel metal2 23240 3024 23240 3024 0 pcpi_rs2[5]
rlabel metal2 23912 3024 23912 3024 0 pcpi_rs2[6]
rlabel metal2 25592 2086 25592 2086 0 pcpi_rs2[7]
rlabel metal2 27608 3472 27608 3472 0 pcpi_rs2[8]
rlabel metal2 29624 2058 29624 2058 0 pcpi_rs2[9]
rlabel metal2 16072 40712 16072 40712 0 picorv32_pcpi_mul_inst_0.instr_any_mul
rlabel metal2 15456 41272 15456 41272 0 picorv32_pcpi_mul_inst_0.instr_mul
rlabel metal3 17472 45304 17472 45304 0 picorv32_pcpi_mul_inst_0.instr_mulh
rlabel metal2 18536 44240 18536 44240 0 picorv32_pcpi_mul_inst_0.instr_mulhsu
rlabel metal3 17528 43512 17528 43512 0 picorv32_pcpi_mul_inst_0.instr_mulhu
rlabel metal3 16072 31864 16072 31864 0 picorv32_pcpi_mul_inst_0.mul_counter\[0\]
rlabel metal2 16632 31416 16632 31416 0 picorv32_pcpi_mul_inst_0.mul_counter\[1\]
rlabel metal2 15624 31584 15624 31584 0 picorv32_pcpi_mul_inst_0.mul_counter\[2\]
rlabel metal2 17304 34888 17304 34888 0 picorv32_pcpi_mul_inst_0.mul_counter\[3\]
rlabel metal2 16520 35616 16520 35616 0 picorv32_pcpi_mul_inst_0.mul_counter\[4\]
rlabel metal2 18424 37744 18424 37744 0 picorv32_pcpi_mul_inst_0.mul_counter\[5\]
rlabel metal2 20160 39032 20160 39032 0 picorv32_pcpi_mul_inst_0.mul_counter\[6\]
rlabel metal2 24248 39536 24248 39536 0 picorv32_pcpi_mul_inst_0.mul_finish
rlabel metal2 20776 40600 20776 40600 0 picorv32_pcpi_mul_inst_0.mul_waiting
rlabel metal3 21392 21448 21392 21448 0 picorv32_pcpi_mul_inst_0.next_rs1\[0\]
rlabel metal2 17752 19376 17752 19376 0 picorv32_pcpi_mul_inst_0.next_rs1\[10\]
rlabel metal3 12320 19208 12320 19208 0 picorv32_pcpi_mul_inst_0.next_rs1\[11\]
rlabel metal3 11592 14504 11592 14504 0 picorv32_pcpi_mul_inst_0.next_rs1\[12\]
rlabel metal2 10360 14616 10360 14616 0 picorv32_pcpi_mul_inst_0.next_rs1\[13\]
rlabel metal3 10248 19880 10248 19880 0 picorv32_pcpi_mul_inst_0.next_rs1\[14\]
rlabel metal3 9688 20888 9688 20888 0 picorv32_pcpi_mul_inst_0.next_rs1\[15\]
rlabel metal2 8008 21952 8008 21952 0 picorv32_pcpi_mul_inst_0.next_rs1\[16\]
rlabel metal2 8120 23856 8120 23856 0 picorv32_pcpi_mul_inst_0.next_rs1\[17\]
rlabel metal3 9744 23912 9744 23912 0 picorv32_pcpi_mul_inst_0.next_rs1\[18\]
rlabel metal2 11256 23408 11256 23408 0 picorv32_pcpi_mul_inst_0.next_rs1\[19\]
rlabel metal2 19992 21000 19992 21000 0 picorv32_pcpi_mul_inst_0.next_rs1\[1\]
rlabel metal2 15848 26544 15848 26544 0 picorv32_pcpi_mul_inst_0.next_rs1\[20\]
rlabel metal2 14056 25788 14056 25788 0 picorv32_pcpi_mul_inst_0.next_rs1\[21\]
rlabel metal2 15176 28560 15176 28560 0 picorv32_pcpi_mul_inst_0.next_rs1\[22\]
rlabel metal2 12264 29344 12264 29344 0 picorv32_pcpi_mul_inst_0.next_rs1\[23\]
rlabel metal2 11928 30856 11928 30856 0 picorv32_pcpi_mul_inst_0.next_rs1\[24\]
rlabel metal2 11144 32872 11144 32872 0 picorv32_pcpi_mul_inst_0.next_rs1\[25\]
rlabel metal2 13048 33320 13048 33320 0 picorv32_pcpi_mul_inst_0.next_rs1\[26\]
rlabel metal2 12712 35560 12712 35560 0 picorv32_pcpi_mul_inst_0.next_rs1\[27\]
rlabel metal2 11928 37688 11928 37688 0 picorv32_pcpi_mul_inst_0.next_rs1\[28\]
rlabel metal3 13384 38696 13384 38696 0 picorv32_pcpi_mul_inst_0.next_rs1\[29\]
rlabel metal3 20440 18424 20440 18424 0 picorv32_pcpi_mul_inst_0.next_rs1\[2\]
rlabel metal3 11816 43736 11816 43736 0 picorv32_pcpi_mul_inst_0.next_rs1\[30\]
rlabel metal2 17416 48720 17416 48720 0 picorv32_pcpi_mul_inst_0.next_rs1\[31\]
rlabel metal3 17136 51464 17136 51464 0 picorv32_pcpi_mul_inst_0.next_rs1\[32\]
rlabel metal2 16016 51800 16016 51800 0 picorv32_pcpi_mul_inst_0.next_rs1\[33\]
rlabel metal2 15288 54992 15288 54992 0 picorv32_pcpi_mul_inst_0.next_rs1\[34\]
rlabel metal2 15176 56336 15176 56336 0 picorv32_pcpi_mul_inst_0.next_rs1\[35\]
rlabel metal2 17920 56952 17920 56952 0 picorv32_pcpi_mul_inst_0.next_rs1\[36\]
rlabel metal2 16856 59472 16856 59472 0 picorv32_pcpi_mul_inst_0.next_rs1\[37\]
rlabel metal2 17528 60704 17528 60704 0 picorv32_pcpi_mul_inst_0.next_rs1\[38\]
rlabel metal2 17528 63728 17528 63728 0 picorv32_pcpi_mul_inst_0.next_rs1\[39\]
rlabel metal2 20496 14504 20496 14504 0 picorv32_pcpi_mul_inst_0.next_rs1\[3\]
rlabel metal2 17472 66360 17472 66360 0 picorv32_pcpi_mul_inst_0.next_rs1\[40\]
rlabel metal2 15960 64680 15960 64680 0 picorv32_pcpi_mul_inst_0.next_rs1\[41\]
rlabel metal2 13944 65576 13944 65576 0 picorv32_pcpi_mul_inst_0.next_rs1\[42\]
rlabel metal2 13384 63728 13384 63728 0 picorv32_pcpi_mul_inst_0.next_rs1\[43\]
rlabel metal3 11256 62216 11256 62216 0 picorv32_pcpi_mul_inst_0.next_rs1\[44\]
rlabel metal2 12488 61208 12488 61208 0 picorv32_pcpi_mul_inst_0.next_rs1\[45\]
rlabel metal2 12488 58856 12488 58856 0 picorv32_pcpi_mul_inst_0.next_rs1\[46\]
rlabel metal2 11256 53984 11256 53984 0 picorv32_pcpi_mul_inst_0.next_rs1\[47\]
rlabel metal2 10360 56560 10360 56560 0 picorv32_pcpi_mul_inst_0.next_rs1\[48\]
rlabel metal2 9016 58296 9016 58296 0 picorv32_pcpi_mul_inst_0.next_rs1\[49\]
rlabel metal2 18984 16632 18984 16632 0 picorv32_pcpi_mul_inst_0.next_rs1\[4\]
rlabel metal2 8512 56168 8512 56168 0 picorv32_pcpi_mul_inst_0.next_rs1\[50\]
rlabel metal2 8008 55272 8008 55272 0 picorv32_pcpi_mul_inst_0.next_rs1\[51\]
rlabel metal2 7672 53704 7672 53704 0 picorv32_pcpi_mul_inst_0.next_rs1\[52\]
rlabel metal2 7784 51632 7784 51632 0 picorv32_pcpi_mul_inst_0.next_rs1\[53\]
rlabel metal2 8512 49112 8512 49112 0 picorv32_pcpi_mul_inst_0.next_rs1\[54\]
rlabel metal2 6328 48048 6328 48048 0 picorv32_pcpi_mul_inst_0.next_rs1\[55\]
rlabel metal2 8120 45248 8120 45248 0 picorv32_pcpi_mul_inst_0.next_rs1\[56\]
rlabel metal2 8624 44408 8624 44408 0 picorv32_pcpi_mul_inst_0.next_rs1\[57\]
rlabel metal2 9576 45360 9576 45360 0 picorv32_pcpi_mul_inst_0.next_rs1\[58\]
rlabel metal2 9576 46480 9576 46480 0 picorv32_pcpi_mul_inst_0.next_rs1\[59\]
rlabel metal2 17416 18088 17416 18088 0 picorv32_pcpi_mul_inst_0.next_rs1\[5\]
rlabel metal2 11816 47880 11816 47880 0 picorv32_pcpi_mul_inst_0.next_rs1\[60\]
rlabel metal2 12376 49756 12376 49756 0 picorv32_pcpi_mul_inst_0.next_rs1\[61\]
rlabel metal2 12936 48552 12936 48552 0 picorv32_pcpi_mul_inst_0.next_rs1\[62\]
rlabel metal2 16184 20272 16184 20272 0 picorv32_pcpi_mul_inst_0.next_rs1\[6\]
rlabel metal2 15792 20776 15792 20776 0 picorv32_pcpi_mul_inst_0.next_rs1\[7\]
rlabel metal2 15512 18648 15512 18648 0 picorv32_pcpi_mul_inst_0.next_rs1\[8\]
rlabel metal2 15064 18760 15064 18760 0 picorv32_pcpi_mul_inst_0.next_rs1\[9\]
rlabel metal3 30016 9800 30016 9800 0 picorv32_pcpi_mul_inst_0.next_rs2\[10\]
rlabel metal2 35112 14112 35112 14112 0 picorv32_pcpi_mul_inst_0.next_rs2\[11\]
rlabel metal2 35000 17920 35000 17920 0 picorv32_pcpi_mul_inst_0.next_rs2\[12\]
rlabel metal2 36456 13608 36456 13608 0 picorv32_pcpi_mul_inst_0.next_rs2\[13\]
rlabel metal2 39928 8372 39928 8372 0 picorv32_pcpi_mul_inst_0.next_rs2\[14\]
rlabel metal2 42168 11256 42168 11256 0 picorv32_pcpi_mul_inst_0.next_rs2\[15\]
rlabel metal2 43064 12544 43064 12544 0 picorv32_pcpi_mul_inst_0.next_rs2\[16\]
rlabel metal2 44520 14000 44520 14000 0 picorv32_pcpi_mul_inst_0.next_rs2\[17\]
rlabel metal2 44744 6664 44744 6664 0 picorv32_pcpi_mul_inst_0.next_rs2\[18\]
rlabel metal3 45752 7560 45752 7560 0 picorv32_pcpi_mul_inst_0.next_rs2\[19\]
rlabel metal3 23352 30184 23352 30184 0 picorv32_pcpi_mul_inst_0.next_rs2\[1\]
rlabel metal2 47320 11032 47320 11032 0 picorv32_pcpi_mul_inst_0.next_rs2\[20\]
rlabel metal3 46536 21560 46536 21560 0 picorv32_pcpi_mul_inst_0.next_rs2\[21\]
rlabel metal2 44408 24696 44408 24696 0 picorv32_pcpi_mul_inst_0.next_rs2\[22\]
rlabel metal3 42784 26264 42784 26264 0 picorv32_pcpi_mul_inst_0.next_rs2\[23\]
rlabel metal2 41496 23912 41496 23912 0 picorv32_pcpi_mul_inst_0.next_rs2\[24\]
rlabel metal3 40432 24024 40432 24024 0 picorv32_pcpi_mul_inst_0.next_rs2\[25\]
rlabel metal2 40488 22680 40488 22680 0 picorv32_pcpi_mul_inst_0.next_rs2\[26\]
rlabel metal2 39928 25312 39928 25312 0 picorv32_pcpi_mul_inst_0.next_rs2\[27\]
rlabel metal2 33488 22456 33488 22456 0 picorv32_pcpi_mul_inst_0.next_rs2\[28\]
rlabel metal2 34888 24752 34888 24752 0 picorv32_pcpi_mul_inst_0.next_rs2\[29\]
rlabel metal2 23240 28616 23240 28616 0 picorv32_pcpi_mul_inst_0.next_rs2\[2\]
rlabel metal3 29568 23016 29568 23016 0 picorv32_pcpi_mul_inst_0.next_rs2\[30\]
rlabel metal2 20216 43960 20216 43960 0 picorv32_pcpi_mul_inst_0.next_rs2\[31\]
rlabel metal2 18312 52080 18312 52080 0 picorv32_pcpi_mul_inst_0.next_rs2\[32\]
rlabel metal3 21672 56056 21672 56056 0 picorv32_pcpi_mul_inst_0.next_rs2\[33\]
rlabel metal2 20664 51240 20664 51240 0 picorv32_pcpi_mul_inst_0.next_rs2\[34\]
rlabel metal2 20216 61320 20216 61320 0 picorv32_pcpi_mul_inst_0.next_rs2\[35\]
rlabel metal3 21560 63112 21560 63112 0 picorv32_pcpi_mul_inst_0.next_rs2\[36\]
rlabel metal2 23576 59948 23576 59948 0 picorv32_pcpi_mul_inst_0.next_rs2\[37\]
rlabel metal3 20888 67816 20888 67816 0 picorv32_pcpi_mul_inst_0.next_rs2\[38\]
rlabel metal2 24696 69160 24696 69160 0 picorv32_pcpi_mul_inst_0.next_rs2\[39\]
rlabel metal2 23576 26852 23576 26852 0 picorv32_pcpi_mul_inst_0.next_rs2\[3\]
rlabel metal3 28784 67144 28784 67144 0 picorv32_pcpi_mul_inst_0.next_rs2\[40\]
rlabel metal2 33432 66752 33432 66752 0 picorv32_pcpi_mul_inst_0.next_rs2\[41\]
rlabel metal2 30912 66136 30912 66136 0 picorv32_pcpi_mul_inst_0.next_rs2\[42\]
rlabel metal2 34104 63280 34104 63280 0 picorv32_pcpi_mul_inst_0.next_rs2\[43\]
rlabel metal2 35896 64512 35896 64512 0 picorv32_pcpi_mul_inst_0.next_rs2\[44\]
rlabel metal2 39424 70056 39424 70056 0 picorv32_pcpi_mul_inst_0.next_rs2\[45\]
rlabel metal2 40264 58576 40264 58576 0 picorv32_pcpi_mul_inst_0.next_rs2\[46\]
rlabel metal2 43848 70112 43848 70112 0 picorv32_pcpi_mul_inst_0.next_rs2\[47\]
rlabel metal2 41496 69160 41496 69160 0 picorv32_pcpi_mul_inst_0.next_rs2\[48\]
rlabel metal2 47936 65464 47936 65464 0 picorv32_pcpi_mul_inst_0.next_rs2\[49\]
rlabel metal2 20776 13664 20776 13664 0 picorv32_pcpi_mul_inst_0.next_rs2\[4\]
rlabel metal2 44688 65576 44688 65576 0 picorv32_pcpi_mul_inst_0.next_rs2\[50\]
rlabel metal3 42336 67144 42336 67144 0 picorv32_pcpi_mul_inst_0.next_rs2\[51\]
rlabel metal2 45920 63784 45920 63784 0 picorv32_pcpi_mul_inst_0.next_rs2\[52\]
rlabel metal2 48104 55216 48104 55216 0 picorv32_pcpi_mul_inst_0.next_rs2\[53\]
rlabel metal2 45976 53144 45976 53144 0 picorv32_pcpi_mul_inst_0.next_rs2\[54\]
rlabel metal3 42280 48776 42280 48776 0 picorv32_pcpi_mul_inst_0.next_rs2\[55\]
rlabel metal2 43848 46368 43848 46368 0 picorv32_pcpi_mul_inst_0.next_rs2\[56\]
rlabel metal2 36792 51184 36792 51184 0 picorv32_pcpi_mul_inst_0.next_rs2\[57\]
rlabel metal2 39480 53704 39480 53704 0 picorv32_pcpi_mul_inst_0.next_rs2\[58\]
rlabel metal2 34664 53760 34664 53760 0 picorv32_pcpi_mul_inst_0.next_rs2\[59\]
rlabel metal2 22680 13944 22680 13944 0 picorv32_pcpi_mul_inst_0.next_rs2\[5\]
rlabel metal3 34552 46760 34552 46760 0 picorv32_pcpi_mul_inst_0.next_rs2\[60\]
rlabel metal2 31360 51240 31360 51240 0 picorv32_pcpi_mul_inst_0.next_rs2\[61\]
rlabel metal2 29400 45808 29400 45808 0 picorv32_pcpi_mul_inst_0.next_rs2\[62\]
rlabel metal2 27216 53144 27216 53144 0 picorv32_pcpi_mul_inst_0.next_rs2\[63\]
rlabel metal2 24696 10976 24696 10976 0 picorv32_pcpi_mul_inst_0.next_rs2\[6\]
rlabel metal2 25480 13496 25480 13496 0 picorv32_pcpi_mul_inst_0.next_rs2\[7\]
rlabel metal2 26264 21392 26264 21392 0 picorv32_pcpi_mul_inst_0.next_rs2\[8\]
rlabel metal2 29960 15260 29960 15260 0 picorv32_pcpi_mul_inst_0.next_rs2\[9\]
rlabel metal2 18984 39760 18984 39760 0 picorv32_pcpi_mul_inst_0.pcpi_wait_q
rlabel metal2 22848 37352 22848 37352 0 picorv32_pcpi_mul_inst_0.rd\[0\]
rlabel metal2 35112 13328 35112 13328 0 picorv32_pcpi_mul_inst_0.rd\[10\]
rlabel metal2 33992 18032 33992 18032 0 picorv32_pcpi_mul_inst_0.rd\[11\]
rlabel metal2 38696 17640 38696 17640 0 picorv32_pcpi_mul_inst_0.rd\[12\]
rlabel metal2 40544 11256 40544 11256 0 picorv32_pcpi_mul_inst_0.rd\[13\]
rlabel metal2 44688 23576 44688 23576 0 picorv32_pcpi_mul_inst_0.rd\[14\]
rlabel metal3 41832 21784 41832 21784 0 picorv32_pcpi_mul_inst_0.rd\[15\]
rlabel metal2 45864 16520 45864 16520 0 picorv32_pcpi_mul_inst_0.rd\[16\]
rlabel metal2 49448 13160 49448 13160 0 picorv32_pcpi_mul_inst_0.rd\[17\]
rlabel metal2 50792 14952 50792 14952 0 picorv32_pcpi_mul_inst_0.rd\[18\]
rlabel metal2 48328 20944 48328 20944 0 picorv32_pcpi_mul_inst_0.rd\[19\]
rlabel metal2 22344 31192 22344 31192 0 picorv32_pcpi_mul_inst_0.rd\[1\]
rlabel metal2 50680 23800 50680 23800 0 picorv32_pcpi_mul_inst_0.rd\[20\]
rlabel metal2 50456 28952 50456 28952 0 picorv32_pcpi_mul_inst_0.rd\[21\]
rlabel metal2 50568 31696 50568 31696 0 picorv32_pcpi_mul_inst_0.rd\[22\]
rlabel metal2 44184 32760 44184 32760 0 picorv32_pcpi_mul_inst_0.rd\[23\]
rlabel metal3 40824 27832 40824 27832 0 picorv32_pcpi_mul_inst_0.rd\[24\]
rlabel metal3 43624 31864 43624 31864 0 picorv32_pcpi_mul_inst_0.rd\[25\]
rlabel metal2 40376 33264 40376 33264 0 picorv32_pcpi_mul_inst_0.rd\[26\]
rlabel metal2 38360 34328 38360 34328 0 picorv32_pcpi_mul_inst_0.rd\[27\]
rlabel metal3 36456 28616 36456 28616 0 picorv32_pcpi_mul_inst_0.rd\[28\]
rlabel metal2 31080 32424 31080 32424 0 picorv32_pcpi_mul_inst_0.rd\[29\]
rlabel metal2 22008 28056 22008 28056 0 picorv32_pcpi_mul_inst_0.rd\[2\]
rlabel metal2 30464 36680 30464 36680 0 picorv32_pcpi_mul_inst_0.rd\[30\]
rlabel metal2 27664 34888 27664 34888 0 picorv32_pcpi_mul_inst_0.rd\[31\]
rlabel metal3 25368 54712 25368 54712 0 picorv32_pcpi_mul_inst_0.rd\[32\]
rlabel metal3 21448 50568 21448 50568 0 picorv32_pcpi_mul_inst_0.rd\[33\]
rlabel metal2 21448 55384 21448 55384 0 picorv32_pcpi_mul_inst_0.rd\[34\]
rlabel metal2 25256 59472 25256 59472 0 picorv32_pcpi_mul_inst_0.rd\[35\]
rlabel metal2 24696 58464 24696 58464 0 picorv32_pcpi_mul_inst_0.rd\[36\]
rlabel metal3 23632 59192 23632 59192 0 picorv32_pcpi_mul_inst_0.rd\[37\]
rlabel metal2 26096 53256 26096 53256 0 picorv32_pcpi_mul_inst_0.rd\[38\]
rlabel metal2 14616 63112 14616 63112 0 picorv32_pcpi_mul_inst_0.rd\[39\]
rlabel metal2 22680 24192 22680 24192 0 picorv32_pcpi_mul_inst_0.rd\[3\]
rlabel metal2 35112 60816 35112 60816 0 picorv32_pcpi_mul_inst_0.rd\[40\]
rlabel metal2 52136 51520 52136 51520 0 picorv32_pcpi_mul_inst_0.rd\[41\]
rlabel metal2 35000 43680 35000 43680 0 picorv32_pcpi_mul_inst_0.rd\[42\]
rlabel metal2 36288 42728 36288 42728 0 picorv32_pcpi_mul_inst_0.rd\[43\]
rlabel metal2 38696 61096 38696 61096 0 picorv32_pcpi_mul_inst_0.rd\[44\]
rlabel metal2 52248 50736 52248 50736 0 picorv32_pcpi_mul_inst_0.rd\[45\]
rlabel metal2 42224 46312 42224 46312 0 picorv32_pcpi_mul_inst_0.rd\[46\]
rlabel metal3 41160 44184 41160 44184 0 picorv32_pcpi_mul_inst_0.rd\[47\]
rlabel metal2 50232 61208 50232 61208 0 picorv32_pcpi_mul_inst_0.rd\[48\]
rlabel metal2 47880 49560 47880 49560 0 picorv32_pcpi_mul_inst_0.rd\[49\]
rlabel metal2 24248 17304 24248 17304 0 picorv32_pcpi_mul_inst_0.rd\[4\]
rlabel metal2 46760 47208 46760 47208 0 picorv32_pcpi_mul_inst_0.rd\[50\]
rlabel metal2 46424 45920 46424 45920 0 picorv32_pcpi_mul_inst_0.rd\[51\]
rlabel metal2 48776 53648 48776 53648 0 picorv32_pcpi_mul_inst_0.rd\[52\]
rlabel metal2 47096 43596 47096 43596 0 picorv32_pcpi_mul_inst_0.rd\[53\]
rlabel metal2 48216 46928 48216 46928 0 picorv32_pcpi_mul_inst_0.rd\[54\]
rlabel metal2 45080 46648 45080 46648 0 picorv32_pcpi_mul_inst_0.rd\[55\]
rlabel metal3 37296 50008 37296 50008 0 picorv32_pcpi_mul_inst_0.rd\[56\]
rlabel metal2 41608 47880 41608 47880 0 picorv32_pcpi_mul_inst_0.rd\[57\]
rlabel metal3 40712 48104 40712 48104 0 picorv32_pcpi_mul_inst_0.rd\[58\]
rlabel metal2 37800 44912 37800 44912 0 picorv32_pcpi_mul_inst_0.rd\[59\]
rlabel metal2 24696 13664 24696 13664 0 picorv32_pcpi_mul_inst_0.rd\[5\]
rlabel metal3 32704 48216 32704 48216 0 picorv32_pcpi_mul_inst_0.rd\[60\]
rlabel metal2 28504 42728 28504 42728 0 picorv32_pcpi_mul_inst_0.rd\[61\]
rlabel metal2 28728 46480 28728 46480 0 picorv32_pcpi_mul_inst_0.rd\[62\]
rlabel metal3 25760 37240 25760 37240 0 picorv32_pcpi_mul_inst_0.rd\[63\]
rlabel metal2 23352 16744 23352 16744 0 picorv32_pcpi_mul_inst_0.rd\[6\]
rlabel metal2 25704 23016 25704 23016 0 picorv32_pcpi_mul_inst_0.rd\[7\]
rlabel metal2 31976 17248 31976 17248 0 picorv32_pcpi_mul_inst_0.rd\[8\]
rlabel metal2 32760 17304 32760 17304 0 picorv32_pcpi_mul_inst_0.rd\[9\]
rlabel metal2 37240 19320 37240 19320 0 picorv32_pcpi_mul_inst_0.rdx\[12\]
rlabel metal2 45640 16352 45640 16352 0 picorv32_pcpi_mul_inst_0.rdx\[16\]
rlabel metal2 50344 23856 50344 23856 0 picorv32_pcpi_mul_inst_0.rdx\[20\]
rlabel metal3 41272 27048 41272 27048 0 picorv32_pcpi_mul_inst_0.rdx\[24\]
rlabel metal3 35280 28616 35280 28616 0 picorv32_pcpi_mul_inst_0.rdx\[28\]
rlabel metal2 29288 55608 29288 55608 0 picorv32_pcpi_mul_inst_0.rdx\[32\]
rlabel metal2 28616 57288 28616 57288 0 picorv32_pcpi_mul_inst_0.rdx\[36\]
rlabel metal2 31976 59136 31976 59136 0 picorv32_pcpi_mul_inst_0.rdx\[40\]
rlabel metal2 36456 57736 36456 57736 0 picorv32_pcpi_mul_inst_0.rdx\[44\]
rlabel metal2 48216 63112 48216 63112 0 picorv32_pcpi_mul_inst_0.rdx\[48\]
rlabel metal2 24696 20720 24696 20720 0 picorv32_pcpi_mul_inst_0.rdx\[4\]
rlabel metal2 50456 49056 50456 49056 0 picorv32_pcpi_mul_inst_0.rdx\[52\]
rlabel metal2 43400 46144 43400 46144 0 picorv32_pcpi_mul_inst_0.rdx\[56\]
rlabel metal3 33768 44408 33768 44408 0 picorv32_pcpi_mul_inst_0.rdx\[60\]
rlabel metal2 30632 21504 30632 21504 0 picorv32_pcpi_mul_inst_0.rdx\[8\]
rlabel metal2 28224 25480 28224 25480 0 picorv32_pcpi_mul_inst_0.rs1\[0\]
rlabel metal2 26544 50568 26544 50568 0 picorv32_pcpi_mul_inst_0.rs2\[63\]
rlabel metal2 1736 40040 1736 40040 0 resetn
<< properties >>
string FIXED_BBOX 0 0 60000 80000
<< end >>

magic
tech gf180mcuD
magscale 1 5
timestamp 1702206233
<< obsm1 >>
rect 672 1538 24304 23158
<< metal2 >>
rect 12096 0 12152 400
rect 12432 0 12488 400
rect 12768 0 12824 400
<< obsm2 >>
rect 2238 430 24122 23147
rect 2238 400 12066 430
rect 12182 400 12402 430
rect 12518 400 12738 430
rect 12854 400 24122 430
<< metal3 >>
rect 24600 12768 25000 12824
rect 0 12432 400 12488
rect 24600 12432 25000 12488
rect 24600 12096 25000 12152
rect 24600 11760 25000 11816
<< obsm3 >>
rect 400 12854 24600 23142
rect 400 12738 24570 12854
rect 400 12518 24600 12738
rect 430 12402 24570 12518
rect 400 12182 24600 12402
rect 400 12066 24570 12182
rect 400 11846 24600 12066
rect 400 11730 24570 11846
rect 400 1554 24600 11730
<< metal4 >>
rect 2224 1538 2384 23158
rect 9904 1538 10064 23158
rect 17584 1538 17744 23158
<< labels >>
rlabel metal3 s 0 12432 400 12488 6 ctrl_in[0]
port 1 nsew signal input
rlabel metal3 s 24600 11760 25000 11816 6 ctrl_in[1]
port 2 nsew signal input
rlabel metal2 s 12432 0 12488 400 6 ctrl_oeb[0]
port 3 nsew signal output
rlabel metal3 s 24600 12768 25000 12824 6 ctrl_oeb[1]
port 4 nsew signal output
rlabel metal2 s 12768 0 12824 400 6 ctrl_out[0]
port 5 nsew signal output
rlabel metal2 s 12096 0 12152 400 6 ctrl_out[1]
port 6 nsew signal output
rlabel metal3 s 24600 12096 25000 12152 6 reset
port 7 nsew signal output
rlabel metal3 s 24600 12432 25000 12488 6 resetn
port 8 nsew signal output
rlabel metal4 s 2224 1538 2384 23158 6 vdd
port 9 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 23158 6 vdd
port 9 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 23158 6 vss
port 10 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 25000 25000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 284648
string GDS_FILE /home/luke/picosoc-w-approximation/openlane/ctrl/runs/23_12_10_12_01/results/signoff/ctrl.magic.gds
string GDS_START 95060
<< end >>


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO spimemio
  CLASS BLOCK ;
  FOREIGN spimemio ;
  ORIGIN 0.000 0.000 ;
  SIZE 250.000 BY 250.000 ;
  PIN addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 127.680 4.000 128.240 ;
    END
  END addr[0]
  PIN addr[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 67.200 246.000 67.760 250.000 ;
    END
  END addr[10]
  PIN addr[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 201.600 4.000 202.160 ;
    END
  END addr[11]
  PIN addr[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 178.080 4.000 178.640 ;
    END
  END addr[12]
  PIN addr[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 161.280 4.000 161.840 ;
    END
  END addr[13]
  PIN addr[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 154.560 4.000 155.120 ;
    END
  END addr[14]
  PIN addr[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 191.520 4.000 192.080 ;
    END
  END addr[15]
  PIN addr[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 198.240 4.000 198.800 ;
    END
  END addr[16]
  PIN addr[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 164.640 4.000 165.200 ;
    END
  END addr[17]
  PIN addr[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 174.720 4.000 175.280 ;
    END
  END addr[18]
  PIN addr[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 124.320 4.000 124.880 ;
    END
  END addr[19]
  PIN addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 117.600 4.000 118.160 ;
    END
  END addr[1]
  PIN addr[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 141.120 4.000 141.680 ;
    END
  END addr[20]
  PIN addr[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 168.000 4.000 168.560 ;
    END
  END addr[21]
  PIN addr[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 157.920 4.000 158.480 ;
    END
  END addr[22]
  PIN addr[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 151.200 4.000 151.760 ;
    END
  END addr[23]
  PIN addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 144.480 4.000 145.040 ;
    END
  END addr[2]
  PIN addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 131.040 4.000 131.600 ;
    END
  END addr[3]
  PIN addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 137.760 4.000 138.320 ;
    END
  END addr[4]
  PIN addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 114.240 246.000 114.800 250.000 ;
    END
  END addr[5]
  PIN addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 90.720 246.000 91.280 250.000 ;
    END
  END addr[6]
  PIN addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 100.800 246.000 101.360 250.000 ;
    END
  END addr[7]
  PIN addr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 188.160 4.000 188.720 ;
    END
  END addr[8]
  PIN addr[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 73.920 246.000 74.480 250.000 ;
    END
  END addr[9]
  PIN cfgreg_di[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 168.000 0.000 168.560 4.000 ;
    END
  END cfgreg_di[0]
  PIN cfgreg_di[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 218.400 0.000 218.960 4.000 ;
    END
  END cfgreg_di[10]
  PIN cfgreg_di[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 225.120 0.000 225.680 4.000 ;
    END
  END cfgreg_di[11]
  PIN cfgreg_di[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 16.800 0.000 17.360 4.000 ;
    END
  END cfgreg_di[12]
  PIN cfgreg_di[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 10.080 0.000 10.640 4.000 ;
    END
  END cfgreg_di[13]
  PIN cfgreg_di[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 13.440 0.000 14.000 4.000 ;
    END
  END cfgreg_di[14]
  PIN cfgreg_di[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 100.800 0.000 101.360 4.000 ;
    END
  END cfgreg_di[15]
  PIN cfgreg_di[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 53.760 0.000 54.320 4.000 ;
    END
  END cfgreg_di[16]
  PIN cfgreg_di[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 63.840 0.000 64.400 4.000 ;
    END
  END cfgreg_di[17]
  PIN cfgreg_di[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 60.480 0.000 61.040 4.000 ;
    END
  END cfgreg_di[18]
  PIN cfgreg_di[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 70.560 0.000 71.120 4.000 ;
    END
  END cfgreg_di[19]
  PIN cfgreg_di[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 110.880 0.000 111.440 4.000 ;
    END
  END cfgreg_di[1]
  PIN cfgreg_di[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 33.600 0.000 34.160 4.000 ;
    END
  END cfgreg_di[20]
  PIN cfgreg_di[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 36.960 0.000 37.520 4.000 ;
    END
  END cfgreg_di[21]
  PIN cfgreg_di[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 84.000 0.000 84.560 4.000 ;
    END
  END cfgreg_di[22]
  PIN cfgreg_di[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 20.160 0.000 20.720 4.000 ;
    END
  END cfgreg_di[23]
  PIN cfgreg_di[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 23.520 0.000 24.080 4.000 ;
    END
  END cfgreg_di[24]
  PIN cfgreg_di[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 26.880 0.000 27.440 4.000 ;
    END
  END cfgreg_di[25]
  PIN cfgreg_di[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 30.240 0.000 30.800 4.000 ;
    END
  END cfgreg_di[26]
  PIN cfgreg_di[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 90.720 0.000 91.280 4.000 ;
    END
  END cfgreg_di[27]
  PIN cfgreg_di[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 40.320 0.000 40.880 4.000 ;
    END
  END cfgreg_di[28]
  PIN cfgreg_di[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3.360 0.000 3.920 4.000 ;
    END
  END cfgreg_di[29]
  PIN cfgreg_di[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 124.320 0.000 124.880 4.000 ;
    END
  END cfgreg_di[2]
  PIN cfgreg_di[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 97.440 0.000 98.000 4.000 ;
    END
  END cfgreg_di[30]
  PIN cfgreg_di[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 117.600 0.000 118.160 4.000 ;
    END
  END cfgreg_di[31]
  PIN cfgreg_di[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 151.200 0.000 151.760 4.000 ;
    END
  END cfgreg_di[3]
  PIN cfgreg_di[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 178.080 0.000 178.640 4.000 ;
    END
  END cfgreg_di[4]
  PIN cfgreg_di[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 157.920 0.000 158.480 4.000 ;
    END
  END cfgreg_di[5]
  PIN cfgreg_di[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 43.680 0.000 44.240 4.000 ;
    END
  END cfgreg_di[6]
  PIN cfgreg_di[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 6.720 0.000 7.280 4.000 ;
    END
  END cfgreg_di[7]
  PIN cfgreg_di[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 215.040 0.000 215.600 4.000 ;
    END
  END cfgreg_di[8]
  PIN cfgreg_di[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 211.680 0.000 212.240 4.000 ;
    END
  END cfgreg_di[9]
  PIN cfgreg_do[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 127.680 250.000 128.240 ;
    END
  END cfgreg_do[0]
  PIN cfgreg_do[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 36.960 250.000 37.520 ;
    END
  END cfgreg_do[10]
  PIN cfgreg_do[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 47.040 250.000 47.600 ;
    END
  END cfgreg_do[11]
  PIN cfgreg_do[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 26.880 4.000 27.440 ;
    END
  END cfgreg_do[12]
  PIN cfgreg_do[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 13.440 4.000 14.000 ;
    END
  END cfgreg_do[13]
  PIN cfgreg_do[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 221.760 250.000 222.320 ;
    END
  END cfgreg_do[14]
  PIN cfgreg_do[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 20.160 4.000 20.720 ;
    END
  END cfgreg_do[15]
  PIN cfgreg_do[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 57.120 0.000 57.680 4.000 ;
    END
  END cfgreg_do[16]
  PIN cfgreg_do[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 73.920 0.000 74.480 4.000 ;
    END
  END cfgreg_do[17]
  PIN cfgreg_do[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 67.200 0.000 67.760 4.000 ;
    END
  END cfgreg_do[18]
  PIN cfgreg_do[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 80.640 0.000 81.200 4.000 ;
    END
  END cfgreg_do[19]
  PIN cfgreg_do[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 117.600 250.000 118.160 ;
    END
  END cfgreg_do[1]
  PIN cfgreg_do[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 87.360 4.000 87.920 ;
    END
  END cfgreg_do[20]
  PIN cfgreg_do[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 47.040 0.000 47.600 4.000 ;
    END
  END cfgreg_do[21]
  PIN cfgreg_do[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 87.360 0.000 87.920 4.000 ;
    END
  END cfgreg_do[22]
  PIN cfgreg_do[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 23.520 250.000 24.080 ;
    END
  END cfgreg_do[23]
  PIN cfgreg_do[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 218.400 250.000 218.960 ;
    END
  END cfgreg_do[24]
  PIN cfgreg_do[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 225.120 250.000 225.680 ;
    END
  END cfgreg_do[25]
  PIN cfgreg_do[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 20.160 250.000 20.720 ;
    END
  END cfgreg_do[26]
  PIN cfgreg_do[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 16.800 250.000 17.360 ;
    END
  END cfgreg_do[27]
  PIN cfgreg_do[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 231.840 250.000 232.400 ;
    END
  END cfgreg_do[28]
  PIN cfgreg_do[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 215.040 250.000 215.600 ;
    END
  END cfgreg_do[29]
  PIN cfgreg_do[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 110.880 250.000 111.440 ;
    END
  END cfgreg_do[2]
  PIN cfgreg_do[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 16.800 4.000 17.360 ;
    END
  END cfgreg_do[30]
  PIN cfgreg_do[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 134.400 0.000 134.960 4.000 ;
    END
  END cfgreg_do[31]
  PIN cfgreg_do[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 100.800 250.000 101.360 ;
    END
  END cfgreg_do[3]
  PIN cfgreg_do[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 184.800 0.000 185.360 4.000 ;
    END
  END cfgreg_do[4]
  PIN cfgreg_do[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 191.520 0.000 192.080 4.000 ;
    END
  END cfgreg_do[5]
  PIN cfgreg_do[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 211.680 250.000 212.240 ;
    END
  END cfgreg_do[6]
  PIN cfgreg_do[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 225.120 4.000 225.680 ;
    END
  END cfgreg_do[7]
  PIN cfgreg_do[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 204.960 0.000 205.520 4.000 ;
    END
  END cfgreg_do[8]
  PIN cfgreg_do[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 208.320 0.000 208.880 4.000 ;
    END
  END cfgreg_do[9]
  PIN cfgreg_we[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 154.560 0.000 155.120 4.000 ;
    END
  END cfgreg_we[0]
  PIN cfgreg_we[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 221.760 0.000 222.320 4.000 ;
    END
  END cfgreg_we[1]
  PIN cfgreg_we[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 50.400 0.000 50.960 4.000 ;
    END
  END cfgreg_we[2]
  PIN cfgreg_we[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 114.240 0.000 114.800 4.000 ;
    END
  END cfgreg_we[3]
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.738000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 221.760 4.000 222.320 ;
    END
  END clk
  PIN flash_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 0.000 0.560 4.000 ;
    END
  END flash_in[0]
  PIN flash_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 77.280 0.000 77.840 4.000 ;
    END
  END flash_in[1]
  PIN flash_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 124.320 250.000 124.880 ;
    END
  END flash_in[2]
  PIN flash_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 120.960 250.000 121.520 ;
    END
  END flash_in[3]
  PIN flash_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 107.520 250.000 108.080 ;
    END
  END flash_in[4]
  PIN flash_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 104.160 250.000 104.720 ;
    END
  END flash_in[5]
  PIN flash_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 228.480 250.000 229.040 ;
    END
  END flash_oeb[0]
  PIN flash_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 23.520 4.000 24.080 ;
    END
  END flash_oeb[1]
  PIN flash_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 201.600 0.000 202.160 4.000 ;
    END
  END flash_oeb[2]
  PIN flash_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 198.240 0.000 198.800 4.000 ;
    END
  END flash_oeb[3]
  PIN flash_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 40.320 250.000 40.880 ;
    END
  END flash_oeb[4]
  PIN flash_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 43.680 250.000 44.240 ;
    END
  END flash_oeb[5]
  PIN flash_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 194.880 0.000 195.440 4.000 ;
    END
  END flash_out[0]
  PIN flash_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 188.160 0.000 188.720 4.000 ;
    END
  END flash_out[1]
  PIN flash_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 164.640 0.000 165.200 4.000 ;
    END
  END flash_out[2]
  PIN flash_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 104.160 0.000 104.720 4.000 ;
    END
  END flash_out[3]
  PIN flash_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 131.040 0.000 131.600 4.000 ;
    END
  END flash_out[4]
  PIN flash_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 147.840 0.000 148.400 4.000 ;
    END
  END flash_out[5]
  PIN rdata[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 117.600 246.000 118.160 250.000 ;
    END
  END rdata[0]
  PIN rdata[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 191.520 246.000 192.080 250.000 ;
    END
  END rdata[10]
  PIN rdata[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 198.240 246.000 198.800 250.000 ;
    END
  END rdata[11]
  PIN rdata[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 198.240 250.000 198.800 ;
    END
  END rdata[12]
  PIN rdata[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 194.880 250.000 195.440 ;
    END
  END rdata[13]
  PIN rdata[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 174.720 246.000 175.280 250.000 ;
    END
  END rdata[14]
  PIN rdata[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 188.160 246.000 188.720 250.000 ;
    END
  END rdata[15]
  PIN rdata[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 168.000 246.000 168.560 250.000 ;
    END
  END rdata[16]
  PIN rdata[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 181.440 246.000 182.000 250.000 ;
    END
  END rdata[17]
  PIN rdata[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 208.320 250.000 208.880 ;
    END
  END rdata[18]
  PIN rdata[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 221.760 246.000 222.320 250.000 ;
    END
  END rdata[19]
  PIN rdata[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 131.040 246.000 131.600 250.000 ;
    END
  END rdata[1]
  PIN rdata[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 201.600 250.000 202.160 ;
    END
  END rdata[20]
  PIN rdata[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 174.720 250.000 175.280 ;
    END
  END rdata[21]
  PIN rdata[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 151.200 246.000 151.760 250.000 ;
    END
  END rdata[22]
  PIN rdata[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 157.920 246.000 158.480 250.000 ;
    END
  END rdata[23]
  PIN rdata[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 164.640 246.000 165.200 250.000 ;
    END
  END rdata[24]
  PIN rdata[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 161.280 246.000 161.840 250.000 ;
    END
  END rdata[25]
  PIN rdata[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 168.000 250.000 168.560 ;
    END
  END rdata[26]
  PIN rdata[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 161.280 250.000 161.840 ;
    END
  END rdata[27]
  PIN rdata[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 157.920 250.000 158.480 ;
    END
  END rdata[28]
  PIN rdata[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 171.360 250.000 171.920 ;
    END
  END rdata[29]
  PIN rdata[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 147.840 250.000 148.400 ;
    END
  END rdata[2]
  PIN rdata[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 154.560 246.000 155.120 250.000 ;
    END
  END rdata[30]
  PIN rdata[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 154.560 250.000 155.120 ;
    END
  END rdata[31]
  PIN rdata[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 144.480 250.000 145.040 ;
    END
  END rdata[3]
  PIN rdata[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 114.240 250.000 114.800 ;
    END
  END rdata[4]
  PIN rdata[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 151.200 250.000 151.760 ;
    END
  END rdata[5]
  PIN rdata[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 137.760 250.000 138.320 ;
    END
  END rdata[6]
  PIN rdata[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 246.000 141.120 250.000 141.680 ;
    END
  END rdata[7]
  PIN rdata[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 127.680 246.000 128.240 250.000 ;
    END
  END rdata[8]
  PIN rdata[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 134.400 246.000 134.960 250.000 ;
    END
  END rdata[9]
  PIN ready
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 147.840 4.000 148.400 ;
    END
  END ready
  PIN resetn
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 94.080 0.000 94.640 4.000 ;
    END
  END resetn
  PIN valid
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 134.400 4.000 134.960 ;
    END
  END valid
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 22.240 15.380 23.840 231.580 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.840 15.380 177.440 231.580 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 99.040 15.380 100.640 231.580 ;
    END
  END vss
  OBS
      LAYER Metal1 ;
        RECT 6.720 15.380 243.040 231.580 ;
      LAYER Metal2 ;
        RECT 6.300 245.700 66.900 246.000 ;
        RECT 68.060 245.700 73.620 246.000 ;
        RECT 74.780 245.700 90.420 246.000 ;
        RECT 91.580 245.700 100.500 246.000 ;
        RECT 101.660 245.700 113.940 246.000 ;
        RECT 115.100 245.700 117.300 246.000 ;
        RECT 118.460 245.700 127.380 246.000 ;
        RECT 128.540 245.700 130.740 246.000 ;
        RECT 131.900 245.700 134.100 246.000 ;
        RECT 135.260 245.700 150.900 246.000 ;
        RECT 152.060 245.700 154.260 246.000 ;
        RECT 155.420 245.700 157.620 246.000 ;
        RECT 158.780 245.700 160.980 246.000 ;
        RECT 162.140 245.700 164.340 246.000 ;
        RECT 165.500 245.700 167.700 246.000 ;
        RECT 168.860 245.700 174.420 246.000 ;
        RECT 175.580 245.700 181.140 246.000 ;
        RECT 182.300 245.700 187.860 246.000 ;
        RECT 189.020 245.700 191.220 246.000 ;
        RECT 192.380 245.700 197.940 246.000 ;
        RECT 199.100 245.700 221.460 246.000 ;
        RECT 222.620 245.700 241.780 246.000 ;
        RECT 6.300 4.300 241.780 245.700 ;
        RECT 6.300 3.500 6.420 4.300 ;
        RECT 7.580 3.500 9.780 4.300 ;
        RECT 10.940 3.500 13.140 4.300 ;
        RECT 14.300 3.500 16.500 4.300 ;
        RECT 17.660 3.500 19.860 4.300 ;
        RECT 21.020 3.500 23.220 4.300 ;
        RECT 24.380 3.500 26.580 4.300 ;
        RECT 27.740 3.500 29.940 4.300 ;
        RECT 31.100 3.500 33.300 4.300 ;
        RECT 34.460 3.500 36.660 4.300 ;
        RECT 37.820 3.500 40.020 4.300 ;
        RECT 41.180 3.500 43.380 4.300 ;
        RECT 44.540 3.500 46.740 4.300 ;
        RECT 47.900 3.500 50.100 4.300 ;
        RECT 51.260 3.500 53.460 4.300 ;
        RECT 54.620 3.500 56.820 4.300 ;
        RECT 57.980 3.500 60.180 4.300 ;
        RECT 61.340 3.500 63.540 4.300 ;
        RECT 64.700 3.500 66.900 4.300 ;
        RECT 68.060 3.500 70.260 4.300 ;
        RECT 71.420 3.500 73.620 4.300 ;
        RECT 74.780 3.500 76.980 4.300 ;
        RECT 78.140 3.500 80.340 4.300 ;
        RECT 81.500 3.500 83.700 4.300 ;
        RECT 84.860 3.500 87.060 4.300 ;
        RECT 88.220 3.500 90.420 4.300 ;
        RECT 91.580 3.500 93.780 4.300 ;
        RECT 94.940 3.500 97.140 4.300 ;
        RECT 98.300 3.500 100.500 4.300 ;
        RECT 101.660 3.500 103.860 4.300 ;
        RECT 105.020 3.500 110.580 4.300 ;
        RECT 111.740 3.500 113.940 4.300 ;
        RECT 115.100 3.500 117.300 4.300 ;
        RECT 118.460 3.500 124.020 4.300 ;
        RECT 125.180 3.500 130.740 4.300 ;
        RECT 131.900 3.500 134.100 4.300 ;
        RECT 135.260 3.500 147.540 4.300 ;
        RECT 148.700 3.500 150.900 4.300 ;
        RECT 152.060 3.500 154.260 4.300 ;
        RECT 155.420 3.500 157.620 4.300 ;
        RECT 158.780 3.500 164.340 4.300 ;
        RECT 165.500 3.500 167.700 4.300 ;
        RECT 168.860 3.500 177.780 4.300 ;
        RECT 178.940 3.500 184.500 4.300 ;
        RECT 185.660 3.500 187.860 4.300 ;
        RECT 189.020 3.500 191.220 4.300 ;
        RECT 192.380 3.500 194.580 4.300 ;
        RECT 195.740 3.500 197.940 4.300 ;
        RECT 199.100 3.500 201.300 4.300 ;
        RECT 202.460 3.500 204.660 4.300 ;
        RECT 205.820 3.500 208.020 4.300 ;
        RECT 209.180 3.500 211.380 4.300 ;
        RECT 212.540 3.500 214.740 4.300 ;
        RECT 215.900 3.500 218.100 4.300 ;
        RECT 219.260 3.500 221.460 4.300 ;
        RECT 222.620 3.500 224.820 4.300 ;
        RECT 225.980 3.500 241.780 4.300 ;
      LAYER Metal3 ;
        RECT 4.000 232.700 246.820 235.060 ;
        RECT 4.000 231.540 245.700 232.700 ;
        RECT 4.000 229.340 246.820 231.540 ;
        RECT 4.000 228.180 245.700 229.340 ;
        RECT 4.000 225.980 246.820 228.180 ;
        RECT 4.300 224.820 245.700 225.980 ;
        RECT 4.000 222.620 246.820 224.820 ;
        RECT 4.300 221.460 245.700 222.620 ;
        RECT 4.000 219.260 246.820 221.460 ;
        RECT 4.000 218.100 245.700 219.260 ;
        RECT 4.000 215.900 246.820 218.100 ;
        RECT 4.000 214.740 245.700 215.900 ;
        RECT 4.000 212.540 246.820 214.740 ;
        RECT 4.000 211.380 245.700 212.540 ;
        RECT 4.000 209.180 246.820 211.380 ;
        RECT 4.000 208.020 245.700 209.180 ;
        RECT 4.000 202.460 246.820 208.020 ;
        RECT 4.300 201.300 245.700 202.460 ;
        RECT 4.000 199.100 246.820 201.300 ;
        RECT 4.300 197.940 245.700 199.100 ;
        RECT 4.000 195.740 246.820 197.940 ;
        RECT 4.000 194.580 245.700 195.740 ;
        RECT 4.000 192.380 246.820 194.580 ;
        RECT 4.300 191.220 246.820 192.380 ;
        RECT 4.000 189.020 246.820 191.220 ;
        RECT 4.300 187.860 246.820 189.020 ;
        RECT 4.000 178.940 246.820 187.860 ;
        RECT 4.300 177.780 246.820 178.940 ;
        RECT 4.000 175.580 246.820 177.780 ;
        RECT 4.300 174.420 245.700 175.580 ;
        RECT 4.000 172.220 246.820 174.420 ;
        RECT 4.000 171.060 245.700 172.220 ;
        RECT 4.000 168.860 246.820 171.060 ;
        RECT 4.300 167.700 245.700 168.860 ;
        RECT 4.000 165.500 246.820 167.700 ;
        RECT 4.300 164.340 246.820 165.500 ;
        RECT 4.000 162.140 246.820 164.340 ;
        RECT 4.300 160.980 245.700 162.140 ;
        RECT 4.000 158.780 246.820 160.980 ;
        RECT 4.300 157.620 245.700 158.780 ;
        RECT 4.000 155.420 246.820 157.620 ;
        RECT 4.300 154.260 245.700 155.420 ;
        RECT 4.000 152.060 246.820 154.260 ;
        RECT 4.300 150.900 245.700 152.060 ;
        RECT 4.000 148.700 246.820 150.900 ;
        RECT 4.300 147.540 245.700 148.700 ;
        RECT 4.000 145.340 246.820 147.540 ;
        RECT 4.300 144.180 245.700 145.340 ;
        RECT 4.000 141.980 246.820 144.180 ;
        RECT 4.300 140.820 245.700 141.980 ;
        RECT 4.000 138.620 246.820 140.820 ;
        RECT 4.300 137.460 245.700 138.620 ;
        RECT 4.000 135.260 246.820 137.460 ;
        RECT 4.300 134.100 246.820 135.260 ;
        RECT 4.000 131.900 246.820 134.100 ;
        RECT 4.300 130.740 246.820 131.900 ;
        RECT 4.000 128.540 246.820 130.740 ;
        RECT 4.300 127.380 245.700 128.540 ;
        RECT 4.000 125.180 246.820 127.380 ;
        RECT 4.300 124.020 245.700 125.180 ;
        RECT 4.000 121.820 246.820 124.020 ;
        RECT 4.000 120.660 245.700 121.820 ;
        RECT 4.000 118.460 246.820 120.660 ;
        RECT 4.300 117.300 245.700 118.460 ;
        RECT 4.000 115.100 246.820 117.300 ;
        RECT 4.000 113.940 245.700 115.100 ;
        RECT 4.000 111.740 246.820 113.940 ;
        RECT 4.000 110.580 245.700 111.740 ;
        RECT 4.000 108.380 246.820 110.580 ;
        RECT 4.000 107.220 245.700 108.380 ;
        RECT 4.000 105.020 246.820 107.220 ;
        RECT 4.000 103.860 245.700 105.020 ;
        RECT 4.000 101.660 246.820 103.860 ;
        RECT 4.000 100.500 245.700 101.660 ;
        RECT 4.000 88.220 246.820 100.500 ;
        RECT 4.300 87.060 246.820 88.220 ;
        RECT 4.000 47.900 246.820 87.060 ;
        RECT 4.000 46.740 245.700 47.900 ;
        RECT 4.000 44.540 246.820 46.740 ;
        RECT 4.000 43.380 245.700 44.540 ;
        RECT 4.000 41.180 246.820 43.380 ;
        RECT 4.000 40.020 245.700 41.180 ;
        RECT 4.000 37.820 246.820 40.020 ;
        RECT 4.000 36.660 245.700 37.820 ;
        RECT 4.000 27.740 246.820 36.660 ;
        RECT 4.300 26.580 246.820 27.740 ;
        RECT 4.000 24.380 246.820 26.580 ;
        RECT 4.300 23.220 245.700 24.380 ;
        RECT 4.000 21.020 246.820 23.220 ;
        RECT 4.300 19.860 245.700 21.020 ;
        RECT 4.000 17.660 246.820 19.860 ;
        RECT 4.300 16.500 245.700 17.660 ;
        RECT 4.000 14.300 246.820 16.500 ;
        RECT 4.300 13.580 246.820 14.300 ;
      LAYER Metal4 ;
        RECT 16.940 16.890 21.940 222.790 ;
        RECT 24.140 16.890 98.740 222.790 ;
        RECT 100.940 16.890 175.540 222.790 ;
        RECT 177.740 16.890 219.380 222.790 ;
  END
END spimemio
END LIBRARY


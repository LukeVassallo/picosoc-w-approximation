magic
tech gf180mcuD
magscale 1 10
timestamp 1702237548
<< metal1 >>
rect 69010 77198 69022 77250
rect 69074 77247 69086 77250
rect 70018 77247 70030 77250
rect 69074 77201 70030 77247
rect 69074 77198 69086 77201
rect 70018 77198 70030 77201
rect 70082 77247 70094 77250
rect 70242 77247 70254 77250
rect 70082 77201 70254 77247
rect 70082 77198 70094 77201
rect 70242 77198 70254 77201
rect 70306 77198 70318 77250
rect 42802 77086 42814 77138
rect 42866 77135 42878 77138
rect 43586 77135 43598 77138
rect 42866 77089 43598 77135
rect 42866 77086 42878 77089
rect 43586 77086 43598 77089
rect 43650 77086 43662 77138
rect 50866 77086 50878 77138
rect 50930 77135 50942 77138
rect 51762 77135 51774 77138
rect 50930 77089 51774 77135
rect 50930 77086 50942 77089
rect 51762 77086 51774 77089
rect 51826 77135 51838 77138
rect 52098 77135 52110 77138
rect 51826 77089 52110 77135
rect 51826 77086 51838 77089
rect 52098 77086 52110 77089
rect 52162 77086 52174 77138
rect 64306 77086 64318 77138
rect 64370 77135 64382 77138
rect 65314 77135 65326 77138
rect 64370 77089 65326 77135
rect 64370 77086 64382 77089
rect 65314 77086 65326 77089
rect 65378 77086 65390 77138
rect 66322 77086 66334 77138
rect 66386 77135 66398 77138
rect 67106 77135 67118 77138
rect 66386 77089 67118 77135
rect 66386 77086 66398 77089
rect 67106 77086 67118 77089
rect 67170 77086 67182 77138
rect 71026 77086 71038 77138
rect 71090 77135 71102 77138
rect 72258 77135 72270 77138
rect 71090 77089 72270 77135
rect 71090 77086 71102 77089
rect 72258 77086 72270 77089
rect 72322 77086 72334 77138
rect 75170 77086 75182 77138
rect 75234 77135 75246 77138
rect 75618 77135 75630 77138
rect 75234 77089 75630 77135
rect 75234 77086 75246 77089
rect 75618 77086 75630 77089
rect 75682 77135 75694 77138
rect 76402 77135 76414 77138
rect 75682 77089 76414 77135
rect 75682 77086 75694 77089
rect 76402 77086 76414 77089
rect 76466 77086 76478 77138
rect 37202 76974 37214 77026
rect 37266 77023 37278 77026
rect 38098 77023 38110 77026
rect 37266 76977 38110 77023
rect 37266 76974 37278 76977
rect 38098 76974 38110 76977
rect 38162 76974 38174 77026
rect 43698 76974 43710 77026
rect 43762 77023 43774 77026
rect 43922 77023 43934 77026
rect 43762 76977 43934 77023
rect 43762 76974 43774 76977
rect 43922 76974 43934 76977
rect 43986 77023 43998 77026
rect 44482 77023 44494 77026
rect 43986 76977 44494 77023
rect 43986 76974 43998 76977
rect 44482 76974 44494 76977
rect 44546 76974 44558 77026
rect 45490 76974 45502 77026
rect 45554 77023 45566 77026
rect 46722 77023 46734 77026
rect 45554 76977 46734 77023
rect 45554 76974 45566 76977
rect 46722 76974 46734 76977
rect 46786 76974 46798 77026
rect 47506 76974 47518 77026
rect 47570 77023 47582 77026
rect 48290 77023 48302 77026
rect 47570 76977 48302 77023
rect 47570 76974 47582 76977
rect 48290 76974 48302 76977
rect 48354 76974 48366 77026
rect 48850 76974 48862 77026
rect 48914 77023 48926 77026
rect 50082 77023 50094 77026
rect 48914 76977 50094 77023
rect 48914 76974 48926 76977
rect 50082 76974 50094 76977
rect 50146 76974 50158 77026
rect 51538 76974 51550 77026
rect 51602 77023 51614 77026
rect 52994 77023 53006 77026
rect 51602 76977 53006 77023
rect 51602 76974 51614 76977
rect 52994 76974 53006 76977
rect 53058 76974 53070 77026
rect 62290 76974 62302 77026
rect 62354 77023 62366 77026
rect 63298 77023 63310 77026
rect 62354 76977 63310 77023
rect 62354 76974 62366 76977
rect 63298 76974 63310 76977
rect 63362 76974 63374 77026
rect 63634 76974 63646 77026
rect 63698 77023 63710 77026
rect 64642 77023 64654 77026
rect 63698 76977 64654 77023
rect 63698 76974 63710 76977
rect 64642 76974 64654 76977
rect 64706 76974 64718 77026
rect 65650 76974 65662 77026
rect 65714 77023 65726 77026
rect 66434 77023 66446 77026
rect 65714 76977 66446 77023
rect 65714 76974 65726 76977
rect 66434 76974 66446 76977
rect 66498 76974 66510 77026
rect 67666 76974 67678 77026
rect 67730 77023 67742 77026
rect 68450 77023 68462 77026
rect 67730 76977 68462 77023
rect 67730 76974 67742 76977
rect 68450 76974 68462 76977
rect 68514 76974 68526 77026
rect 69010 76974 69022 77026
rect 69074 77023 69086 77026
rect 70130 77023 70142 77026
rect 69074 76977 70142 77023
rect 69074 76974 69086 76977
rect 70130 76974 70142 76977
rect 70194 76974 70206 77026
rect 74386 76974 74398 77026
rect 74450 77023 74462 77026
rect 74946 77023 74958 77026
rect 74450 76977 74958 77023
rect 74450 76974 74462 76977
rect 74946 76974 74958 76977
rect 75010 77023 75022 77026
rect 75730 77023 75742 77026
rect 75010 76977 75742 77023
rect 75010 76974 75022 76977
rect 75730 76974 75742 76977
rect 75794 76974 75806 77026
rect 1344 76858 78624 76892
rect 1344 76806 19838 76858
rect 19890 76806 19942 76858
rect 19994 76806 20046 76858
rect 20098 76806 50558 76858
rect 50610 76806 50662 76858
rect 50714 76806 50766 76858
rect 50818 76806 78624 76858
rect 1344 76772 78624 76806
rect 4622 76690 4674 76702
rect 4622 76626 4674 76638
rect 15374 76690 15426 76702
rect 15374 76626 15426 76638
rect 21086 76690 21138 76702
rect 21086 76626 21138 76638
rect 24894 76690 24946 76702
rect 24894 76626 24946 76638
rect 25566 76690 25618 76702
rect 25566 76626 25618 76638
rect 26238 76690 26290 76702
rect 26238 76626 26290 76638
rect 26910 76690 26962 76702
rect 26910 76626 26962 76638
rect 27582 76690 27634 76702
rect 27582 76626 27634 76638
rect 28366 76690 28418 76702
rect 28366 76626 28418 76638
rect 28926 76690 28978 76702
rect 28926 76626 28978 76638
rect 29598 76690 29650 76702
rect 29598 76626 29650 76638
rect 30270 76690 30322 76702
rect 30270 76626 30322 76638
rect 30942 76690 30994 76702
rect 30942 76626 30994 76638
rect 31502 76690 31554 76702
rect 31502 76626 31554 76638
rect 32286 76690 32338 76702
rect 32286 76626 32338 76638
rect 36878 76690 36930 76702
rect 36878 76626 36930 76638
rect 38334 76690 38386 76702
rect 38334 76626 38386 76638
rect 39230 76690 39282 76702
rect 39230 76626 39282 76638
rect 40126 76690 40178 76702
rect 40126 76626 40178 76638
rect 41022 76690 41074 76702
rect 41022 76626 41074 76638
rect 42030 76690 42082 76702
rect 42030 76626 42082 76638
rect 42366 76690 42418 76702
rect 42366 76626 42418 76638
rect 43598 76690 43650 76702
rect 43598 76626 43650 76638
rect 44494 76690 44546 76702
rect 44494 76626 44546 76638
rect 48302 76690 48354 76702
rect 48302 76626 48354 76638
rect 49198 76690 49250 76702
rect 49198 76626 49250 76638
rect 50094 76690 50146 76702
rect 50094 76626 50146 76638
rect 51214 76690 51266 76702
rect 51214 76626 51266 76638
rect 52110 76690 52162 76702
rect 52110 76626 52162 76638
rect 53006 76690 53058 76702
rect 53006 76626 53058 76638
rect 53902 76690 53954 76702
rect 53902 76626 53954 76638
rect 55134 76690 55186 76702
rect 55134 76626 55186 76638
rect 59838 76690 59890 76702
rect 59838 76626 59890 76638
rect 63310 76690 63362 76702
rect 63310 76626 63362 76638
rect 63982 76690 64034 76702
rect 63982 76626 64034 76638
rect 64654 76690 64706 76702
rect 64654 76626 64706 76638
rect 65326 76690 65378 76702
rect 65326 76626 65378 76638
rect 66446 76690 66498 76702
rect 66446 76626 66498 76638
rect 67118 76690 67170 76702
rect 67118 76626 67170 76638
rect 67790 76690 67842 76702
rect 67790 76626 67842 76638
rect 68462 76690 68514 76702
rect 68462 76626 68514 76638
rect 69358 76690 69410 76702
rect 69358 76626 69410 76638
rect 70254 76690 70306 76702
rect 70254 76626 70306 76638
rect 72270 76690 72322 76702
rect 72270 76626 72322 76638
rect 76078 76690 76130 76702
rect 76078 76626 76130 76638
rect 77310 76690 77362 76702
rect 77310 76626 77362 76638
rect 4958 76578 5010 76590
rect 4958 76514 5010 76526
rect 5518 76578 5570 76590
rect 45950 76578 46002 76590
rect 62638 76578 62690 76590
rect 70926 76578 70978 76590
rect 19282 76526 19294 76578
rect 19346 76526 19358 76578
rect 36194 76526 36206 76578
rect 36258 76526 36270 76578
rect 61730 76526 61742 76578
rect 61794 76526 61806 76578
rect 63634 76526 63646 76578
rect 63698 76526 63710 76578
rect 64306 76526 64318 76578
rect 64370 76526 64382 76578
rect 64978 76526 64990 76578
rect 65042 76526 65054 76578
rect 65650 76526 65662 76578
rect 65714 76526 65726 76578
rect 66770 76526 66782 76578
rect 66834 76526 66846 76578
rect 67442 76526 67454 76578
rect 67506 76526 67518 76578
rect 68114 76526 68126 76578
rect 68178 76526 68190 76578
rect 69682 76526 69694 76578
rect 69746 76526 69758 76578
rect 70578 76526 70590 76578
rect 70642 76526 70654 76578
rect 5518 76514 5570 76526
rect 45950 76514 46002 76526
rect 62638 76514 62690 76526
rect 70926 76514 70978 76526
rect 71262 76578 71314 76590
rect 71262 76514 71314 76526
rect 71598 76578 71650 76590
rect 71598 76514 71650 76526
rect 71934 76578 71986 76590
rect 72942 76578 72994 76590
rect 74734 76578 74786 76590
rect 72594 76526 72606 76578
rect 72658 76526 72670 76578
rect 74050 76526 74062 76578
rect 74114 76526 74126 76578
rect 71934 76514 71986 76526
rect 72942 76514 72994 76526
rect 74734 76514 74786 76526
rect 75070 76578 75122 76590
rect 75070 76514 75122 76526
rect 75406 76578 75458 76590
rect 75406 76514 75458 76526
rect 75742 76578 75794 76590
rect 75742 76514 75794 76526
rect 76414 76578 76466 76590
rect 78194 76526 78206 76578
rect 78258 76526 78270 76578
rect 76414 76514 76466 76526
rect 62078 76466 62130 76478
rect 77870 76466 77922 76478
rect 4274 76414 4286 76466
rect 4338 76414 4350 76466
rect 5730 76414 5742 76466
rect 5794 76414 5806 76466
rect 12450 76414 12462 76466
rect 12514 76414 12526 76466
rect 16370 76414 16382 76466
rect 16434 76414 16446 76466
rect 18050 76414 18062 76466
rect 18114 76414 18126 76466
rect 23762 76414 23774 76466
rect 23826 76414 23838 76466
rect 35074 76414 35086 76466
rect 35138 76414 35150 76466
rect 36418 76414 36430 76466
rect 36482 76414 36494 76466
rect 46722 76414 46734 76466
rect 46786 76414 46798 76466
rect 47842 76414 47854 76466
rect 47906 76414 47918 76466
rect 58258 76414 58270 76466
rect 58322 76414 58334 76466
rect 58818 76414 58830 76466
rect 58882 76414 58894 76466
rect 62850 76414 62862 76466
rect 62914 76414 62926 76466
rect 73154 76414 73166 76466
rect 73218 76414 73230 76466
rect 74274 76414 74286 76466
rect 74338 76414 74350 76466
rect 62078 76402 62130 76414
rect 77870 76402 77922 76414
rect 13358 76354 13410 76366
rect 13358 76290 13410 76302
rect 17166 76354 17218 76366
rect 17166 76290 17218 76302
rect 21646 76354 21698 76366
rect 37438 76354 37490 76366
rect 40686 76354 40738 76366
rect 33394 76302 33406 76354
rect 33458 76302 33470 76354
rect 37874 76302 37886 76354
rect 37938 76302 37950 76354
rect 38770 76302 38782 76354
rect 38834 76302 38846 76354
rect 21646 76290 21698 76302
rect 37438 76290 37490 76302
rect 40686 76290 40738 76302
rect 41582 76354 41634 76366
rect 41582 76290 41634 76302
rect 42926 76354 42978 76366
rect 46286 76354 46338 76366
rect 44034 76302 44046 76354
rect 44098 76302 44110 76354
rect 44930 76302 44942 76354
rect 44994 76302 45006 76354
rect 45490 76302 45502 76354
rect 45554 76302 45566 76354
rect 42926 76290 42978 76302
rect 46286 76290 46338 76302
rect 47406 76354 47458 76366
rect 47406 76290 47458 76302
rect 48862 76354 48914 76366
rect 54462 76354 54514 76366
rect 49634 76302 49646 76354
rect 49698 76302 49710 76354
rect 50530 76302 50542 76354
rect 50594 76302 50606 76354
rect 51650 76302 51662 76354
rect 51714 76302 51726 76354
rect 52546 76302 52558 76354
rect 52610 76302 52622 76354
rect 53442 76302 53454 76354
rect 53506 76302 53518 76354
rect 48862 76290 48914 76302
rect 54462 76290 54514 76302
rect 55918 76354 55970 76366
rect 55918 76290 55970 76302
rect 69022 76354 69074 76366
rect 69022 76290 69074 76302
rect 76750 76354 76802 76366
rect 76750 76290 76802 76302
rect 1934 76242 1986 76254
rect 1934 76178 1986 76190
rect 11566 76242 11618 76254
rect 11566 76178 11618 76190
rect 1344 76074 78624 76108
rect 1344 76022 4478 76074
rect 4530 76022 4582 76074
rect 4634 76022 4686 76074
rect 4738 76022 35198 76074
rect 35250 76022 35302 76074
rect 35354 76022 35406 76074
rect 35458 76022 65918 76074
rect 65970 76022 66022 76074
rect 66074 76022 66126 76074
rect 66178 76022 78624 76074
rect 1344 75988 78624 76022
rect 11902 75906 11954 75918
rect 11902 75842 11954 75854
rect 16830 75906 16882 75918
rect 56702 75906 56754 75918
rect 21970 75854 21982 75906
rect 22034 75854 22046 75906
rect 45826 75854 45838 75906
rect 45890 75903 45902 75906
rect 46498 75903 46510 75906
rect 45890 75857 46510 75903
rect 45890 75854 45902 75857
rect 46498 75854 46510 75857
rect 46562 75854 46574 75906
rect 63298 75854 63310 75906
rect 63362 75903 63374 75906
rect 63746 75903 63758 75906
rect 63362 75857 63758 75903
rect 63362 75854 63374 75857
rect 63746 75854 63758 75857
rect 63810 75854 63822 75906
rect 16830 75842 16882 75854
rect 56702 75842 56754 75854
rect 1934 75794 1986 75806
rect 32734 75794 32786 75806
rect 37214 75794 37266 75806
rect 18610 75742 18622 75794
rect 18674 75742 18686 75794
rect 35186 75742 35198 75794
rect 35250 75742 35262 75794
rect 1934 75730 1986 75742
rect 32734 75730 32786 75742
rect 37214 75730 37266 75742
rect 39454 75794 39506 75806
rect 39454 75730 39506 75742
rect 41470 75794 41522 75806
rect 41470 75730 41522 75742
rect 42478 75794 42530 75806
rect 42478 75730 42530 75742
rect 43374 75794 43426 75806
rect 43374 75730 43426 75742
rect 43934 75794 43986 75806
rect 43934 75730 43986 75742
rect 44382 75794 44434 75806
rect 44382 75730 44434 75742
rect 46062 75794 46114 75806
rect 46062 75730 46114 75742
rect 46622 75794 46674 75806
rect 46622 75730 46674 75742
rect 48078 75794 48130 75806
rect 48078 75730 48130 75742
rect 48526 75794 48578 75806
rect 48526 75730 48578 75742
rect 49086 75794 49138 75806
rect 49086 75730 49138 75742
rect 49534 75794 49586 75806
rect 49534 75730 49586 75742
rect 50766 75794 50818 75806
rect 50766 75730 50818 75742
rect 51214 75794 51266 75806
rect 51214 75730 51266 75742
rect 51774 75794 51826 75806
rect 51774 75730 51826 75742
rect 52222 75794 52274 75806
rect 52222 75730 52274 75742
rect 63758 75794 63810 75806
rect 63758 75730 63810 75742
rect 64206 75794 64258 75806
rect 64206 75730 64258 75742
rect 64990 75794 65042 75806
rect 64990 75730 65042 75742
rect 65998 75794 66050 75806
rect 65998 75730 66050 75742
rect 66446 75794 66498 75806
rect 66446 75730 66498 75742
rect 67006 75794 67058 75806
rect 67006 75730 67058 75742
rect 67566 75794 67618 75806
rect 67566 75730 67618 75742
rect 68462 75794 68514 75806
rect 68462 75730 68514 75742
rect 69134 75794 69186 75806
rect 69134 75730 69186 75742
rect 70030 75794 70082 75806
rect 70030 75730 70082 75742
rect 70702 75794 70754 75806
rect 70702 75730 70754 75742
rect 71374 75794 71426 75806
rect 71374 75730 71426 75742
rect 71934 75794 71986 75806
rect 71934 75730 71986 75742
rect 72382 75794 72434 75806
rect 72382 75730 72434 75742
rect 73390 75794 73442 75806
rect 73390 75730 73442 75742
rect 73950 75794 74002 75806
rect 73950 75730 74002 75742
rect 74510 75794 74562 75806
rect 74510 75730 74562 75742
rect 75070 75794 75122 75806
rect 77746 75742 77758 75794
rect 77810 75742 77822 75794
rect 75070 75730 75122 75742
rect 4958 75682 5010 75694
rect 13582 75682 13634 75694
rect 4274 75630 4286 75682
rect 4338 75630 4350 75682
rect 12562 75630 12574 75682
rect 12626 75630 12638 75682
rect 4958 75618 5010 75630
rect 13582 75618 13634 75630
rect 14702 75682 14754 75694
rect 24782 75682 24834 75694
rect 17826 75630 17838 75682
rect 17890 75630 17902 75682
rect 20290 75630 20302 75682
rect 20354 75630 20366 75682
rect 23874 75630 23886 75682
rect 23938 75630 23950 75682
rect 14702 75618 14754 75630
rect 24782 75618 24834 75630
rect 25230 75682 25282 75694
rect 25230 75618 25282 75630
rect 32958 75682 33010 75694
rect 32958 75618 33010 75630
rect 33518 75682 33570 75694
rect 34414 75682 34466 75694
rect 33954 75630 33966 75682
rect 34018 75630 34030 75682
rect 33518 75618 33570 75630
rect 34414 75618 34466 75630
rect 34750 75682 34802 75694
rect 34750 75618 34802 75630
rect 35646 75682 35698 75694
rect 35646 75618 35698 75630
rect 36206 75682 36258 75694
rect 36206 75618 36258 75630
rect 37438 75682 37490 75694
rect 37438 75618 37490 75630
rect 37998 75682 38050 75694
rect 37998 75618 38050 75630
rect 38334 75682 38386 75694
rect 38334 75618 38386 75630
rect 38894 75682 38946 75694
rect 38894 75618 38946 75630
rect 40910 75682 40962 75694
rect 40910 75618 40962 75630
rect 41694 75682 41746 75694
rect 41694 75618 41746 75630
rect 45054 75682 45106 75694
rect 45054 75618 45106 75630
rect 47070 75682 47122 75694
rect 47070 75618 47122 75630
rect 47630 75682 47682 75694
rect 47630 75618 47682 75630
rect 49758 75682 49810 75694
rect 49758 75618 49810 75630
rect 50318 75682 50370 75694
rect 50318 75618 50370 75630
rect 52670 75682 52722 75694
rect 52670 75618 52722 75630
rect 53230 75682 53282 75694
rect 53230 75618 53282 75630
rect 53790 75682 53842 75694
rect 53790 75618 53842 75630
rect 54350 75682 54402 75694
rect 54350 75618 54402 75630
rect 54686 75682 54738 75694
rect 54686 75618 54738 75630
rect 55246 75682 55298 75694
rect 56142 75682 56194 75694
rect 61742 75682 61794 75694
rect 55682 75630 55694 75682
rect 55746 75630 55758 75682
rect 59042 75630 59054 75682
rect 59106 75630 59118 75682
rect 55246 75618 55298 75630
rect 56142 75618 56194 75630
rect 61742 75618 61794 75630
rect 63310 75682 63362 75694
rect 63310 75618 63362 75630
rect 65214 75682 65266 75694
rect 65214 75618 65266 75630
rect 72606 75682 72658 75694
rect 76190 75682 76242 75694
rect 75394 75630 75406 75682
rect 75458 75630 75470 75682
rect 72606 75618 72658 75630
rect 76190 75618 76242 75630
rect 76862 75682 76914 75694
rect 76862 75618 76914 75630
rect 4622 75570 4674 75582
rect 4622 75506 4674 75518
rect 24222 75570 24274 75582
rect 24222 75506 24274 75518
rect 45614 75570 45666 75582
rect 45614 75506 45666 75518
rect 61182 75570 61234 75582
rect 61182 75506 61234 75518
rect 62078 75570 62130 75582
rect 62078 75506 62130 75518
rect 75630 75570 75682 75582
rect 77198 75570 77250 75582
rect 76514 75518 76526 75570
rect 76578 75518 76590 75570
rect 75630 75506 75682 75518
rect 77198 75506 77250 75518
rect 78206 75570 78258 75582
rect 78206 75506 78258 75518
rect 14254 75458 14306 75470
rect 59390 75458 59442 75470
rect 60510 75458 60562 75470
rect 62414 75458 62466 75470
rect 42018 75406 42030 75458
rect 42082 75406 42094 75458
rect 59714 75406 59726 75458
rect 59778 75406 59790 75458
rect 60834 75406 60846 75458
rect 60898 75406 60910 75458
rect 14254 75394 14306 75406
rect 59390 75394 59442 75406
rect 60510 75394 60562 75406
rect 62414 75394 62466 75406
rect 62862 75458 62914 75470
rect 65538 75406 65550 75458
rect 65602 75406 65614 75458
rect 72930 75406 72942 75458
rect 72994 75406 73006 75458
rect 62862 75394 62914 75406
rect 1344 75290 78624 75324
rect 1344 75238 19838 75290
rect 19890 75238 19942 75290
rect 19994 75238 20046 75290
rect 20098 75238 50558 75290
rect 50610 75238 50662 75290
rect 50714 75238 50766 75290
rect 50818 75238 78624 75290
rect 1344 75204 78624 75238
rect 4622 75122 4674 75134
rect 4622 75058 4674 75070
rect 12910 75122 12962 75134
rect 12910 75058 12962 75070
rect 23102 75122 23154 75134
rect 23102 75058 23154 75070
rect 23550 75122 23602 75134
rect 23550 75058 23602 75070
rect 34638 75122 34690 75134
rect 34638 75058 34690 75070
rect 35534 75122 35586 75134
rect 35534 75058 35586 75070
rect 35982 75122 36034 75134
rect 35982 75058 36034 75070
rect 36766 75122 36818 75134
rect 36766 75058 36818 75070
rect 37662 75122 37714 75134
rect 37662 75058 37714 75070
rect 46846 75122 46898 75134
rect 46846 75058 46898 75070
rect 52782 75122 52834 75134
rect 52782 75058 52834 75070
rect 53566 75122 53618 75134
rect 53566 75058 53618 75070
rect 54462 75122 54514 75134
rect 54462 75058 54514 75070
rect 55358 75122 55410 75134
rect 55358 75058 55410 75070
rect 57598 75122 57650 75134
rect 57598 75058 57650 75070
rect 61294 75122 61346 75134
rect 61294 75058 61346 75070
rect 61742 75122 61794 75134
rect 61742 75058 61794 75070
rect 62190 75122 62242 75134
rect 62190 75058 62242 75070
rect 64654 75122 64706 75134
rect 64654 75058 64706 75070
rect 74062 75122 74114 75134
rect 74062 75058 74114 75070
rect 74510 75122 74562 75134
rect 74510 75058 74562 75070
rect 74958 75122 75010 75134
rect 74958 75058 75010 75070
rect 76862 75122 76914 75134
rect 76862 75058 76914 75070
rect 78206 75122 78258 75134
rect 78206 75058 78258 75070
rect 75406 75010 75458 75022
rect 15250 74958 15262 75010
rect 15314 74958 15326 75010
rect 75406 74946 75458 74958
rect 75630 75010 75682 75022
rect 75630 74946 75682 74958
rect 75966 75010 76018 75022
rect 75966 74946 76018 74958
rect 60846 74898 60898 74910
rect 4162 74846 4174 74898
rect 4226 74846 4238 74898
rect 4834 74846 4846 74898
rect 4898 74846 4910 74898
rect 13458 74846 13470 74898
rect 13522 74846 13534 74898
rect 16482 74846 16494 74898
rect 16546 74846 16558 74898
rect 22754 74846 22766 74898
rect 22818 74846 22830 74898
rect 60386 74846 60398 74898
rect 60450 74846 60462 74898
rect 77298 74846 77310 74898
rect 77362 74846 77374 74898
rect 60846 74834 60898 74846
rect 17950 74786 18002 74798
rect 2146 74734 2158 74786
rect 2210 74734 2222 74786
rect 17950 74722 18002 74734
rect 18286 74786 18338 74798
rect 18286 74722 18338 74734
rect 19406 74786 19458 74798
rect 19406 74722 19458 74734
rect 19854 74786 19906 74798
rect 19854 74722 19906 74734
rect 20414 74786 20466 74798
rect 20414 74722 20466 74734
rect 35086 74786 35138 74798
rect 35086 74722 35138 74734
rect 38222 74786 38274 74798
rect 38222 74722 38274 74734
rect 38782 74786 38834 74798
rect 38782 74722 38834 74734
rect 58046 74786 58098 74798
rect 77758 74786 77810 74798
rect 76402 74734 76414 74786
rect 76466 74734 76478 74786
rect 58046 74722 58098 74734
rect 77758 74722 77810 74734
rect 37426 74622 37438 74674
rect 37490 74671 37502 74674
rect 38210 74671 38222 74674
rect 37490 74625 38222 74671
rect 37490 74622 37502 74625
rect 38210 74622 38222 74625
rect 38274 74622 38286 74674
rect 1344 74506 78624 74540
rect 1344 74454 4478 74506
rect 4530 74454 4582 74506
rect 4634 74454 4686 74506
rect 4738 74454 35198 74506
rect 35250 74454 35302 74506
rect 35354 74454 35406 74506
rect 35458 74454 65918 74506
rect 65970 74454 66022 74506
rect 66074 74454 66126 74506
rect 66178 74454 78624 74506
rect 1344 74420 78624 74454
rect 19182 74338 19234 74350
rect 15922 74286 15934 74338
rect 15986 74286 15998 74338
rect 76066 74286 76078 74338
rect 76130 74335 76142 74338
rect 76402 74335 76414 74338
rect 76130 74289 76414 74335
rect 76130 74286 76142 74289
rect 76402 74286 76414 74289
rect 76466 74286 76478 74338
rect 19182 74274 19234 74286
rect 1934 74226 1986 74238
rect 58494 74226 58546 74238
rect 11218 74174 11230 74226
rect 11282 74174 11294 74226
rect 1934 74162 1986 74174
rect 58494 74162 58546 74174
rect 59166 74226 59218 74238
rect 59166 74162 59218 74174
rect 59502 74226 59554 74238
rect 59502 74162 59554 74174
rect 75742 74226 75794 74238
rect 75742 74162 75794 74174
rect 76414 74226 76466 74238
rect 76414 74162 76466 74174
rect 75294 74114 75346 74126
rect 4274 74062 4286 74114
rect 4338 74062 4350 74114
rect 4834 74062 4846 74114
rect 4898 74062 4910 74114
rect 12674 74062 12686 74114
rect 12738 74062 12750 74114
rect 17602 74062 17614 74114
rect 17666 74062 17678 74114
rect 18162 74062 18174 74114
rect 18226 74062 18238 74114
rect 75294 74050 75346 74062
rect 76974 74114 77026 74126
rect 76974 74050 77026 74062
rect 77534 74114 77586 74126
rect 78082 74062 78094 74114
rect 78146 74062 78158 74114
rect 77534 74050 77586 74062
rect 4622 74002 4674 74014
rect 4622 73938 4674 73950
rect 14030 74002 14082 74014
rect 14030 73938 14082 73950
rect 14366 74002 14418 74014
rect 14366 73938 14418 73950
rect 22990 74002 23042 74014
rect 22990 73938 23042 73950
rect 77870 74002 77922 74014
rect 77870 73938 77922 73950
rect 1344 73722 78624 73756
rect 1344 73670 19838 73722
rect 19890 73670 19942 73722
rect 19994 73670 20046 73722
rect 20098 73670 50558 73722
rect 50610 73670 50662 73722
rect 50714 73670 50766 73722
rect 50818 73670 78624 73722
rect 1344 73636 78624 73670
rect 76190 73554 76242 73566
rect 76190 73490 76242 73502
rect 76638 73554 76690 73566
rect 76638 73490 76690 73502
rect 77198 73554 77250 73566
rect 77198 73490 77250 73502
rect 77646 73554 77698 73566
rect 77646 73490 77698 73502
rect 78206 73554 78258 73566
rect 78206 73490 78258 73502
rect 4622 73442 4674 73454
rect 12114 73390 12126 73442
rect 12178 73390 12190 73442
rect 77858 73390 77870 73442
rect 77922 73390 77934 73442
rect 4622 73378 4674 73390
rect 4274 73278 4286 73330
rect 4338 73278 4350 73330
rect 4834 73278 4846 73330
rect 4898 73278 4910 73330
rect 13906 73278 13918 73330
rect 13970 73278 13982 73330
rect 16370 73278 16382 73330
rect 16434 73278 16446 73330
rect 18062 73218 18114 73230
rect 14578 73166 14590 73218
rect 14642 73166 14654 73218
rect 18062 73154 18114 73166
rect 1934 73106 1986 73118
rect 1934 73042 1986 73054
rect 1344 72938 78624 72972
rect 1344 72886 4478 72938
rect 4530 72886 4582 72938
rect 4634 72886 4686 72938
rect 4738 72886 35198 72938
rect 35250 72886 35302 72938
rect 35354 72886 35406 72938
rect 35458 72886 65918 72938
rect 65970 72886 66022 72938
rect 66074 72886 66126 72938
rect 66178 72886 78624 72938
rect 1344 72852 78624 72886
rect 1934 72658 1986 72670
rect 1934 72594 1986 72606
rect 77198 72658 77250 72670
rect 77198 72594 77250 72606
rect 3826 72494 3838 72546
rect 3890 72494 3902 72546
rect 77646 72434 77698 72446
rect 77646 72370 77698 72382
rect 78206 72434 78258 72446
rect 78206 72370 78258 72382
rect 14142 72322 14194 72334
rect 14142 72258 14194 72270
rect 77870 72322 77922 72334
rect 77870 72258 77922 72270
rect 1344 72154 78624 72188
rect 1344 72102 19838 72154
rect 19890 72102 19942 72154
rect 19994 72102 20046 72154
rect 20098 72102 50558 72154
rect 50610 72102 50662 72154
rect 50714 72102 50766 72154
rect 50818 72102 78624 72154
rect 1344 72068 78624 72102
rect 3166 71986 3218 71998
rect 3166 71922 3218 71934
rect 3502 71986 3554 71998
rect 3502 71922 3554 71934
rect 4174 71986 4226 71998
rect 4174 71922 4226 71934
rect 2494 71874 2546 71886
rect 2494 71810 2546 71822
rect 3838 71874 3890 71886
rect 3838 71810 3890 71822
rect 4510 71874 4562 71886
rect 4510 71810 4562 71822
rect 77870 71874 77922 71886
rect 77870 71810 77922 71822
rect 2158 71762 2210 71774
rect 78206 71762 78258 71774
rect 2930 71710 2942 71762
rect 2994 71710 3006 71762
rect 2158 71698 2210 71710
rect 78206 71698 78258 71710
rect 1934 71650 1986 71662
rect 1934 71586 1986 71598
rect 77646 71650 77698 71662
rect 77646 71586 77698 71598
rect 1344 71370 78624 71404
rect 1344 71318 4478 71370
rect 4530 71318 4582 71370
rect 4634 71318 4686 71370
rect 4738 71318 35198 71370
rect 35250 71318 35302 71370
rect 35354 71318 35406 71370
rect 35458 71318 65918 71370
rect 65970 71318 66022 71370
rect 66074 71318 66126 71370
rect 66178 71318 78624 71370
rect 1344 71284 78624 71318
rect 1934 71090 1986 71102
rect 1934 71026 1986 71038
rect 77646 70978 77698 70990
rect 3938 70926 3950 70978
rect 4002 70926 4014 70978
rect 77646 70914 77698 70926
rect 77422 70754 77474 70766
rect 77422 70690 77474 70702
rect 78206 70754 78258 70766
rect 78206 70690 78258 70702
rect 1344 70586 78624 70620
rect 1344 70534 19838 70586
rect 19890 70534 19942 70586
rect 19994 70534 20046 70586
rect 20098 70534 50558 70586
rect 50610 70534 50662 70586
rect 50714 70534 50766 70586
rect 50818 70534 78624 70586
rect 1344 70500 78624 70534
rect 3826 70142 3838 70194
rect 3890 70142 3902 70194
rect 1934 69970 1986 69982
rect 1934 69906 1986 69918
rect 1344 69802 78624 69836
rect 1344 69750 4478 69802
rect 4530 69750 4582 69802
rect 4634 69750 4686 69802
rect 4738 69750 35198 69802
rect 35250 69750 35302 69802
rect 35354 69750 35406 69802
rect 35458 69750 65918 69802
rect 65970 69750 66022 69802
rect 66074 69750 66126 69802
rect 66178 69750 78624 69802
rect 1344 69716 78624 69750
rect 2930 69358 2942 69410
rect 2994 69358 3006 69410
rect 2382 69298 2434 69310
rect 2382 69234 2434 69246
rect 2718 69298 2770 69310
rect 2718 69234 2770 69246
rect 2046 69186 2098 69198
rect 2046 69122 2098 69134
rect 77646 69186 77698 69198
rect 78206 69186 78258 69198
rect 77858 69134 77870 69186
rect 77922 69134 77934 69186
rect 77646 69122 77698 69134
rect 78206 69122 78258 69134
rect 1344 69018 78624 69052
rect 1344 68966 19838 69018
rect 19890 68966 19942 69018
rect 19994 68966 20046 69018
rect 20098 68966 50558 69018
rect 50610 68966 50662 69018
rect 50714 68966 50766 69018
rect 50818 68966 78624 69018
rect 1344 68932 78624 68966
rect 77422 68626 77474 68638
rect 2034 68574 2046 68626
rect 2098 68574 2110 68626
rect 77422 68562 77474 68574
rect 78206 68626 78258 68638
rect 78206 68562 78258 68574
rect 77646 68514 77698 68526
rect 77646 68450 77698 68462
rect 2718 68402 2770 68414
rect 2718 68338 2770 68350
rect 1344 68234 78624 68268
rect 1344 68182 4478 68234
rect 4530 68182 4582 68234
rect 4634 68182 4686 68234
rect 4738 68182 35198 68234
rect 35250 68182 35302 68234
rect 35354 68182 35406 68234
rect 35458 68182 65918 68234
rect 65970 68182 66022 68234
rect 66074 68182 66126 68234
rect 66178 68182 78624 68234
rect 1344 68148 78624 68182
rect 1934 67954 1986 67966
rect 1934 67890 1986 67902
rect 3826 67790 3838 67842
rect 3890 67790 3902 67842
rect 1344 67450 78624 67484
rect 1344 67398 19838 67450
rect 19890 67398 19942 67450
rect 19994 67398 20046 67450
rect 20098 67398 50558 67450
rect 50610 67398 50662 67450
rect 50714 67398 50766 67450
rect 50818 67398 78624 67450
rect 1344 67364 78624 67398
rect 3390 67282 3442 67294
rect 3390 67218 3442 67230
rect 2046 67170 2098 67182
rect 2046 67106 2098 67118
rect 2382 67170 2434 67182
rect 2382 67106 2434 67118
rect 3054 67170 3106 67182
rect 77858 67118 77870 67170
rect 77922 67118 77934 67170
rect 3054 67106 3106 67118
rect 2718 67058 2770 67070
rect 78206 67058 78258 67070
rect 3602 67006 3614 67058
rect 3666 67006 3678 67058
rect 2718 66994 2770 67006
rect 78206 66994 78258 67006
rect 77646 66946 77698 66958
rect 77646 66882 77698 66894
rect 1344 66666 78624 66700
rect 1344 66614 4478 66666
rect 4530 66614 4582 66666
rect 4634 66614 4686 66666
rect 4738 66614 35198 66666
rect 35250 66614 35302 66666
rect 35354 66614 35406 66666
rect 35458 66614 65918 66666
rect 65970 66614 66022 66666
rect 66074 66614 66126 66666
rect 66178 66614 78624 66666
rect 1344 66580 78624 66614
rect 2034 66222 2046 66274
rect 2098 66222 2110 66274
rect 2718 66050 2770 66062
rect 2718 65986 2770 65998
rect 77646 66050 77698 66062
rect 78206 66050 78258 66062
rect 77858 65998 77870 66050
rect 77922 65998 77934 66050
rect 77646 65986 77698 65998
rect 78206 65986 78258 65998
rect 1344 65882 78624 65916
rect 1344 65830 19838 65882
rect 19890 65830 19942 65882
rect 19994 65830 20046 65882
rect 20098 65830 50558 65882
rect 50610 65830 50662 65882
rect 50714 65830 50766 65882
rect 50818 65830 78624 65882
rect 1344 65796 78624 65830
rect 4274 65438 4286 65490
rect 4338 65438 4350 65490
rect 1934 65266 1986 65278
rect 1934 65202 1986 65214
rect 1344 65098 78624 65132
rect 1344 65046 4478 65098
rect 4530 65046 4582 65098
rect 4634 65046 4686 65098
rect 4738 65046 35198 65098
rect 35250 65046 35302 65098
rect 35354 65046 35406 65098
rect 35458 65046 65918 65098
rect 65970 65046 66022 65098
rect 66074 65046 66126 65098
rect 66178 65046 78624 65098
rect 1344 65012 78624 65046
rect 1934 64818 1986 64830
rect 1934 64754 1986 64766
rect 77646 64706 77698 64718
rect 3826 64654 3838 64706
rect 3890 64654 3902 64706
rect 77646 64642 77698 64654
rect 4622 64594 4674 64606
rect 4622 64530 4674 64542
rect 4958 64594 5010 64606
rect 4958 64530 5010 64542
rect 77422 64594 77474 64606
rect 77422 64530 77474 64542
rect 78206 64594 78258 64606
rect 78206 64530 78258 64542
rect 1344 64314 78624 64348
rect 1344 64262 19838 64314
rect 19890 64262 19942 64314
rect 19994 64262 20046 64314
rect 20098 64262 50558 64314
rect 50610 64262 50662 64314
rect 50714 64262 50766 64314
rect 50818 64262 78624 64314
rect 1344 64228 78624 64262
rect 3838 64146 3890 64158
rect 3838 64082 3890 64094
rect 2494 64034 2546 64046
rect 2494 63970 2546 63982
rect 3166 64034 3218 64046
rect 3166 63970 3218 63982
rect 77422 63922 77474 63934
rect 2258 63870 2270 63922
rect 2322 63870 2334 63922
rect 2930 63870 2942 63922
rect 2994 63870 3006 63922
rect 3602 63870 3614 63922
rect 3666 63870 3678 63922
rect 77422 63858 77474 63870
rect 77646 63922 77698 63934
rect 77646 63858 77698 63870
rect 78206 63922 78258 63934
rect 78206 63858 78258 63870
rect 1344 63530 78624 63564
rect 1344 63478 4478 63530
rect 4530 63478 4582 63530
rect 4634 63478 4686 63530
rect 4738 63478 35198 63530
rect 35250 63478 35302 63530
rect 35354 63478 35406 63530
rect 35458 63478 65918 63530
rect 65970 63478 66022 63530
rect 66074 63478 66126 63530
rect 66178 63478 78624 63530
rect 1344 63444 78624 63478
rect 1934 63250 1986 63262
rect 1934 63186 1986 63198
rect 3826 63086 3838 63138
rect 3890 63086 3902 63138
rect 78206 63026 78258 63038
rect 78206 62962 78258 62974
rect 77646 62914 77698 62926
rect 77646 62850 77698 62862
rect 77870 62914 77922 62926
rect 77870 62850 77922 62862
rect 1344 62746 78624 62780
rect 1344 62694 19838 62746
rect 19890 62694 19942 62746
rect 19994 62694 20046 62746
rect 20098 62694 50558 62746
rect 50610 62694 50662 62746
rect 50714 62694 50766 62746
rect 50818 62694 78624 62746
rect 1344 62660 78624 62694
rect 3826 62302 3838 62354
rect 3890 62302 3902 62354
rect 1934 62130 1986 62142
rect 1934 62066 1986 62078
rect 1344 61962 78624 61996
rect 1344 61910 4478 61962
rect 4530 61910 4582 61962
rect 4634 61910 4686 61962
rect 4738 61910 35198 61962
rect 35250 61910 35302 61962
rect 35354 61910 35406 61962
rect 35458 61910 65918 61962
rect 65970 61910 66022 61962
rect 66074 61910 66126 61962
rect 66178 61910 78624 61962
rect 1344 61876 78624 61910
rect 77646 61570 77698 61582
rect 2258 61518 2270 61570
rect 2322 61518 2334 61570
rect 3602 61518 3614 61570
rect 3666 61518 3678 61570
rect 77646 61506 77698 61518
rect 2718 61458 2770 61470
rect 2718 61394 2770 61406
rect 3054 61458 3106 61470
rect 3054 61394 3106 61406
rect 3390 61458 3442 61470
rect 3390 61394 3442 61406
rect 2046 61346 2098 61358
rect 2046 61282 2098 61294
rect 4286 61346 4338 61358
rect 4286 61282 4338 61294
rect 77422 61346 77474 61358
rect 77422 61282 77474 61294
rect 78206 61346 78258 61358
rect 78206 61282 78258 61294
rect 1344 61178 78624 61212
rect 1344 61126 19838 61178
rect 19890 61126 19942 61178
rect 19994 61126 20046 61178
rect 20098 61126 50558 61178
rect 50610 61126 50662 61178
rect 50714 61126 50766 61178
rect 50818 61126 78624 61178
rect 1344 61092 78624 61126
rect 77870 60898 77922 60910
rect 77870 60834 77922 60846
rect 77646 60786 77698 60798
rect 2034 60734 2046 60786
rect 2098 60734 2110 60786
rect 77646 60722 77698 60734
rect 78206 60786 78258 60798
rect 78206 60722 78258 60734
rect 2718 60562 2770 60574
rect 2718 60498 2770 60510
rect 1344 60394 78624 60428
rect 1344 60342 4478 60394
rect 4530 60342 4582 60394
rect 4634 60342 4686 60394
rect 4738 60342 35198 60394
rect 35250 60342 35302 60394
rect 35354 60342 35406 60394
rect 35458 60342 65918 60394
rect 65970 60342 66022 60394
rect 66074 60342 66126 60394
rect 66178 60342 78624 60394
rect 1344 60308 78624 60342
rect 1934 60114 1986 60126
rect 1934 60050 1986 60062
rect 3826 59950 3838 60002
rect 3890 59950 3902 60002
rect 1344 59610 78624 59644
rect 1344 59558 19838 59610
rect 19890 59558 19942 59610
rect 19994 59558 20046 59610
rect 20098 59558 50558 59610
rect 50610 59558 50662 59610
rect 50714 59558 50766 59610
rect 50818 59558 78624 59610
rect 1344 59524 78624 59558
rect 2718 59442 2770 59454
rect 2718 59378 2770 59390
rect 2046 59330 2098 59342
rect 2046 59266 2098 59278
rect 2382 59218 2434 59230
rect 3502 59218 3554 59230
rect 2930 59166 2942 59218
rect 2994 59166 3006 59218
rect 2382 59154 2434 59166
rect 3502 59154 3554 59166
rect 78206 59218 78258 59230
rect 78206 59154 78258 59166
rect 77422 59106 77474 59118
rect 77422 59042 77474 59054
rect 77646 59106 77698 59118
rect 77646 59042 77698 59054
rect 1344 58826 78624 58860
rect 1344 58774 4478 58826
rect 4530 58774 4582 58826
rect 4634 58774 4686 58826
rect 4738 58774 35198 58826
rect 35250 58774 35302 58826
rect 35354 58774 35406 58826
rect 35458 58774 65918 58826
rect 65970 58774 66022 58826
rect 66074 58774 66126 58826
rect 66178 58774 78624 58826
rect 1344 58740 78624 58774
rect 2034 58382 2046 58434
rect 2098 58382 2110 58434
rect 2718 58210 2770 58222
rect 2718 58146 2770 58158
rect 77646 58210 77698 58222
rect 78206 58210 78258 58222
rect 77858 58158 77870 58210
rect 77922 58158 77934 58210
rect 77646 58146 77698 58158
rect 78206 58146 78258 58158
rect 1344 58042 78624 58076
rect 1344 57990 19838 58042
rect 19890 57990 19942 58042
rect 19994 57990 20046 58042
rect 20098 57990 50558 58042
rect 50610 57990 50662 58042
rect 50714 57990 50766 58042
rect 50818 57990 78624 58042
rect 1344 57956 78624 57990
rect 4274 57598 4286 57650
rect 4338 57598 4350 57650
rect 1934 57426 1986 57438
rect 1934 57362 1986 57374
rect 1344 57258 78624 57292
rect 1344 57206 4478 57258
rect 4530 57206 4582 57258
rect 4634 57206 4686 57258
rect 4738 57206 35198 57258
rect 35250 57206 35302 57258
rect 35354 57206 35406 57258
rect 35458 57206 65918 57258
rect 65970 57206 66022 57258
rect 66074 57206 66126 57258
rect 66178 57206 78624 57258
rect 1344 57172 78624 57206
rect 1934 56978 1986 56990
rect 1934 56914 1986 56926
rect 3826 56814 3838 56866
rect 3890 56814 3902 56866
rect 4834 56814 4846 56866
rect 4898 56814 4910 56866
rect 4622 56754 4674 56766
rect 4622 56690 4674 56702
rect 77646 56754 77698 56766
rect 77646 56690 77698 56702
rect 78206 56754 78258 56766
rect 78206 56690 78258 56702
rect 77870 56642 77922 56654
rect 77870 56578 77922 56590
rect 1344 56474 78624 56508
rect 1344 56422 19838 56474
rect 19890 56422 19942 56474
rect 19994 56422 20046 56474
rect 20098 56422 50558 56474
rect 50610 56422 50662 56474
rect 50714 56422 50766 56474
rect 50818 56422 78624 56474
rect 1344 56388 78624 56422
rect 2718 56306 2770 56318
rect 2718 56242 2770 56254
rect 3726 56306 3778 56318
rect 3726 56242 3778 56254
rect 2046 56194 2098 56206
rect 2046 56130 2098 56142
rect 2382 56194 2434 56206
rect 2382 56130 2434 56142
rect 3390 56194 3442 56206
rect 77858 56142 77870 56194
rect 77922 56142 77934 56194
rect 3390 56130 3442 56142
rect 78206 56082 78258 56094
rect 2930 56030 2942 56082
rect 2994 56030 3006 56082
rect 78206 56018 78258 56030
rect 77646 55970 77698 55982
rect 77646 55906 77698 55918
rect 1344 55690 78624 55724
rect 1344 55638 4478 55690
rect 4530 55638 4582 55690
rect 4634 55638 4686 55690
rect 4738 55638 35198 55690
rect 35250 55638 35302 55690
rect 35354 55638 35406 55690
rect 35458 55638 65918 55690
rect 65970 55638 66022 55690
rect 66074 55638 66126 55690
rect 66178 55638 78624 55690
rect 1344 55604 78624 55638
rect 2034 55246 2046 55298
rect 2098 55246 2110 55298
rect 78206 55186 78258 55198
rect 78206 55122 78258 55134
rect 2718 55074 2770 55086
rect 2718 55010 2770 55022
rect 77646 55074 77698 55086
rect 77646 55010 77698 55022
rect 77870 55074 77922 55086
rect 77870 55010 77922 55022
rect 1344 54906 78624 54940
rect 1344 54854 19838 54906
rect 19890 54854 19942 54906
rect 19994 54854 20046 54906
rect 20098 54854 50558 54906
rect 50610 54854 50662 54906
rect 50714 54854 50766 54906
rect 50818 54854 78624 54906
rect 1344 54820 78624 54854
rect 3826 54462 3838 54514
rect 3890 54462 3902 54514
rect 1934 54290 1986 54302
rect 1934 54226 1986 54238
rect 1344 54122 78624 54156
rect 1344 54070 4478 54122
rect 4530 54070 4582 54122
rect 4634 54070 4686 54122
rect 4738 54070 35198 54122
rect 35250 54070 35302 54122
rect 35354 54070 35406 54122
rect 35458 54070 65918 54122
rect 65970 54070 66022 54122
rect 66074 54070 66126 54122
rect 66178 54070 78624 54122
rect 1344 54036 78624 54070
rect 2930 53678 2942 53730
rect 2994 53678 3006 53730
rect 2158 53618 2210 53630
rect 2158 53554 2210 53566
rect 3166 53618 3218 53630
rect 3166 53554 3218 53566
rect 3502 53618 3554 53630
rect 3502 53554 3554 53566
rect 3838 53618 3890 53630
rect 3838 53554 3890 53566
rect 77870 53618 77922 53630
rect 77870 53554 77922 53566
rect 78206 53618 78258 53630
rect 78206 53554 78258 53566
rect 1934 53506 1986 53518
rect 1934 53442 1986 53454
rect 2494 53506 2546 53518
rect 2494 53442 2546 53454
rect 77646 53506 77698 53518
rect 77646 53442 77698 53454
rect 1344 53338 78624 53372
rect 1344 53286 19838 53338
rect 19890 53286 19942 53338
rect 19994 53286 20046 53338
rect 20098 53286 50558 53338
rect 50610 53286 50662 53338
rect 50714 53286 50766 53338
rect 50818 53286 78624 53338
rect 1344 53252 78624 53286
rect 77870 53058 77922 53070
rect 77870 52994 77922 53006
rect 78206 52946 78258 52958
rect 3938 52894 3950 52946
rect 4002 52894 4014 52946
rect 78206 52882 78258 52894
rect 77646 52834 77698 52846
rect 77646 52770 77698 52782
rect 1934 52722 1986 52734
rect 1934 52658 1986 52670
rect 1344 52554 78624 52588
rect 1344 52502 4478 52554
rect 4530 52502 4582 52554
rect 4634 52502 4686 52554
rect 4738 52502 35198 52554
rect 35250 52502 35302 52554
rect 35354 52502 35406 52554
rect 35458 52502 65918 52554
rect 65970 52502 66022 52554
rect 66074 52502 66126 52554
rect 66178 52502 78624 52554
rect 1344 52468 78624 52502
rect 1934 52274 1986 52286
rect 1934 52210 1986 52222
rect 3826 52110 3838 52162
rect 3890 52110 3902 52162
rect 1344 51770 78624 51804
rect 1344 51718 19838 51770
rect 19890 51718 19942 51770
rect 19994 51718 20046 51770
rect 20098 51718 50558 51770
rect 50610 51718 50662 51770
rect 50714 51718 50766 51770
rect 50818 51718 78624 51770
rect 1344 51684 78624 51718
rect 2494 51602 2546 51614
rect 2494 51538 2546 51550
rect 3502 51602 3554 51614
rect 3502 51538 3554 51550
rect 2830 51490 2882 51502
rect 2830 51426 2882 51438
rect 3838 51490 3890 51502
rect 3838 51426 3890 51438
rect 77870 51490 77922 51502
rect 77870 51426 77922 51438
rect 3166 51378 3218 51390
rect 2258 51326 2270 51378
rect 2322 51326 2334 51378
rect 3166 51314 3218 51326
rect 78206 51378 78258 51390
rect 78206 51314 78258 51326
rect 77646 51266 77698 51278
rect 77646 51202 77698 51214
rect 1344 50986 78624 51020
rect 1344 50934 4478 50986
rect 4530 50934 4582 50986
rect 4634 50934 4686 50986
rect 4738 50934 35198 50986
rect 35250 50934 35302 50986
rect 35354 50934 35406 50986
rect 35458 50934 65918 50986
rect 65970 50934 66022 50986
rect 66074 50934 66126 50986
rect 66178 50934 78624 50986
rect 1344 50900 78624 50934
rect 1934 50706 1986 50718
rect 1934 50642 1986 50654
rect 3826 50542 3838 50594
rect 3890 50542 3902 50594
rect 77646 50482 77698 50494
rect 77646 50418 77698 50430
rect 78206 50482 78258 50494
rect 78206 50418 78258 50430
rect 77870 50370 77922 50382
rect 77870 50306 77922 50318
rect 1344 50202 78624 50236
rect 1344 50150 19838 50202
rect 19890 50150 19942 50202
rect 19994 50150 20046 50202
rect 20098 50150 50558 50202
rect 50610 50150 50662 50202
rect 50714 50150 50766 50202
rect 50818 50150 78624 50202
rect 1344 50116 78624 50150
rect 3826 49758 3838 49810
rect 3890 49758 3902 49810
rect 1934 49586 1986 49598
rect 1934 49522 1986 49534
rect 1344 49418 78624 49452
rect 1344 49366 4478 49418
rect 4530 49366 4582 49418
rect 4634 49366 4686 49418
rect 4738 49366 35198 49418
rect 35250 49366 35302 49418
rect 35354 49366 35406 49418
rect 35458 49366 65918 49418
rect 65970 49366 66022 49418
rect 66074 49366 66126 49418
rect 66178 49366 78624 49418
rect 1344 49332 78624 49366
rect 1934 49138 1986 49150
rect 1934 49074 1986 49086
rect 3826 48974 3838 49026
rect 3890 48974 3902 49026
rect 77646 48914 77698 48926
rect 77646 48850 77698 48862
rect 78206 48914 78258 48926
rect 78206 48850 78258 48862
rect 77870 48802 77922 48814
rect 77870 48738 77922 48750
rect 1344 48634 78624 48668
rect 1344 48582 19838 48634
rect 19890 48582 19942 48634
rect 19994 48582 20046 48634
rect 20098 48582 50558 48634
rect 50610 48582 50662 48634
rect 50714 48582 50766 48634
rect 50818 48582 78624 48634
rect 1344 48548 78624 48582
rect 2718 48466 2770 48478
rect 2718 48402 2770 48414
rect 3390 48466 3442 48478
rect 3390 48402 3442 48414
rect 2046 48354 2098 48366
rect 2046 48290 2098 48302
rect 77870 48354 77922 48366
rect 77870 48290 77922 48302
rect 2382 48242 2434 48254
rect 78206 48242 78258 48254
rect 2930 48190 2942 48242
rect 2994 48190 3006 48242
rect 3602 48190 3614 48242
rect 3666 48190 3678 48242
rect 2382 48178 2434 48190
rect 78206 48178 78258 48190
rect 77646 48130 77698 48142
rect 77646 48066 77698 48078
rect 1344 47850 78624 47884
rect 1344 47798 4478 47850
rect 4530 47798 4582 47850
rect 4634 47798 4686 47850
rect 4738 47798 35198 47850
rect 35250 47798 35302 47850
rect 35354 47798 35406 47850
rect 35458 47798 65918 47850
rect 65970 47798 66022 47850
rect 66074 47798 66126 47850
rect 66178 47798 78624 47850
rect 1344 47764 78624 47798
rect 2034 47406 2046 47458
rect 2098 47406 2110 47458
rect 77646 47346 77698 47358
rect 77646 47282 77698 47294
rect 78206 47346 78258 47358
rect 78206 47282 78258 47294
rect 2718 47234 2770 47246
rect 2718 47170 2770 47182
rect 77870 47234 77922 47246
rect 77870 47170 77922 47182
rect 1344 47066 78624 47100
rect 1344 47014 19838 47066
rect 19890 47014 19942 47066
rect 19994 47014 20046 47066
rect 20098 47014 50558 47066
rect 50610 47014 50662 47066
rect 50714 47014 50766 47066
rect 50818 47014 78624 47066
rect 1344 46980 78624 47014
rect 3826 46622 3838 46674
rect 3890 46622 3902 46674
rect 1934 46450 1986 46462
rect 1934 46386 1986 46398
rect 1344 46282 78624 46316
rect 1344 46230 4478 46282
rect 4530 46230 4582 46282
rect 4634 46230 4686 46282
rect 4738 46230 35198 46282
rect 35250 46230 35302 46282
rect 35354 46230 35406 46282
rect 35458 46230 65918 46282
rect 65970 46230 66022 46282
rect 66074 46230 66126 46282
rect 66178 46230 78624 46282
rect 1344 46196 78624 46230
rect 2382 45890 2434 45902
rect 2818 45838 2830 45890
rect 2882 45838 2894 45890
rect 3602 45838 3614 45890
rect 3666 45838 3678 45890
rect 2382 45826 2434 45838
rect 3054 45778 3106 45790
rect 3054 45714 3106 45726
rect 3390 45778 3442 45790
rect 3390 45714 3442 45726
rect 4286 45778 4338 45790
rect 4286 45714 4338 45726
rect 78206 45778 78258 45790
rect 78206 45714 78258 45726
rect 2046 45666 2098 45678
rect 2046 45602 2098 45614
rect 77646 45666 77698 45678
rect 77646 45602 77698 45614
rect 77870 45666 77922 45678
rect 77870 45602 77922 45614
rect 1344 45498 78624 45532
rect 1344 45446 19838 45498
rect 19890 45446 19942 45498
rect 19994 45446 20046 45498
rect 20098 45446 50558 45498
rect 50610 45446 50662 45498
rect 50714 45446 50766 45498
rect 50818 45446 78624 45498
rect 1344 45412 78624 45446
rect 77870 45218 77922 45230
rect 77870 45154 77922 45166
rect 78206 45106 78258 45118
rect 2034 45054 2046 45106
rect 2098 45054 2110 45106
rect 78206 45042 78258 45054
rect 77646 44994 77698 45006
rect 77646 44930 77698 44942
rect 2718 44882 2770 44894
rect 2718 44818 2770 44830
rect 1344 44714 78624 44748
rect 1344 44662 4478 44714
rect 4530 44662 4582 44714
rect 4634 44662 4686 44714
rect 4738 44662 35198 44714
rect 35250 44662 35302 44714
rect 35354 44662 35406 44714
rect 35458 44662 65918 44714
rect 65970 44662 66022 44714
rect 66074 44662 66126 44714
rect 66178 44662 78624 44714
rect 1344 44628 78624 44662
rect 2034 44270 2046 44322
rect 2098 44270 2110 44322
rect 2718 44098 2770 44110
rect 2718 44034 2770 44046
rect 77982 44098 78034 44110
rect 77982 44034 78034 44046
rect 1344 43930 78624 43964
rect 1344 43878 19838 43930
rect 19890 43878 19942 43930
rect 19994 43878 20046 43930
rect 20098 43878 50558 43930
rect 50610 43878 50662 43930
rect 50714 43878 50766 43930
rect 50818 43878 78624 43930
rect 1344 43844 78624 43878
rect 2046 43762 2098 43774
rect 2046 43698 2098 43710
rect 2718 43650 2770 43662
rect 2718 43586 2770 43598
rect 77870 43650 77922 43662
rect 77870 43586 77922 43598
rect 77086 43538 77138 43550
rect 2258 43486 2270 43538
rect 2322 43486 2334 43538
rect 2930 43486 2942 43538
rect 2994 43486 3006 43538
rect 77086 43474 77138 43486
rect 78206 43538 78258 43550
rect 78206 43474 78258 43486
rect 77646 43426 77698 43438
rect 77646 43362 77698 43374
rect 1344 43146 78624 43180
rect 1344 43094 4478 43146
rect 4530 43094 4582 43146
rect 4634 43094 4686 43146
rect 4738 43094 35198 43146
rect 35250 43094 35302 43146
rect 35354 43094 35406 43146
rect 35458 43094 65918 43146
rect 65970 43094 66022 43146
rect 66074 43094 66126 43146
rect 66178 43094 78624 43146
rect 1344 43060 78624 43094
rect 1934 42866 1986 42878
rect 1934 42802 1986 42814
rect 55806 42866 55858 42878
rect 55806 42802 55858 42814
rect 56702 42866 56754 42878
rect 56702 42802 56754 42814
rect 57598 42866 57650 42878
rect 57598 42802 57650 42814
rect 58494 42866 58546 42878
rect 58494 42802 58546 42814
rect 62414 42866 62466 42878
rect 62414 42802 62466 42814
rect 75294 42866 75346 42878
rect 75294 42802 75346 42814
rect 76526 42866 76578 42878
rect 76526 42802 76578 42814
rect 76750 42754 76802 42766
rect 3826 42702 3838 42754
rect 3890 42702 3902 42754
rect 57138 42702 57150 42754
rect 57202 42702 57214 42754
rect 58034 42702 58046 42754
rect 58098 42702 58110 42754
rect 76750 42690 76802 42702
rect 77086 42754 77138 42766
rect 77086 42690 77138 42702
rect 77422 42642 77474 42654
rect 77422 42578 77474 42590
rect 77758 42642 77810 42654
rect 77758 42578 77810 42590
rect 55246 42530 55298 42542
rect 55246 42466 55298 42478
rect 56142 42530 56194 42542
rect 56142 42466 56194 42478
rect 77086 42530 77138 42542
rect 77086 42466 77138 42478
rect 78094 42530 78146 42542
rect 78094 42466 78146 42478
rect 1344 42362 78624 42396
rect 1344 42310 19838 42362
rect 19890 42310 19942 42362
rect 19994 42310 20046 42362
rect 20098 42310 50558 42362
rect 50610 42310 50662 42362
rect 50714 42310 50766 42362
rect 50818 42310 78624 42362
rect 1344 42276 78624 42310
rect 55010 42142 55022 42194
rect 55074 42142 55086 42194
rect 57138 42142 57150 42194
rect 57202 42142 57214 42194
rect 58034 42142 58046 42194
rect 58098 42142 58110 42194
rect 62862 42082 62914 42094
rect 62862 42018 62914 42030
rect 75294 42082 75346 42094
rect 75294 42018 75346 42030
rect 4734 41970 4786 41982
rect 3826 41918 3838 41970
rect 3890 41918 3902 41970
rect 4734 41906 4786 41918
rect 61630 41970 61682 41982
rect 61630 41906 61682 41918
rect 62750 41970 62802 41982
rect 62750 41906 62802 41918
rect 63310 41970 63362 41982
rect 63310 41906 63362 41918
rect 64542 41970 64594 41982
rect 64542 41906 64594 41918
rect 73950 41970 74002 41982
rect 73950 41906 74002 41918
rect 74958 41970 75010 41982
rect 75618 41918 75630 41970
rect 75682 41918 75694 41970
rect 74958 41906 75010 41918
rect 55582 41858 55634 41870
rect 55582 41794 55634 41806
rect 56142 41858 56194 41870
rect 56142 41794 56194 41806
rect 56590 41858 56642 41870
rect 56590 41794 56642 41806
rect 57486 41858 57538 41870
rect 57486 41794 57538 41806
rect 62190 41858 62242 41870
rect 62190 41794 62242 41806
rect 63086 41858 63138 41870
rect 63086 41794 63138 41806
rect 63646 41858 63698 41870
rect 63646 41794 63698 41806
rect 70590 41858 70642 41870
rect 70590 41794 70642 41806
rect 71038 41858 71090 41870
rect 71038 41794 71090 41806
rect 74734 41858 74786 41870
rect 74734 41794 74786 41806
rect 77982 41858 78034 41870
rect 77982 41794 78034 41806
rect 1934 41746 1986 41758
rect 1934 41682 1986 41694
rect 55358 41746 55410 41758
rect 56814 41746 56866 41758
rect 55794 41694 55806 41746
rect 55858 41743 55870 41746
rect 56018 41743 56030 41746
rect 55858 41697 56030 41743
rect 55858 41694 55870 41697
rect 56018 41694 56030 41697
rect 56082 41694 56094 41746
rect 55358 41682 55410 41694
rect 56814 41682 56866 41694
rect 57710 41746 57762 41758
rect 57710 41682 57762 41694
rect 1344 41578 78624 41612
rect 1344 41526 4478 41578
rect 4530 41526 4582 41578
rect 4634 41526 4686 41578
rect 4738 41526 35198 41578
rect 35250 41526 35302 41578
rect 35354 41526 35406 41578
rect 35458 41526 65918 41578
rect 65970 41526 66022 41578
rect 66074 41526 66126 41578
rect 66178 41526 78624 41578
rect 1344 41492 78624 41526
rect 55470 41410 55522 41422
rect 71374 41410 71426 41422
rect 55794 41358 55806 41410
rect 55858 41358 55870 41410
rect 74610 41358 74622 41410
rect 74674 41358 74686 41410
rect 75506 41358 75518 41410
rect 75570 41358 75582 41410
rect 55470 41346 55522 41358
rect 71374 41346 71426 41358
rect 1934 41298 1986 41310
rect 1934 41234 1986 41246
rect 4734 41298 4786 41310
rect 4734 41234 4786 41246
rect 57150 41298 57202 41310
rect 57150 41234 57202 41246
rect 61518 41298 61570 41310
rect 61518 41234 61570 41246
rect 65326 41298 65378 41310
rect 71486 41298 71538 41310
rect 70802 41246 70814 41298
rect 70866 41246 70878 41298
rect 65326 41234 65378 41246
rect 71486 41234 71538 41246
rect 71934 41298 71986 41310
rect 71934 41234 71986 41246
rect 72046 41298 72098 41310
rect 72046 41234 72098 41246
rect 75182 41298 75234 41310
rect 75182 41234 75234 41246
rect 78094 41298 78146 41310
rect 78094 41234 78146 41246
rect 55246 41186 55298 41198
rect 4050 41134 4062 41186
rect 4114 41134 4126 41186
rect 55246 41122 55298 41134
rect 60510 41186 60562 41198
rect 60510 41122 60562 41134
rect 61854 41186 61906 41198
rect 61854 41122 61906 41134
rect 62190 41186 62242 41198
rect 62190 41122 62242 41134
rect 62414 41186 62466 41198
rect 64878 41186 64930 41198
rect 71710 41186 71762 41198
rect 62962 41134 62974 41186
rect 63026 41134 63038 41186
rect 63298 41134 63310 41186
rect 63362 41134 63374 41186
rect 64418 41134 64430 41186
rect 64482 41134 64494 41186
rect 65650 41134 65662 41186
rect 65714 41134 65726 41186
rect 66770 41134 66782 41186
rect 66834 41134 66846 41186
rect 62414 41122 62466 41134
rect 64878 41122 64930 41134
rect 71710 41122 71762 41134
rect 73502 41186 73554 41198
rect 73502 41122 73554 41134
rect 74062 41186 74114 41198
rect 74062 41122 74114 41134
rect 74286 41186 74338 41198
rect 74286 41122 74338 41134
rect 74958 41186 75010 41198
rect 74958 41122 75010 41134
rect 76414 41186 76466 41198
rect 76414 41122 76466 41134
rect 76750 41186 76802 41198
rect 76750 41122 76802 41134
rect 77422 41186 77474 41198
rect 77422 41122 77474 41134
rect 58382 41074 58434 41086
rect 58382 41010 58434 41022
rect 58718 41074 58770 41086
rect 58718 41010 58770 41022
rect 61070 41074 61122 41086
rect 73166 41074 73218 41086
rect 63410 41022 63422 41074
rect 63474 41022 63486 41074
rect 65762 41022 65774 41074
rect 65826 41022 65838 41074
rect 69570 41022 69582 41074
rect 69634 41022 69646 41074
rect 61070 41010 61122 41022
rect 73166 41010 73218 41022
rect 73726 41074 73778 41086
rect 73726 41010 73778 41022
rect 76190 41074 76242 41086
rect 76190 41010 76242 41022
rect 77086 41074 77138 41086
rect 77086 41010 77138 41022
rect 77646 41074 77698 41086
rect 77646 41010 77698 41022
rect 54910 40962 54962 40974
rect 54910 40898 54962 40910
rect 56254 40962 56306 40974
rect 56254 40898 56306 40910
rect 62078 40962 62130 40974
rect 69022 40962 69074 40974
rect 62962 40910 62974 40962
rect 63026 40910 63038 40962
rect 66658 40910 66670 40962
rect 66722 40910 66734 40962
rect 62078 40898 62130 40910
rect 69022 40898 69074 40910
rect 69246 40962 69298 40974
rect 69246 40898 69298 40910
rect 70030 40962 70082 40974
rect 70030 40898 70082 40910
rect 70366 40962 70418 40974
rect 70366 40898 70418 40910
rect 73390 40962 73442 40974
rect 73390 40898 73442 40910
rect 76638 40962 76690 40974
rect 76638 40898 76690 40910
rect 77198 40962 77250 40974
rect 77198 40898 77250 40910
rect 1344 40794 78624 40828
rect 1344 40742 19838 40794
rect 19890 40742 19942 40794
rect 19994 40742 20046 40794
rect 20098 40742 50558 40794
rect 50610 40742 50662 40794
rect 50714 40742 50766 40794
rect 50818 40742 78624 40794
rect 1344 40708 78624 40742
rect 2270 40626 2322 40638
rect 67454 40626 67506 40638
rect 69582 40626 69634 40638
rect 63522 40574 63534 40626
rect 63586 40574 63598 40626
rect 68338 40574 68350 40626
rect 68402 40574 68414 40626
rect 2270 40562 2322 40574
rect 67454 40562 67506 40574
rect 69582 40562 69634 40574
rect 70254 40626 70306 40638
rect 74610 40574 74622 40626
rect 74674 40574 74686 40626
rect 70254 40562 70306 40574
rect 4062 40514 4114 40526
rect 4062 40450 4114 40462
rect 4510 40514 4562 40526
rect 67902 40514 67954 40526
rect 59826 40462 59838 40514
rect 59890 40462 59902 40514
rect 61506 40462 61518 40514
rect 61570 40462 61582 40514
rect 62514 40462 62526 40514
rect 62578 40462 62590 40514
rect 65090 40462 65102 40514
rect 65154 40462 65166 40514
rect 66322 40462 66334 40514
rect 66386 40462 66398 40514
rect 4510 40450 4562 40462
rect 67902 40450 67954 40462
rect 75294 40514 75346 40526
rect 76514 40462 76526 40514
rect 76578 40462 76590 40514
rect 75294 40450 75346 40462
rect 1710 40402 1762 40414
rect 1710 40338 1762 40350
rect 2606 40402 2658 40414
rect 2606 40338 2658 40350
rect 3166 40402 3218 40414
rect 3166 40338 3218 40350
rect 3502 40402 3554 40414
rect 3502 40338 3554 40350
rect 4958 40402 5010 40414
rect 4958 40338 5010 40350
rect 5406 40402 5458 40414
rect 69134 40402 69186 40414
rect 74286 40402 74338 40414
rect 60050 40350 60062 40402
rect 60114 40350 60126 40402
rect 60722 40350 60734 40402
rect 60786 40350 60798 40402
rect 61058 40350 61070 40402
rect 61122 40350 61134 40402
rect 62178 40350 62190 40402
rect 62242 40350 62254 40402
rect 63074 40350 63086 40402
rect 63138 40350 63150 40402
rect 63410 40350 63422 40402
rect 63474 40350 63486 40402
rect 64418 40350 64430 40402
rect 64482 40350 64494 40402
rect 65538 40350 65550 40402
rect 65602 40350 65614 40402
rect 65874 40350 65886 40402
rect 65938 40350 65950 40402
rect 66770 40350 66782 40402
rect 66834 40350 66846 40402
rect 68562 40350 68574 40402
rect 68626 40350 68638 40402
rect 73154 40350 73166 40402
rect 73218 40350 73230 40402
rect 73602 40350 73614 40402
rect 73666 40350 73678 40402
rect 75058 40350 75070 40402
rect 75122 40350 75134 40402
rect 78194 40350 78206 40402
rect 78258 40350 78270 40402
rect 5406 40338 5458 40350
rect 69134 40338 69186 40350
rect 74286 40338 74338 40350
rect 70702 40290 70754 40302
rect 60162 40238 60174 40290
rect 60226 40238 60238 40290
rect 61394 40238 61406 40290
rect 61458 40238 61470 40290
rect 64866 40238 64878 40290
rect 64930 40238 64942 40290
rect 66434 40238 66446 40290
rect 66498 40238 66510 40290
rect 73378 40238 73390 40290
rect 73442 40238 73454 40290
rect 70702 40226 70754 40238
rect 72930 40126 72942 40178
rect 72994 40126 73006 40178
rect 1344 40010 78624 40044
rect 1344 39958 4478 40010
rect 4530 39958 4582 40010
rect 4634 39958 4686 40010
rect 4738 39958 35198 40010
rect 35250 39958 35302 40010
rect 35354 39958 35406 40010
rect 35458 39958 65918 40010
rect 65970 39958 66022 40010
rect 66074 39958 66126 40010
rect 66178 39958 78624 40010
rect 1344 39924 78624 39958
rect 1934 39730 1986 39742
rect 1934 39666 1986 39678
rect 62302 39730 62354 39742
rect 62302 39666 62354 39678
rect 62638 39730 62690 39742
rect 67118 39730 67170 39742
rect 71374 39730 71426 39742
rect 63186 39678 63198 39730
rect 63250 39678 63262 39730
rect 66210 39678 66222 39730
rect 66274 39678 66286 39730
rect 69010 39678 69022 39730
rect 69074 39678 69086 39730
rect 62638 39666 62690 39678
rect 67118 39666 67170 39678
rect 71374 39666 71426 39678
rect 71822 39730 71874 39742
rect 71822 39666 71874 39678
rect 73166 39730 73218 39742
rect 73166 39666 73218 39678
rect 74622 39730 74674 39742
rect 77982 39730 78034 39742
rect 76738 39678 76750 39730
rect 76802 39678 76814 39730
rect 74622 39666 74674 39678
rect 77982 39666 78034 39678
rect 4734 39618 4786 39630
rect 70254 39618 70306 39630
rect 3826 39566 3838 39618
rect 3890 39566 3902 39618
rect 60722 39566 60734 39618
rect 60786 39566 60798 39618
rect 61058 39566 61070 39618
rect 61122 39566 61134 39618
rect 65650 39566 65662 39618
rect 65714 39566 65726 39618
rect 66098 39566 66110 39618
rect 66162 39566 66174 39618
rect 68562 39566 68574 39618
rect 68626 39566 68638 39618
rect 69570 39566 69582 39618
rect 69634 39566 69646 39618
rect 4734 39554 4786 39566
rect 70254 39554 70306 39566
rect 70702 39618 70754 39630
rect 70702 39554 70754 39566
rect 72830 39618 72882 39630
rect 72830 39554 72882 39566
rect 72942 39618 72994 39630
rect 72942 39554 72994 39566
rect 74958 39618 75010 39630
rect 74958 39554 75010 39566
rect 75406 39618 75458 39630
rect 75406 39554 75458 39566
rect 75630 39618 75682 39630
rect 76514 39566 76526 39618
rect 76578 39566 76590 39618
rect 77298 39566 77310 39618
rect 77362 39566 77374 39618
rect 75630 39554 75682 39566
rect 70926 39506 70978 39518
rect 61170 39454 61182 39506
rect 61234 39454 61246 39506
rect 63970 39454 63982 39506
rect 64034 39454 64046 39506
rect 66546 39454 66558 39506
rect 66610 39454 66622 39506
rect 69234 39454 69246 39506
rect 69298 39454 69310 39506
rect 70926 39442 70978 39454
rect 73278 39506 73330 39518
rect 73278 39442 73330 39454
rect 73838 39506 73890 39518
rect 73838 39442 73890 39454
rect 74174 39506 74226 39518
rect 77870 39506 77922 39518
rect 76178 39454 76190 39506
rect 76242 39454 76254 39506
rect 74174 39442 74226 39454
rect 77870 39442 77922 39454
rect 78094 39506 78146 39518
rect 78094 39442 78146 39454
rect 63646 39394 63698 39406
rect 60610 39342 60622 39394
rect 60674 39342 60686 39394
rect 63646 39330 63698 39342
rect 64318 39394 64370 39406
rect 64318 39330 64370 39342
rect 67566 39394 67618 39406
rect 67566 39330 67618 39342
rect 70478 39394 70530 39406
rect 70478 39330 70530 39342
rect 72382 39394 72434 39406
rect 72382 39330 72434 39342
rect 75294 39394 75346 39406
rect 75294 39330 75346 39342
rect 1344 39226 78624 39260
rect 1344 39174 19838 39226
rect 19890 39174 19942 39226
rect 19994 39174 20046 39226
rect 20098 39174 50558 39226
rect 50610 39174 50662 39226
rect 50714 39174 50766 39226
rect 50818 39174 78624 39226
rect 1344 39140 78624 39174
rect 41134 39058 41186 39070
rect 41134 38994 41186 39006
rect 42926 39058 42978 39070
rect 42926 38994 42978 39006
rect 43262 39058 43314 39070
rect 43262 38994 43314 39006
rect 60958 39058 61010 39070
rect 60958 38994 61010 39006
rect 63310 39058 63362 39070
rect 63310 38994 63362 39006
rect 72830 39058 72882 39070
rect 72830 38994 72882 39006
rect 75966 39058 76018 39070
rect 75966 38994 76018 39006
rect 78206 39058 78258 39070
rect 78206 38994 78258 39006
rect 41246 38946 41298 38958
rect 42702 38946 42754 38958
rect 71374 38946 71426 38958
rect 42242 38894 42254 38946
rect 42306 38894 42318 38946
rect 66994 38894 67006 38946
rect 67058 38894 67070 38946
rect 67666 38894 67678 38946
rect 67730 38894 67742 38946
rect 69906 38894 69918 38946
rect 69970 38894 69982 38946
rect 41246 38882 41298 38894
rect 42702 38882 42754 38894
rect 71374 38882 71426 38894
rect 72494 38946 72546 38958
rect 72494 38882 72546 38894
rect 73166 38946 73218 38958
rect 73166 38882 73218 38894
rect 73502 38946 73554 38958
rect 73502 38882 73554 38894
rect 74510 38946 74562 38958
rect 74510 38882 74562 38894
rect 75406 38946 75458 38958
rect 75406 38882 75458 38894
rect 76526 38946 76578 38958
rect 76526 38882 76578 38894
rect 77534 38946 77586 38958
rect 77534 38882 77586 38894
rect 40910 38834 40962 38846
rect 42590 38834 42642 38846
rect 2034 38782 2046 38834
rect 2098 38782 2110 38834
rect 41682 38782 41694 38834
rect 41746 38782 41758 38834
rect 40910 38770 40962 38782
rect 42590 38770 42642 38782
rect 43710 38834 43762 38846
rect 65214 38834 65266 38846
rect 63522 38782 63534 38834
rect 63586 38782 63598 38834
rect 43710 38770 43762 38782
rect 65214 38770 65266 38782
rect 65774 38834 65826 38846
rect 70366 38834 70418 38846
rect 66098 38782 66110 38834
rect 66162 38782 66174 38834
rect 67218 38782 67230 38834
rect 67282 38782 67294 38834
rect 68114 38782 68126 38834
rect 68178 38782 68190 38834
rect 68562 38782 68574 38834
rect 68626 38782 68638 38834
rect 69010 38782 69022 38834
rect 69074 38782 69086 38834
rect 69570 38782 69582 38834
rect 69634 38782 69646 38834
rect 65774 38770 65826 38782
rect 70366 38770 70418 38782
rect 70702 38834 70754 38846
rect 70702 38770 70754 38782
rect 70926 38834 70978 38846
rect 74174 38834 74226 38846
rect 71586 38782 71598 38834
rect 71650 38782 71662 38834
rect 70926 38770 70978 38782
rect 74174 38770 74226 38782
rect 74734 38834 74786 38846
rect 74734 38770 74786 38782
rect 75070 38834 75122 38846
rect 75070 38770 75122 38782
rect 76302 38834 76354 38846
rect 76302 38770 76354 38782
rect 76974 38834 77026 38846
rect 76974 38770 77026 38782
rect 77086 38834 77138 38846
rect 77086 38770 77138 38782
rect 77646 38834 77698 38846
rect 77646 38770 77698 38782
rect 62974 38722 63026 38734
rect 70590 38722 70642 38734
rect 3378 38670 3390 38722
rect 3442 38670 3454 38722
rect 41570 38670 41582 38722
rect 41634 38670 41646 38722
rect 66546 38670 66558 38722
rect 66610 38670 66622 38722
rect 67666 38670 67678 38722
rect 67730 38670 67742 38722
rect 69458 38670 69470 38722
rect 69522 38670 69534 38722
rect 62974 38658 63026 38670
rect 70590 38658 70642 38670
rect 74958 38722 75010 38734
rect 74958 38658 75010 38670
rect 76750 38722 76802 38734
rect 76750 38658 76802 38670
rect 77310 38722 77362 38734
rect 77310 38658 77362 38670
rect 1344 38442 78624 38476
rect 1344 38390 4478 38442
rect 4530 38390 4582 38442
rect 4634 38390 4686 38442
rect 4738 38390 35198 38442
rect 35250 38390 35302 38442
rect 35354 38390 35406 38442
rect 35458 38390 65918 38442
rect 65970 38390 66022 38442
rect 66074 38390 66126 38442
rect 66178 38390 78624 38442
rect 1344 38356 78624 38390
rect 77310 38274 77362 38286
rect 72706 38222 72718 38274
rect 72770 38271 72782 38274
rect 73266 38271 73278 38274
rect 72770 38225 73278 38271
rect 72770 38222 72782 38225
rect 73266 38222 73278 38225
rect 73330 38222 73342 38274
rect 77310 38210 77362 38222
rect 2942 38162 2994 38174
rect 2034 38110 2046 38162
rect 2098 38110 2110 38162
rect 2942 38098 2994 38110
rect 41470 38162 41522 38174
rect 69918 38162 69970 38174
rect 67330 38110 67342 38162
rect 67394 38110 67406 38162
rect 41470 38098 41522 38110
rect 69918 38098 69970 38110
rect 72158 38162 72210 38174
rect 72158 38098 72210 38110
rect 72606 38162 72658 38174
rect 72606 38098 72658 38110
rect 75742 38162 75794 38174
rect 77982 38162 78034 38174
rect 76402 38110 76414 38162
rect 76466 38110 76478 38162
rect 75742 38098 75794 38110
rect 77982 38098 78034 38110
rect 2494 38050 2546 38062
rect 66558 38050 66610 38062
rect 70254 38050 70306 38062
rect 66098 37998 66110 38050
rect 66162 37998 66174 38050
rect 68338 37998 68350 38050
rect 68402 37998 68414 38050
rect 69346 37998 69358 38050
rect 69410 37998 69422 38050
rect 2494 37986 2546 37998
rect 66558 37986 66610 37998
rect 70254 37986 70306 37998
rect 70590 38050 70642 38062
rect 70590 37986 70642 37998
rect 70814 38050 70866 38062
rect 70814 37986 70866 37998
rect 71150 38050 71202 38062
rect 71150 37986 71202 37998
rect 71374 38050 71426 38062
rect 71374 37986 71426 37998
rect 73054 38050 73106 38062
rect 73054 37986 73106 37998
rect 74510 38050 74562 38062
rect 74510 37986 74562 37998
rect 74846 38050 74898 38062
rect 74846 37986 74898 37998
rect 75070 38050 75122 38062
rect 77186 37998 77198 38050
rect 77250 37998 77262 38050
rect 77522 37998 77534 38050
rect 77586 37998 77598 38050
rect 75070 37986 75122 37998
rect 71710 37938 71762 37950
rect 69234 37886 69246 37938
rect 69298 37886 69310 37938
rect 71710 37874 71762 37886
rect 73838 37938 73890 37950
rect 73838 37874 73890 37886
rect 74174 37938 74226 37950
rect 74174 37874 74226 37886
rect 76190 37938 76242 37950
rect 76190 37874 76242 37886
rect 67790 37826 67842 37838
rect 70366 37826 70418 37838
rect 68562 37774 68574 37826
rect 68626 37774 68638 37826
rect 67790 37762 67842 37774
rect 70366 37762 70418 37774
rect 71598 37826 71650 37838
rect 71598 37762 71650 37774
rect 73502 37826 73554 37838
rect 73502 37762 73554 37774
rect 74622 37826 74674 37838
rect 74622 37762 74674 37774
rect 76414 37826 76466 37838
rect 76414 37762 76466 37774
rect 1344 37658 78624 37692
rect 1344 37606 19838 37658
rect 19890 37606 19942 37658
rect 19994 37606 20046 37658
rect 20098 37606 50558 37658
rect 50610 37606 50662 37658
rect 50714 37606 50766 37658
rect 50818 37606 78624 37658
rect 1344 37572 78624 37606
rect 68462 37490 68514 37502
rect 68462 37426 68514 37438
rect 69470 37490 69522 37502
rect 71150 37490 71202 37502
rect 76414 37490 76466 37502
rect 69794 37438 69806 37490
rect 69858 37438 69870 37490
rect 70802 37438 70814 37490
rect 70866 37438 70878 37490
rect 71474 37438 71486 37490
rect 71538 37438 71550 37490
rect 69470 37426 69522 37438
rect 71150 37426 71202 37438
rect 76414 37426 76466 37438
rect 72270 37378 72322 37390
rect 2034 37326 2046 37378
rect 2098 37326 2110 37378
rect 72270 37314 72322 37326
rect 72830 37378 72882 37390
rect 72830 37314 72882 37326
rect 73726 37378 73778 37390
rect 73726 37314 73778 37326
rect 74062 37378 74114 37390
rect 74062 37314 74114 37326
rect 75630 37378 75682 37390
rect 75630 37314 75682 37326
rect 76190 37378 76242 37390
rect 76190 37314 76242 37326
rect 1710 37266 1762 37278
rect 69134 37266 69186 37278
rect 72494 37266 72546 37278
rect 68674 37214 68686 37266
rect 68738 37214 68750 37266
rect 70018 37214 70030 37266
rect 70082 37214 70094 37266
rect 70578 37214 70590 37266
rect 70642 37214 70654 37266
rect 1710 37202 1762 37214
rect 69134 37202 69186 37214
rect 72494 37202 72546 37214
rect 73054 37266 73106 37278
rect 73054 37202 73106 37214
rect 73390 37266 73442 37278
rect 73390 37202 73442 37214
rect 74286 37266 74338 37278
rect 74286 37202 74338 37214
rect 74622 37266 74674 37278
rect 74622 37202 74674 37214
rect 75070 37266 75122 37278
rect 75070 37202 75122 37214
rect 75406 37266 75458 37278
rect 75406 37202 75458 37214
rect 76078 37266 76130 37278
rect 76078 37202 76130 37214
rect 76526 37266 76578 37278
rect 77298 37214 77310 37266
rect 77362 37214 77374 37266
rect 77858 37214 77870 37266
rect 77922 37214 77934 37266
rect 76526 37202 76578 37214
rect 2494 37154 2546 37166
rect 2494 37090 2546 37102
rect 68126 37154 68178 37166
rect 68126 37090 68178 37102
rect 72382 37154 72434 37166
rect 72382 37090 72434 37102
rect 73278 37154 73330 37166
rect 73278 37090 73330 37102
rect 74510 37154 74562 37166
rect 74510 37090 74562 37102
rect 75182 37154 75234 37166
rect 77410 37102 77422 37154
rect 77474 37102 77486 37154
rect 75182 37090 75234 37102
rect 77522 36990 77534 37042
rect 77586 36990 77598 37042
rect 1344 36874 78624 36908
rect 1344 36822 4478 36874
rect 4530 36822 4582 36874
rect 4634 36822 4686 36874
rect 4738 36822 35198 36874
rect 35250 36822 35302 36874
rect 35354 36822 35406 36874
rect 35458 36822 65918 36874
rect 65970 36822 66022 36874
rect 66074 36822 66126 36874
rect 66178 36822 78624 36874
rect 1344 36788 78624 36822
rect 76302 36706 76354 36718
rect 76302 36642 76354 36654
rect 68798 36594 68850 36606
rect 68798 36530 68850 36542
rect 71262 36594 71314 36606
rect 71262 36530 71314 36542
rect 71710 36594 71762 36606
rect 71710 36530 71762 36542
rect 72606 36594 72658 36606
rect 72606 36530 72658 36542
rect 73838 36594 73890 36606
rect 73838 36530 73890 36542
rect 74398 36594 74450 36606
rect 74398 36530 74450 36542
rect 75518 36594 75570 36606
rect 77074 36542 77086 36594
rect 77138 36542 77150 36594
rect 75518 36530 75570 36542
rect 69694 36482 69746 36494
rect 69694 36418 69746 36430
rect 72158 36482 72210 36494
rect 72158 36418 72210 36430
rect 72830 36482 72882 36494
rect 72830 36418 72882 36430
rect 73166 36482 73218 36494
rect 73166 36418 73218 36430
rect 73390 36482 73442 36494
rect 74722 36430 74734 36482
rect 74786 36430 74798 36482
rect 75282 36430 75294 36482
rect 75346 36430 75358 36482
rect 76514 36430 76526 36482
rect 76578 36430 76590 36482
rect 76850 36430 76862 36482
rect 76914 36430 76926 36482
rect 73390 36418 73442 36430
rect 1710 36370 1762 36382
rect 1710 36306 1762 36318
rect 45054 36370 45106 36382
rect 45054 36306 45106 36318
rect 45614 36370 45666 36382
rect 45614 36306 45666 36318
rect 74958 36370 75010 36382
rect 74958 36306 75010 36318
rect 75630 36370 75682 36382
rect 75630 36306 75682 36318
rect 77870 36370 77922 36382
rect 77870 36306 77922 36318
rect 78206 36370 78258 36382
rect 78206 36306 78258 36318
rect 2046 36258 2098 36270
rect 2046 36194 2098 36206
rect 2494 36258 2546 36270
rect 2494 36194 2546 36206
rect 45166 36258 45218 36270
rect 45166 36194 45218 36206
rect 73054 36258 73106 36270
rect 73054 36194 73106 36206
rect 1344 36090 78624 36124
rect 1344 36038 19838 36090
rect 19890 36038 19942 36090
rect 19994 36038 20046 36090
rect 20098 36038 50558 36090
rect 50610 36038 50662 36090
rect 50714 36038 50766 36090
rect 50818 36038 78624 36090
rect 1344 36004 78624 36038
rect 44718 35922 44770 35934
rect 44718 35858 44770 35870
rect 56814 35922 56866 35934
rect 56814 35858 56866 35870
rect 71374 35922 71426 35934
rect 71374 35858 71426 35870
rect 72606 35922 72658 35934
rect 72606 35858 72658 35870
rect 74286 35922 74338 35934
rect 74286 35858 74338 35870
rect 77310 35922 77362 35934
rect 77310 35858 77362 35870
rect 77982 35922 78034 35934
rect 77982 35858 78034 35870
rect 45054 35810 45106 35822
rect 74174 35810 74226 35822
rect 54226 35758 54238 35810
rect 54290 35758 54302 35810
rect 55346 35758 55358 35810
rect 55410 35758 55422 35810
rect 72930 35758 72942 35810
rect 72994 35758 73006 35810
rect 45054 35746 45106 35758
rect 74174 35746 74226 35758
rect 75182 35810 75234 35822
rect 75182 35746 75234 35758
rect 76302 35810 76354 35822
rect 76302 35746 76354 35758
rect 76974 35810 77026 35822
rect 76974 35746 77026 35758
rect 77534 35810 77586 35822
rect 77534 35746 77586 35758
rect 78094 35810 78146 35822
rect 78094 35746 78146 35758
rect 45726 35698 45778 35710
rect 45726 35634 45778 35646
rect 45950 35698 46002 35710
rect 45950 35634 46002 35646
rect 46174 35698 46226 35710
rect 46174 35634 46226 35646
rect 46398 35698 46450 35710
rect 72270 35698 72322 35710
rect 74062 35698 74114 35710
rect 54002 35646 54014 35698
rect 54066 35646 54078 35698
rect 55010 35646 55022 35698
rect 55074 35646 55086 35698
rect 73154 35646 73166 35698
rect 73218 35646 73230 35698
rect 46398 35634 46450 35646
rect 72270 35634 72322 35646
rect 74062 35634 74114 35646
rect 74622 35698 74674 35710
rect 74622 35634 74674 35646
rect 74734 35698 74786 35710
rect 74734 35634 74786 35646
rect 75406 35698 75458 35710
rect 75406 35634 75458 35646
rect 76078 35698 76130 35710
rect 76078 35634 76130 35646
rect 76750 35698 76802 35710
rect 76750 35634 76802 35646
rect 77310 35698 77362 35710
rect 77310 35634 77362 35646
rect 71710 35586 71762 35598
rect 54674 35534 54686 35586
rect 54738 35534 54750 35586
rect 55682 35534 55694 35586
rect 55746 35534 55758 35586
rect 71710 35522 71762 35534
rect 74958 35586 75010 35598
rect 74958 35522 75010 35534
rect 76526 35586 76578 35598
rect 76526 35522 76578 35534
rect 45166 35474 45218 35486
rect 45166 35410 45218 35422
rect 77870 35474 77922 35486
rect 77870 35410 77922 35422
rect 1344 35306 78624 35340
rect 1344 35254 4478 35306
rect 4530 35254 4582 35306
rect 4634 35254 4686 35306
rect 4738 35254 35198 35306
rect 35250 35254 35302 35306
rect 35354 35254 35406 35306
rect 35458 35254 65918 35306
rect 65970 35254 66022 35306
rect 66074 35254 66126 35306
rect 66178 35254 78624 35306
rect 1344 35220 78624 35254
rect 55022 35026 55074 35038
rect 55022 34962 55074 34974
rect 55358 35026 55410 35038
rect 55358 34962 55410 34974
rect 72606 35026 72658 35038
rect 76290 34974 76302 35026
rect 76354 34974 76366 35026
rect 77186 34974 77198 35026
rect 77250 34974 77262 35026
rect 72606 34962 72658 34974
rect 45726 34914 45778 34926
rect 45726 34850 45778 34862
rect 46174 34914 46226 34926
rect 46174 34850 46226 34862
rect 46622 34914 46674 34926
rect 46622 34850 46674 34862
rect 46846 34914 46898 34926
rect 46846 34850 46898 34862
rect 46958 34914 47010 34926
rect 46958 34850 47010 34862
rect 47182 34914 47234 34926
rect 72830 34914 72882 34926
rect 53890 34862 53902 34914
rect 53954 34862 53966 34914
rect 47182 34850 47234 34862
rect 72830 34850 72882 34862
rect 73278 34914 73330 34926
rect 77870 34914 77922 34926
rect 73938 34862 73950 34914
rect 74002 34862 74014 34914
rect 74834 34862 74846 34914
rect 74898 34862 74910 34914
rect 75394 34862 75406 34914
rect 75458 34862 75470 34914
rect 76178 34862 76190 34914
rect 76242 34862 76254 34914
rect 76850 34862 76862 34914
rect 76914 34862 76926 34914
rect 73278 34850 73330 34862
rect 77870 34850 77922 34862
rect 1710 34802 1762 34814
rect 1710 34738 1762 34750
rect 2494 34802 2546 34814
rect 2494 34738 2546 34750
rect 45166 34802 45218 34814
rect 45166 34738 45218 34750
rect 45278 34802 45330 34814
rect 45278 34738 45330 34750
rect 46398 34802 46450 34814
rect 73502 34802 73554 34814
rect 78206 34802 78258 34814
rect 53778 34750 53790 34802
rect 53842 34750 53854 34802
rect 75618 34750 75630 34802
rect 75682 34750 75694 34802
rect 46398 34738 46450 34750
rect 73502 34738 73554 34750
rect 78206 34738 78258 34750
rect 2046 34690 2098 34702
rect 2046 34626 2098 34638
rect 44382 34690 44434 34702
rect 44382 34626 44434 34638
rect 46062 34690 46114 34702
rect 71822 34690 71874 34702
rect 54002 34638 54014 34690
rect 54066 34638 54078 34690
rect 46062 34626 46114 34638
rect 71822 34626 71874 34638
rect 72158 34690 72210 34702
rect 72158 34626 72210 34638
rect 73054 34690 73106 34702
rect 73054 34626 73106 34638
rect 74174 34690 74226 34702
rect 74610 34638 74622 34690
rect 74674 34638 74686 34690
rect 74174 34626 74226 34638
rect 1344 34522 78624 34556
rect 1344 34470 19838 34522
rect 19890 34470 19942 34522
rect 19994 34470 20046 34522
rect 20098 34470 50558 34522
rect 50610 34470 50662 34522
rect 50714 34470 50766 34522
rect 50818 34470 78624 34522
rect 1344 34436 78624 34470
rect 78206 34354 78258 34366
rect 78206 34290 78258 34302
rect 46286 34242 46338 34254
rect 2034 34190 2046 34242
rect 2098 34190 2110 34242
rect 46286 34178 46338 34190
rect 71150 34242 71202 34254
rect 71150 34178 71202 34190
rect 71486 34242 71538 34254
rect 71486 34178 71538 34190
rect 72606 34242 72658 34254
rect 72606 34178 72658 34190
rect 73166 34242 73218 34254
rect 73166 34178 73218 34190
rect 73502 34242 73554 34254
rect 73502 34178 73554 34190
rect 74622 34242 74674 34254
rect 74622 34178 74674 34190
rect 75294 34242 75346 34254
rect 75294 34178 75346 34190
rect 75966 34242 76018 34254
rect 75966 34178 76018 34190
rect 77534 34242 77586 34254
rect 77534 34178 77586 34190
rect 1710 34130 1762 34142
rect 1710 34066 1762 34078
rect 45838 34130 45890 34142
rect 45838 34066 45890 34078
rect 46510 34130 46562 34142
rect 46510 34066 46562 34078
rect 71710 34130 71762 34142
rect 71710 34066 71762 34078
rect 72158 34130 72210 34142
rect 72158 34066 72210 34078
rect 72718 34130 72770 34142
rect 72718 34066 72770 34078
rect 73726 34130 73778 34142
rect 73726 34066 73778 34078
rect 74286 34130 74338 34142
rect 76302 34130 76354 34142
rect 75058 34078 75070 34130
rect 75122 34078 75134 34130
rect 75730 34078 75742 34130
rect 75794 34078 75806 34130
rect 74286 34066 74338 34078
rect 76302 34066 76354 34078
rect 76526 34130 76578 34142
rect 76526 34066 76578 34078
rect 76862 34130 76914 34142
rect 76862 34066 76914 34078
rect 77086 34130 77138 34142
rect 77086 34066 77138 34078
rect 77646 34130 77698 34142
rect 77646 34066 77698 34078
rect 2494 34018 2546 34030
rect 2494 33954 2546 33966
rect 46062 34018 46114 34030
rect 46062 33954 46114 33966
rect 70926 34018 70978 34030
rect 70926 33954 70978 33966
rect 71262 34018 71314 34030
rect 71262 33954 71314 33966
rect 72382 34018 72434 34030
rect 72382 33954 72434 33966
rect 73278 34018 73330 34030
rect 73278 33954 73330 33966
rect 76414 34018 76466 34030
rect 76414 33954 76466 33966
rect 77310 34018 77362 34030
rect 77310 33954 77362 33966
rect 1344 33738 78624 33772
rect 1344 33686 4478 33738
rect 4530 33686 4582 33738
rect 4634 33686 4686 33738
rect 4738 33686 35198 33738
rect 35250 33686 35302 33738
rect 35354 33686 35406 33738
rect 35458 33686 65918 33738
rect 65970 33686 66022 33738
rect 66074 33686 66126 33738
rect 66178 33686 78624 33738
rect 1344 33652 78624 33686
rect 45278 33570 45330 33582
rect 73950 33570 74002 33582
rect 71474 33518 71486 33570
rect 71538 33567 71550 33570
rect 72034 33567 72046 33570
rect 71538 33521 72046 33567
rect 71538 33518 71550 33521
rect 72034 33518 72046 33521
rect 72098 33518 72110 33570
rect 45278 33506 45330 33518
rect 73950 33506 74002 33518
rect 54126 33458 54178 33470
rect 53106 33406 53118 33458
rect 53170 33406 53182 33458
rect 54126 33394 54178 33406
rect 71150 33458 71202 33470
rect 71150 33394 71202 33406
rect 72046 33458 72098 33470
rect 72046 33394 72098 33406
rect 73838 33458 73890 33470
rect 78318 33458 78370 33470
rect 74386 33406 74398 33458
rect 74450 33406 74462 33458
rect 74834 33406 74846 33458
rect 74898 33406 74910 33458
rect 73838 33394 73890 33406
rect 78318 33394 78370 33406
rect 76862 33346 76914 33358
rect 46834 33294 46846 33346
rect 46898 33294 46910 33346
rect 52994 33294 53006 33346
rect 53058 33294 53070 33346
rect 72706 33294 72718 33346
rect 72770 33294 72782 33346
rect 74498 33294 74510 33346
rect 74562 33294 74574 33346
rect 75282 33294 75294 33346
rect 75346 33294 75358 33346
rect 76862 33282 76914 33294
rect 77086 33346 77138 33358
rect 77086 33282 77138 33294
rect 77758 33346 77810 33358
rect 77758 33282 77810 33294
rect 45166 33234 45218 33246
rect 45166 33170 45218 33182
rect 45726 33234 45778 33246
rect 47070 33234 47122 33246
rect 76526 33234 76578 33246
rect 46386 33182 46398 33234
rect 46450 33182 46462 33234
rect 53330 33182 53342 33234
rect 53394 33182 53406 33234
rect 77410 33182 77422 33234
rect 77474 33182 77486 33234
rect 45726 33170 45778 33182
rect 47070 33170 47122 33182
rect 76526 33170 76578 33182
rect 1710 33122 1762 33134
rect 2494 33122 2546 33134
rect 2034 33070 2046 33122
rect 2098 33070 2110 33122
rect 1710 33058 1762 33070
rect 2494 33058 2546 33070
rect 46062 33122 46114 33134
rect 46062 33058 46114 33070
rect 71598 33122 71650 33134
rect 71598 33058 71650 33070
rect 72942 33122 72994 33134
rect 72942 33058 72994 33070
rect 73726 33122 73778 33134
rect 73726 33058 73778 33070
rect 76638 33122 76690 33134
rect 76638 33058 76690 33070
rect 1344 32954 78624 32988
rect 1344 32902 19838 32954
rect 19890 32902 19942 32954
rect 19994 32902 20046 32954
rect 20098 32902 50558 32954
rect 50610 32902 50662 32954
rect 50714 32902 50766 32954
rect 50818 32902 78624 32954
rect 1344 32868 78624 32902
rect 70926 32786 70978 32798
rect 70926 32722 70978 32734
rect 74174 32786 74226 32798
rect 74174 32722 74226 32734
rect 77758 32786 77810 32798
rect 77758 32722 77810 32734
rect 45502 32674 45554 32686
rect 45502 32610 45554 32622
rect 45838 32674 45890 32686
rect 45838 32610 45890 32622
rect 46174 32674 46226 32686
rect 46174 32610 46226 32622
rect 71710 32674 71762 32686
rect 71710 32610 71762 32622
rect 72382 32674 72434 32686
rect 72382 32610 72434 32622
rect 72718 32674 72770 32686
rect 77534 32674 77586 32686
rect 76738 32622 76750 32674
rect 76802 32622 76814 32674
rect 72718 32610 72770 32622
rect 77534 32610 77586 32622
rect 71038 32562 71090 32574
rect 71038 32498 71090 32510
rect 71374 32562 71426 32574
rect 71374 32498 71426 32510
rect 73726 32562 73778 32574
rect 73726 32498 73778 32510
rect 74398 32562 74450 32574
rect 76414 32562 76466 32574
rect 74946 32510 74958 32562
rect 75010 32510 75022 32562
rect 75506 32510 75518 32562
rect 75570 32510 75582 32562
rect 74398 32498 74450 32510
rect 76414 32498 76466 32510
rect 77310 32562 77362 32574
rect 77310 32498 77362 32510
rect 71262 32450 71314 32462
rect 71262 32386 71314 32398
rect 73502 32450 73554 32462
rect 73502 32386 73554 32398
rect 74286 32450 74338 32462
rect 75394 32398 75406 32450
rect 75458 32398 75470 32450
rect 77858 32398 77870 32450
rect 77922 32398 77934 32450
rect 74286 32386 74338 32398
rect 74846 32338 74898 32350
rect 74846 32274 74898 32286
rect 1344 32170 78624 32204
rect 1344 32118 4478 32170
rect 4530 32118 4582 32170
rect 4634 32118 4686 32170
rect 4738 32118 35198 32170
rect 35250 32118 35302 32170
rect 35354 32118 35406 32170
rect 35458 32118 65918 32170
rect 65970 32118 66022 32170
rect 66074 32118 66126 32170
rect 66178 32118 78624 32170
rect 1344 32084 78624 32118
rect 77534 32002 77586 32014
rect 77534 31938 77586 31950
rect 52782 31890 52834 31902
rect 52782 31826 52834 31838
rect 75294 31890 75346 31902
rect 75294 31826 75346 31838
rect 75742 31890 75794 31902
rect 75742 31826 75794 31838
rect 77646 31890 77698 31902
rect 77646 31826 77698 31838
rect 44942 31778 44994 31790
rect 44942 31714 44994 31726
rect 45950 31778 46002 31790
rect 45950 31714 46002 31726
rect 46174 31778 46226 31790
rect 70926 31778 70978 31790
rect 51090 31726 51102 31778
rect 51154 31726 51166 31778
rect 46174 31714 46226 31726
rect 70926 31714 70978 31726
rect 71710 31778 71762 31790
rect 71710 31714 71762 31726
rect 72270 31778 72322 31790
rect 72270 31714 72322 31726
rect 72606 31778 72658 31790
rect 72606 31714 72658 31726
rect 73054 31778 73106 31790
rect 73054 31714 73106 31726
rect 73726 31778 73778 31790
rect 73726 31714 73778 31726
rect 74062 31778 74114 31790
rect 74062 31714 74114 31726
rect 76526 31778 76578 31790
rect 76526 31714 76578 31726
rect 76862 31778 76914 31790
rect 77858 31726 77870 31778
rect 77922 31726 77934 31778
rect 76862 31714 76914 31726
rect 1710 31666 1762 31678
rect 1710 31602 1762 31614
rect 45054 31666 45106 31678
rect 45054 31602 45106 31614
rect 46398 31666 46450 31678
rect 46398 31602 46450 31614
rect 46622 31666 46674 31678
rect 71262 31666 71314 31678
rect 51426 31614 51438 31666
rect 51490 31614 51502 31666
rect 46622 31602 46674 31614
rect 71262 31602 71314 31614
rect 71486 31666 71538 31678
rect 71486 31602 71538 31614
rect 72158 31666 72210 31678
rect 72158 31602 72210 31614
rect 73278 31666 73330 31678
rect 73278 31602 73330 31614
rect 74622 31666 74674 31678
rect 74622 31602 74674 31614
rect 77086 31666 77138 31678
rect 77086 31602 77138 31614
rect 2046 31554 2098 31566
rect 2046 31490 2098 31502
rect 2494 31554 2546 31566
rect 2494 31490 2546 31502
rect 45502 31554 45554 31566
rect 71150 31554 71202 31566
rect 51650 31502 51662 31554
rect 51714 31502 51726 31554
rect 45502 31490 45554 31502
rect 71150 31490 71202 31502
rect 72046 31554 72098 31566
rect 72046 31490 72098 31502
rect 72830 31554 72882 31566
rect 72830 31490 72882 31502
rect 74510 31554 74562 31566
rect 74510 31490 74562 31502
rect 74734 31554 74786 31566
rect 74734 31490 74786 31502
rect 76638 31554 76690 31566
rect 76638 31490 76690 31502
rect 1344 31386 78624 31420
rect 1344 31334 19838 31386
rect 19890 31334 19942 31386
rect 19994 31334 20046 31386
rect 20098 31334 50558 31386
rect 50610 31334 50662 31386
rect 50714 31334 50766 31386
rect 50818 31334 78624 31386
rect 1344 31300 78624 31334
rect 44270 31218 44322 31230
rect 44270 31154 44322 31166
rect 52334 31218 52386 31230
rect 52334 31154 52386 31166
rect 52782 31218 52834 31230
rect 52782 31154 52834 31166
rect 71822 31218 71874 31230
rect 71822 31154 71874 31166
rect 72718 31218 72770 31230
rect 72718 31154 72770 31166
rect 73502 31218 73554 31230
rect 73502 31154 73554 31166
rect 75854 31218 75906 31230
rect 75854 31154 75906 31166
rect 44606 31106 44658 31118
rect 46398 31106 46450 31118
rect 2034 31054 2046 31106
rect 2098 31054 2110 31106
rect 45714 31054 45726 31106
rect 45778 31054 45790 31106
rect 44606 31042 44658 31054
rect 46398 31042 46450 31054
rect 46622 31106 46674 31118
rect 46622 31042 46674 31054
rect 47294 31106 47346 31118
rect 70926 31106 70978 31118
rect 50306 31054 50318 31106
rect 50370 31054 50382 31106
rect 51426 31054 51438 31106
rect 51490 31054 51502 31106
rect 47294 31042 47346 31054
rect 70926 31042 70978 31054
rect 74510 31106 74562 31118
rect 74510 31042 74562 31054
rect 75182 31106 75234 31118
rect 75182 31042 75234 31054
rect 75518 31106 75570 31118
rect 75518 31042 75570 31054
rect 76190 31106 76242 31118
rect 76190 31042 76242 31054
rect 77422 31106 77474 31118
rect 77422 31042 77474 31054
rect 1710 30994 1762 31006
rect 1710 30930 1762 30942
rect 44718 30994 44770 31006
rect 45950 30994 46002 31006
rect 45490 30942 45502 30994
rect 45554 30942 45566 30994
rect 44718 30930 44770 30942
rect 45950 30930 46002 30942
rect 46174 30994 46226 31006
rect 46174 30930 46226 30942
rect 46958 30994 47010 31006
rect 46958 30930 47010 30942
rect 47406 30994 47458 31006
rect 73838 30994 73890 31006
rect 50530 30942 50542 30994
rect 50594 30942 50606 30994
rect 51090 30942 51102 30994
rect 51154 30942 51166 30994
rect 47406 30930 47458 30942
rect 73838 30930 73890 30942
rect 74174 30994 74226 31006
rect 74174 30930 74226 30942
rect 74846 30994 74898 31006
rect 74846 30930 74898 30942
rect 76526 30994 76578 31006
rect 76526 30930 76578 30942
rect 76638 30994 76690 31006
rect 76638 30930 76690 30942
rect 76974 30994 77026 31006
rect 76974 30930 77026 30942
rect 77646 30994 77698 31006
rect 77646 30930 77698 30942
rect 2494 30882 2546 30894
rect 2494 30818 2546 30830
rect 47070 30882 47122 30894
rect 71374 30882 71426 30894
rect 50754 30830 50766 30882
rect 50818 30830 50830 30882
rect 47070 30818 47122 30830
rect 71374 30818 71426 30830
rect 76302 30882 76354 30894
rect 76302 30818 76354 30830
rect 77198 30882 77250 30894
rect 77198 30818 77250 30830
rect 78206 30882 78258 30894
rect 78206 30818 78258 30830
rect 51214 30770 51266 30782
rect 71250 30718 71262 30770
rect 71314 30767 71326 30770
rect 71810 30767 71822 30770
rect 71314 30721 71822 30767
rect 71314 30718 71326 30721
rect 71810 30718 71822 30721
rect 71874 30718 71886 30770
rect 51214 30706 51266 30718
rect 1344 30602 78624 30636
rect 1344 30550 4478 30602
rect 4530 30550 4582 30602
rect 4634 30550 4686 30602
rect 4738 30550 35198 30602
rect 35250 30550 35302 30602
rect 35354 30550 35406 30602
rect 35458 30550 65918 30602
rect 65970 30550 66022 30602
rect 66074 30550 66126 30602
rect 66178 30550 78624 30602
rect 1344 30516 78624 30550
rect 77534 30434 77586 30446
rect 45490 30382 45502 30434
rect 45554 30431 45566 30434
rect 45826 30431 45838 30434
rect 45554 30385 45838 30431
rect 45554 30382 45566 30385
rect 45826 30382 45838 30385
rect 45890 30382 45902 30434
rect 77534 30370 77586 30382
rect 77646 30322 77698 30334
rect 74050 30270 74062 30322
rect 74114 30270 74126 30322
rect 77646 30258 77698 30270
rect 44942 30210 44994 30222
rect 44942 30146 44994 30158
rect 46174 30210 46226 30222
rect 46174 30146 46226 30158
rect 46398 30210 46450 30222
rect 46398 30146 46450 30158
rect 46622 30210 46674 30222
rect 51774 30210 51826 30222
rect 73278 30210 73330 30222
rect 76638 30210 76690 30222
rect 47058 30158 47070 30210
rect 47122 30158 47134 30210
rect 50642 30158 50654 30210
rect 50706 30158 50718 30210
rect 71810 30158 71822 30210
rect 71874 30158 71886 30210
rect 73938 30158 73950 30210
rect 74002 30158 74014 30210
rect 74946 30158 74958 30210
rect 75010 30158 75022 30210
rect 75170 30158 75182 30210
rect 75234 30158 75246 30210
rect 46622 30146 46674 30158
rect 51774 30146 51826 30158
rect 73278 30146 73330 30158
rect 76638 30146 76690 30158
rect 76750 30210 76802 30222
rect 77858 30158 77870 30210
rect 77922 30158 77934 30210
rect 76750 30146 76802 30158
rect 44830 30098 44882 30110
rect 44830 30034 44882 30046
rect 46062 30098 46114 30110
rect 46062 30034 46114 30046
rect 47294 30098 47346 30110
rect 72494 30098 72546 30110
rect 50754 30046 50766 30098
rect 50818 30046 50830 30098
rect 51314 30046 51326 30098
rect 51378 30046 51390 30098
rect 71586 30046 71598 30098
rect 71650 30046 71662 30098
rect 47294 30034 47346 30046
rect 72494 30034 72546 30046
rect 72718 30098 72770 30110
rect 72718 30034 72770 30046
rect 73054 30098 73106 30110
rect 73054 30034 73106 30046
rect 76302 30098 76354 30110
rect 76302 30034 76354 30046
rect 45390 29986 45442 29998
rect 45390 29922 45442 29934
rect 72830 29986 72882 29998
rect 72830 29922 72882 29934
rect 76414 29986 76466 29998
rect 76414 29922 76466 29934
rect 1344 29818 78624 29852
rect 1344 29766 19838 29818
rect 19890 29766 19942 29818
rect 19994 29766 20046 29818
rect 20098 29766 50558 29818
rect 50610 29766 50662 29818
rect 50714 29766 50766 29818
rect 50818 29766 78624 29818
rect 1344 29732 78624 29766
rect 45166 29650 45218 29662
rect 45166 29586 45218 29598
rect 72382 29650 72434 29662
rect 72382 29586 72434 29598
rect 72606 29650 72658 29662
rect 72606 29586 72658 29598
rect 73278 29650 73330 29662
rect 73278 29586 73330 29598
rect 73502 29650 73554 29662
rect 73502 29586 73554 29598
rect 77870 29650 77922 29662
rect 77870 29586 77922 29598
rect 2046 29538 2098 29550
rect 2046 29474 2098 29486
rect 44830 29538 44882 29550
rect 44830 29474 44882 29486
rect 45054 29538 45106 29550
rect 45054 29474 45106 29486
rect 71710 29538 71762 29550
rect 71710 29474 71762 29486
rect 74398 29538 74450 29550
rect 74398 29474 74450 29486
rect 74958 29538 75010 29550
rect 74958 29474 75010 29486
rect 75518 29538 75570 29550
rect 75518 29474 75570 29486
rect 76078 29538 76130 29550
rect 76078 29474 76130 29486
rect 78206 29538 78258 29550
rect 78206 29474 78258 29486
rect 1710 29426 1762 29438
rect 1710 29362 1762 29374
rect 71038 29426 71090 29438
rect 71038 29362 71090 29374
rect 71374 29426 71426 29438
rect 71374 29362 71426 29374
rect 72830 29426 72882 29438
rect 72830 29362 72882 29374
rect 73726 29426 73778 29438
rect 73726 29362 73778 29374
rect 74622 29426 74674 29438
rect 74622 29362 74674 29374
rect 76414 29426 76466 29438
rect 76414 29362 76466 29374
rect 76638 29426 76690 29438
rect 77522 29374 77534 29426
rect 77586 29374 77598 29426
rect 76638 29362 76690 29374
rect 2494 29314 2546 29326
rect 2494 29250 2546 29262
rect 72718 29314 72770 29326
rect 72718 29250 72770 29262
rect 73614 29314 73666 29326
rect 76190 29314 76242 29326
rect 75394 29262 75406 29314
rect 75458 29262 75470 29314
rect 77410 29262 77422 29314
rect 77474 29262 77486 29314
rect 73614 29250 73666 29262
rect 76190 29250 76242 29262
rect 75742 29202 75794 29214
rect 75742 29138 75794 29150
rect 77198 29202 77250 29214
rect 77198 29138 77250 29150
rect 1344 29034 78624 29068
rect 1344 28982 4478 29034
rect 4530 28982 4582 29034
rect 4634 28982 4686 29034
rect 4738 28982 35198 29034
rect 35250 28982 35302 29034
rect 35354 28982 35406 29034
rect 35458 28982 65918 29034
rect 65970 28982 66022 29034
rect 66074 28982 66126 29034
rect 66178 28982 78624 29034
rect 1344 28948 78624 28982
rect 77198 28866 77250 28878
rect 77198 28802 77250 28814
rect 37550 28754 37602 28766
rect 37550 28690 37602 28702
rect 40910 28754 40962 28766
rect 40910 28690 40962 28702
rect 71262 28754 71314 28766
rect 71262 28690 71314 28702
rect 71710 28754 71762 28766
rect 71710 28690 71762 28702
rect 72158 28754 72210 28766
rect 72158 28690 72210 28702
rect 73390 28754 73442 28766
rect 73390 28690 73442 28702
rect 73726 28754 73778 28766
rect 73726 28690 73778 28702
rect 77310 28754 77362 28766
rect 77310 28690 77362 28702
rect 1710 28642 1762 28654
rect 1710 28578 1762 28590
rect 2494 28642 2546 28654
rect 72382 28642 72434 28654
rect 75406 28642 75458 28654
rect 37874 28590 37886 28642
rect 37938 28590 37950 28642
rect 38322 28590 38334 28642
rect 38386 28590 38398 28642
rect 74274 28590 74286 28642
rect 74338 28590 74350 28642
rect 2494 28578 2546 28590
rect 72382 28578 72434 28590
rect 75406 28578 75458 28590
rect 75630 28642 75682 28654
rect 75630 28578 75682 28590
rect 76526 28642 76578 28654
rect 76526 28578 76578 28590
rect 76638 28642 76690 28654
rect 78206 28642 78258 28654
rect 77522 28590 77534 28642
rect 77586 28590 77598 28642
rect 76638 28578 76690 28590
rect 78206 28578 78258 28590
rect 72718 28530 72770 28542
rect 2034 28478 2046 28530
rect 2098 28478 2110 28530
rect 38770 28478 38782 28530
rect 38834 28478 38846 28530
rect 72718 28466 72770 28478
rect 75070 28530 75122 28542
rect 75070 28466 75122 28478
rect 75182 28530 75234 28542
rect 75182 28466 75234 28478
rect 76190 28530 76242 28542
rect 76190 28466 76242 28478
rect 77870 28530 77922 28542
rect 77870 28466 77922 28478
rect 76302 28418 76354 28430
rect 37986 28366 37998 28418
rect 38050 28366 38062 28418
rect 74498 28366 74510 28418
rect 74562 28366 74574 28418
rect 76302 28354 76354 28366
rect 1344 28250 78624 28284
rect 1344 28198 19838 28250
rect 19890 28198 19942 28250
rect 19994 28198 20046 28250
rect 20098 28198 50558 28250
rect 50610 28198 50662 28250
rect 50714 28198 50766 28250
rect 50818 28198 78624 28250
rect 1344 28164 78624 28198
rect 34750 28082 34802 28094
rect 34750 28018 34802 28030
rect 37102 28082 37154 28094
rect 37102 28018 37154 28030
rect 37662 28082 37714 28094
rect 37662 28018 37714 28030
rect 39902 28082 39954 28094
rect 39902 28018 39954 28030
rect 40350 28082 40402 28094
rect 40350 28018 40402 28030
rect 42478 28082 42530 28094
rect 42478 28018 42530 28030
rect 44606 28082 44658 28094
rect 44606 28018 44658 28030
rect 70702 28082 70754 28094
rect 70702 28018 70754 28030
rect 71822 28082 71874 28094
rect 71822 28018 71874 28030
rect 75966 28082 76018 28094
rect 75966 28018 76018 28030
rect 76750 28082 76802 28094
rect 76750 28018 76802 28030
rect 77870 28082 77922 28094
rect 77870 28018 77922 28030
rect 44942 27970 44994 27982
rect 35074 27918 35086 27970
rect 35138 27918 35150 27970
rect 38770 27918 38782 27970
rect 38834 27918 38846 27970
rect 41906 27918 41918 27970
rect 41970 27918 41982 27970
rect 44942 27906 44994 27918
rect 72718 27970 72770 27982
rect 72718 27906 72770 27918
rect 72942 27970 72994 27982
rect 72942 27906 72994 27918
rect 73278 27970 73330 27982
rect 73278 27906 73330 27918
rect 74174 27970 74226 27982
rect 74174 27906 74226 27918
rect 74958 27970 75010 27982
rect 74958 27906 75010 27918
rect 75854 27970 75906 27982
rect 75854 27906 75906 27918
rect 76190 27970 76242 27982
rect 76190 27906 76242 27918
rect 76414 27970 76466 27982
rect 76414 27906 76466 27918
rect 78206 27970 78258 27982
rect 78206 27906 78258 27918
rect 36654 27858 36706 27870
rect 39454 27858 39506 27870
rect 70254 27858 70306 27870
rect 35298 27806 35310 27858
rect 35362 27806 35374 27858
rect 36194 27806 36206 27858
rect 36258 27806 36270 27858
rect 37874 27806 37886 27858
rect 37938 27806 37950 27858
rect 38994 27806 39006 27858
rect 39058 27806 39070 27858
rect 41010 27806 41022 27858
rect 41074 27806 41086 27858
rect 41458 27806 41470 27858
rect 41522 27806 41534 27858
rect 36654 27794 36706 27806
rect 39454 27794 39506 27806
rect 70254 27794 70306 27806
rect 70926 27858 70978 27870
rect 70926 27794 70978 27806
rect 73502 27858 73554 27870
rect 73502 27794 73554 27806
rect 73726 27858 73778 27870
rect 73726 27794 73778 27806
rect 74286 27858 74338 27870
rect 74286 27794 74338 27806
rect 74734 27858 74786 27870
rect 74734 27794 74786 27806
rect 75294 27858 75346 27870
rect 75294 27794 75346 27806
rect 77086 27858 77138 27870
rect 77086 27794 77138 27806
rect 77646 27858 77698 27870
rect 77646 27794 77698 27806
rect 70814 27746 70866 27758
rect 35522 27694 35534 27746
rect 35586 27694 35598 27746
rect 38546 27694 38558 27746
rect 38610 27694 38622 27746
rect 41346 27694 41358 27746
rect 41410 27694 41422 27746
rect 70814 27682 70866 27694
rect 73054 27746 73106 27758
rect 73054 27682 73106 27694
rect 73950 27746 74002 27758
rect 73950 27682 74002 27694
rect 75182 27746 75234 27758
rect 75182 27682 75234 27694
rect 45054 27634 45106 27646
rect 45054 27570 45106 27582
rect 1344 27466 78624 27500
rect 1344 27414 4478 27466
rect 4530 27414 4582 27466
rect 4634 27414 4686 27466
rect 4738 27414 35198 27466
rect 35250 27414 35302 27466
rect 35354 27414 35406 27466
rect 35458 27414 65918 27466
rect 65970 27414 66022 27466
rect 66074 27414 66126 27466
rect 66178 27414 78624 27466
rect 1344 27380 78624 27414
rect 76190 27298 76242 27310
rect 76190 27234 76242 27246
rect 76862 27298 76914 27310
rect 76862 27234 76914 27246
rect 43822 27186 43874 27198
rect 43822 27122 43874 27134
rect 44830 27186 44882 27198
rect 44830 27122 44882 27134
rect 45390 27186 45442 27198
rect 45390 27122 45442 27134
rect 46398 27186 46450 27198
rect 46398 27122 46450 27134
rect 50318 27186 50370 27198
rect 50318 27122 50370 27134
rect 50766 27186 50818 27198
rect 50766 27122 50818 27134
rect 71934 27186 71986 27198
rect 76974 27186 77026 27198
rect 75394 27134 75406 27186
rect 75458 27134 75470 27186
rect 71934 27122 71986 27134
rect 76974 27122 77026 27134
rect 36990 27074 37042 27086
rect 43038 27074 43090 27086
rect 34066 27022 34078 27074
rect 34130 27022 34142 27074
rect 34738 27022 34750 27074
rect 34802 27022 34814 27074
rect 35746 27022 35758 27074
rect 35810 27022 35822 27074
rect 36194 27022 36206 27074
rect 36258 27022 36270 27074
rect 37426 27022 37438 27074
rect 37490 27022 37502 27074
rect 38098 27022 38110 27074
rect 38162 27022 38174 27074
rect 38658 27022 38670 27074
rect 38722 27022 38734 27074
rect 39778 27022 39790 27074
rect 39842 27022 39854 27074
rect 40674 27022 40686 27074
rect 40738 27022 40750 27074
rect 41010 27022 41022 27074
rect 41074 27022 41086 27074
rect 42130 27022 42142 27074
rect 42194 27022 42206 27074
rect 36990 27010 37042 27022
rect 43038 27010 43090 27022
rect 46174 27074 46226 27086
rect 46174 27010 46226 27022
rect 47070 27074 47122 27086
rect 47070 27010 47122 27022
rect 47294 27074 47346 27086
rect 47294 27010 47346 27022
rect 49086 27074 49138 27086
rect 49086 27010 49138 27022
rect 49646 27074 49698 27086
rect 49646 27010 49698 27022
rect 70590 27074 70642 27086
rect 70590 27010 70642 27022
rect 71038 27074 71090 27086
rect 71038 27010 71090 27022
rect 72382 27074 72434 27086
rect 72382 27010 72434 27022
rect 73390 27074 73442 27086
rect 73390 27010 73442 27022
rect 73502 27074 73554 27086
rect 75282 27022 75294 27074
rect 75346 27022 75358 27074
rect 77186 27022 77198 27074
rect 77250 27022 77262 27074
rect 73502 27010 73554 27022
rect 1710 26962 1762 26974
rect 1710 26898 1762 26910
rect 2046 26962 2098 26974
rect 2046 26898 2098 26910
rect 2494 26962 2546 26974
rect 44942 26962 44994 26974
rect 34962 26910 34974 26962
rect 35026 26910 35038 26962
rect 35634 26910 35646 26962
rect 35698 26910 35710 26962
rect 38770 26910 38782 26962
rect 38834 26910 38846 26962
rect 40562 26910 40574 26962
rect 40626 26910 40638 26962
rect 41682 26910 41694 26962
rect 41746 26910 41758 26962
rect 2494 26898 2546 26910
rect 44942 26898 44994 26910
rect 46622 26962 46674 26974
rect 46622 26898 46674 26910
rect 46846 26962 46898 26974
rect 46846 26898 46898 26910
rect 47518 26962 47570 26974
rect 47518 26898 47570 26910
rect 47742 26962 47794 26974
rect 47742 26898 47794 26910
rect 49758 26962 49810 26974
rect 49758 26898 49810 26910
rect 73054 26962 73106 26974
rect 73054 26898 73106 26910
rect 74286 26962 74338 26974
rect 74286 26898 74338 26910
rect 74622 26962 74674 26974
rect 74622 26898 74674 26910
rect 75630 26962 75682 26974
rect 75630 26898 75682 26910
rect 76526 26962 76578 26974
rect 76526 26898 76578 26910
rect 77534 26962 77586 26974
rect 77534 26898 77586 26910
rect 77870 26962 77922 26974
rect 77870 26898 77922 26910
rect 42478 26850 42530 26862
rect 33954 26798 33966 26850
rect 34018 26798 34030 26850
rect 36194 26798 36206 26850
rect 36258 26798 36270 26850
rect 38322 26798 38334 26850
rect 38386 26798 38398 26850
rect 39778 26798 39790 26850
rect 39842 26798 39854 26850
rect 41122 26798 41134 26850
rect 41186 26798 41198 26850
rect 42478 26786 42530 26798
rect 44382 26850 44434 26862
rect 44382 26786 44434 26798
rect 49198 26850 49250 26862
rect 49198 26786 49250 26798
rect 49422 26850 49474 26862
rect 49422 26786 49474 26798
rect 49982 26850 50034 26862
rect 49982 26786 50034 26798
rect 71150 26850 71202 26862
rect 71150 26786 71202 26798
rect 71262 26850 71314 26862
rect 71262 26786 71314 26798
rect 72830 26850 72882 26862
rect 72830 26786 72882 26798
rect 73166 26850 73218 26862
rect 73166 26786 73218 26798
rect 76302 26850 76354 26862
rect 76302 26786 76354 26798
rect 1344 26682 78624 26716
rect 1344 26630 19838 26682
rect 19890 26630 19942 26682
rect 19994 26630 20046 26682
rect 20098 26630 50558 26682
rect 50610 26630 50662 26682
rect 50714 26630 50766 26682
rect 50818 26630 78624 26682
rect 1344 26596 78624 26630
rect 35198 26514 35250 26526
rect 35198 26450 35250 26462
rect 42590 26514 42642 26526
rect 44606 26514 44658 26526
rect 44034 26462 44046 26514
rect 44098 26462 44110 26514
rect 42590 26450 42642 26462
rect 44606 26450 44658 26462
rect 47518 26514 47570 26526
rect 47518 26450 47570 26462
rect 50094 26514 50146 26526
rect 50094 26450 50146 26462
rect 50542 26514 50594 26526
rect 50542 26450 50594 26462
rect 70926 26514 70978 26526
rect 70926 26450 70978 26462
rect 76974 26514 77026 26526
rect 76974 26450 77026 26462
rect 77198 26514 77250 26526
rect 77198 26450 77250 26462
rect 77870 26514 77922 26526
rect 77870 26450 77922 26462
rect 2046 26402 2098 26414
rect 44942 26402 44994 26414
rect 46734 26402 46786 26414
rect 35858 26350 35870 26402
rect 35922 26350 35934 26402
rect 38770 26350 38782 26402
rect 38834 26350 38846 26402
rect 41682 26350 41694 26402
rect 41746 26350 41758 26402
rect 43026 26350 43038 26402
rect 43090 26350 43102 26402
rect 46050 26350 46062 26402
rect 46114 26350 46126 26402
rect 2046 26338 2098 26350
rect 44942 26338 44994 26350
rect 46734 26338 46786 26350
rect 47630 26402 47682 26414
rect 47630 26338 47682 26350
rect 48862 26402 48914 26414
rect 48862 26338 48914 26350
rect 49310 26402 49362 26414
rect 49310 26338 49362 26350
rect 49422 26402 49474 26414
rect 76302 26402 76354 26414
rect 75618 26350 75630 26402
rect 75682 26350 75694 26402
rect 49422 26338 49474 26350
rect 76302 26338 76354 26350
rect 77534 26402 77586 26414
rect 77534 26338 77586 26350
rect 1710 26290 1762 26302
rect 37774 26290 37826 26302
rect 40350 26290 40402 26302
rect 45054 26290 45106 26302
rect 46286 26290 46338 26302
rect 35970 26238 35982 26290
rect 36034 26238 36046 26290
rect 36306 26238 36318 26290
rect 36370 26238 36382 26290
rect 37314 26238 37326 26290
rect 37378 26238 37390 26290
rect 38098 26238 38110 26290
rect 38162 26238 38174 26290
rect 39218 26238 39230 26290
rect 39282 26238 39294 26290
rect 41010 26238 41022 26290
rect 41074 26238 41086 26290
rect 41794 26238 41806 26290
rect 41858 26238 41870 26290
rect 43586 26238 43598 26290
rect 43650 26238 43662 26290
rect 44146 26238 44158 26290
rect 44210 26238 44222 26290
rect 45826 26238 45838 26290
rect 45890 26238 45902 26290
rect 1710 26226 1762 26238
rect 37774 26226 37826 26238
rect 40350 26226 40402 26238
rect 45054 26226 45106 26238
rect 46286 26226 46338 26238
rect 46510 26290 46562 26302
rect 46510 26226 46562 26238
rect 46846 26290 46898 26302
rect 46846 26226 46898 26238
rect 47182 26290 47234 26302
rect 47182 26226 47234 26238
rect 47742 26290 47794 26302
rect 47742 26226 47794 26238
rect 48750 26290 48802 26302
rect 48750 26226 48802 26238
rect 71150 26290 71202 26302
rect 71150 26226 71202 26238
rect 71374 26290 71426 26302
rect 71374 26226 71426 26238
rect 72382 26290 72434 26302
rect 75966 26290 76018 26302
rect 73490 26238 73502 26290
rect 73554 26238 73566 26290
rect 74274 26238 74286 26290
rect 74338 26238 74350 26290
rect 74834 26238 74846 26290
rect 74898 26238 74910 26290
rect 75394 26238 75406 26290
rect 75458 26238 75470 26290
rect 72382 26226 72434 26238
rect 75966 26226 76018 26238
rect 78206 26290 78258 26302
rect 78206 26226 78258 26238
rect 2494 26178 2546 26190
rect 71262 26178 71314 26190
rect 35746 26126 35758 26178
rect 35810 26126 35822 26178
rect 38546 26126 38558 26178
rect 38610 26126 38622 26178
rect 39890 26126 39902 26178
rect 39954 26126 39966 26178
rect 41458 26126 41470 26178
rect 41522 26126 41534 26178
rect 70802 26175 70814 26178
rect 70593 26129 70814 26175
rect 2494 26114 2546 26126
rect 48862 26066 48914 26078
rect 48862 26002 48914 26014
rect 49422 26066 49474 26078
rect 70593 26066 70639 26129
rect 70802 26126 70814 26129
rect 70866 26126 70878 26178
rect 71262 26114 71314 26126
rect 72942 26178 72994 26190
rect 72942 26114 72994 26126
rect 73278 26178 73330 26190
rect 73278 26114 73330 26126
rect 74062 26066 74114 26078
rect 70578 26014 70590 26066
rect 70642 26014 70654 26066
rect 49422 26002 49474 26014
rect 74062 26002 74114 26014
rect 1344 25898 78624 25932
rect 1344 25846 4478 25898
rect 4530 25846 4582 25898
rect 4634 25846 4686 25898
rect 4738 25846 35198 25898
rect 35250 25846 35302 25898
rect 35354 25846 35406 25898
rect 35458 25846 65918 25898
rect 65970 25846 66022 25898
rect 66074 25846 66126 25898
rect 66178 25846 78624 25898
rect 1344 25812 78624 25846
rect 47070 25730 47122 25742
rect 47070 25666 47122 25678
rect 72718 25730 72770 25742
rect 72718 25666 72770 25678
rect 74398 25730 74450 25742
rect 74398 25666 74450 25678
rect 77758 25730 77810 25742
rect 77758 25666 77810 25678
rect 78094 25730 78146 25742
rect 78094 25666 78146 25678
rect 35870 25618 35922 25630
rect 35870 25554 35922 25566
rect 37774 25618 37826 25630
rect 37774 25554 37826 25566
rect 44046 25618 44098 25630
rect 44046 25554 44098 25566
rect 46958 25618 47010 25630
rect 46958 25554 47010 25566
rect 47518 25618 47570 25630
rect 47518 25554 47570 25566
rect 47966 25618 48018 25630
rect 47966 25554 48018 25566
rect 63310 25618 63362 25630
rect 71026 25566 71038 25618
rect 71090 25566 71102 25618
rect 63310 25554 63362 25566
rect 38110 25506 38162 25518
rect 63198 25506 63250 25518
rect 76750 25506 76802 25518
rect 37314 25454 37326 25506
rect 37378 25454 37390 25506
rect 38322 25454 38334 25506
rect 38386 25454 38398 25506
rect 40338 25454 40350 25506
rect 40402 25454 40414 25506
rect 42466 25454 42478 25506
rect 42530 25454 42542 25506
rect 43362 25454 43374 25506
rect 43426 25454 43438 25506
rect 44818 25454 44830 25506
rect 44882 25454 44894 25506
rect 45714 25454 45726 25506
rect 45778 25454 45790 25506
rect 62850 25454 62862 25506
rect 62914 25454 62926 25506
rect 70802 25454 70814 25506
rect 70866 25454 70878 25506
rect 71810 25454 71822 25506
rect 71874 25454 71886 25506
rect 72146 25454 72158 25506
rect 72210 25454 72222 25506
rect 72482 25454 72494 25506
rect 72546 25454 72558 25506
rect 73266 25454 73278 25506
rect 73330 25454 73342 25506
rect 73826 25454 73838 25506
rect 73890 25454 73902 25506
rect 74162 25454 74174 25506
rect 74226 25454 74238 25506
rect 74946 25454 74958 25506
rect 75010 25454 75022 25506
rect 75506 25454 75518 25506
rect 75570 25454 75582 25506
rect 38110 25442 38162 25454
rect 63198 25442 63250 25454
rect 76750 25442 76802 25454
rect 77422 25506 77474 25518
rect 77422 25442 77474 25454
rect 23998 25394 24050 25406
rect 2034 25342 2046 25394
rect 2098 25342 2110 25394
rect 23998 25330 24050 25342
rect 27134 25394 27186 25406
rect 27134 25330 27186 25342
rect 36430 25394 36482 25406
rect 42142 25394 42194 25406
rect 46286 25394 46338 25406
rect 40450 25342 40462 25394
rect 40514 25342 40526 25394
rect 42578 25342 42590 25394
rect 42642 25342 42654 25394
rect 44930 25342 44942 25394
rect 44994 25342 45006 25394
rect 36430 25330 36482 25342
rect 42142 25330 42194 25342
rect 46286 25330 46338 25342
rect 46622 25394 46674 25406
rect 46622 25330 46674 25342
rect 70702 25394 70754 25406
rect 70702 25330 70754 25342
rect 76414 25394 76466 25406
rect 76414 25330 76466 25342
rect 77086 25394 77138 25406
rect 77086 25330 77138 25342
rect 1710 25282 1762 25294
rect 1710 25218 1762 25230
rect 2494 25282 2546 25294
rect 2494 25218 2546 25230
rect 23662 25282 23714 25294
rect 23662 25218 23714 25230
rect 24110 25282 24162 25294
rect 24110 25218 24162 25230
rect 24334 25282 24386 25294
rect 24334 25218 24386 25230
rect 27022 25282 27074 25294
rect 27022 25218 27074 25230
rect 35534 25282 35586 25294
rect 41806 25282 41858 25294
rect 63422 25282 63474 25294
rect 40002 25230 40014 25282
rect 40066 25230 40078 25282
rect 43474 25230 43486 25282
rect 43538 25230 43550 25282
rect 45826 25230 45838 25282
rect 45890 25230 45902 25282
rect 35534 25218 35586 25230
rect 41806 25218 41858 25230
rect 63422 25218 63474 25230
rect 77982 25282 78034 25294
rect 77982 25218 78034 25230
rect 1344 25114 78624 25148
rect 1344 25062 19838 25114
rect 19890 25062 19942 25114
rect 19994 25062 20046 25114
rect 20098 25062 50558 25114
rect 50610 25062 50662 25114
rect 50714 25062 50766 25114
rect 50818 25062 78624 25114
rect 1344 25028 78624 25062
rect 25342 24946 25394 24958
rect 25342 24882 25394 24894
rect 34974 24946 35026 24958
rect 34974 24882 35026 24894
rect 35310 24946 35362 24958
rect 39454 24946 39506 24958
rect 37426 24894 37438 24946
rect 37490 24894 37502 24946
rect 35310 24882 35362 24894
rect 39454 24882 39506 24894
rect 40350 24946 40402 24958
rect 48190 24946 48242 24958
rect 44370 24894 44382 24946
rect 44434 24894 44446 24946
rect 45938 24894 45950 24946
rect 46002 24894 46014 24946
rect 40350 24882 40402 24894
rect 48190 24882 48242 24894
rect 63198 24946 63250 24958
rect 63198 24882 63250 24894
rect 63982 24946 64034 24958
rect 63982 24882 64034 24894
rect 71710 24946 71762 24958
rect 71710 24882 71762 24894
rect 74174 24946 74226 24958
rect 74174 24882 74226 24894
rect 74958 24946 75010 24958
rect 74958 24882 75010 24894
rect 75406 24946 75458 24958
rect 75406 24882 75458 24894
rect 76190 24946 76242 24958
rect 76190 24882 76242 24894
rect 77646 24946 77698 24958
rect 77646 24882 77698 24894
rect 46958 24834 47010 24846
rect 35746 24782 35758 24834
rect 35810 24782 35822 24834
rect 41682 24782 41694 24834
rect 41746 24782 41758 24834
rect 44930 24782 44942 24834
rect 44994 24782 45006 24834
rect 46610 24782 46622 24834
rect 46674 24782 46686 24834
rect 46958 24770 47010 24782
rect 47294 24834 47346 24846
rect 47294 24770 47346 24782
rect 76078 24834 76130 24846
rect 76078 24770 76130 24782
rect 77086 24834 77138 24846
rect 77086 24770 77138 24782
rect 77534 24834 77586 24846
rect 77534 24770 77586 24782
rect 77758 24834 77810 24846
rect 77758 24770 77810 24782
rect 25566 24722 25618 24734
rect 17490 24670 17502 24722
rect 17554 24670 17566 24722
rect 20626 24670 20638 24722
rect 20690 24670 20702 24722
rect 25566 24658 25618 24670
rect 25790 24722 25842 24734
rect 30382 24722 30434 24734
rect 27234 24670 27246 24722
rect 27298 24670 27310 24722
rect 25790 24658 25842 24670
rect 30382 24658 30434 24670
rect 30494 24722 30546 24734
rect 30494 24658 30546 24670
rect 35086 24722 35138 24734
rect 35086 24658 35138 24670
rect 35422 24722 35474 24734
rect 39342 24722 39394 24734
rect 45614 24722 45666 24734
rect 48862 24722 48914 24734
rect 35970 24670 35982 24722
rect 36034 24670 36046 24722
rect 37538 24670 37550 24722
rect 37602 24670 37614 24722
rect 37874 24670 37886 24722
rect 37938 24670 37950 24722
rect 40114 24670 40126 24722
rect 40178 24670 40190 24722
rect 40898 24670 40910 24722
rect 40962 24670 40974 24722
rect 44146 24670 44158 24722
rect 44210 24670 44222 24722
rect 45266 24670 45278 24722
rect 45330 24670 45342 24722
rect 46386 24670 46398 24722
rect 46450 24670 46462 24722
rect 35422 24658 35474 24670
rect 39342 24658 39394 24670
rect 45614 24658 45666 24670
rect 48862 24658 48914 24670
rect 62750 24722 62802 24734
rect 62750 24658 62802 24670
rect 63422 24722 63474 24734
rect 74622 24722 74674 24734
rect 72146 24670 72158 24722
rect 72210 24670 72222 24722
rect 73042 24670 73054 24722
rect 73106 24670 73118 24722
rect 73490 24670 73502 24722
rect 73554 24670 73566 24722
rect 75618 24670 75630 24722
rect 75682 24670 75694 24722
rect 63422 24658 63474 24670
rect 74622 24658 74674 24670
rect 23886 24610 23938 24622
rect 25678 24610 25730 24622
rect 47854 24610 47906 24622
rect 18162 24558 18174 24610
rect 18226 24558 18238 24610
rect 20290 24558 20302 24610
rect 20354 24558 20366 24610
rect 21410 24558 21422 24610
rect 21474 24558 21486 24610
rect 23538 24558 23550 24610
rect 23602 24558 23614 24610
rect 24210 24558 24222 24610
rect 24274 24558 24286 24610
rect 27906 24558 27918 24610
rect 27970 24558 27982 24610
rect 30034 24558 30046 24610
rect 30098 24558 30110 24610
rect 43810 24558 43822 24610
rect 43874 24558 43886 24610
rect 23886 24546 23938 24558
rect 25678 24546 25730 24558
rect 47854 24546 47906 24558
rect 63310 24610 63362 24622
rect 63310 24546 63362 24558
rect 71374 24610 71426 24622
rect 77186 24558 77198 24610
rect 77250 24558 77262 24610
rect 71374 24546 71426 24558
rect 39454 24498 39506 24510
rect 39454 24434 39506 24446
rect 72382 24498 72434 24510
rect 72382 24434 72434 24446
rect 75294 24498 75346 24510
rect 75294 24434 75346 24446
rect 76302 24498 76354 24510
rect 76302 24434 76354 24446
rect 76862 24498 76914 24510
rect 76862 24434 76914 24446
rect 1344 24330 78624 24364
rect 1344 24278 4478 24330
rect 4530 24278 4582 24330
rect 4634 24278 4686 24330
rect 4738 24278 35198 24330
rect 35250 24278 35302 24330
rect 35354 24278 35406 24330
rect 35458 24278 65918 24330
rect 65970 24278 66022 24330
rect 66074 24278 66126 24330
rect 66178 24278 78624 24330
rect 1344 24244 78624 24278
rect 35982 24162 36034 24174
rect 35982 24098 36034 24110
rect 75294 24162 75346 24174
rect 75294 24098 75346 24110
rect 76190 24162 76242 24174
rect 76190 24098 76242 24110
rect 76526 24162 76578 24174
rect 76526 24098 76578 24110
rect 17166 24050 17218 24062
rect 17166 23986 17218 23998
rect 17614 24050 17666 24062
rect 20078 24050 20130 24062
rect 19730 23998 19742 24050
rect 19794 23998 19806 24050
rect 17614 23986 17666 23998
rect 20078 23986 20130 23998
rect 21758 24050 21810 24062
rect 21758 23986 21810 23998
rect 23326 24050 23378 24062
rect 28030 24050 28082 24062
rect 24994 23998 25006 24050
rect 25058 23998 25070 24050
rect 27122 23998 27134 24050
rect 27186 23998 27198 24050
rect 23326 23986 23378 23998
rect 28030 23986 28082 23998
rect 42366 24050 42418 24062
rect 42366 23986 42418 23998
rect 43262 24050 43314 24062
rect 43262 23986 43314 23998
rect 44158 24050 44210 24062
rect 44158 23986 44210 23998
rect 48302 24050 48354 24062
rect 48302 23986 48354 23998
rect 74286 24050 74338 24062
rect 74286 23986 74338 23998
rect 17726 23938 17778 23950
rect 17726 23874 17778 23886
rect 18174 23938 18226 23950
rect 18174 23874 18226 23886
rect 18286 23938 18338 23950
rect 18286 23874 18338 23886
rect 18622 23938 18674 23950
rect 18622 23874 18674 23886
rect 20750 23938 20802 23950
rect 20750 23874 20802 23886
rect 21198 23938 21250 23950
rect 21198 23874 21250 23886
rect 23662 23938 23714 23950
rect 23662 23874 23714 23886
rect 23998 23938 24050 23950
rect 27470 23938 27522 23950
rect 24322 23886 24334 23938
rect 24386 23886 24398 23938
rect 23998 23874 24050 23886
rect 27470 23874 27522 23886
rect 34750 23938 34802 23950
rect 34750 23874 34802 23886
rect 35870 23938 35922 23950
rect 35870 23874 35922 23886
rect 38222 23938 38274 23950
rect 41806 23938 41858 23950
rect 39442 23886 39454 23938
rect 39506 23886 39518 23938
rect 40338 23886 40350 23938
rect 40402 23886 40414 23938
rect 38222 23874 38274 23886
rect 41806 23874 41858 23886
rect 42702 23938 42754 23950
rect 42702 23874 42754 23886
rect 46062 23938 46114 23950
rect 46062 23874 46114 23886
rect 46510 23938 46562 23950
rect 46510 23874 46562 23886
rect 46734 23938 46786 23950
rect 75406 23938 75458 23950
rect 72258 23886 72270 23938
rect 72322 23886 72334 23938
rect 73266 23886 73278 23938
rect 73330 23886 73342 23938
rect 73602 23886 73614 23938
rect 73666 23886 73678 23938
rect 46734 23874 46786 23886
rect 75406 23874 75458 23886
rect 1710 23826 1762 23838
rect 1710 23762 1762 23774
rect 2046 23826 2098 23838
rect 2046 23762 2098 23774
rect 18510 23826 18562 23838
rect 18510 23762 18562 23774
rect 20414 23826 20466 23838
rect 20414 23762 20466 23774
rect 27918 23826 27970 23838
rect 27918 23762 27970 23774
rect 35646 23826 35698 23838
rect 35646 23762 35698 23774
rect 37102 23826 37154 23838
rect 37102 23762 37154 23774
rect 37214 23826 37266 23838
rect 37214 23762 37266 23774
rect 37662 23826 37714 23838
rect 37662 23762 37714 23774
rect 37774 23826 37826 23838
rect 43598 23826 43650 23838
rect 40450 23774 40462 23826
rect 40514 23774 40526 23826
rect 37774 23762 37826 23774
rect 43598 23762 43650 23774
rect 43710 23826 43762 23838
rect 43710 23762 43762 23774
rect 44830 23826 44882 23838
rect 44830 23762 44882 23774
rect 45390 23826 45442 23838
rect 45390 23762 45442 23774
rect 47070 23826 47122 23838
rect 47070 23762 47122 23774
rect 47182 23826 47234 23838
rect 47182 23762 47234 23774
rect 47630 23826 47682 23838
rect 47630 23762 47682 23774
rect 47742 23826 47794 23838
rect 47742 23762 47794 23774
rect 48750 23826 48802 23838
rect 74622 23826 74674 23838
rect 73714 23774 73726 23826
rect 73778 23774 73790 23826
rect 48750 23762 48802 23774
rect 74622 23762 74674 23774
rect 74958 23826 75010 23838
rect 74958 23762 75010 23774
rect 76862 23826 76914 23838
rect 76862 23762 76914 23774
rect 77198 23826 77250 23838
rect 77198 23762 77250 23774
rect 77870 23826 77922 23838
rect 77870 23762 77922 23774
rect 78206 23826 78258 23838
rect 78206 23762 78258 23774
rect 2494 23714 2546 23726
rect 2494 23650 2546 23662
rect 17502 23714 17554 23726
rect 17502 23650 17554 23662
rect 19406 23714 19458 23726
rect 19406 23650 19458 23662
rect 20526 23714 20578 23726
rect 20526 23650 20578 23662
rect 21646 23714 21698 23726
rect 21646 23650 21698 23662
rect 21870 23714 21922 23726
rect 21870 23650 21922 23662
rect 22318 23714 22370 23726
rect 22318 23650 22370 23662
rect 23774 23714 23826 23726
rect 23774 23650 23826 23662
rect 28142 23714 28194 23726
rect 28142 23650 28194 23662
rect 34302 23714 34354 23726
rect 34302 23650 34354 23662
rect 35086 23714 35138 23726
rect 35086 23650 35138 23662
rect 35982 23714 36034 23726
rect 35982 23650 36034 23662
rect 37438 23714 37490 23726
rect 37438 23650 37490 23662
rect 37998 23714 38050 23726
rect 43934 23714 43986 23726
rect 39330 23662 39342 23714
rect 39394 23662 39406 23714
rect 37998 23650 38050 23662
rect 43934 23650 43986 23662
rect 44270 23714 44322 23726
rect 44270 23650 44322 23662
rect 44942 23714 44994 23726
rect 44942 23650 44994 23662
rect 45166 23714 45218 23726
rect 45166 23650 45218 23662
rect 45502 23714 45554 23726
rect 45502 23650 45554 23662
rect 46398 23714 46450 23726
rect 46398 23650 46450 23662
rect 47406 23714 47458 23726
rect 47406 23650 47458 23662
rect 47966 23714 48018 23726
rect 47966 23650 48018 23662
rect 49310 23714 49362 23726
rect 49310 23650 49362 23662
rect 49646 23714 49698 23726
rect 49646 23650 49698 23662
rect 72158 23714 72210 23726
rect 72158 23650 72210 23662
rect 75518 23714 75570 23726
rect 75518 23650 75570 23662
rect 76414 23714 76466 23726
rect 76414 23650 76466 23662
rect 1344 23546 78624 23580
rect 1344 23494 19838 23546
rect 19890 23494 19942 23546
rect 19994 23494 20046 23546
rect 20098 23494 50558 23546
rect 50610 23494 50662 23546
rect 50714 23494 50766 23546
rect 50818 23494 78624 23546
rect 1344 23460 78624 23494
rect 18398 23378 18450 23390
rect 18398 23314 18450 23326
rect 24222 23378 24274 23390
rect 24222 23314 24274 23326
rect 25790 23378 25842 23390
rect 25790 23314 25842 23326
rect 27582 23378 27634 23390
rect 27582 23314 27634 23326
rect 33742 23378 33794 23390
rect 33742 23314 33794 23326
rect 34526 23378 34578 23390
rect 34526 23314 34578 23326
rect 35086 23378 35138 23390
rect 43374 23378 43426 23390
rect 47182 23378 47234 23390
rect 36642 23326 36654 23378
rect 36706 23326 36718 23378
rect 45714 23326 45726 23378
rect 45778 23326 45790 23378
rect 35086 23314 35138 23326
rect 43374 23314 43426 23326
rect 47182 23314 47234 23326
rect 51102 23378 51154 23390
rect 51102 23314 51154 23326
rect 71710 23378 71762 23390
rect 71710 23314 71762 23326
rect 74398 23378 74450 23390
rect 74398 23314 74450 23326
rect 17502 23266 17554 23278
rect 2034 23214 2046 23266
rect 2098 23214 2110 23266
rect 17502 23202 17554 23214
rect 17614 23266 17666 23278
rect 17614 23202 17666 23214
rect 19518 23266 19570 23278
rect 19518 23202 19570 23214
rect 19630 23266 19682 23278
rect 19630 23202 19682 23214
rect 23886 23266 23938 23278
rect 23886 23202 23938 23214
rect 23998 23266 24050 23278
rect 41246 23266 41298 23278
rect 35858 23214 35870 23266
rect 35922 23214 35934 23266
rect 23998 23202 24050 23214
rect 41246 23202 41298 23214
rect 41694 23266 41746 23278
rect 47966 23266 48018 23278
rect 42802 23214 42814 23266
rect 42866 23214 42878 23266
rect 44482 23214 44494 23266
rect 44546 23214 44558 23266
rect 46498 23214 46510 23266
rect 46562 23214 46574 23266
rect 47506 23214 47518 23266
rect 47570 23214 47582 23266
rect 41694 23202 41746 23214
rect 47966 23202 48018 23214
rect 76862 23266 76914 23278
rect 76862 23202 76914 23214
rect 77086 23266 77138 23278
rect 77086 23202 77138 23214
rect 77534 23266 77586 23278
rect 77534 23202 77586 23214
rect 77758 23266 77810 23278
rect 77758 23202 77810 23214
rect 1710 23154 1762 23166
rect 1710 23090 1762 23102
rect 19854 23154 19906 23166
rect 25118 23154 25170 23166
rect 20290 23102 20302 23154
rect 20354 23102 20366 23154
rect 19854 23090 19906 23102
rect 25118 23090 25170 23102
rect 25566 23154 25618 23166
rect 25566 23090 25618 23102
rect 26910 23154 26962 23166
rect 26910 23090 26962 23102
rect 27358 23154 27410 23166
rect 34190 23154 34242 23166
rect 27906 23102 27918 23154
rect 27970 23102 27982 23154
rect 27358 23090 27410 23102
rect 34190 23090 34242 23102
rect 34302 23154 34354 23166
rect 34302 23090 34354 23102
rect 34638 23154 34690 23166
rect 34638 23090 34690 23102
rect 35198 23154 35250 23166
rect 40910 23154 40962 23166
rect 35746 23102 35758 23154
rect 35810 23102 35822 23154
rect 37314 23102 37326 23154
rect 37378 23102 37390 23154
rect 37650 23102 37662 23154
rect 37714 23102 37726 23154
rect 39778 23102 39790 23154
rect 39842 23102 39854 23154
rect 35198 23090 35250 23102
rect 40910 23090 40962 23102
rect 41582 23154 41634 23166
rect 47854 23154 47906 23166
rect 42354 23102 42366 23154
rect 42418 23102 42430 23154
rect 44146 23102 44158 23154
rect 44210 23102 44222 23154
rect 45602 23102 45614 23154
rect 45666 23102 45678 23154
rect 41582 23090 41634 23102
rect 47854 23090 47906 23102
rect 48190 23154 48242 23166
rect 48190 23090 48242 23102
rect 48862 23154 48914 23166
rect 72146 23102 72158 23154
rect 72210 23102 72222 23154
rect 72930 23102 72942 23154
rect 72994 23102 73006 23154
rect 73490 23102 73502 23154
rect 73554 23102 73566 23154
rect 74498 23102 74510 23154
rect 74562 23102 74574 23154
rect 74834 23102 74846 23154
rect 74898 23102 74910 23154
rect 75954 23102 75966 23154
rect 76018 23102 76030 23154
rect 76178 23102 76190 23154
rect 76242 23102 76254 23154
rect 48862 23090 48914 23102
rect 2494 23042 2546 23054
rect 2494 22978 2546 22990
rect 16830 23042 16882 23054
rect 16830 22978 16882 22990
rect 19182 23042 19234 23054
rect 24558 23042 24610 23054
rect 21074 22990 21086 23042
rect 21138 22990 21150 23042
rect 23202 22990 23214 23042
rect 23266 22990 23278 23042
rect 19182 22978 19234 22990
rect 24558 22978 24610 22990
rect 25678 23042 25730 23054
rect 25678 22978 25730 22990
rect 27470 23042 27522 23054
rect 40350 23042 40402 23054
rect 49310 23042 49362 23054
rect 28690 22990 28702 23042
rect 28754 22990 28766 23042
rect 30818 22990 30830 23042
rect 30882 22990 30894 23042
rect 39442 22990 39454 23042
rect 39506 22990 39518 23042
rect 42242 22990 42254 23042
rect 42306 22990 42318 23042
rect 49186 22990 49198 23042
rect 49250 22990 49262 23042
rect 27470 22978 27522 22990
rect 40350 22978 40402 22990
rect 17502 22930 17554 22942
rect 17502 22866 17554 22878
rect 35086 22930 35138 22942
rect 35086 22866 35138 22878
rect 41694 22930 41746 22942
rect 48738 22878 48750 22930
rect 48802 22927 48814 22930
rect 49201 22927 49247 22990
rect 49310 22978 49362 22990
rect 49870 23042 49922 23054
rect 49870 22978 49922 22990
rect 50206 23042 50258 23054
rect 74513 23039 74559 23102
rect 74834 23039 74846 23042
rect 74513 22993 74846 23039
rect 74834 22990 74846 22993
rect 74898 22990 74910 23042
rect 77186 22990 77198 23042
rect 77250 22990 77262 23042
rect 77858 22990 77870 23042
rect 77922 22990 77934 23042
rect 50206 22978 50258 22990
rect 72382 22930 72434 22942
rect 50194 22927 50206 22930
rect 48802 22881 50206 22927
rect 48802 22878 48814 22881
rect 50194 22878 50206 22881
rect 50258 22878 50270 22930
rect 41694 22866 41746 22878
rect 72382 22866 72434 22878
rect 75070 22930 75122 22942
rect 76402 22878 76414 22930
rect 76466 22927 76478 22930
rect 76626 22927 76638 22930
rect 76466 22881 76638 22927
rect 76466 22878 76478 22881
rect 76626 22878 76638 22881
rect 76690 22878 76702 22930
rect 75070 22866 75122 22878
rect 1344 22762 78624 22796
rect 1344 22710 4478 22762
rect 4530 22710 4582 22762
rect 4634 22710 4686 22762
rect 4738 22710 35198 22762
rect 35250 22710 35302 22762
rect 35354 22710 35406 22762
rect 35458 22710 65918 22762
rect 65970 22710 66022 22762
rect 66074 22710 66126 22762
rect 66178 22710 78624 22762
rect 1344 22676 78624 22710
rect 74174 22594 74226 22606
rect 50530 22542 50542 22594
rect 50594 22591 50606 22594
rect 51090 22591 51102 22594
rect 50594 22545 51102 22591
rect 50594 22542 50606 22545
rect 51090 22542 51102 22545
rect 51154 22542 51166 22594
rect 51314 22542 51326 22594
rect 51378 22591 51390 22594
rect 51762 22591 51774 22594
rect 51378 22545 51774 22591
rect 51378 22542 51390 22545
rect 51762 22542 51774 22545
rect 51826 22542 51838 22594
rect 74174 22530 74226 22542
rect 77534 22594 77586 22606
rect 77534 22530 77586 22542
rect 77870 22594 77922 22606
rect 77870 22530 77922 22542
rect 20414 22482 20466 22494
rect 19394 22430 19406 22482
rect 19458 22430 19470 22482
rect 20414 22418 20466 22430
rect 21758 22482 21810 22494
rect 21758 22418 21810 22430
rect 23102 22482 23154 22494
rect 42030 22482 42082 22494
rect 44830 22482 44882 22494
rect 50430 22482 50482 22494
rect 25106 22430 25118 22482
rect 25170 22430 25182 22482
rect 27234 22430 27246 22482
rect 27298 22430 27310 22482
rect 37314 22430 37326 22482
rect 37378 22430 37390 22482
rect 43362 22430 43374 22482
rect 43426 22430 43438 22482
rect 48626 22430 48638 22482
rect 48690 22430 48702 22482
rect 23102 22418 23154 22430
rect 42030 22418 42082 22430
rect 44830 22418 44882 22430
rect 50430 22418 50482 22430
rect 51774 22482 51826 22494
rect 51774 22418 51826 22430
rect 53790 22482 53842 22494
rect 53790 22418 53842 22430
rect 54238 22482 54290 22494
rect 54238 22418 54290 22430
rect 71710 22482 71762 22494
rect 71710 22418 71762 22430
rect 72158 22482 72210 22494
rect 76526 22482 76578 22494
rect 72482 22430 72494 22482
rect 72546 22430 72558 22482
rect 75058 22430 75070 22482
rect 75122 22430 75134 22482
rect 72158 22418 72210 22430
rect 76526 22418 76578 22430
rect 21198 22370 21250 22382
rect 27582 22370 27634 22382
rect 16594 22318 16606 22370
rect 16658 22318 16670 22370
rect 19954 22318 19966 22370
rect 20018 22318 20030 22370
rect 23538 22318 23550 22370
rect 23602 22318 23614 22370
rect 24322 22318 24334 22370
rect 24386 22318 24398 22370
rect 21198 22306 21250 22318
rect 27582 22306 27634 22318
rect 30830 22370 30882 22382
rect 30830 22306 30882 22318
rect 30942 22370 30994 22382
rect 37774 22370 37826 22382
rect 43822 22370 43874 22382
rect 46062 22370 46114 22382
rect 34290 22318 34302 22370
rect 34354 22318 34366 22370
rect 35298 22318 35310 22370
rect 35362 22318 35374 22370
rect 38994 22318 39006 22370
rect 39058 22318 39070 22370
rect 41346 22318 41358 22370
rect 41410 22318 41422 22370
rect 42466 22318 42478 22370
rect 42530 22318 42542 22370
rect 45378 22318 45390 22370
rect 45442 22318 45454 22370
rect 30942 22306 30994 22318
rect 37774 22306 37826 22318
rect 43822 22306 43874 22318
rect 46062 22306 46114 22318
rect 46510 22370 46562 22382
rect 46510 22306 46562 22318
rect 46734 22370 46786 22382
rect 46734 22306 46786 22318
rect 47406 22370 47458 22382
rect 47406 22306 47458 22318
rect 47518 22370 47570 22382
rect 47518 22306 47570 22318
rect 49422 22370 49474 22382
rect 49422 22306 49474 22318
rect 49982 22370 50034 22382
rect 49982 22306 50034 22318
rect 52782 22370 52834 22382
rect 52782 22306 52834 22318
rect 53342 22370 53394 22382
rect 72258 22318 72270 22370
rect 72322 22318 72334 22370
rect 73266 22318 73278 22370
rect 73330 22318 73342 22370
rect 73602 22318 73614 22370
rect 73666 22318 73678 22370
rect 73938 22318 73950 22370
rect 74002 22318 74014 22370
rect 74946 22318 74958 22370
rect 75010 22318 75022 22370
rect 53342 22306 53394 22318
rect 44942 22258 44994 22270
rect 17266 22206 17278 22258
rect 17330 22206 17342 22258
rect 19730 22206 19742 22258
rect 19794 22206 19806 22258
rect 20738 22206 20750 22258
rect 20802 22206 20814 22258
rect 23762 22206 23774 22258
rect 23826 22206 23838 22258
rect 33506 22206 33518 22258
rect 33570 22206 33582 22258
rect 35746 22206 35758 22258
rect 35810 22206 35822 22258
rect 39442 22206 39454 22258
rect 39506 22206 39518 22258
rect 41234 22206 41246 22258
rect 41298 22206 41310 22258
rect 44942 22194 44994 22206
rect 47070 22258 47122 22270
rect 47070 22194 47122 22206
rect 47966 22258 48018 22270
rect 47966 22194 48018 22206
rect 48078 22258 48130 22270
rect 48078 22194 48130 22206
rect 76750 22258 76802 22270
rect 76750 22194 76802 22206
rect 21646 22146 21698 22158
rect 21646 22082 21698 22094
rect 21870 22146 21922 22158
rect 21870 22082 21922 22094
rect 22990 22146 23042 22158
rect 22990 22082 23042 22094
rect 27694 22146 27746 22158
rect 44270 22146 44322 22158
rect 34290 22094 34302 22146
rect 34354 22094 34366 22146
rect 40562 22094 40574 22146
rect 40626 22094 40638 22146
rect 27694 22082 27746 22094
rect 44270 22082 44322 22094
rect 45614 22146 45666 22158
rect 45614 22082 45666 22094
rect 46398 22146 46450 22158
rect 46398 22082 46450 22094
rect 47294 22146 47346 22158
rect 47294 22082 47346 22094
rect 48302 22146 48354 22158
rect 48302 22082 48354 22094
rect 49086 22146 49138 22158
rect 49086 22082 49138 22094
rect 50878 22146 50930 22158
rect 50878 22082 50930 22094
rect 51438 22146 51490 22158
rect 51438 22082 51490 22094
rect 77086 22146 77138 22158
rect 77086 22082 77138 22094
rect 77758 22146 77810 22158
rect 77758 22082 77810 22094
rect 1344 21978 78624 22012
rect 1344 21926 19838 21978
rect 19890 21926 19942 21978
rect 19994 21926 20046 21978
rect 20098 21926 50558 21978
rect 50610 21926 50662 21978
rect 50714 21926 50766 21978
rect 50818 21926 78624 21978
rect 1344 21892 78624 21926
rect 17502 21810 17554 21822
rect 2034 21758 2046 21810
rect 2098 21758 2110 21810
rect 17502 21746 17554 21758
rect 17838 21810 17890 21822
rect 17838 21746 17890 21758
rect 24222 21810 24274 21822
rect 35422 21810 35474 21822
rect 26226 21758 26238 21810
rect 26290 21758 26302 21810
rect 24222 21746 24274 21758
rect 35422 21746 35474 21758
rect 36206 21810 36258 21822
rect 41246 21810 41298 21822
rect 38210 21758 38222 21810
rect 38274 21758 38286 21810
rect 36206 21746 36258 21758
rect 41246 21746 41298 21758
rect 47742 21810 47794 21822
rect 56030 21810 56082 21822
rect 48850 21758 48862 21810
rect 48914 21758 48926 21810
rect 55010 21758 55022 21810
rect 55074 21758 55086 21810
rect 47742 21746 47794 21758
rect 56030 21746 56082 21758
rect 70030 21810 70082 21822
rect 70030 21746 70082 21758
rect 74622 21810 74674 21822
rect 74622 21746 74674 21758
rect 75854 21810 75906 21822
rect 75854 21746 75906 21758
rect 77310 21810 77362 21822
rect 77310 21746 77362 21758
rect 77870 21810 77922 21822
rect 77870 21746 77922 21758
rect 23886 21698 23938 21710
rect 22306 21646 22318 21698
rect 22370 21646 22382 21698
rect 23886 21634 23938 21646
rect 23998 21698 24050 21710
rect 23998 21634 24050 21646
rect 25678 21698 25730 21710
rect 42478 21698 42530 21710
rect 55582 21698 55634 21710
rect 75182 21698 75234 21710
rect 37426 21646 37438 21698
rect 37490 21646 37502 21698
rect 39442 21646 39454 21698
rect 39506 21646 39518 21698
rect 44034 21646 44046 21698
rect 44098 21646 44110 21698
rect 46162 21646 46174 21698
rect 46226 21646 46238 21698
rect 49858 21646 49870 21698
rect 49922 21646 49934 21698
rect 50866 21646 50878 21698
rect 50930 21646 50942 21698
rect 51762 21646 51774 21698
rect 51826 21646 51838 21698
rect 54450 21646 54462 21698
rect 54514 21646 54526 21698
rect 72258 21646 72270 21698
rect 72322 21646 72334 21698
rect 25678 21634 25730 21646
rect 42478 21634 42530 21646
rect 55582 21634 55634 21646
rect 75182 21634 75234 21646
rect 76638 21698 76690 21710
rect 76638 21634 76690 21646
rect 77198 21698 77250 21710
rect 77198 21634 77250 21646
rect 78206 21698 78258 21710
rect 78206 21634 78258 21646
rect 1710 21586 1762 21598
rect 1710 21522 1762 21534
rect 17726 21586 17778 21598
rect 17726 21522 17778 21534
rect 17950 21586 18002 21598
rect 35086 21586 35138 21598
rect 19170 21534 19182 21586
rect 19234 21534 19246 21586
rect 22530 21534 22542 21586
rect 22594 21534 22606 21586
rect 26450 21534 26462 21586
rect 26514 21534 26526 21586
rect 17950 21522 18002 21534
rect 35086 21522 35138 21534
rect 35534 21586 35586 21598
rect 35534 21522 35586 21534
rect 35758 21586 35810 21598
rect 35758 21522 35810 21534
rect 35982 21586 36034 21598
rect 35982 21522 36034 21534
rect 36430 21586 36482 21598
rect 36430 21522 36482 21534
rect 36542 21586 36594 21598
rect 47406 21586 47458 21598
rect 37538 21534 37550 21586
rect 37602 21534 37614 21586
rect 39218 21534 39230 21586
rect 39282 21534 39294 21586
rect 44930 21534 44942 21586
rect 44994 21534 45006 21586
rect 45826 21534 45838 21586
rect 45890 21534 45902 21586
rect 36542 21522 36594 21534
rect 47406 21522 47458 21534
rect 47630 21586 47682 21598
rect 47630 21522 47682 21534
rect 47966 21586 48018 21598
rect 53118 21586 53170 21598
rect 74062 21586 74114 21598
rect 48738 21534 48750 21586
rect 48802 21534 48814 21586
rect 49410 21534 49422 21586
rect 49474 21534 49486 21586
rect 50194 21534 50206 21586
rect 50258 21534 50270 21586
rect 51314 21534 51326 21586
rect 51378 21534 51390 21586
rect 52210 21534 52222 21586
rect 52274 21534 52286 21586
rect 52770 21534 52782 21586
rect 52834 21534 52846 21586
rect 54338 21534 54350 21586
rect 54402 21534 54414 21586
rect 54898 21534 54910 21586
rect 54962 21534 54974 21586
rect 70242 21534 70254 21586
rect 70306 21534 70318 21586
rect 71362 21534 71374 21586
rect 71426 21534 71438 21586
rect 71586 21534 71598 21586
rect 71650 21534 71662 21586
rect 72594 21534 72606 21586
rect 72658 21534 72670 21586
rect 73266 21534 73278 21586
rect 73330 21534 73342 21586
rect 47966 21522 48018 21534
rect 53118 21522 53170 21534
rect 74062 21522 74114 21534
rect 74846 21586 74898 21598
rect 74846 21522 74898 21534
rect 75518 21586 75570 21598
rect 75518 21522 75570 21534
rect 76862 21586 76914 21598
rect 77522 21534 77534 21586
rect 77586 21534 77598 21586
rect 76862 21522 76914 21534
rect 2494 21474 2546 21486
rect 2494 21410 2546 21422
rect 18398 21474 18450 21486
rect 23550 21474 23602 21486
rect 33630 21474 33682 21486
rect 19842 21422 19854 21474
rect 19906 21422 19918 21474
rect 21970 21422 21982 21474
rect 22034 21422 22046 21474
rect 33282 21422 33294 21474
rect 33346 21422 33358 21474
rect 18398 21410 18450 21422
rect 23550 21410 23602 21422
rect 33630 21410 33682 21422
rect 34526 21474 34578 21486
rect 34526 21410 34578 21422
rect 34862 21474 34914 21486
rect 46622 21474 46674 21486
rect 53678 21474 53730 21486
rect 43250 21422 43262 21474
rect 43314 21422 43326 21474
rect 50866 21422 50878 21474
rect 50930 21422 50942 21474
rect 52322 21422 52334 21474
rect 52386 21422 52398 21474
rect 70578 21422 70590 21474
rect 70642 21422 70654 21474
rect 73042 21422 73054 21474
rect 73106 21422 73118 21474
rect 76514 21422 76526 21474
rect 76578 21422 76590 21474
rect 34862 21410 34914 21422
rect 46622 21410 46674 21422
rect 53678 21410 53730 21422
rect 42030 21362 42082 21374
rect 42030 21298 42082 21310
rect 1344 21194 78624 21228
rect 1344 21142 4478 21194
rect 4530 21142 4582 21194
rect 4634 21142 4686 21194
rect 4738 21142 35198 21194
rect 35250 21142 35302 21194
rect 35354 21142 35406 21194
rect 35458 21142 65918 21194
rect 65970 21142 66022 21194
rect 66074 21142 66126 21194
rect 66178 21142 78624 21194
rect 1344 21108 78624 21142
rect 75294 21026 75346 21038
rect 75294 20962 75346 20974
rect 77086 21026 77138 21038
rect 77086 20962 77138 20974
rect 77422 21026 77474 21038
rect 77422 20962 77474 20974
rect 21758 20914 21810 20926
rect 34414 20914 34466 20926
rect 24994 20862 25006 20914
rect 25058 20862 25070 20914
rect 30146 20862 30158 20914
rect 30210 20862 30222 20914
rect 33618 20862 33630 20914
rect 33682 20862 33694 20914
rect 21758 20850 21810 20862
rect 34414 20850 34466 20862
rect 35310 20914 35362 20926
rect 35310 20850 35362 20862
rect 38110 20914 38162 20926
rect 57150 20914 57202 20926
rect 46162 20862 46174 20914
rect 46226 20862 46238 20914
rect 47058 20862 47070 20914
rect 47122 20862 47134 20914
rect 51314 20862 51326 20914
rect 51378 20862 51390 20914
rect 38110 20850 38162 20862
rect 57150 20850 57202 20862
rect 70926 20914 70978 20926
rect 74734 20914 74786 20926
rect 71250 20862 71262 20914
rect 71314 20862 71326 20914
rect 72146 20862 72158 20914
rect 72210 20862 72222 20914
rect 72930 20862 72942 20914
rect 72994 20862 73006 20914
rect 73826 20862 73838 20914
rect 73890 20862 73902 20914
rect 70926 20850 70978 20862
rect 74734 20850 74786 20862
rect 77534 20914 77586 20926
rect 77534 20850 77586 20862
rect 78318 20914 78370 20926
rect 78318 20850 78370 20862
rect 18622 20802 18674 20814
rect 25342 20802 25394 20814
rect 22082 20750 22094 20802
rect 22146 20750 22158 20802
rect 18622 20738 18674 20750
rect 25342 20738 25394 20750
rect 26014 20802 26066 20814
rect 26014 20738 26066 20750
rect 27246 20802 27298 20814
rect 27246 20738 27298 20750
rect 29038 20802 29090 20814
rect 29038 20738 29090 20750
rect 29486 20802 29538 20814
rect 34190 20802 34242 20814
rect 30818 20750 30830 20802
rect 30882 20750 30894 20802
rect 29486 20738 29538 20750
rect 34190 20738 34242 20750
rect 34862 20802 34914 20814
rect 34862 20738 34914 20750
rect 35758 20802 35810 20814
rect 35758 20738 35810 20750
rect 36430 20802 36482 20814
rect 36430 20738 36482 20750
rect 37886 20802 37938 20814
rect 37886 20738 37938 20750
rect 39342 20802 39394 20814
rect 42926 20802 42978 20814
rect 44830 20802 44882 20814
rect 45726 20802 45778 20814
rect 41234 20750 41246 20802
rect 41298 20750 41310 20802
rect 43250 20750 43262 20802
rect 43314 20750 43326 20802
rect 45266 20750 45278 20802
rect 45330 20750 45342 20802
rect 46610 20750 46622 20802
rect 46674 20750 46686 20802
rect 47170 20750 47182 20802
rect 47234 20750 47246 20802
rect 48290 20750 48302 20802
rect 48354 20750 48366 20802
rect 49410 20750 49422 20802
rect 49474 20750 49486 20802
rect 49746 20750 49758 20802
rect 49810 20750 49822 20802
rect 50418 20750 50430 20802
rect 50482 20750 50494 20802
rect 51650 20750 51662 20802
rect 51714 20750 51726 20802
rect 52770 20750 52782 20802
rect 52834 20750 52846 20802
rect 53218 20750 53230 20802
rect 53282 20750 53294 20802
rect 54114 20750 54126 20802
rect 54178 20750 54190 20802
rect 54674 20750 54686 20802
rect 54738 20750 54750 20802
rect 55570 20750 55582 20802
rect 55634 20750 55646 20802
rect 56130 20750 56142 20802
rect 56194 20750 56206 20802
rect 71026 20750 71038 20802
rect 71090 20750 71102 20802
rect 72034 20750 72046 20802
rect 72098 20750 72110 20802
rect 72706 20750 72718 20802
rect 72770 20750 72782 20802
rect 73490 20750 73502 20802
rect 73554 20750 73566 20802
rect 76738 20750 76750 20802
rect 76802 20750 76814 20802
rect 77746 20750 77758 20802
rect 77810 20750 77822 20802
rect 39342 20738 39394 20750
rect 42926 20738 42978 20750
rect 44830 20738 44882 20750
rect 45726 20738 45778 20750
rect 18958 20690 19010 20702
rect 2034 20638 2046 20690
rect 2098 20638 2110 20690
rect 18958 20626 19010 20638
rect 19070 20690 19122 20702
rect 25678 20690 25730 20702
rect 22866 20638 22878 20690
rect 22930 20638 22942 20690
rect 19070 20626 19122 20638
rect 25678 20626 25730 20638
rect 26350 20690 26402 20702
rect 26350 20626 26402 20638
rect 30382 20690 30434 20702
rect 34638 20690 34690 20702
rect 31490 20638 31502 20690
rect 31554 20638 31566 20690
rect 30382 20626 30434 20638
rect 34638 20626 34690 20638
rect 35198 20690 35250 20702
rect 35198 20626 35250 20638
rect 35534 20690 35586 20702
rect 35534 20626 35586 20638
rect 36094 20690 36146 20702
rect 38334 20690 38386 20702
rect 36978 20638 36990 20690
rect 37042 20638 37054 20690
rect 36094 20626 36146 20638
rect 38334 20626 38386 20638
rect 38558 20690 38610 20702
rect 38558 20626 38610 20638
rect 39006 20690 39058 20702
rect 39006 20626 39058 20638
rect 40014 20690 40066 20702
rect 75630 20690 75682 20702
rect 40338 20638 40350 20690
rect 40402 20638 40414 20690
rect 41122 20638 41134 20690
rect 41186 20638 41198 20690
rect 47730 20638 47742 20690
rect 47794 20638 47806 20690
rect 48626 20638 48638 20690
rect 48690 20638 48702 20690
rect 50642 20638 50654 20690
rect 50706 20638 50718 20690
rect 53442 20638 53454 20690
rect 53506 20638 53518 20690
rect 55234 20638 55246 20690
rect 55298 20638 55310 20690
rect 56242 20638 56254 20690
rect 56306 20638 56318 20690
rect 40014 20626 40066 20638
rect 75630 20626 75682 20638
rect 1710 20578 1762 20590
rect 1710 20514 1762 20526
rect 2494 20578 2546 20590
rect 2494 20514 2546 20526
rect 19294 20578 19346 20590
rect 19294 20514 19346 20526
rect 20638 20578 20690 20590
rect 20638 20514 20690 20526
rect 21646 20578 21698 20590
rect 21646 20514 21698 20526
rect 26126 20578 26178 20590
rect 26126 20514 26178 20526
rect 26574 20578 26626 20590
rect 27358 20578 27410 20590
rect 26898 20526 26910 20578
rect 26962 20526 26974 20578
rect 26574 20514 26626 20526
rect 27358 20514 27410 20526
rect 27582 20578 27634 20590
rect 27582 20514 27634 20526
rect 27918 20578 27970 20590
rect 27918 20514 27970 20526
rect 29598 20578 29650 20590
rect 29598 20514 29650 20526
rect 29710 20578 29762 20590
rect 29710 20514 29762 20526
rect 37326 20578 37378 20590
rect 37326 20514 37378 20526
rect 39678 20578 39730 20590
rect 39678 20514 39730 20526
rect 40686 20578 40738 20590
rect 75406 20578 75458 20590
rect 43026 20526 43038 20578
rect 43090 20526 43102 20578
rect 49186 20526 49198 20578
rect 49250 20526 49262 20578
rect 49858 20526 49870 20578
rect 49922 20526 49934 20578
rect 52882 20526 52894 20578
rect 52946 20526 52958 20578
rect 54226 20526 54238 20578
rect 54290 20526 54302 20578
rect 55682 20526 55694 20578
rect 55746 20526 55758 20578
rect 40686 20514 40738 20526
rect 75406 20514 75458 20526
rect 76302 20578 76354 20590
rect 76302 20514 76354 20526
rect 76974 20578 77026 20590
rect 76974 20514 77026 20526
rect 1344 20410 78624 20444
rect 1344 20358 19838 20410
rect 19890 20358 19942 20410
rect 19994 20358 20046 20410
rect 20098 20358 50558 20410
rect 50610 20358 50662 20410
rect 50714 20358 50766 20410
rect 50818 20358 78624 20410
rect 1344 20324 78624 20358
rect 18734 20242 18786 20254
rect 18734 20178 18786 20190
rect 31502 20242 31554 20254
rect 31502 20178 31554 20190
rect 33966 20242 34018 20254
rect 33966 20178 34018 20190
rect 34414 20242 34466 20254
rect 34414 20178 34466 20190
rect 39678 20242 39730 20254
rect 48078 20242 48130 20254
rect 72606 20242 72658 20254
rect 42802 20190 42814 20242
rect 42866 20190 42878 20242
rect 46498 20190 46510 20242
rect 46562 20190 46574 20242
rect 52882 20190 52894 20242
rect 52946 20190 52958 20242
rect 54338 20190 54350 20242
rect 54402 20190 54414 20242
rect 39678 20178 39730 20190
rect 48078 20178 48130 20190
rect 72606 20178 72658 20190
rect 74622 20242 74674 20254
rect 74622 20178 74674 20190
rect 25230 20130 25282 20142
rect 18386 20078 18398 20130
rect 18450 20078 18462 20130
rect 25230 20066 25282 20078
rect 26238 20130 26290 20142
rect 26238 20066 26290 20078
rect 26350 20130 26402 20142
rect 26350 20066 26402 20078
rect 26910 20130 26962 20142
rect 31390 20130 31442 20142
rect 28466 20078 28478 20130
rect 28530 20078 28542 20130
rect 26910 20066 26962 20078
rect 31390 20066 31442 20078
rect 33518 20130 33570 20142
rect 33518 20066 33570 20078
rect 34862 20130 34914 20142
rect 34862 20066 34914 20078
rect 35534 20130 35586 20142
rect 38782 20130 38834 20142
rect 52110 20130 52162 20142
rect 56702 20130 56754 20142
rect 36306 20078 36318 20130
rect 36370 20078 36382 20130
rect 41346 20078 41358 20130
rect 41410 20078 41422 20130
rect 42914 20078 42926 20130
rect 42978 20078 42990 20130
rect 44482 20078 44494 20130
rect 44546 20078 44558 20130
rect 46946 20078 46958 20130
rect 47010 20078 47022 20130
rect 49410 20078 49422 20130
rect 49474 20078 49486 20130
rect 53442 20078 53454 20130
rect 53506 20078 53518 20130
rect 55234 20078 55246 20130
rect 55298 20078 55310 20130
rect 35534 20066 35586 20078
rect 38782 20066 38834 20078
rect 52110 20066 52162 20078
rect 56702 20066 56754 20078
rect 75182 20130 75234 20142
rect 75182 20066 75234 20078
rect 76190 20130 76242 20142
rect 76190 20066 76242 20078
rect 76302 20130 76354 20142
rect 76302 20066 76354 20078
rect 76750 20130 76802 20142
rect 76750 20066 76802 20078
rect 77086 20130 77138 20142
rect 77086 20066 77138 20078
rect 77870 20130 77922 20142
rect 77870 20066 77922 20078
rect 26574 20018 26626 20030
rect 30942 20018 30994 20030
rect 24658 19966 24670 20018
rect 24722 19966 24734 20018
rect 27794 19966 27806 20018
rect 27858 19966 27870 20018
rect 26574 19954 26626 19966
rect 30942 19954 30994 19966
rect 31614 20018 31666 20030
rect 31614 19954 31666 19966
rect 35422 20018 35474 20030
rect 39342 20018 39394 20030
rect 36194 19966 36206 20018
rect 36258 19966 36270 20018
rect 37650 19966 37662 20018
rect 37714 19966 37726 20018
rect 37986 19966 37998 20018
rect 38050 19966 38062 20018
rect 35422 19954 35474 19966
rect 39342 19954 39394 19966
rect 39678 20018 39730 20030
rect 39678 19954 39730 19966
rect 39902 20018 39954 20030
rect 48862 20018 48914 20030
rect 51102 20018 51154 20030
rect 55806 20018 55858 20030
rect 41122 19966 41134 20018
rect 41186 19966 41198 20018
rect 43026 19966 43038 20018
rect 43090 19966 43102 20018
rect 44706 19966 44718 20018
rect 44770 19966 44782 20018
rect 46610 19966 46622 20018
rect 46674 19966 46686 20018
rect 50082 19966 50094 20018
rect 50146 19966 50158 20018
rect 51426 19966 51438 20018
rect 51490 19966 51502 20018
rect 52770 19966 52782 20018
rect 52834 19966 52846 20018
rect 53330 19966 53342 20018
rect 53394 19966 53406 20018
rect 54450 19966 54462 20018
rect 54514 19966 54526 20018
rect 54786 19966 54798 20018
rect 54850 19966 54862 20018
rect 39902 19954 39954 19966
rect 48862 19954 48914 19966
rect 51102 19954 51154 19966
rect 55806 19954 55858 19966
rect 76078 20018 76130 20030
rect 78082 19966 78094 20018
rect 78146 19966 78158 20018
rect 76078 19954 76130 19966
rect 27470 19906 27522 19918
rect 32174 19906 32226 19918
rect 19618 19854 19630 19906
rect 19682 19854 19694 19906
rect 25554 19854 25566 19906
rect 25618 19854 25630 19906
rect 30594 19854 30606 19906
rect 30658 19854 30670 19906
rect 27470 19842 27522 19854
rect 32174 19842 32226 19854
rect 32622 19906 32674 19918
rect 32622 19842 32674 19854
rect 33406 19906 33458 19918
rect 33406 19842 33458 19854
rect 33854 19906 33906 19918
rect 33854 19842 33906 19854
rect 34302 19906 34354 19918
rect 34302 19842 34354 19854
rect 34750 19906 34802 19918
rect 34750 19842 34802 19854
rect 48190 19906 48242 19918
rect 48190 19842 48242 19854
rect 77646 19906 77698 19918
rect 77646 19842 77698 19854
rect 1344 19626 78624 19660
rect 1344 19574 4478 19626
rect 4530 19574 4582 19626
rect 4634 19574 4686 19626
rect 4738 19574 35198 19626
rect 35250 19574 35302 19626
rect 35354 19574 35406 19626
rect 35458 19574 65918 19626
rect 65970 19574 66022 19626
rect 66074 19574 66126 19626
rect 66178 19574 78624 19626
rect 1344 19540 78624 19574
rect 76750 19458 76802 19470
rect 76750 19394 76802 19406
rect 77422 19458 77474 19470
rect 77422 19394 77474 19406
rect 18846 19346 18898 19358
rect 18846 19282 18898 19294
rect 20302 19346 20354 19358
rect 20302 19282 20354 19294
rect 21758 19346 21810 19358
rect 21758 19282 21810 19294
rect 22766 19346 22818 19358
rect 22766 19282 22818 19294
rect 24446 19346 24498 19358
rect 24446 19282 24498 19294
rect 35534 19346 35586 19358
rect 35534 19282 35586 19294
rect 36430 19346 36482 19358
rect 36430 19282 36482 19294
rect 38110 19346 38162 19358
rect 38110 19282 38162 19294
rect 43934 19346 43986 19358
rect 43934 19282 43986 19294
rect 48526 19346 48578 19358
rect 48526 19282 48578 19294
rect 51774 19346 51826 19358
rect 51774 19282 51826 19294
rect 78318 19346 78370 19358
rect 78318 19282 78370 19294
rect 19742 19234 19794 19246
rect 19742 19170 19794 19182
rect 20414 19234 20466 19246
rect 20414 19170 20466 19182
rect 22318 19234 22370 19246
rect 22318 19170 22370 19182
rect 22654 19234 22706 19246
rect 22654 19170 22706 19182
rect 26350 19234 26402 19246
rect 26350 19170 26402 19182
rect 26686 19234 26738 19246
rect 26686 19170 26738 19182
rect 27022 19234 27074 19246
rect 27022 19170 27074 19182
rect 27694 19234 27746 19246
rect 35646 19234 35698 19246
rect 34402 19182 34414 19234
rect 34466 19182 34478 19234
rect 27694 19170 27746 19182
rect 35646 19170 35698 19182
rect 35870 19234 35922 19246
rect 35870 19170 35922 19182
rect 38334 19234 38386 19246
rect 38334 19170 38386 19182
rect 38558 19234 38610 19246
rect 38558 19170 38610 19182
rect 38782 19234 38834 19246
rect 38782 19170 38834 19182
rect 39230 19234 39282 19246
rect 39230 19170 39282 19182
rect 39342 19234 39394 19246
rect 39342 19170 39394 19182
rect 40798 19234 40850 19246
rect 44830 19234 44882 19246
rect 52670 19234 52722 19246
rect 42242 19182 42254 19234
rect 42306 19182 42318 19234
rect 43362 19182 43374 19234
rect 43426 19182 43438 19234
rect 45378 19182 45390 19234
rect 45442 19182 45454 19234
rect 47058 19182 47070 19234
rect 47122 19182 47134 19234
rect 49858 19182 49870 19234
rect 49922 19182 49934 19234
rect 50978 19182 50990 19234
rect 51042 19182 51054 19234
rect 40798 19170 40850 19182
rect 44830 19170 44882 19182
rect 52670 19170 52722 19182
rect 53230 19234 53282 19246
rect 76862 19234 76914 19246
rect 53890 19182 53902 19234
rect 53954 19182 53966 19234
rect 55458 19182 55470 19234
rect 55522 19182 55534 19234
rect 56130 19182 56142 19234
rect 56194 19182 56206 19234
rect 77746 19182 77758 19234
rect 77810 19182 77822 19234
rect 53230 19170 53282 19182
rect 76862 19170 76914 19182
rect 1710 19122 1762 19134
rect 1710 19058 1762 19070
rect 2046 19122 2098 19134
rect 2046 19058 2098 19070
rect 2494 19122 2546 19134
rect 2494 19058 2546 19070
rect 19182 19122 19234 19134
rect 19182 19058 19234 19070
rect 19294 19122 19346 19134
rect 22878 19122 22930 19134
rect 21970 19070 21982 19122
rect 22034 19070 22046 19122
rect 19294 19058 19346 19070
rect 22878 19058 22930 19070
rect 23550 19122 23602 19134
rect 24782 19122 24834 19134
rect 23874 19070 23886 19122
rect 23938 19070 23950 19122
rect 23550 19058 23602 19070
rect 24782 19058 24834 19070
rect 25118 19122 25170 19134
rect 25118 19058 25170 19070
rect 25454 19122 25506 19134
rect 25454 19058 25506 19070
rect 25790 19122 25842 19134
rect 25790 19058 25842 19070
rect 29150 19122 29202 19134
rect 35422 19122 35474 19134
rect 37998 19122 38050 19134
rect 29474 19070 29486 19122
rect 29538 19070 29550 19122
rect 30258 19070 30270 19122
rect 30322 19070 30334 19122
rect 37650 19070 37662 19122
rect 37714 19070 37726 19122
rect 29150 19058 29202 19070
rect 35422 19058 35474 19070
rect 37998 19058 38050 19070
rect 40126 19122 40178 19134
rect 40126 19058 40178 19070
rect 40462 19122 40514 19134
rect 57374 19122 57426 19134
rect 41234 19070 41246 19122
rect 41298 19070 41310 19122
rect 42914 19070 42926 19122
rect 42978 19070 42990 19122
rect 46946 19070 46958 19122
rect 47010 19070 47022 19122
rect 49298 19070 49310 19122
rect 49362 19070 49374 19122
rect 51090 19070 51102 19122
rect 51154 19070 51166 19122
rect 54114 19070 54126 19122
rect 54178 19070 54190 19122
rect 40462 19058 40514 19070
rect 57374 19058 57426 19070
rect 19518 19010 19570 19022
rect 19518 18946 19570 18958
rect 20190 19010 20242 19022
rect 20190 18946 20242 18958
rect 23102 19010 23154 19022
rect 23102 18946 23154 18958
rect 26462 19010 26514 19022
rect 26462 18946 26514 18958
rect 27470 19010 27522 19022
rect 27470 18946 27522 18958
rect 27582 19010 27634 19022
rect 27582 18946 27634 18958
rect 28142 19010 28194 19022
rect 28142 18946 28194 18958
rect 28590 19010 28642 19022
rect 28590 18946 28642 18958
rect 37326 19010 37378 19022
rect 37326 18946 37378 18958
rect 39118 19010 39170 19022
rect 39118 18946 39170 18958
rect 39790 19010 39842 19022
rect 39790 18946 39842 18958
rect 40574 19010 40626 19022
rect 76526 19010 76578 19022
rect 46834 18958 46846 19010
rect 46898 18958 46910 19010
rect 55346 18958 55358 19010
rect 55410 18958 55422 19010
rect 40574 18946 40626 18958
rect 76526 18946 76578 18958
rect 76974 19010 77026 19022
rect 76974 18946 77026 18958
rect 77534 19010 77586 19022
rect 77534 18946 77586 18958
rect 1344 18842 78624 18876
rect 1344 18790 19838 18842
rect 19890 18790 19942 18842
rect 19994 18790 20046 18842
rect 20098 18790 50558 18842
rect 50610 18790 50662 18842
rect 50714 18790 50766 18842
rect 50818 18790 78624 18842
rect 1344 18756 78624 18790
rect 17614 18674 17666 18686
rect 17614 18610 17666 18622
rect 18062 18674 18114 18686
rect 18062 18610 18114 18622
rect 40014 18674 40066 18686
rect 40014 18610 40066 18622
rect 41694 18674 41746 18686
rect 77534 18674 77586 18686
rect 46946 18622 46958 18674
rect 47010 18622 47022 18674
rect 49858 18622 49870 18674
rect 49922 18622 49934 18674
rect 54002 18622 54014 18674
rect 54066 18622 54078 18674
rect 41694 18610 41746 18622
rect 77534 18610 77586 18622
rect 77870 18674 77922 18686
rect 77870 18610 77922 18622
rect 2046 18562 2098 18574
rect 2046 18498 2098 18510
rect 18174 18562 18226 18574
rect 41582 18562 41634 18574
rect 27122 18510 27134 18562
rect 27186 18510 27198 18562
rect 40898 18510 40910 18562
rect 40962 18510 40974 18562
rect 42130 18510 42142 18562
rect 42194 18510 42206 18562
rect 44034 18510 44046 18562
rect 44098 18510 44110 18562
rect 47506 18510 47518 18562
rect 47570 18510 47582 18562
rect 48850 18510 48862 18562
rect 48914 18510 48926 18562
rect 51090 18510 51102 18562
rect 51154 18510 51166 18562
rect 53442 18510 53454 18562
rect 53506 18510 53518 18562
rect 55682 18510 55694 18562
rect 55746 18510 55758 18562
rect 18174 18498 18226 18510
rect 41582 18498 41634 18510
rect 1710 18450 1762 18462
rect 41918 18450 41970 18462
rect 18610 18398 18622 18450
rect 18674 18398 18686 18450
rect 21858 18398 21870 18450
rect 21922 18398 21934 18450
rect 26450 18398 26462 18450
rect 26514 18398 26526 18450
rect 29698 18398 29710 18450
rect 29762 18398 29774 18450
rect 34402 18398 34414 18450
rect 34466 18398 34478 18450
rect 40226 18398 40238 18450
rect 40290 18398 40302 18450
rect 41122 18398 41134 18450
rect 41186 18398 41198 18450
rect 1710 18386 1762 18398
rect 41918 18386 41970 18398
rect 42478 18450 42530 18462
rect 44830 18450 44882 18462
rect 57150 18450 57202 18462
rect 78206 18450 78258 18462
rect 43922 18398 43934 18450
rect 43986 18398 43998 18450
rect 45266 18398 45278 18450
rect 45330 18398 45342 18450
rect 46834 18398 46846 18450
rect 46898 18398 46910 18450
rect 47394 18398 47406 18450
rect 47458 18398 47470 18450
rect 48962 18398 48974 18450
rect 49026 18398 49038 18450
rect 51314 18398 51326 18450
rect 51378 18398 51390 18450
rect 53666 18398 53678 18450
rect 53730 18398 53742 18450
rect 55122 18398 55134 18450
rect 55186 18398 55198 18450
rect 77298 18398 77310 18450
rect 77362 18398 77374 18450
rect 42478 18386 42530 18398
rect 44830 18386 44882 18398
rect 57150 18386 57202 18398
rect 78206 18386 78258 18398
rect 2494 18338 2546 18350
rect 25342 18338 25394 18350
rect 33182 18338 33234 18350
rect 19282 18286 19294 18338
rect 19346 18286 19358 18338
rect 21410 18286 21422 18338
rect 21474 18286 21486 18338
rect 22530 18286 22542 18338
rect 22594 18286 22606 18338
rect 24658 18286 24670 18338
rect 24722 18286 24734 18338
rect 25666 18286 25678 18338
rect 25730 18286 25742 18338
rect 29250 18286 29262 18338
rect 29314 18286 29326 18338
rect 30370 18286 30382 18338
rect 30434 18286 30446 18338
rect 32498 18286 32510 18338
rect 32562 18286 32574 18338
rect 2494 18274 2546 18286
rect 25342 18274 25394 18286
rect 33182 18274 33234 18286
rect 33518 18338 33570 18350
rect 52446 18338 52498 18350
rect 33730 18286 33742 18338
rect 33794 18286 33806 18338
rect 38434 18286 38446 18338
rect 38498 18286 38510 18338
rect 33518 18274 33570 18286
rect 52446 18274 52498 18286
rect 56702 18338 56754 18350
rect 56702 18274 56754 18286
rect 76974 18338 77026 18350
rect 76974 18274 77026 18286
rect 18062 18226 18114 18238
rect 43698 18174 43710 18226
rect 43762 18174 43774 18226
rect 18062 18162 18114 18174
rect 1344 18058 78624 18092
rect 1344 18006 4478 18058
rect 4530 18006 4582 18058
rect 4634 18006 4686 18058
rect 4738 18006 35198 18058
rect 35250 18006 35302 18058
rect 35354 18006 35406 18058
rect 35458 18006 65918 18058
rect 65970 18006 66022 18058
rect 66074 18006 66126 18058
rect 66178 18006 78624 18058
rect 1344 17972 78624 18006
rect 33854 17890 33906 17902
rect 33854 17826 33906 17838
rect 37998 17890 38050 17902
rect 37998 17826 38050 17838
rect 20638 17778 20690 17790
rect 20638 17714 20690 17726
rect 21422 17778 21474 17790
rect 21422 17714 21474 17726
rect 22430 17778 22482 17790
rect 22430 17714 22482 17726
rect 28590 17778 28642 17790
rect 28590 17714 28642 17726
rect 33406 17778 33458 17790
rect 33406 17714 33458 17726
rect 33742 17778 33794 17790
rect 33742 17714 33794 17726
rect 34750 17778 34802 17790
rect 34750 17714 34802 17726
rect 35310 17778 35362 17790
rect 50206 17778 50258 17790
rect 52110 17778 52162 17790
rect 46050 17726 46062 17778
rect 46114 17726 46126 17778
rect 50754 17726 50766 17778
rect 50818 17726 50830 17778
rect 35310 17714 35362 17726
rect 50206 17714 50258 17726
rect 52110 17714 52162 17726
rect 19070 17666 19122 17678
rect 19070 17602 19122 17614
rect 19406 17666 19458 17678
rect 20526 17666 20578 17678
rect 20178 17614 20190 17666
rect 20242 17614 20254 17666
rect 19406 17602 19458 17614
rect 20526 17602 20578 17614
rect 20750 17666 20802 17678
rect 22318 17666 22370 17678
rect 30718 17666 30770 17678
rect 21970 17614 21982 17666
rect 22034 17614 22046 17666
rect 28130 17614 28142 17666
rect 28194 17614 28206 17666
rect 20750 17602 20802 17614
rect 22318 17602 22370 17614
rect 30718 17602 30770 17614
rect 31166 17666 31218 17678
rect 31166 17602 31218 17614
rect 31390 17666 31442 17678
rect 31390 17602 31442 17614
rect 35086 17666 35138 17678
rect 35086 17602 35138 17614
rect 35534 17666 35586 17678
rect 35534 17602 35586 17614
rect 35758 17666 35810 17678
rect 35758 17602 35810 17614
rect 36430 17666 36482 17678
rect 36430 17602 36482 17614
rect 37886 17666 37938 17678
rect 37886 17602 37938 17614
rect 39006 17666 39058 17678
rect 39006 17602 39058 17614
rect 39790 17666 39842 17678
rect 39790 17602 39842 17614
rect 40574 17666 40626 17678
rect 42926 17666 42978 17678
rect 56590 17666 56642 17678
rect 41682 17614 41694 17666
rect 41746 17614 41758 17666
rect 43138 17614 43150 17666
rect 43202 17614 43214 17666
rect 45266 17614 45278 17666
rect 45330 17614 45342 17666
rect 45938 17614 45950 17666
rect 46002 17614 46014 17666
rect 47282 17614 47294 17666
rect 47346 17614 47358 17666
rect 48738 17614 48750 17666
rect 48802 17614 48814 17666
rect 50978 17614 50990 17666
rect 51042 17614 51054 17666
rect 51650 17614 51662 17666
rect 51714 17614 51726 17666
rect 53218 17614 53230 17666
rect 53282 17614 53294 17666
rect 54786 17614 54798 17666
rect 54850 17614 54862 17666
rect 55682 17614 55694 17666
rect 55746 17614 55758 17666
rect 56802 17614 56814 17666
rect 56866 17614 56878 17666
rect 58706 17614 58718 17666
rect 58770 17614 58782 17666
rect 40574 17602 40626 17614
rect 42926 17602 42978 17614
rect 56590 17602 56642 17614
rect 1710 17554 1762 17566
rect 1710 17490 1762 17502
rect 18734 17554 18786 17566
rect 18734 17490 18786 17502
rect 22542 17554 22594 17566
rect 31278 17554 31330 17566
rect 25106 17502 25118 17554
rect 25170 17502 25182 17554
rect 22542 17490 22594 17502
rect 31278 17490 31330 17502
rect 34190 17554 34242 17566
rect 34190 17490 34242 17502
rect 34302 17554 34354 17566
rect 34302 17490 34354 17502
rect 34638 17554 34690 17566
rect 34638 17490 34690 17502
rect 36990 17554 37042 17566
rect 36990 17490 37042 17502
rect 37326 17554 37378 17566
rect 37326 17490 37378 17502
rect 37550 17554 37602 17566
rect 37550 17490 37602 17502
rect 38446 17554 38498 17566
rect 38446 17490 38498 17502
rect 38782 17554 38834 17566
rect 38782 17490 38834 17502
rect 39342 17554 39394 17566
rect 39342 17490 39394 17502
rect 39678 17554 39730 17566
rect 39678 17490 39730 17502
rect 40238 17554 40290 17566
rect 77646 17554 77698 17566
rect 41458 17502 41470 17554
rect 41522 17502 41534 17554
rect 46162 17502 46174 17554
rect 46226 17502 46238 17554
rect 46946 17502 46958 17554
rect 47010 17502 47022 17554
rect 48850 17502 48862 17554
rect 48914 17502 48926 17554
rect 50866 17502 50878 17554
rect 50930 17502 50942 17554
rect 53442 17502 53454 17554
rect 53506 17502 53518 17554
rect 58818 17502 58830 17554
rect 58882 17502 58894 17554
rect 70802 17502 70814 17554
rect 70866 17502 70878 17554
rect 40238 17490 40290 17502
rect 77646 17490 77698 17502
rect 77870 17554 77922 17566
rect 77870 17490 77922 17502
rect 78206 17554 78258 17566
rect 78206 17490 78258 17502
rect 2046 17442 2098 17454
rect 2046 17378 2098 17390
rect 2494 17442 2546 17454
rect 2494 17378 2546 17390
rect 19182 17442 19234 17454
rect 19182 17378 19234 17390
rect 29262 17442 29314 17454
rect 29262 17378 29314 17390
rect 32734 17442 32786 17454
rect 37214 17442 37266 17454
rect 36082 17390 36094 17442
rect 36146 17390 36158 17442
rect 32734 17378 32786 17390
rect 37214 17378 37266 17390
rect 38558 17442 38610 17454
rect 38558 17378 38610 17390
rect 39566 17442 39618 17454
rect 39566 17378 39618 17390
rect 40350 17442 40402 17454
rect 70254 17442 70306 17454
rect 43026 17390 43038 17442
rect 43090 17390 43102 17442
rect 48402 17390 48414 17442
rect 48466 17390 48478 17442
rect 55010 17390 55022 17442
rect 55074 17390 55086 17442
rect 58370 17390 58382 17442
rect 58434 17390 58446 17442
rect 40350 17378 40402 17390
rect 70254 17378 70306 17390
rect 70478 17442 70530 17454
rect 70478 17378 70530 17390
rect 1344 17274 78624 17308
rect 1344 17222 19838 17274
rect 19890 17222 19942 17274
rect 19994 17222 20046 17274
rect 20098 17222 50558 17274
rect 50610 17222 50662 17274
rect 50714 17222 50766 17274
rect 50818 17222 78624 17274
rect 1344 17188 78624 17222
rect 22766 17106 22818 17118
rect 22766 17042 22818 17054
rect 33406 17106 33458 17118
rect 33406 17042 33458 17054
rect 35422 17106 35474 17118
rect 35422 17042 35474 17054
rect 35982 17106 36034 17118
rect 35982 17042 36034 17054
rect 37774 17106 37826 17118
rect 37774 17042 37826 17054
rect 38670 17106 38722 17118
rect 38670 17042 38722 17054
rect 39454 17106 39506 17118
rect 39454 17042 39506 17054
rect 40462 17106 40514 17118
rect 40462 17042 40514 17054
rect 41694 17106 41746 17118
rect 41694 17042 41746 17054
rect 42030 17106 42082 17118
rect 42030 17042 42082 17054
rect 42254 17106 42306 17118
rect 42254 17042 42306 17054
rect 43934 17106 43986 17118
rect 56814 17106 56866 17118
rect 50418 17054 50430 17106
rect 50482 17054 50494 17106
rect 53442 17054 53454 17106
rect 53506 17054 53518 17106
rect 43934 17042 43986 17054
rect 56814 17042 56866 17054
rect 57150 17106 57202 17118
rect 57150 17042 57202 17054
rect 77870 17106 77922 17118
rect 77870 17042 77922 17054
rect 36094 16994 36146 17006
rect 32274 16942 32286 16994
rect 32338 16942 32350 16994
rect 36094 16930 36146 16942
rect 36990 16994 37042 17006
rect 36990 16930 37042 16942
rect 37326 16994 37378 17006
rect 37326 16930 37378 16942
rect 38782 16994 38834 17006
rect 38782 16930 38834 16942
rect 39678 16994 39730 17006
rect 39678 16930 39730 16942
rect 41134 16994 41186 17006
rect 41134 16930 41186 16942
rect 41358 16994 41410 17006
rect 41358 16930 41410 16942
rect 41470 16994 41522 17006
rect 45278 16994 45330 17006
rect 42578 16942 42590 16994
rect 42642 16942 42654 16994
rect 47506 16942 47518 16994
rect 47570 16942 47582 16994
rect 49074 16942 49086 16994
rect 49138 16942 49150 16994
rect 51090 16942 51102 16994
rect 51154 16942 51166 16994
rect 52322 16942 52334 16994
rect 52386 16942 52398 16994
rect 54562 16942 54574 16994
rect 54626 16942 54638 16994
rect 41470 16930 41522 16942
rect 45278 16930 45330 16942
rect 33854 16882 33906 16894
rect 25330 16830 25342 16882
rect 25394 16830 25406 16882
rect 28690 16830 28702 16882
rect 28754 16830 28766 16882
rect 29474 16830 29486 16882
rect 29538 16830 29550 16882
rect 33854 16818 33906 16830
rect 34302 16882 34354 16894
rect 34302 16818 34354 16830
rect 35646 16882 35698 16894
rect 35646 16818 35698 16830
rect 36206 16882 36258 16894
rect 36206 16818 36258 16830
rect 37662 16882 37714 16894
rect 37662 16818 37714 16830
rect 38222 16882 38274 16894
rect 38222 16818 38274 16830
rect 39230 16882 39282 16894
rect 39230 16818 39282 16830
rect 39790 16882 39842 16894
rect 39790 16818 39842 16830
rect 41918 16882 41970 16894
rect 41918 16818 41970 16830
rect 42702 16882 42754 16894
rect 56030 16882 56082 16894
rect 46386 16830 46398 16882
rect 46450 16830 46462 16882
rect 46722 16830 46734 16882
rect 46786 16830 46798 16882
rect 47282 16830 47294 16882
rect 47346 16830 47358 16882
rect 49298 16830 49310 16882
rect 49362 16830 49374 16882
rect 51426 16830 51438 16882
rect 51490 16830 51502 16882
rect 52546 16830 52558 16882
rect 52610 16830 52622 16882
rect 54674 16830 54686 16882
rect 54738 16830 54750 16882
rect 42702 16818 42754 16830
rect 56030 16818 56082 16830
rect 77646 16882 77698 16894
rect 77646 16818 77698 16830
rect 78206 16882 78258 16894
rect 78206 16818 78258 16830
rect 31950 16770 32002 16782
rect 26114 16718 26126 16770
rect 26178 16718 26190 16770
rect 28242 16718 28254 16770
rect 28306 16718 28318 16770
rect 31602 16718 31614 16770
rect 31666 16718 31678 16770
rect 47730 16718 47742 16770
rect 47794 16718 47806 16770
rect 31950 16706 32002 16718
rect 38334 16658 38386 16670
rect 38334 16594 38386 16606
rect 1344 16490 78624 16524
rect 1344 16438 4478 16490
rect 4530 16438 4582 16490
rect 4634 16438 4686 16490
rect 4738 16438 35198 16490
rect 35250 16438 35302 16490
rect 35354 16438 35406 16490
rect 35458 16438 65918 16490
rect 65970 16438 66022 16490
rect 66074 16438 66126 16490
rect 66178 16438 78624 16490
rect 1344 16404 78624 16438
rect 37438 16322 37490 16334
rect 37986 16270 37998 16322
rect 38050 16319 38062 16322
rect 38322 16319 38334 16322
rect 38050 16273 38334 16319
rect 38050 16270 38062 16273
rect 38322 16270 38334 16273
rect 38386 16270 38398 16322
rect 37438 16258 37490 16270
rect 25566 16210 25618 16222
rect 25566 16146 25618 16158
rect 26686 16210 26738 16222
rect 26686 16146 26738 16158
rect 28142 16210 28194 16222
rect 35646 16210 35698 16222
rect 32050 16158 32062 16210
rect 32114 16158 32126 16210
rect 35298 16158 35310 16210
rect 35362 16158 35374 16210
rect 28142 16146 28194 16158
rect 35646 16146 35698 16158
rect 36542 16210 36594 16222
rect 36542 16146 36594 16158
rect 37326 16210 37378 16222
rect 37326 16146 37378 16158
rect 37886 16210 37938 16222
rect 37886 16146 37938 16158
rect 38334 16210 38386 16222
rect 38334 16146 38386 16158
rect 38782 16210 38834 16222
rect 38782 16146 38834 16158
rect 40686 16210 40738 16222
rect 40686 16146 40738 16158
rect 41134 16210 41186 16222
rect 41134 16146 41186 16158
rect 41582 16210 41634 16222
rect 41582 16146 41634 16158
rect 43934 16210 43986 16222
rect 43934 16146 43986 16158
rect 45054 16210 45106 16222
rect 45054 16146 45106 16158
rect 45502 16210 45554 16222
rect 45502 16146 45554 16158
rect 45838 16210 45890 16222
rect 52110 16210 52162 16222
rect 51090 16158 51102 16210
rect 51154 16158 51166 16210
rect 45838 16146 45890 16158
rect 52110 16146 52162 16158
rect 26574 16098 26626 16110
rect 26574 16034 26626 16046
rect 28254 16098 28306 16110
rect 28254 16034 28306 16046
rect 28702 16098 28754 16110
rect 39230 16098 39282 16110
rect 29138 16046 29150 16098
rect 29202 16046 29214 16098
rect 32498 16046 32510 16098
rect 32562 16046 32574 16098
rect 28702 16034 28754 16046
rect 39230 16034 39282 16046
rect 39678 16098 39730 16110
rect 39678 16034 39730 16046
rect 39790 16098 39842 16110
rect 39790 16034 39842 16046
rect 43374 16098 43426 16110
rect 43374 16034 43426 16046
rect 43710 16098 43762 16110
rect 43710 16034 43762 16046
rect 46174 16098 46226 16110
rect 52670 16098 52722 16110
rect 54574 16098 54626 16110
rect 47842 16046 47854 16098
rect 47906 16046 47918 16098
rect 48962 16046 48974 16098
rect 49026 16046 49038 16098
rect 53666 16046 53678 16098
rect 53730 16046 53742 16098
rect 54786 16046 54798 16098
rect 54850 16046 54862 16098
rect 46174 16034 46226 16046
rect 52670 16034 52722 16046
rect 54574 16034 54626 16046
rect 1710 15986 1762 15998
rect 1710 15922 1762 15934
rect 2046 15986 2098 15998
rect 41918 15986 41970 15998
rect 29922 15934 29934 15986
rect 29986 15934 29998 15986
rect 33170 15934 33182 15986
rect 33234 15934 33246 15986
rect 35970 15934 35982 15986
rect 36034 15934 36046 15986
rect 2046 15922 2098 15934
rect 41918 15922 41970 15934
rect 42478 15986 42530 15998
rect 42478 15922 42530 15934
rect 43486 15986 43538 15998
rect 77870 15986 77922 15998
rect 47170 15934 47182 15986
rect 47234 15934 47246 15986
rect 49410 15934 49422 15986
rect 49474 15934 49486 15986
rect 43486 15922 43538 15934
rect 77870 15922 77922 15934
rect 78206 15986 78258 15998
rect 78206 15922 78258 15934
rect 2494 15874 2546 15886
rect 2494 15810 2546 15822
rect 26014 15874 26066 15886
rect 26014 15810 26066 15822
rect 26350 15874 26402 15886
rect 26350 15810 26402 15822
rect 26798 15874 26850 15886
rect 26798 15810 26850 15822
rect 27246 15874 27298 15886
rect 27246 15810 27298 15822
rect 27470 15874 27522 15886
rect 27470 15810 27522 15822
rect 27582 15874 27634 15886
rect 27582 15810 27634 15822
rect 27694 15874 27746 15886
rect 27694 15810 27746 15822
rect 28030 15874 28082 15886
rect 28030 15810 28082 15822
rect 39566 15874 39618 15886
rect 39566 15810 39618 15822
rect 41806 15874 41858 15886
rect 41806 15810 41858 15822
rect 42814 15874 42866 15886
rect 42814 15810 42866 15822
rect 44046 15874 44098 15886
rect 50430 15874 50482 15886
rect 46498 15822 46510 15874
rect 46562 15822 46574 15874
rect 47954 15822 47966 15874
rect 48018 15822 48030 15874
rect 44046 15810 44098 15822
rect 50430 15810 50482 15822
rect 51662 15874 51714 15886
rect 77646 15874 77698 15886
rect 53778 15822 53790 15874
rect 53842 15822 53854 15874
rect 51662 15810 51714 15822
rect 77646 15810 77698 15822
rect 1344 15706 78624 15740
rect 1344 15654 19838 15706
rect 19890 15654 19942 15706
rect 19994 15654 20046 15706
rect 20098 15654 50558 15706
rect 50610 15654 50662 15706
rect 50714 15654 50766 15706
rect 50818 15654 78624 15706
rect 1344 15620 78624 15654
rect 33406 15538 33458 15550
rect 33406 15474 33458 15486
rect 33518 15538 33570 15550
rect 33518 15474 33570 15486
rect 38558 15538 38610 15550
rect 38558 15474 38610 15486
rect 41134 15538 41186 15550
rect 41134 15474 41186 15486
rect 41582 15538 41634 15550
rect 41582 15474 41634 15486
rect 46174 15538 46226 15550
rect 46174 15474 46226 15486
rect 46622 15538 46674 15550
rect 46622 15474 46674 15486
rect 47182 15538 47234 15550
rect 47182 15474 47234 15486
rect 47966 15538 48018 15550
rect 53442 15486 53454 15538
rect 53506 15486 53518 15538
rect 47966 15474 48018 15486
rect 2046 15426 2098 15438
rect 31950 15426 32002 15438
rect 27906 15374 27918 15426
rect 27970 15374 27982 15426
rect 31602 15374 31614 15426
rect 31666 15374 31678 15426
rect 39218 15374 39230 15426
rect 39282 15374 39294 15426
rect 48738 15374 48750 15426
rect 48802 15374 48814 15426
rect 50642 15374 50654 15426
rect 50706 15374 50718 15426
rect 52770 15374 52782 15426
rect 52834 15374 52846 15426
rect 54562 15374 54574 15426
rect 54626 15374 54638 15426
rect 2046 15362 2098 15374
rect 31950 15362 32002 15374
rect 1710 15314 1762 15326
rect 32958 15314 33010 15326
rect 31042 15262 31054 15314
rect 31106 15262 31118 15314
rect 1710 15250 1762 15262
rect 32958 15250 33010 15262
rect 33630 15314 33682 15326
rect 39454 15314 39506 15326
rect 35074 15262 35086 15314
rect 35138 15262 35150 15314
rect 33630 15250 33682 15262
rect 39454 15250 39506 15262
rect 39902 15314 39954 15326
rect 39902 15250 39954 15262
rect 40126 15314 40178 15326
rect 45390 15314 45442 15326
rect 42130 15262 42142 15314
rect 42194 15262 42206 15314
rect 40126 15250 40178 15262
rect 45390 15250 45442 15262
rect 45502 15314 45554 15326
rect 49746 15262 49758 15314
rect 49810 15262 49822 15314
rect 50866 15262 50878 15314
rect 50930 15262 50942 15314
rect 52546 15262 52558 15314
rect 52610 15262 52622 15314
rect 54450 15262 54462 15314
rect 54514 15262 54526 15314
rect 45502 15250 45554 15262
rect 2494 15202 2546 15214
rect 38446 15202 38498 15214
rect 35858 15150 35870 15202
rect 35922 15150 35934 15202
rect 37986 15150 37998 15202
rect 38050 15150 38062 15202
rect 2494 15138 2546 15150
rect 38446 15138 38498 15150
rect 38894 15202 38946 15214
rect 38894 15138 38946 15150
rect 40014 15202 40066 15214
rect 51662 15202 51714 15214
rect 42914 15150 42926 15202
rect 42978 15150 42990 15202
rect 45042 15150 45054 15202
rect 45106 15150 45118 15202
rect 40014 15138 40066 15150
rect 51662 15138 51714 15150
rect 1344 14922 78624 14956
rect 1344 14870 4478 14922
rect 4530 14870 4582 14922
rect 4634 14870 4686 14922
rect 4738 14870 35198 14922
rect 35250 14870 35302 14922
rect 35354 14870 35406 14922
rect 35458 14870 65918 14922
rect 65970 14870 66022 14922
rect 66074 14870 66126 14922
rect 66178 14870 78624 14922
rect 1344 14836 78624 14870
rect 52110 14754 52162 14766
rect 30818 14702 30830 14754
rect 30882 14751 30894 14754
rect 31490 14751 31502 14754
rect 30882 14705 31502 14751
rect 30882 14702 30894 14705
rect 31490 14702 31502 14705
rect 31554 14702 31566 14754
rect 52110 14690 52162 14702
rect 29598 14642 29650 14654
rect 25666 14590 25678 14642
rect 25730 14590 25742 14642
rect 27794 14590 27806 14642
rect 27858 14590 27870 14642
rect 28466 14590 28478 14642
rect 28530 14590 28542 14642
rect 29598 14578 29650 14590
rect 30830 14642 30882 14654
rect 35198 14642 35250 14654
rect 34626 14590 34638 14642
rect 34690 14590 34702 14642
rect 30830 14578 30882 14590
rect 35198 14578 35250 14590
rect 35870 14642 35922 14654
rect 35870 14578 35922 14590
rect 37214 14642 37266 14654
rect 37214 14578 37266 14590
rect 38334 14642 38386 14654
rect 38334 14578 38386 14590
rect 38670 14642 38722 14654
rect 42814 14642 42866 14654
rect 39778 14590 39790 14642
rect 39842 14590 39854 14642
rect 41906 14590 41918 14642
rect 41970 14590 41982 14642
rect 38670 14578 38722 14590
rect 42814 14578 42866 14590
rect 43374 14642 43426 14654
rect 43374 14578 43426 14590
rect 43934 14642 43986 14654
rect 43934 14578 43986 14590
rect 44270 14642 44322 14654
rect 44270 14578 44322 14590
rect 46286 14642 46338 14654
rect 46286 14578 46338 14590
rect 51102 14642 51154 14654
rect 53106 14590 53118 14642
rect 53170 14590 53182 14642
rect 51102 14578 51154 14590
rect 19966 14530 20018 14542
rect 29038 14530 29090 14542
rect 24882 14478 24894 14530
rect 24946 14478 24958 14530
rect 28242 14478 28254 14530
rect 28306 14478 28318 14530
rect 19966 14466 20018 14478
rect 29038 14466 29090 14478
rect 29486 14530 29538 14542
rect 29486 14466 29538 14478
rect 29710 14530 29762 14542
rect 35758 14530 35810 14542
rect 42702 14530 42754 14542
rect 31826 14478 31838 14530
rect 31890 14478 31902 14530
rect 38994 14478 39006 14530
rect 39058 14478 39070 14530
rect 29710 14466 29762 14478
rect 35758 14466 35810 14478
rect 42702 14466 42754 14478
rect 46510 14530 46562 14542
rect 51326 14530 51378 14542
rect 47730 14478 47742 14530
rect 47794 14478 47806 14530
rect 48738 14478 48750 14530
rect 48802 14478 48814 14530
rect 46510 14466 46562 14478
rect 51326 14466 51378 14478
rect 52670 14530 52722 14542
rect 52670 14466 52722 14478
rect 19854 14418 19906 14430
rect 43262 14418 43314 14430
rect 77870 14418 77922 14430
rect 30034 14366 30046 14418
rect 30098 14366 30110 14418
rect 32498 14366 32510 14418
rect 32562 14366 32574 14418
rect 48962 14366 48974 14418
rect 49026 14366 49038 14418
rect 19854 14354 19906 14366
rect 43262 14354 43314 14366
rect 77870 14354 77922 14366
rect 78206 14418 78258 14430
rect 78206 14354 78258 14366
rect 20078 14306 20130 14318
rect 20078 14242 20130 14254
rect 20302 14306 20354 14318
rect 20302 14242 20354 14254
rect 21422 14306 21474 14318
rect 21422 14242 21474 14254
rect 30382 14306 30434 14318
rect 30382 14242 30434 14254
rect 31278 14306 31330 14318
rect 31278 14242 31330 14254
rect 35534 14306 35586 14318
rect 35534 14242 35586 14254
rect 35982 14306 36034 14318
rect 35982 14242 36034 14254
rect 42478 14306 42530 14318
rect 42478 14242 42530 14254
rect 42926 14306 42978 14318
rect 77646 14306 77698 14318
rect 48178 14254 48190 14306
rect 48242 14254 48254 14306
rect 42926 14242 42978 14254
rect 77646 14242 77698 14254
rect 1344 14138 78624 14172
rect 1344 14086 19838 14138
rect 19890 14086 19942 14138
rect 19994 14086 20046 14138
rect 20098 14086 50558 14138
rect 50610 14086 50662 14138
rect 50714 14086 50766 14138
rect 50818 14086 78624 14138
rect 1344 14052 78624 14086
rect 2046 13970 2098 13982
rect 2046 13906 2098 13918
rect 19182 13970 19234 13982
rect 26238 13970 26290 13982
rect 22866 13918 22878 13970
rect 22930 13918 22942 13970
rect 19182 13906 19234 13918
rect 26238 13906 26290 13918
rect 27246 13970 27298 13982
rect 27246 13906 27298 13918
rect 28814 13970 28866 13982
rect 28814 13906 28866 13918
rect 29598 13970 29650 13982
rect 29598 13906 29650 13918
rect 30942 13970 30994 13982
rect 30942 13906 30994 13918
rect 33406 13970 33458 13982
rect 33406 13906 33458 13918
rect 33518 13970 33570 13982
rect 33518 13906 33570 13918
rect 33630 13970 33682 13982
rect 33630 13906 33682 13918
rect 34078 13970 34130 13982
rect 38558 13970 38610 13982
rect 39342 13970 39394 13982
rect 35298 13918 35310 13970
rect 35362 13918 35374 13970
rect 39106 13918 39118 13970
rect 39170 13918 39182 13970
rect 34078 13906 34130 13918
rect 38558 13906 38610 13918
rect 39342 13906 39394 13918
rect 41246 13970 41298 13982
rect 41246 13906 41298 13918
rect 41470 13970 41522 13982
rect 41470 13906 41522 13918
rect 45390 13970 45442 13982
rect 45390 13906 45442 13918
rect 48078 13970 48130 13982
rect 48078 13906 48130 13918
rect 48862 13970 48914 13982
rect 55134 13970 55186 13982
rect 52658 13918 52670 13970
rect 52722 13918 52734 13970
rect 48862 13906 48914 13918
rect 55134 13906 55186 13918
rect 77870 13970 77922 13982
rect 77870 13906 77922 13918
rect 18622 13858 18674 13870
rect 18622 13794 18674 13806
rect 26462 13858 26514 13870
rect 26462 13794 26514 13806
rect 26574 13858 26626 13870
rect 26574 13794 26626 13806
rect 27022 13858 27074 13870
rect 28478 13858 28530 13870
rect 28018 13806 28030 13858
rect 28082 13806 28094 13858
rect 27022 13794 27074 13806
rect 28478 13794 28530 13806
rect 28590 13858 28642 13870
rect 29822 13858 29874 13870
rect 29026 13806 29038 13858
rect 29090 13806 29102 13858
rect 28590 13794 28642 13806
rect 29822 13794 29874 13806
rect 29934 13858 29986 13870
rect 29934 13794 29986 13806
rect 31166 13858 31218 13870
rect 31166 13794 31218 13806
rect 31726 13858 31778 13870
rect 31726 13794 31778 13806
rect 32286 13858 32338 13870
rect 32286 13794 32338 13806
rect 34638 13858 34690 13870
rect 37774 13858 37826 13870
rect 34962 13806 34974 13858
rect 35026 13806 35038 13858
rect 34638 13794 34690 13806
rect 37774 13794 37826 13806
rect 38222 13858 38274 13870
rect 38222 13794 38274 13806
rect 38334 13858 38386 13870
rect 38334 13794 38386 13806
rect 38782 13858 38834 13870
rect 38782 13794 38834 13806
rect 39566 13858 39618 13870
rect 54226 13806 54238 13858
rect 54290 13806 54302 13858
rect 39566 13794 39618 13806
rect 1710 13746 1762 13758
rect 1710 13682 1762 13694
rect 18958 13746 19010 13758
rect 26910 13746 26962 13758
rect 29374 13746 29426 13758
rect 19506 13694 19518 13746
rect 19570 13694 19582 13746
rect 19842 13694 19854 13746
rect 19906 13694 19918 13746
rect 27794 13694 27806 13746
rect 27858 13694 27870 13746
rect 18958 13682 19010 13694
rect 26910 13682 26962 13694
rect 29374 13682 29426 13694
rect 31278 13746 31330 13758
rect 31278 13682 31330 13694
rect 31614 13746 31666 13758
rect 31614 13682 31666 13694
rect 31950 13746 32002 13758
rect 31950 13682 32002 13694
rect 32174 13746 32226 13758
rect 32174 13682 32226 13694
rect 32958 13746 33010 13758
rect 32958 13682 33010 13694
rect 35646 13746 35698 13758
rect 35646 13682 35698 13694
rect 37662 13746 37714 13758
rect 37662 13682 37714 13694
rect 37998 13746 38050 13758
rect 37998 13682 38050 13694
rect 39678 13746 39730 13758
rect 39678 13682 39730 13694
rect 40798 13746 40850 13758
rect 45278 13746 45330 13758
rect 78206 13746 78258 13758
rect 42130 13694 42142 13746
rect 42194 13694 42206 13746
rect 52210 13694 52222 13746
rect 52274 13694 52286 13746
rect 52882 13694 52894 13746
rect 52946 13694 52958 13746
rect 53890 13694 53902 13746
rect 53954 13694 53966 13746
rect 40798 13682 40850 13694
rect 45278 13682 45330 13694
rect 78206 13682 78258 13694
rect 2494 13634 2546 13646
rect 2494 13570 2546 13582
rect 19070 13634 19122 13646
rect 41358 13634 41410 13646
rect 46622 13634 46674 13646
rect 20626 13582 20638 13634
rect 20690 13582 20702 13634
rect 42802 13582 42814 13634
rect 42866 13582 42878 13634
rect 44930 13582 44942 13634
rect 44994 13582 45006 13634
rect 19070 13570 19122 13582
rect 41358 13570 41410 13582
rect 46622 13570 46674 13582
rect 77646 13634 77698 13646
rect 77646 13570 77698 13582
rect 32286 13522 32338 13534
rect 32286 13458 32338 13470
rect 1344 13354 78624 13388
rect 1344 13302 4478 13354
rect 4530 13302 4582 13354
rect 4634 13302 4686 13354
rect 4738 13302 35198 13354
rect 35250 13302 35302 13354
rect 35354 13302 35406 13354
rect 35458 13302 65918 13354
rect 65970 13302 66022 13354
rect 66074 13302 66126 13354
rect 66178 13302 78624 13354
rect 1344 13268 78624 13302
rect 20078 13186 20130 13198
rect 20078 13122 20130 13134
rect 20414 13186 20466 13198
rect 20414 13122 20466 13134
rect 12462 13074 12514 13086
rect 12462 13010 12514 13022
rect 19518 13074 19570 13086
rect 37774 13074 37826 13086
rect 43150 13074 43202 13086
rect 25442 13022 25454 13074
rect 25506 13022 25518 13074
rect 36418 13022 36430 13074
rect 36482 13022 36494 13074
rect 40226 13022 40238 13074
rect 40290 13022 40302 13074
rect 42354 13022 42366 13074
rect 42418 13022 42430 13074
rect 19518 13010 19570 13022
rect 37774 13010 37826 13022
rect 43150 13010 43202 13022
rect 74510 13074 74562 13086
rect 74510 13010 74562 13022
rect 74734 13074 74786 13086
rect 74734 13010 74786 13022
rect 74958 13074 75010 13086
rect 74958 13010 75010 13022
rect 76302 13074 76354 13086
rect 76302 13010 76354 13022
rect 32174 12962 32226 12974
rect 38446 12962 38498 12974
rect 42590 12962 42642 12974
rect 16594 12910 16606 12962
rect 16658 12910 16670 12962
rect 22530 12910 22542 12962
rect 22594 12910 22606 12962
rect 28354 12910 28366 12962
rect 28418 12910 28430 12962
rect 31602 12910 31614 12962
rect 31666 12910 31678 12962
rect 33618 12910 33630 12962
rect 33682 12910 33694 12962
rect 39554 12910 39566 12962
rect 39618 12910 39630 12962
rect 32174 12898 32226 12910
rect 38446 12898 38498 12910
rect 42590 12898 42642 12910
rect 43038 12962 43090 12974
rect 43038 12898 43090 12910
rect 43262 12962 43314 12974
rect 43262 12898 43314 12910
rect 1710 12850 1762 12862
rect 1710 12786 1762 12798
rect 2046 12850 2098 12862
rect 29486 12850 29538 12862
rect 17378 12798 17390 12850
rect 17442 12798 17454 12850
rect 23314 12798 23326 12850
rect 23378 12798 23390 12850
rect 31826 12798 31838 12850
rect 31890 12798 31902 12850
rect 34290 12798 34302 12850
rect 34354 12798 34366 12850
rect 37426 12798 37438 12850
rect 37490 12798 37502 12850
rect 2046 12786 2098 12798
rect 29486 12786 29538 12798
rect 2494 12738 2546 12750
rect 2494 12674 2546 12686
rect 20302 12738 20354 12750
rect 20302 12674 20354 12686
rect 28590 12738 28642 12750
rect 28590 12674 28642 12686
rect 29822 12738 29874 12750
rect 29822 12674 29874 12686
rect 32286 12738 32338 12750
rect 32286 12674 32338 12686
rect 32510 12738 32562 12750
rect 32510 12674 32562 12686
rect 37102 12738 37154 12750
rect 37102 12674 37154 12686
rect 37886 12738 37938 12750
rect 38770 12686 38782 12738
rect 38834 12686 38846 12738
rect 75282 12686 75294 12738
rect 75346 12686 75358 12738
rect 37886 12674 37938 12686
rect 1344 12570 78624 12604
rect 1344 12518 19838 12570
rect 19890 12518 19942 12570
rect 19994 12518 20046 12570
rect 20098 12518 50558 12570
rect 50610 12518 50662 12570
rect 50714 12518 50766 12570
rect 50818 12518 78624 12570
rect 1344 12484 78624 12518
rect 11902 12402 11954 12414
rect 18510 12402 18562 12414
rect 15586 12350 15598 12402
rect 15650 12350 15662 12402
rect 17378 12350 17390 12402
rect 17442 12350 17454 12402
rect 11902 12338 11954 12350
rect 17393 12287 17439 12350
rect 18510 12338 18562 12350
rect 25454 12402 25506 12414
rect 25454 12338 25506 12350
rect 35086 12402 35138 12414
rect 35086 12338 35138 12350
rect 35198 12402 35250 12414
rect 35198 12338 35250 12350
rect 35310 12402 35362 12414
rect 35310 12338 35362 12350
rect 35758 12402 35810 12414
rect 35758 12338 35810 12350
rect 41246 12402 41298 12414
rect 41246 12338 41298 12350
rect 41582 12402 41634 12414
rect 41582 12338 41634 12350
rect 17838 12290 17890 12302
rect 17602 12287 17614 12290
rect 17393 12241 17614 12287
rect 17602 12238 17614 12241
rect 17666 12238 17678 12290
rect 17838 12226 17890 12238
rect 18062 12290 18114 12302
rect 18062 12226 18114 12238
rect 25678 12290 25730 12302
rect 25678 12226 25730 12238
rect 26462 12290 26514 12302
rect 26462 12226 26514 12238
rect 35646 12290 35698 12302
rect 35646 12226 35698 12238
rect 36206 12290 36258 12302
rect 36206 12226 36258 12238
rect 40910 12290 40962 12302
rect 40910 12226 40962 12238
rect 41022 12290 41074 12302
rect 77522 12238 77534 12290
rect 77586 12238 77598 12290
rect 41022 12226 41074 12238
rect 11678 12178 11730 12190
rect 9538 12126 9550 12178
rect 9602 12126 9614 12178
rect 11678 12114 11730 12126
rect 12350 12178 12402 12190
rect 25230 12178 25282 12190
rect 34638 12178 34690 12190
rect 12674 12126 12686 12178
rect 12738 12126 12750 12178
rect 21858 12126 21870 12178
rect 21922 12126 21934 12178
rect 29698 12126 29710 12178
rect 29762 12126 29774 12178
rect 37538 12126 37550 12178
rect 37602 12126 37614 12178
rect 77746 12126 77758 12178
rect 77810 12126 77822 12178
rect 12350 12114 12402 12126
rect 25230 12114 25282 12126
rect 34638 12114 34690 12126
rect 9774 12066 9826 12078
rect 9774 12002 9826 12014
rect 9886 12066 9938 12078
rect 9886 12002 9938 12014
rect 11790 12066 11842 12078
rect 25342 12066 25394 12078
rect 37214 12066 37266 12078
rect 13346 12014 13358 12066
rect 13410 12014 13422 12066
rect 17714 12014 17726 12066
rect 17778 12014 17790 12066
rect 22530 12014 22542 12066
rect 22594 12014 22606 12066
rect 24658 12014 24670 12066
rect 24722 12014 24734 12066
rect 26450 12014 26462 12066
rect 26514 12014 26526 12066
rect 30370 12014 30382 12066
rect 30434 12014 30446 12066
rect 32498 12014 32510 12066
rect 32562 12014 32574 12066
rect 38210 12014 38222 12066
rect 38274 12014 38286 12066
rect 40338 12014 40350 12066
rect 40402 12014 40414 12066
rect 11790 12002 11842 12014
rect 25342 12002 25394 12014
rect 37214 12002 37266 12014
rect 26238 11954 26290 11966
rect 26238 11890 26290 11902
rect 1344 11786 78624 11820
rect 1344 11734 4478 11786
rect 4530 11734 4582 11786
rect 4634 11734 4686 11786
rect 4738 11734 35198 11786
rect 35250 11734 35302 11786
rect 35354 11734 35406 11786
rect 35458 11734 65918 11786
rect 65970 11734 66022 11786
rect 66074 11734 66126 11786
rect 66178 11734 78624 11786
rect 1344 11700 78624 11734
rect 37774 11618 37826 11630
rect 37774 11554 37826 11566
rect 11902 11506 11954 11518
rect 9762 11454 9774 11506
rect 9826 11454 9838 11506
rect 11902 11442 11954 11454
rect 14478 11506 14530 11518
rect 20750 11506 20802 11518
rect 18274 11454 18286 11506
rect 18338 11454 18350 11506
rect 14478 11442 14530 11454
rect 20750 11442 20802 11454
rect 22542 11506 22594 11518
rect 22542 11442 22594 11454
rect 23214 11506 23266 11518
rect 76526 11506 76578 11518
rect 26450 11454 26462 11506
rect 26514 11454 26526 11506
rect 28578 11454 28590 11506
rect 28642 11454 28654 11506
rect 30146 11454 30158 11506
rect 30210 11454 30222 11506
rect 32386 11454 32398 11506
rect 32450 11503 32462 11506
rect 32610 11503 32622 11506
rect 32450 11457 32622 11503
rect 32450 11454 32462 11457
rect 32610 11454 32622 11457
rect 32674 11454 32686 11506
rect 36418 11454 36430 11506
rect 36482 11454 36494 11506
rect 23214 11442 23266 11454
rect 76526 11442 76578 11454
rect 13694 11394 13746 11406
rect 19406 11394 19458 11406
rect 9090 11342 9102 11394
rect 9154 11342 9166 11394
rect 15362 11342 15374 11394
rect 15426 11342 15438 11394
rect 13694 11330 13746 11342
rect 19406 11330 19458 11342
rect 19854 11394 19906 11406
rect 19854 11330 19906 11342
rect 19966 11394 20018 11406
rect 19966 11330 20018 11342
rect 20414 11394 20466 11406
rect 25006 11394 25058 11406
rect 22306 11342 22318 11394
rect 22370 11342 22382 11394
rect 22978 11342 22990 11394
rect 23042 11342 23054 11394
rect 20414 11330 20466 11342
rect 25006 11330 25058 11342
rect 25454 11394 25506 11406
rect 31950 11394 32002 11406
rect 25778 11342 25790 11394
rect 25842 11342 25854 11394
rect 25454 11330 25506 11342
rect 31950 11330 32002 11342
rect 32398 11394 32450 11406
rect 32958 11394 33010 11406
rect 78206 11394 78258 11406
rect 32610 11342 32622 11394
rect 32674 11342 32686 11394
rect 33618 11342 33630 11394
rect 33682 11342 33694 11394
rect 37090 11342 37102 11394
rect 37154 11342 37166 11394
rect 38658 11342 38670 11394
rect 38722 11342 38734 11394
rect 32398 11330 32450 11342
rect 32958 11330 33010 11342
rect 78206 11330 78258 11342
rect 1710 11282 1762 11294
rect 1710 11218 1762 11230
rect 2494 11282 2546 11294
rect 22654 11282 22706 11294
rect 16034 11230 16046 11282
rect 16098 11230 16110 11282
rect 2494 11218 2546 11230
rect 22654 11218 22706 11230
rect 23326 11282 23378 11294
rect 23326 11218 23378 11230
rect 24894 11282 24946 11294
rect 24894 11218 24946 11230
rect 30382 11282 30434 11294
rect 30382 11218 30434 11230
rect 31838 11282 31890 11294
rect 37662 11282 37714 11294
rect 44830 11282 44882 11294
rect 34290 11230 34302 11282
rect 34354 11230 34366 11282
rect 41346 11230 41358 11282
rect 41410 11230 41422 11282
rect 31838 11218 31890 11230
rect 37662 11218 37714 11230
rect 44830 11218 44882 11230
rect 77198 11282 77250 11294
rect 77198 11218 77250 11230
rect 77534 11282 77586 11294
rect 77534 11218 77586 11230
rect 77870 11282 77922 11294
rect 77870 11218 77922 11230
rect 2046 11170 2098 11182
rect 2046 11106 2098 11118
rect 13470 11170 13522 11182
rect 13470 11106 13522 11118
rect 13582 11170 13634 11182
rect 13582 11106 13634 11118
rect 13918 11170 13970 11182
rect 13918 11106 13970 11118
rect 19182 11170 19234 11182
rect 19182 11106 19234 11118
rect 19294 11170 19346 11182
rect 19294 11106 19346 11118
rect 19742 11170 19794 11182
rect 19742 11106 19794 11118
rect 24782 11170 24834 11182
rect 24782 11106 24834 11118
rect 30158 11170 30210 11182
rect 30158 11106 30210 11118
rect 31726 11170 31778 11182
rect 31726 11106 31778 11118
rect 33070 11170 33122 11182
rect 33070 11106 33122 11118
rect 33182 11170 33234 11182
rect 33182 11106 33234 11118
rect 37326 11170 37378 11182
rect 37326 11106 37378 11118
rect 38334 11170 38386 11182
rect 38334 11106 38386 11118
rect 44942 11170 44994 11182
rect 44942 11106 44994 11118
rect 76974 11170 77026 11182
rect 76974 11106 77026 11118
rect 1344 11002 78624 11036
rect 1344 10950 19838 11002
rect 19890 10950 19942 11002
rect 19994 10950 20046 11002
rect 20098 10950 50558 11002
rect 50610 10950 50662 11002
rect 50714 10950 50766 11002
rect 50818 10950 78624 11002
rect 1344 10916 78624 10950
rect 2046 10834 2098 10846
rect 2046 10770 2098 10782
rect 13246 10834 13298 10846
rect 13246 10770 13298 10782
rect 17950 10834 18002 10846
rect 25230 10834 25282 10846
rect 21634 10782 21646 10834
rect 21698 10782 21710 10834
rect 17950 10770 18002 10782
rect 25230 10770 25282 10782
rect 26462 10834 26514 10846
rect 26462 10770 26514 10782
rect 26574 10834 26626 10846
rect 26574 10770 26626 10782
rect 32510 10834 32562 10846
rect 32510 10770 32562 10782
rect 39342 10834 39394 10846
rect 39342 10770 39394 10782
rect 39454 10834 39506 10846
rect 39454 10770 39506 10782
rect 39566 10834 39618 10846
rect 39566 10770 39618 10782
rect 40238 10834 40290 10846
rect 40238 10770 40290 10782
rect 13134 10722 13186 10734
rect 13134 10658 13186 10670
rect 13358 10722 13410 10734
rect 25678 10722 25730 10734
rect 19394 10670 19406 10722
rect 19458 10670 19470 10722
rect 13358 10658 13410 10670
rect 25678 10658 25730 10670
rect 40350 10722 40402 10734
rect 40350 10658 40402 10670
rect 1710 10610 1762 10622
rect 17726 10610 17778 10622
rect 9538 10558 9550 10610
rect 9602 10558 9614 10610
rect 1710 10546 1762 10558
rect 17726 10546 17778 10558
rect 17838 10610 17890 10622
rect 17838 10546 17890 10558
rect 18398 10610 18450 10622
rect 25454 10610 25506 10622
rect 18722 10558 18734 10610
rect 18786 10558 18798 10610
rect 22642 10558 22654 10610
rect 22706 10558 22718 10610
rect 18398 10546 18450 10558
rect 25454 10546 25506 10558
rect 26014 10610 26066 10622
rect 26014 10546 26066 10558
rect 26686 10610 26738 10622
rect 38894 10610 38946 10622
rect 28466 10558 28478 10610
rect 28530 10558 28542 10610
rect 36978 10558 36990 10610
rect 37042 10558 37054 10610
rect 41346 10558 41358 10610
rect 41410 10558 41422 10610
rect 78194 10558 78206 10610
rect 78258 10558 78270 10610
rect 26686 10546 26738 10558
rect 38894 10546 38946 10558
rect 2494 10498 2546 10510
rect 12462 10498 12514 10510
rect 10322 10446 10334 10498
rect 10386 10446 10398 10498
rect 2494 10434 2546 10446
rect 12462 10434 12514 10446
rect 14142 10498 14194 10510
rect 14142 10434 14194 10446
rect 14478 10498 14530 10510
rect 14478 10434 14530 10446
rect 15150 10498 15202 10510
rect 15150 10434 15202 10446
rect 15598 10498 15650 10510
rect 15598 10434 15650 10446
rect 16046 10498 16098 10510
rect 16046 10434 16098 10446
rect 22878 10498 22930 10510
rect 22878 10434 22930 10446
rect 22990 10498 23042 10510
rect 22990 10434 23042 10446
rect 25342 10498 25394 10510
rect 41022 10498 41074 10510
rect 25778 10446 25790 10498
rect 25842 10495 25854 10498
rect 26002 10495 26014 10498
rect 25842 10449 26014 10495
rect 25842 10446 25854 10449
rect 26002 10446 26014 10449
rect 26066 10446 26078 10498
rect 29138 10446 29150 10498
rect 29202 10446 29214 10498
rect 31266 10446 31278 10498
rect 31330 10446 31342 10498
rect 34066 10446 34078 10498
rect 34130 10446 34142 10498
rect 42130 10446 42142 10498
rect 42194 10446 42206 10498
rect 44258 10446 44270 10498
rect 44322 10446 44334 10498
rect 76514 10446 76526 10498
rect 76578 10446 76590 10498
rect 25342 10434 25394 10446
rect 41022 10434 41074 10446
rect 1344 10218 78624 10252
rect 1344 10166 4478 10218
rect 4530 10166 4582 10218
rect 4634 10166 4686 10218
rect 4738 10166 35198 10218
rect 35250 10166 35302 10218
rect 35354 10166 35406 10218
rect 35458 10166 65918 10218
rect 65970 10166 66022 10218
rect 66074 10166 66126 10218
rect 66178 10166 78624 10218
rect 1344 10132 78624 10166
rect 29150 10050 29202 10062
rect 29150 9986 29202 9998
rect 33966 10050 34018 10062
rect 33966 9986 34018 9998
rect 35758 10050 35810 10062
rect 35758 9986 35810 9998
rect 37438 10050 37490 10062
rect 37438 9986 37490 9998
rect 9438 9938 9490 9950
rect 27806 9938 27858 9950
rect 40350 9938 40402 9950
rect 44942 9938 44994 9950
rect 12450 9886 12462 9938
rect 12514 9935 12526 9938
rect 12674 9935 12686 9938
rect 12514 9889 12686 9935
rect 12514 9886 12526 9889
rect 12674 9886 12686 9889
rect 12738 9886 12750 9938
rect 15362 9886 15374 9938
rect 15426 9886 15438 9938
rect 34178 9886 34190 9938
rect 34242 9886 34254 9938
rect 34962 9886 34974 9938
rect 35026 9886 35038 9938
rect 41010 9886 41022 9938
rect 41074 9886 41086 9938
rect 44258 9886 44270 9938
rect 44322 9886 44334 9938
rect 9438 9874 9490 9886
rect 27806 9874 27858 9886
rect 40350 9874 40402 9886
rect 44942 9874 44994 9886
rect 11790 9826 11842 9838
rect 11790 9762 11842 9774
rect 12014 9826 12066 9838
rect 12798 9826 12850 9838
rect 20862 9826 20914 9838
rect 32398 9826 32450 9838
rect 12338 9774 12350 9826
rect 12402 9774 12414 9826
rect 20290 9774 20302 9826
rect 20354 9774 20366 9826
rect 22754 9774 22766 9826
rect 22818 9774 22830 9826
rect 12014 9762 12066 9774
rect 12798 9762 12850 9774
rect 20862 9762 20914 9774
rect 32398 9762 32450 9774
rect 33070 9826 33122 9838
rect 33070 9762 33122 9774
rect 33294 9826 33346 9838
rect 33294 9762 33346 9774
rect 35870 9826 35922 9838
rect 35870 9762 35922 9774
rect 36206 9826 36258 9838
rect 36206 9762 36258 9774
rect 37326 9826 37378 9838
rect 38670 9826 38722 9838
rect 39454 9826 39506 9838
rect 38098 9774 38110 9826
rect 38162 9774 38174 9826
rect 39218 9774 39230 9826
rect 39282 9774 39294 9826
rect 37326 9762 37378 9774
rect 38670 9762 38722 9774
rect 39454 9762 39506 9774
rect 39790 9826 39842 9838
rect 41346 9774 41358 9826
rect 41410 9774 41422 9826
rect 39790 9762 39842 9774
rect 1710 9714 1762 9726
rect 1710 9650 1762 9662
rect 2046 9714 2098 9726
rect 2046 9650 2098 9662
rect 9550 9714 9602 9726
rect 9550 9650 9602 9662
rect 11902 9714 11954 9726
rect 14702 9714 14754 9726
rect 29486 9714 29538 9726
rect 13458 9662 13470 9714
rect 13522 9662 13534 9714
rect 23650 9662 23662 9714
rect 23714 9662 23726 9714
rect 26898 9662 26910 9714
rect 26962 9662 26974 9714
rect 11902 9650 11954 9662
rect 14702 9650 14754 9662
rect 29486 9650 29538 9662
rect 32622 9714 32674 9726
rect 32622 9650 32674 9662
rect 33182 9714 33234 9726
rect 33182 9650 33234 9662
rect 33518 9714 33570 9726
rect 33518 9650 33570 9662
rect 34638 9714 34690 9726
rect 34638 9650 34690 9662
rect 36542 9714 36594 9726
rect 36542 9650 36594 9662
rect 40686 9714 40738 9726
rect 77646 9714 77698 9726
rect 42130 9662 42142 9714
rect 42194 9662 42206 9714
rect 45266 9662 45278 9714
rect 45330 9662 45342 9714
rect 40686 9650 40738 9662
rect 77646 9650 77698 9662
rect 78206 9714 78258 9726
rect 78206 9650 78258 9662
rect 2494 9602 2546 9614
rect 2494 9538 2546 9550
rect 9326 9602 9378 9614
rect 9326 9538 9378 9550
rect 13806 9602 13858 9614
rect 13806 9538 13858 9550
rect 14478 9602 14530 9614
rect 14478 9538 14530 9550
rect 14590 9602 14642 9614
rect 14590 9538 14642 9550
rect 27246 9602 27298 9614
rect 27246 9538 27298 9550
rect 28590 9602 28642 9614
rect 28590 9538 28642 9550
rect 29262 9602 29314 9614
rect 29262 9538 29314 9550
rect 29934 9602 29986 9614
rect 29934 9538 29986 9550
rect 30382 9602 30434 9614
rect 30382 9538 30434 9550
rect 31838 9602 31890 9614
rect 31838 9538 31890 9550
rect 32174 9602 32226 9614
rect 32174 9538 32226 9550
rect 32286 9602 32338 9614
rect 32286 9538 32338 9550
rect 34190 9602 34242 9614
rect 34190 9538 34242 9550
rect 34862 9602 34914 9614
rect 34862 9538 34914 9550
rect 35758 9602 35810 9614
rect 35758 9538 35810 9550
rect 36318 9602 36370 9614
rect 36318 9538 36370 9550
rect 37438 9602 37490 9614
rect 37438 9538 37490 9550
rect 37886 9602 37938 9614
rect 37886 9538 37938 9550
rect 38782 9602 38834 9614
rect 38782 9538 38834 9550
rect 38894 9602 38946 9614
rect 38894 9538 38946 9550
rect 39678 9602 39730 9614
rect 39678 9538 39730 9550
rect 75294 9602 75346 9614
rect 75294 9538 75346 9550
rect 75742 9602 75794 9614
rect 75742 9538 75794 9550
rect 76302 9602 76354 9614
rect 76302 9538 76354 9550
rect 76974 9602 77026 9614
rect 76974 9538 77026 9550
rect 77870 9602 77922 9614
rect 77870 9538 77922 9550
rect 1344 9434 78624 9468
rect 1344 9382 19838 9434
rect 19890 9382 19942 9434
rect 19994 9382 20046 9434
rect 20098 9382 50558 9434
rect 50610 9382 50662 9434
rect 50714 9382 50766 9434
rect 50818 9382 78624 9434
rect 1344 9348 78624 9382
rect 13358 9266 13410 9278
rect 17614 9266 17666 9278
rect 12562 9214 12574 9266
rect 12626 9214 12638 9266
rect 13010 9214 13022 9266
rect 13074 9214 13086 9266
rect 16706 9214 16718 9266
rect 16770 9214 16782 9266
rect 13358 9202 13410 9214
rect 17614 9202 17666 9214
rect 18510 9266 18562 9278
rect 18510 9202 18562 9214
rect 18622 9266 18674 9278
rect 18622 9202 18674 9214
rect 18846 9266 18898 9278
rect 24670 9266 24722 9278
rect 22306 9214 22318 9266
rect 22370 9214 22382 9266
rect 18846 9202 18898 9214
rect 24670 9202 24722 9214
rect 25230 9266 25282 9278
rect 43374 9266 43426 9278
rect 25554 9214 25566 9266
rect 25618 9214 25630 9266
rect 33506 9214 33518 9266
rect 33570 9214 33582 9266
rect 25230 9202 25282 9214
rect 43374 9202 43426 9214
rect 43486 9266 43538 9278
rect 43486 9202 43538 9214
rect 43598 9266 43650 9278
rect 43598 9202 43650 9214
rect 43934 9266 43986 9278
rect 43934 9202 43986 9214
rect 44046 9266 44098 9278
rect 44046 9202 44098 9214
rect 44158 9266 44210 9278
rect 44158 9202 44210 9214
rect 44382 9266 44434 9278
rect 44382 9202 44434 9214
rect 45614 9266 45666 9278
rect 45614 9202 45666 9214
rect 46062 9266 46114 9278
rect 46062 9202 46114 9214
rect 17726 9154 17778 9166
rect 42702 9154 42754 9166
rect 14466 9102 14478 9154
rect 14530 9102 14542 9154
rect 34962 9102 34974 9154
rect 35026 9102 35038 9154
rect 38210 9102 38222 9154
rect 38274 9102 38286 9154
rect 17726 9090 17778 9102
rect 42702 9090 42754 9102
rect 44942 9154 44994 9166
rect 44942 9090 44994 9102
rect 45054 9154 45106 9166
rect 45054 9090 45106 9102
rect 18398 9042 18450 9054
rect 33182 9042 33234 9054
rect 41022 9042 41074 9054
rect 9650 8990 9662 9042
rect 9714 8990 9726 9042
rect 13682 8990 13694 9042
rect 13746 8990 13758 9042
rect 17378 8990 17390 9042
rect 17442 8990 17454 9042
rect 19394 8990 19406 9042
rect 19458 8990 19470 9042
rect 25890 8990 25902 9042
rect 25954 8990 25966 9042
rect 29586 8990 29598 9042
rect 29650 8990 29662 9042
rect 34178 8990 34190 9042
rect 34242 8990 34254 9042
rect 37426 8990 37438 9042
rect 37490 8990 37502 9042
rect 18398 8978 18450 8990
rect 33182 8978 33234 8990
rect 41022 8978 41074 8990
rect 41134 9042 41186 9054
rect 41134 8978 41186 8990
rect 41246 9042 41298 9054
rect 41918 9042 41970 9054
rect 41458 8990 41470 9042
rect 41522 8990 41534 9042
rect 41246 8978 41298 8990
rect 41918 8978 41970 8990
rect 42142 9042 42194 9054
rect 42142 8978 42194 8990
rect 42926 9042 42978 9054
rect 75282 8990 75294 9042
rect 75346 8990 75358 9042
rect 77746 8990 77758 9042
rect 77810 8990 77822 9042
rect 42926 8978 42978 8990
rect 22990 8930 23042 8942
rect 10322 8878 10334 8930
rect 10386 8878 10398 8930
rect 20066 8878 20078 8930
rect 20130 8878 20142 8930
rect 22990 8866 23042 8878
rect 23550 8930 23602 8942
rect 23550 8866 23602 8878
rect 24334 8930 24386 8942
rect 26674 8878 26686 8930
rect 26738 8878 26750 8930
rect 28802 8878 28814 8930
rect 28866 8878 28878 8930
rect 30258 8878 30270 8930
rect 30322 8878 30334 8930
rect 32386 8878 32398 8930
rect 32450 8878 32462 8930
rect 37090 8878 37102 8930
rect 37154 8878 37166 8930
rect 40338 8878 40350 8930
rect 40402 8878 40414 8930
rect 24334 8866 24386 8878
rect 44942 8818 44994 8830
rect 75854 8818 75906 8830
rect 73378 8766 73390 8818
rect 73442 8766 73454 8818
rect 44942 8754 44994 8766
rect 75854 8754 75906 8766
rect 1344 8650 78624 8684
rect 1344 8598 4478 8650
rect 4530 8598 4582 8650
rect 4634 8598 4686 8650
rect 4738 8598 35198 8650
rect 35250 8598 35302 8650
rect 35354 8598 35406 8650
rect 35458 8598 65918 8650
rect 65970 8598 66022 8650
rect 66074 8598 66126 8650
rect 66178 8598 78624 8650
rect 1344 8564 78624 8598
rect 28142 8482 28194 8494
rect 28142 8418 28194 8430
rect 9326 8370 9378 8382
rect 9326 8306 9378 8318
rect 17838 8370 17890 8382
rect 17838 8306 17890 8318
rect 19966 8370 20018 8382
rect 26910 8370 26962 8382
rect 22866 8318 22878 8370
rect 22930 8318 22942 8370
rect 24994 8318 25006 8370
rect 25058 8318 25070 8370
rect 19966 8306 20018 8318
rect 26910 8306 26962 8318
rect 27358 8370 27410 8382
rect 27358 8306 27410 8318
rect 27470 8370 27522 8382
rect 27470 8306 27522 8318
rect 30158 8370 30210 8382
rect 30158 8306 30210 8318
rect 30270 8370 30322 8382
rect 30270 8306 30322 8318
rect 31166 8370 31218 8382
rect 31166 8306 31218 8318
rect 34638 8370 34690 8382
rect 36418 8318 36430 8370
rect 36482 8318 36494 8370
rect 38770 8318 38782 8370
rect 38834 8318 38846 8370
rect 40114 8318 40126 8370
rect 40178 8318 40190 8370
rect 42578 8318 42590 8370
rect 42642 8318 42654 8370
rect 45266 8318 45278 8370
rect 45330 8318 45342 8370
rect 74274 8318 74286 8370
rect 74338 8318 74350 8370
rect 34638 8306 34690 8318
rect 11006 8258 11058 8270
rect 11006 8194 11058 8206
rect 11790 8258 11842 8270
rect 11790 8194 11842 8206
rect 12014 8258 12066 8270
rect 18622 8258 18674 8270
rect 12338 8206 12350 8258
rect 12402 8206 12414 8258
rect 14914 8206 14926 8258
rect 14978 8206 14990 8258
rect 12014 8194 12066 8206
rect 18622 8194 18674 8206
rect 19854 8258 19906 8270
rect 19854 8194 19906 8206
rect 20078 8258 20130 8270
rect 20078 8194 20130 8206
rect 20526 8258 20578 8270
rect 25566 8258 25618 8270
rect 22082 8206 22094 8258
rect 22146 8206 22158 8258
rect 20526 8194 20578 8206
rect 25566 8194 25618 8206
rect 25790 8258 25842 8270
rect 25790 8194 25842 8206
rect 26238 8258 26290 8270
rect 26238 8194 26290 8206
rect 26798 8258 26850 8270
rect 32958 8258 33010 8270
rect 29922 8206 29934 8258
rect 29986 8206 29998 8258
rect 32162 8206 32174 8258
rect 32226 8206 32238 8258
rect 26798 8194 26850 8206
rect 32958 8194 33010 8206
rect 33854 8258 33906 8270
rect 33854 8194 33906 8206
rect 34750 8258 34802 8270
rect 34750 8194 34802 8206
rect 38894 8258 38946 8270
rect 38894 8194 38946 8206
rect 40686 8258 40738 8270
rect 40686 8194 40738 8206
rect 40798 8258 40850 8270
rect 76862 8258 76914 8270
rect 41794 8206 41806 8258
rect 41858 8206 41870 8258
rect 43026 8206 43038 8258
rect 43090 8206 43102 8258
rect 43586 8206 43598 8258
rect 43650 8206 43662 8258
rect 75506 8206 75518 8258
rect 75570 8206 75582 8258
rect 78082 8206 78094 8258
rect 78146 8206 78158 8258
rect 40798 8194 40850 8206
rect 76862 8194 76914 8206
rect 1710 8146 1762 8158
rect 1710 8082 1762 8094
rect 2046 8146 2098 8158
rect 2046 8082 2098 8094
rect 9438 8146 9490 8158
rect 9438 8082 9490 8094
rect 11902 8146 11954 8158
rect 11902 8082 11954 8094
rect 13022 8146 13074 8158
rect 13022 8082 13074 8094
rect 14254 8146 14306 8158
rect 14254 8082 14306 8094
rect 14590 8146 14642 8158
rect 18846 8146 18898 8158
rect 26574 8146 26626 8158
rect 15698 8094 15710 8146
rect 15762 8094 15774 8146
rect 21298 8094 21310 8146
rect 21362 8094 21374 8146
rect 14590 8082 14642 8094
rect 18846 8082 18898 8094
rect 26574 8082 26626 8094
rect 28142 8146 28194 8158
rect 28142 8082 28194 8094
rect 28254 8146 28306 8158
rect 34302 8146 34354 8158
rect 31938 8094 31950 8146
rect 32002 8094 32014 8146
rect 28254 8082 28306 8094
rect 34302 8082 34354 8094
rect 35422 8146 35474 8158
rect 35422 8082 35474 8094
rect 36094 8146 36146 8158
rect 36094 8082 36146 8094
rect 37102 8146 37154 8158
rect 37102 8082 37154 8094
rect 37774 8146 37826 8158
rect 37774 8082 37826 8094
rect 39230 8146 39282 8158
rect 44270 8146 44322 8158
rect 41122 8094 41134 8146
rect 41186 8094 41198 8146
rect 42914 8094 42926 8146
rect 42978 8094 42990 8146
rect 39230 8082 39282 8094
rect 44270 8082 44322 8094
rect 77198 8146 77250 8158
rect 77198 8082 77250 8094
rect 77534 8146 77586 8158
rect 77534 8082 77586 8094
rect 77870 8146 77922 8158
rect 77870 8082 77922 8094
rect 2494 8034 2546 8046
rect 2494 7970 2546 7982
rect 9214 8034 9266 8046
rect 9214 7970 9266 7982
rect 10670 8034 10722 8046
rect 10670 7970 10722 7982
rect 11454 8034 11506 8046
rect 11454 7970 11506 7982
rect 14030 8034 14082 8046
rect 14030 7970 14082 7982
rect 18398 8034 18450 8046
rect 18398 7970 18450 7982
rect 18510 8034 18562 8046
rect 18510 7970 18562 7982
rect 19630 8034 19682 8046
rect 19630 7970 19682 7982
rect 21646 8034 21698 8046
rect 21646 7970 21698 7982
rect 25678 8034 25730 8046
rect 25678 7970 25730 7982
rect 27022 8034 27074 8046
rect 27022 7970 27074 7982
rect 27582 8034 27634 8046
rect 27582 7970 27634 7982
rect 29710 8034 29762 8046
rect 29710 7970 29762 7982
rect 30830 8034 30882 8046
rect 30830 7970 30882 7982
rect 31726 8034 31778 8046
rect 34526 8034 34578 8046
rect 33282 7982 33294 8034
rect 33346 7982 33358 8034
rect 31726 7970 31778 7982
rect 34526 7970 34578 7982
rect 34974 8034 35026 8046
rect 34974 7970 35026 7982
rect 35758 8034 35810 8046
rect 35758 7970 35810 7982
rect 36318 8034 36370 8046
rect 36318 7970 36370 7982
rect 37438 8034 37490 8046
rect 37438 7970 37490 7982
rect 38110 8034 38162 8046
rect 38110 7970 38162 7982
rect 44158 8034 44210 8046
rect 44158 7970 44210 7982
rect 44830 8034 44882 8046
rect 44830 7970 44882 7982
rect 45950 8034 46002 8046
rect 45950 7970 46002 7982
rect 46286 8034 46338 8046
rect 46286 7970 46338 7982
rect 76302 8034 76354 8046
rect 76302 7970 76354 7982
rect 1344 7866 78624 7900
rect 1344 7814 19838 7866
rect 19890 7814 19942 7866
rect 19994 7814 20046 7866
rect 20098 7814 50558 7866
rect 50610 7814 50662 7866
rect 50714 7814 50766 7866
rect 50818 7814 78624 7866
rect 1344 7780 78624 7814
rect 2046 7698 2098 7710
rect 2046 7634 2098 7646
rect 15710 7698 15762 7710
rect 15710 7634 15762 7646
rect 16494 7698 16546 7710
rect 16494 7634 16546 7646
rect 16942 7698 16994 7710
rect 16942 7634 16994 7646
rect 17950 7698 18002 7710
rect 17950 7634 18002 7646
rect 18398 7698 18450 7710
rect 18398 7634 18450 7646
rect 19406 7698 19458 7710
rect 20638 7698 20690 7710
rect 25342 7698 25394 7710
rect 20290 7646 20302 7698
rect 20354 7646 20366 7698
rect 21410 7646 21422 7698
rect 21474 7646 21486 7698
rect 19406 7634 19458 7646
rect 20638 7634 20690 7646
rect 25342 7634 25394 7646
rect 26350 7698 26402 7710
rect 26350 7634 26402 7646
rect 26574 7698 26626 7710
rect 38222 7698 38274 7710
rect 66670 7698 66722 7710
rect 28130 7646 28142 7698
rect 28194 7646 28206 7698
rect 29026 7646 29038 7698
rect 29090 7646 29102 7698
rect 33394 7646 33406 7698
rect 33458 7646 33470 7698
rect 42914 7646 42926 7698
rect 42978 7646 42990 7698
rect 26574 7634 26626 7646
rect 38222 7634 38274 7646
rect 66670 7634 66722 7646
rect 15822 7586 15874 7598
rect 15822 7522 15874 7534
rect 19742 7586 19794 7598
rect 19742 7522 19794 7534
rect 19966 7586 20018 7598
rect 27694 7586 27746 7598
rect 26898 7534 26910 7586
rect 26962 7534 26974 7586
rect 19966 7522 20018 7534
rect 27694 7522 27746 7534
rect 30270 7586 30322 7598
rect 30270 7522 30322 7534
rect 31278 7586 31330 7598
rect 31278 7522 31330 7534
rect 32062 7586 32114 7598
rect 32062 7522 32114 7534
rect 32286 7586 32338 7598
rect 32286 7522 32338 7534
rect 34078 7586 34130 7598
rect 43038 7586 43090 7598
rect 38770 7534 38782 7586
rect 38834 7534 38846 7586
rect 39330 7534 39342 7586
rect 39394 7534 39406 7586
rect 41234 7534 41246 7586
rect 41298 7534 41310 7586
rect 34078 7522 34130 7534
rect 43038 7522 43090 7534
rect 44494 7586 44546 7598
rect 44494 7522 44546 7534
rect 46062 7586 46114 7598
rect 46062 7522 46114 7534
rect 71710 7586 71762 7598
rect 71710 7522 71762 7534
rect 1710 7474 1762 7486
rect 14030 7474 14082 7486
rect 10546 7422 10558 7474
rect 10610 7422 10622 7474
rect 1710 7410 1762 7422
rect 14030 7410 14082 7422
rect 14254 7474 14306 7486
rect 14254 7410 14306 7422
rect 14702 7474 14754 7486
rect 18174 7474 18226 7486
rect 15474 7422 15486 7474
rect 15538 7422 15550 7474
rect 14702 7410 14754 7422
rect 18174 7410 18226 7422
rect 18846 7474 18898 7486
rect 27806 7474 27858 7486
rect 21186 7422 21198 7474
rect 21250 7422 21262 7474
rect 21858 7422 21870 7474
rect 21922 7422 21934 7474
rect 18846 7410 18898 7422
rect 27806 7410 27858 7422
rect 29598 7474 29650 7486
rect 29598 7410 29650 7422
rect 29934 7474 29986 7486
rect 29934 7410 29986 7422
rect 30942 7474 30994 7486
rect 30942 7410 30994 7422
rect 33070 7474 33122 7486
rect 33070 7410 33122 7422
rect 33742 7474 33794 7486
rect 46846 7474 46898 7486
rect 34514 7422 34526 7474
rect 34578 7422 34590 7474
rect 35298 7422 35310 7474
rect 35362 7422 35374 7474
rect 40226 7422 40238 7474
rect 40290 7422 40302 7474
rect 41570 7422 41582 7474
rect 41634 7422 41646 7474
rect 41906 7422 41918 7474
rect 41970 7422 41982 7474
rect 43922 7422 43934 7474
rect 43986 7422 43998 7474
rect 46274 7422 46286 7474
rect 46338 7422 46350 7474
rect 66994 7422 67006 7474
rect 67058 7422 67070 7474
rect 72370 7422 72382 7474
rect 72434 7422 72446 7474
rect 75282 7422 75294 7474
rect 75346 7422 75358 7474
rect 33742 7410 33794 7422
rect 46846 7410 46898 7422
rect 2494 7362 2546 7374
rect 2494 7298 2546 7310
rect 9886 7362 9938 7374
rect 9886 7298 9938 7310
rect 10334 7362 10386 7374
rect 13470 7362 13522 7374
rect 11330 7310 11342 7362
rect 11394 7310 11406 7362
rect 10334 7298 10386 7310
rect 13470 7298 13522 7310
rect 14142 7362 14194 7374
rect 14142 7298 14194 7310
rect 15262 7362 15314 7374
rect 15262 7298 15314 7310
rect 18286 7362 18338 7374
rect 25790 7362 25842 7374
rect 19618 7310 19630 7362
rect 19682 7310 19694 7362
rect 22530 7310 22542 7362
rect 22594 7310 22606 7362
rect 24658 7310 24670 7362
rect 24722 7310 24734 7362
rect 18286 7298 18338 7310
rect 25790 7298 25842 7310
rect 28478 7362 28530 7374
rect 28478 7298 28530 7310
rect 28702 7362 28754 7374
rect 28702 7298 28754 7310
rect 29374 7362 29426 7374
rect 29374 7298 29426 7310
rect 31838 7362 31890 7374
rect 47518 7362 47570 7374
rect 32386 7310 32398 7362
rect 32450 7310 32462 7362
rect 37426 7310 37438 7362
rect 37490 7310 37502 7362
rect 39890 7310 39902 7362
rect 39954 7310 39966 7362
rect 41458 7310 41470 7362
rect 41522 7310 41534 7362
rect 31838 7298 31890 7310
rect 47518 7298 47570 7310
rect 48078 7362 48130 7374
rect 48078 7298 48130 7310
rect 60174 7362 60226 7374
rect 68562 7310 68574 7362
rect 68626 7310 68638 7362
rect 73938 7310 73950 7362
rect 74002 7310 74014 7362
rect 60174 7298 60226 7310
rect 27694 7250 27746 7262
rect 27694 7186 27746 7198
rect 38558 7250 38610 7262
rect 38558 7186 38610 7198
rect 76302 7250 76354 7262
rect 76302 7186 76354 7198
rect 1344 7082 78624 7116
rect 1344 7030 4478 7082
rect 4530 7030 4582 7082
rect 4634 7030 4686 7082
rect 4738 7030 35198 7082
rect 35250 7030 35302 7082
rect 35354 7030 35406 7082
rect 35458 7030 65918 7082
rect 65970 7030 66022 7082
rect 66074 7030 66126 7082
rect 66178 7030 78624 7082
rect 1344 6996 78624 7030
rect 9438 6914 9490 6926
rect 9438 6850 9490 6862
rect 11230 6914 11282 6926
rect 11230 6850 11282 6862
rect 8318 6802 8370 6814
rect 8318 6738 8370 6750
rect 8430 6802 8482 6814
rect 8430 6738 8482 6750
rect 8990 6802 9042 6814
rect 8990 6738 9042 6750
rect 9102 6802 9154 6814
rect 9102 6738 9154 6750
rect 9774 6802 9826 6814
rect 9774 6738 9826 6750
rect 11118 6802 11170 6814
rect 11118 6738 11170 6750
rect 19294 6802 19346 6814
rect 19294 6738 19346 6750
rect 20750 6802 20802 6814
rect 20750 6738 20802 6750
rect 23886 6802 23938 6814
rect 23886 6738 23938 6750
rect 26126 6802 26178 6814
rect 42254 6802 42306 6814
rect 33282 6750 33294 6802
rect 33346 6750 33358 6802
rect 40114 6750 40126 6802
rect 40178 6750 40190 6802
rect 26126 6738 26178 6750
rect 42254 6738 42306 6750
rect 13806 6690 13858 6702
rect 10322 6638 10334 6690
rect 10386 6638 10398 6690
rect 10882 6638 10894 6690
rect 10946 6638 10958 6690
rect 13806 6626 13858 6638
rect 15038 6690 15090 6702
rect 26014 6690 26066 6702
rect 16370 6638 16382 6690
rect 16434 6638 16446 6690
rect 17154 6638 17166 6690
rect 17218 6638 17230 6690
rect 20066 6638 20078 6690
rect 20130 6638 20142 6690
rect 22418 6638 22430 6690
rect 22482 6638 22494 6690
rect 15038 6626 15090 6638
rect 26014 6626 26066 6638
rect 26238 6690 26290 6702
rect 26238 6626 26290 6638
rect 26686 6690 26738 6702
rect 26686 6626 26738 6638
rect 27246 6690 27298 6702
rect 27246 6626 27298 6638
rect 28366 6690 28418 6702
rect 28366 6626 28418 6638
rect 28590 6690 28642 6702
rect 34414 6690 34466 6702
rect 29810 6638 29822 6690
rect 29874 6638 29886 6690
rect 30482 6638 30494 6690
rect 30546 6638 30558 6690
rect 28590 6626 28642 6638
rect 34414 6626 34466 6638
rect 34638 6690 34690 6702
rect 34638 6626 34690 6638
rect 34862 6690 34914 6702
rect 34862 6626 34914 6638
rect 35870 6690 35922 6702
rect 46510 6690 46562 6702
rect 50206 6690 50258 6702
rect 37314 6638 37326 6690
rect 37378 6638 37390 6690
rect 37986 6638 37998 6690
rect 38050 6638 38062 6690
rect 40450 6638 40462 6690
rect 40514 6638 40526 6690
rect 44258 6638 44270 6690
rect 44322 6638 44334 6690
rect 47058 6638 47070 6690
rect 47122 6638 47134 6690
rect 35870 6626 35922 6638
rect 46510 6626 46562 6638
rect 50206 6626 50258 6638
rect 51102 6690 51154 6702
rect 59502 6690 59554 6702
rect 51538 6638 51550 6690
rect 51602 6638 51614 6690
rect 51102 6626 51154 6638
rect 59502 6626 59554 6638
rect 60062 6690 60114 6702
rect 67902 6690 67954 6702
rect 74510 6690 74562 6702
rect 60498 6638 60510 6690
rect 60562 6638 60574 6690
rect 63410 6638 63422 6690
rect 63474 6638 63486 6690
rect 68338 6638 68350 6690
rect 68402 6638 68414 6690
rect 71250 6638 71262 6690
rect 71314 6638 71326 6690
rect 60062 6626 60114 6638
rect 67902 6626 67954 6638
rect 74510 6626 74562 6638
rect 74734 6690 74786 6702
rect 74734 6626 74786 6638
rect 76190 6690 76242 6702
rect 76190 6626 76242 6638
rect 76414 6690 76466 6702
rect 76414 6626 76466 6638
rect 10110 6578 10162 6590
rect 10110 6514 10162 6526
rect 16158 6578 16210 6590
rect 23214 6578 23266 6590
rect 19842 6526 19854 6578
rect 19906 6526 19918 6578
rect 16158 6514 16210 6526
rect 23214 6514 23266 6526
rect 23326 6578 23378 6590
rect 23326 6514 23378 6526
rect 23438 6578 23490 6590
rect 23438 6514 23490 6526
rect 23774 6578 23826 6590
rect 23774 6514 23826 6526
rect 25342 6578 25394 6590
rect 25342 6514 25394 6526
rect 25678 6578 25730 6590
rect 29262 6578 29314 6590
rect 28018 6526 28030 6578
rect 28082 6526 28094 6578
rect 25678 6514 25730 6526
rect 29262 6514 29314 6526
rect 29374 6578 29426 6590
rect 33742 6578 33794 6590
rect 31154 6526 31166 6578
rect 31218 6526 31230 6578
rect 29374 6514 29426 6526
rect 33742 6514 33794 6526
rect 33966 6578 34018 6590
rect 33966 6514 34018 6526
rect 35086 6578 35138 6590
rect 35086 6514 35138 6526
rect 36094 6578 36146 6590
rect 36094 6514 36146 6526
rect 41582 6578 41634 6590
rect 46062 6578 46114 6590
rect 50766 6578 50818 6590
rect 44146 6526 44158 6578
rect 44210 6526 44222 6578
rect 48626 6526 48638 6578
rect 48690 6526 48702 6578
rect 41582 6514 41634 6526
rect 46062 6514 46114 6526
rect 50766 6514 50818 6526
rect 77198 6578 77250 6590
rect 77198 6514 77250 6526
rect 77534 6578 77586 6590
rect 77534 6514 77586 6526
rect 77870 6578 77922 6590
rect 77870 6514 77922 6526
rect 78206 6578 78258 6590
rect 78206 6514 78258 6526
rect 7422 6466 7474 6478
rect 7422 6402 7474 6414
rect 7870 6466 7922 6478
rect 7870 6402 7922 6414
rect 8206 6466 8258 6478
rect 8206 6402 8258 6414
rect 8878 6466 8930 6478
rect 8878 6402 8930 6414
rect 9550 6466 9602 6478
rect 9550 6402 9602 6414
rect 12126 6466 12178 6478
rect 12126 6402 12178 6414
rect 12574 6466 12626 6478
rect 12574 6402 12626 6414
rect 13022 6466 13074 6478
rect 14478 6466 14530 6478
rect 15710 6466 15762 6478
rect 13458 6414 13470 6466
rect 13522 6414 13534 6466
rect 14690 6414 14702 6466
rect 14754 6414 14766 6466
rect 13022 6402 13074 6414
rect 14478 6402 14530 6414
rect 15710 6402 15762 6414
rect 21534 6466 21586 6478
rect 21534 6402 21586 6414
rect 21982 6466 22034 6478
rect 21982 6402 22034 6414
rect 22206 6466 22258 6478
rect 22206 6402 22258 6414
rect 23998 6466 24050 6478
rect 23998 6402 24050 6414
rect 24670 6466 24722 6478
rect 24670 6402 24722 6414
rect 25118 6466 25170 6478
rect 27806 6466 27858 6478
rect 26898 6414 26910 6466
rect 26962 6414 26974 6466
rect 25118 6402 25170 6414
rect 27806 6402 27858 6414
rect 29038 6466 29090 6478
rect 29038 6402 29090 6414
rect 30046 6466 30098 6478
rect 30046 6402 30098 6414
rect 33854 6466 33906 6478
rect 33854 6402 33906 6414
rect 34750 6466 34802 6478
rect 34750 6402 34802 6414
rect 36430 6466 36482 6478
rect 49086 6466 49138 6478
rect 46610 6414 46622 6466
rect 46674 6414 46686 6466
rect 36430 6402 36482 6414
rect 49086 6402 49138 6414
rect 52110 6466 52162 6478
rect 52110 6402 52162 6414
rect 56814 6466 56866 6478
rect 56814 6402 56866 6414
rect 61518 6466 61570 6478
rect 61518 6402 61570 6414
rect 64430 6466 64482 6478
rect 64430 6402 64482 6414
rect 67342 6466 67394 6478
rect 67342 6402 67394 6414
rect 69358 6466 69410 6478
rect 69358 6402 69410 6414
rect 72270 6466 72322 6478
rect 75518 6466 75570 6478
rect 75058 6414 75070 6466
rect 75122 6414 75134 6466
rect 76738 6414 76750 6466
rect 76802 6414 76814 6466
rect 72270 6402 72322 6414
rect 75518 6402 75570 6414
rect 1344 6298 78624 6332
rect 1344 6246 19838 6298
rect 19890 6246 19942 6298
rect 19994 6246 20046 6298
rect 20098 6246 50558 6298
rect 50610 6246 50662 6298
rect 50714 6246 50766 6298
rect 50818 6246 78624 6298
rect 1344 6212 78624 6246
rect 14254 6130 14306 6142
rect 2034 6078 2046 6130
rect 2098 6078 2110 6130
rect 14254 6066 14306 6078
rect 15598 6130 15650 6142
rect 18846 6130 18898 6142
rect 20190 6130 20242 6142
rect 18050 6078 18062 6130
rect 18114 6078 18126 6130
rect 19842 6078 19854 6130
rect 19906 6078 19918 6130
rect 15598 6066 15650 6078
rect 8990 6018 9042 6030
rect 8990 5954 9042 5966
rect 13582 6018 13634 6030
rect 13582 5954 13634 5966
rect 13918 6018 13970 6030
rect 13918 5954 13970 5966
rect 14702 6018 14754 6030
rect 14702 5954 14754 5966
rect 17502 6018 17554 6030
rect 17826 5966 17838 6018
rect 17890 6015 17902 6018
rect 18065 6015 18111 6078
rect 18846 6066 18898 6078
rect 20190 6066 20242 6078
rect 22094 6130 22146 6142
rect 22094 6066 22146 6078
rect 22654 6130 22706 6142
rect 22654 6066 22706 6078
rect 23550 6130 23602 6142
rect 23550 6066 23602 6078
rect 24782 6130 24834 6142
rect 24782 6066 24834 6078
rect 25902 6130 25954 6142
rect 25902 6066 25954 6078
rect 26350 6130 26402 6142
rect 26350 6066 26402 6078
rect 26798 6130 26850 6142
rect 26798 6066 26850 6078
rect 27582 6130 27634 6142
rect 29262 6130 29314 6142
rect 28018 6078 28030 6130
rect 28082 6078 28094 6130
rect 27582 6066 27634 6078
rect 29038 6074 29090 6086
rect 17890 5969 18111 6015
rect 22206 6018 22258 6030
rect 17890 5966 17902 5969
rect 17502 5954 17554 5966
rect 22206 5954 22258 5966
rect 22766 6018 22818 6030
rect 22766 5954 22818 5966
rect 23886 6018 23938 6030
rect 23886 5954 23938 5966
rect 24110 6018 24162 6030
rect 24110 5954 24162 5966
rect 27470 6018 27522 6030
rect 27470 5954 27522 5966
rect 28926 6018 28978 6030
rect 29262 6066 29314 6078
rect 29822 6130 29874 6142
rect 33182 6130 33234 6142
rect 31378 6078 31390 6130
rect 31442 6078 31454 6130
rect 29822 6066 29874 6078
rect 33182 6066 33234 6078
rect 33294 6130 33346 6142
rect 44942 6130 44994 6142
rect 35186 6078 35198 6130
rect 35250 6078 35262 6130
rect 33294 6066 33346 6078
rect 44942 6066 44994 6078
rect 56030 6130 56082 6142
rect 56030 6066 56082 6078
rect 63198 6130 63250 6142
rect 63198 6066 63250 6078
rect 63870 6130 63922 6142
rect 63870 6066 63922 6078
rect 78318 6130 78370 6142
rect 78318 6066 78370 6078
rect 29038 6010 29090 6022
rect 30494 6018 30546 6030
rect 29474 5966 29486 6018
rect 29538 5966 29550 6018
rect 28926 5954 28978 5966
rect 30494 5954 30546 5966
rect 31838 6018 31890 6030
rect 31838 5954 31890 5966
rect 32062 6018 32114 6030
rect 32062 5954 32114 5966
rect 34750 6018 34802 6030
rect 34750 5954 34802 5966
rect 35646 6018 35698 6030
rect 35646 5954 35698 5966
rect 37662 6018 37714 6030
rect 45614 6018 45666 6030
rect 39330 5966 39342 6018
rect 39394 5966 39406 6018
rect 40114 5966 40126 6018
rect 40178 5966 40190 6018
rect 42578 5966 42590 6018
rect 42642 5966 42654 6018
rect 37662 5954 37714 5966
rect 45614 5954 45666 5966
rect 47742 6018 47794 6030
rect 47742 5954 47794 5966
rect 1710 5906 1762 5918
rect 9886 5906 9938 5918
rect 14478 5906 14530 5918
rect 17726 5906 17778 5918
rect 21534 5906 21586 5918
rect 22542 5906 22594 5918
rect 26574 5906 26626 5918
rect 8642 5854 8654 5906
rect 8706 5854 8718 5906
rect 10210 5854 10222 5906
rect 10274 5854 10286 5906
rect 15362 5854 15374 5906
rect 15426 5854 15438 5906
rect 21186 5854 21198 5906
rect 21250 5854 21262 5906
rect 21858 5854 21870 5906
rect 21922 5854 21934 5906
rect 25666 5854 25678 5906
rect 25730 5854 25742 5906
rect 1710 5842 1762 5854
rect 9886 5842 9938 5854
rect 14478 5842 14530 5854
rect 17726 5842 17778 5854
rect 21534 5842 21586 5854
rect 22542 5842 22594 5854
rect 26574 5842 26626 5854
rect 28366 5906 28418 5918
rect 28366 5842 28418 5854
rect 28590 5906 28642 5918
rect 30830 5906 30882 5918
rect 30146 5854 30158 5906
rect 30210 5854 30222 5906
rect 28590 5842 28642 5854
rect 30830 5842 30882 5854
rect 31054 5906 31106 5918
rect 31054 5842 31106 5854
rect 32622 5906 32674 5918
rect 32622 5842 32674 5854
rect 33070 5906 33122 5918
rect 33070 5842 33122 5854
rect 33742 5906 33794 5918
rect 48750 5906 48802 5918
rect 71038 5906 71090 5918
rect 34402 5854 34414 5906
rect 34466 5854 34478 5906
rect 35074 5854 35086 5906
rect 35138 5854 35150 5906
rect 37090 5854 37102 5906
rect 37154 5854 37166 5906
rect 39218 5854 39230 5906
rect 39282 5854 39294 5906
rect 42466 5854 42478 5906
rect 42530 5854 42542 5906
rect 44482 5854 44494 5906
rect 44546 5854 44558 5906
rect 46946 5854 46958 5906
rect 47010 5854 47022 5906
rect 47954 5854 47966 5906
rect 48018 5854 48030 5906
rect 49186 5854 49198 5906
rect 49250 5854 49262 5906
rect 56914 5854 56926 5906
rect 56978 5854 56990 5906
rect 59826 5854 59838 5906
rect 59890 5854 59902 5906
rect 64418 5854 64430 5906
rect 64482 5854 64494 5906
rect 67330 5854 67342 5906
rect 67394 5854 67406 5906
rect 72258 5854 72270 5906
rect 72322 5854 72334 5906
rect 75170 5854 75182 5906
rect 75234 5854 75246 5906
rect 33742 5842 33794 5854
rect 48750 5842 48802 5854
rect 71038 5842 71090 5854
rect 2494 5794 2546 5806
rect 2494 5730 2546 5742
rect 6190 5794 6242 5806
rect 6190 5730 6242 5742
rect 6638 5794 6690 5806
rect 6638 5730 6690 5742
rect 7086 5794 7138 5806
rect 7086 5730 7138 5742
rect 7534 5794 7586 5806
rect 7534 5730 7586 5742
rect 7982 5794 8034 5806
rect 7982 5730 8034 5742
rect 8430 5794 8482 5806
rect 13022 5794 13074 5806
rect 8754 5742 8766 5794
rect 8818 5742 8830 5794
rect 10882 5742 10894 5794
rect 10946 5742 10958 5794
rect 8430 5730 8482 5742
rect 13022 5730 13074 5742
rect 14366 5794 14418 5806
rect 14366 5730 14418 5742
rect 16494 5794 16546 5806
rect 16494 5730 16546 5742
rect 16942 5794 16994 5806
rect 18398 5794 18450 5806
rect 17378 5742 17390 5794
rect 17442 5742 17454 5794
rect 16942 5730 16994 5742
rect 18398 5730 18450 5742
rect 19294 5794 19346 5806
rect 19294 5730 19346 5742
rect 20974 5794 21026 5806
rect 23998 5794 24050 5806
rect 21298 5742 21310 5794
rect 21362 5742 21374 5794
rect 20974 5730 21026 5742
rect 23998 5730 24050 5742
rect 25454 5794 25506 5806
rect 25454 5730 25506 5742
rect 26462 5794 26514 5806
rect 34190 5794 34242 5806
rect 40462 5794 40514 5806
rect 30258 5742 30270 5794
rect 30322 5742 30334 5794
rect 34514 5742 34526 5794
rect 34578 5742 34590 5794
rect 26462 5730 26514 5742
rect 34190 5730 34242 5742
rect 40462 5730 40514 5742
rect 41022 5794 41074 5806
rect 41022 5730 41074 5742
rect 41470 5794 41522 5806
rect 41470 5730 41522 5742
rect 42254 5794 42306 5806
rect 49758 5794 49810 5806
rect 46722 5742 46734 5794
rect 46786 5742 46798 5794
rect 42254 5730 42306 5742
rect 49758 5730 49810 5742
rect 50206 5794 50258 5806
rect 50206 5730 50258 5742
rect 50990 5794 51042 5806
rect 50990 5730 51042 5742
rect 51438 5794 51490 5806
rect 51438 5730 51490 5742
rect 52558 5794 52610 5806
rect 70478 5794 70530 5806
rect 65538 5742 65550 5794
rect 65602 5742 65614 5794
rect 68898 5742 68910 5794
rect 68962 5742 68974 5794
rect 52558 5730 52610 5742
rect 70478 5730 70530 5742
rect 71710 5794 71762 5806
rect 71710 5730 71762 5742
rect 15710 5682 15762 5694
rect 7410 5630 7422 5682
rect 7474 5679 7486 5682
rect 8082 5679 8094 5682
rect 7474 5633 8094 5679
rect 7474 5630 7486 5633
rect 8082 5630 8094 5633
rect 8146 5630 8158 5682
rect 15710 5618 15762 5630
rect 26014 5682 26066 5694
rect 26014 5618 26066 5630
rect 27694 5682 27746 5694
rect 27694 5618 27746 5630
rect 31726 5682 31778 5694
rect 57934 5682 57986 5694
rect 47282 5630 47294 5682
rect 47346 5630 47358 5682
rect 31726 5618 31778 5630
rect 57934 5618 57986 5630
rect 60846 5682 60898 5694
rect 60846 5618 60898 5630
rect 73278 5682 73330 5694
rect 73278 5618 73330 5630
rect 76190 5682 76242 5694
rect 76190 5618 76242 5630
rect 1344 5514 78624 5548
rect 1344 5462 4478 5514
rect 4530 5462 4582 5514
rect 4634 5462 4686 5514
rect 4738 5462 35198 5514
rect 35250 5462 35302 5514
rect 35354 5462 35406 5514
rect 35458 5462 65918 5514
rect 65970 5462 66022 5514
rect 66074 5462 66126 5514
rect 66178 5462 78624 5514
rect 1344 5428 78624 5462
rect 21758 5346 21810 5358
rect 7186 5294 7198 5346
rect 7250 5343 7262 5346
rect 7858 5343 7870 5346
rect 7250 5297 7870 5343
rect 7250 5294 7262 5297
rect 7858 5294 7870 5297
rect 7922 5294 7934 5346
rect 21758 5282 21810 5294
rect 22094 5346 22146 5358
rect 22094 5282 22146 5294
rect 27246 5346 27298 5358
rect 27246 5282 27298 5294
rect 29598 5346 29650 5358
rect 29598 5282 29650 5294
rect 30270 5346 30322 5358
rect 30270 5282 30322 5294
rect 30942 5346 30994 5358
rect 74846 5346 74898 5358
rect 37090 5294 37102 5346
rect 37154 5343 37166 5346
rect 37426 5343 37438 5346
rect 37154 5297 37438 5343
rect 37154 5294 37166 5297
rect 37426 5294 37438 5297
rect 37490 5294 37502 5346
rect 50306 5294 50318 5346
rect 50370 5343 50382 5346
rect 50978 5343 50990 5346
rect 50370 5297 50990 5343
rect 50370 5294 50382 5297
rect 50978 5294 50990 5297
rect 51042 5343 51054 5346
rect 51986 5343 51998 5346
rect 51042 5297 51998 5343
rect 51042 5294 51054 5297
rect 51986 5294 51998 5297
rect 52050 5294 52062 5346
rect 67330 5294 67342 5346
rect 67394 5343 67406 5346
rect 67554 5343 67566 5346
rect 67394 5297 67566 5343
rect 67394 5294 67406 5297
rect 67554 5294 67566 5297
rect 67618 5294 67630 5346
rect 30942 5282 30994 5294
rect 74846 5282 74898 5294
rect 7422 5234 7474 5246
rect 7422 5170 7474 5182
rect 7870 5234 7922 5246
rect 7870 5170 7922 5182
rect 8318 5234 8370 5246
rect 10782 5234 10834 5246
rect 10210 5182 10222 5234
rect 10274 5182 10286 5234
rect 8318 5170 8370 5182
rect 10782 5170 10834 5182
rect 10894 5234 10946 5246
rect 10894 5170 10946 5182
rect 13582 5234 13634 5246
rect 17278 5234 17330 5246
rect 18622 5234 18674 5246
rect 15138 5182 15150 5234
rect 15202 5182 15214 5234
rect 17938 5182 17950 5234
rect 18002 5182 18014 5234
rect 13582 5170 13634 5182
rect 17278 5170 17330 5182
rect 18622 5170 18674 5182
rect 19966 5234 20018 5246
rect 19966 5170 20018 5182
rect 21534 5234 21586 5246
rect 26686 5234 26738 5246
rect 23986 5182 23998 5234
rect 24050 5182 24062 5234
rect 26114 5182 26126 5234
rect 26178 5182 26190 5234
rect 21534 5170 21586 5182
rect 26686 5170 26738 5182
rect 27134 5234 27186 5246
rect 27134 5170 27186 5182
rect 31838 5234 31890 5246
rect 50878 5234 50930 5246
rect 46946 5182 46958 5234
rect 47010 5182 47022 5234
rect 31838 5170 31890 5182
rect 50878 5170 50930 5182
rect 51326 5234 51378 5246
rect 51326 5170 51378 5182
rect 54014 5234 54066 5246
rect 54014 5170 54066 5182
rect 55246 5234 55298 5246
rect 55246 5170 55298 5182
rect 58158 5234 58210 5246
rect 58158 5170 58210 5182
rect 64430 5234 64482 5246
rect 64430 5170 64482 5182
rect 66446 5234 66498 5246
rect 66446 5170 66498 5182
rect 67118 5234 67170 5246
rect 67118 5170 67170 5182
rect 69358 5234 69410 5246
rect 69358 5170 69410 5182
rect 74398 5234 74450 5246
rect 74398 5170 74450 5182
rect 74622 5234 74674 5246
rect 76626 5182 76638 5234
rect 76690 5182 76702 5234
rect 74622 5170 74674 5182
rect 1710 5122 1762 5134
rect 1710 5058 1762 5070
rect 2494 5122 2546 5134
rect 2494 5058 2546 5070
rect 6190 5122 6242 5134
rect 8766 5122 8818 5134
rect 6514 5070 6526 5122
rect 6578 5070 6590 5122
rect 6190 5058 6242 5070
rect 8766 5058 8818 5070
rect 8878 5122 8930 5134
rect 8878 5058 8930 5070
rect 9550 5122 9602 5134
rect 11902 5122 11954 5134
rect 11554 5070 11566 5122
rect 11618 5070 11630 5122
rect 9550 5058 9602 5070
rect 11902 5058 11954 5070
rect 12462 5122 12514 5134
rect 12462 5058 12514 5070
rect 13022 5122 13074 5134
rect 13022 5058 13074 5070
rect 13470 5122 13522 5134
rect 13470 5058 13522 5070
rect 14142 5122 14194 5134
rect 19518 5122 19570 5134
rect 14354 5070 14366 5122
rect 14418 5070 14430 5122
rect 17826 5070 17838 5122
rect 17890 5070 17902 5122
rect 18834 5070 18846 5122
rect 18898 5070 18910 5122
rect 14142 5058 14194 5070
rect 19518 5058 19570 5070
rect 22878 5122 22930 5134
rect 27918 5122 27970 5134
rect 29486 5122 29538 5134
rect 23202 5070 23214 5122
rect 23266 5070 23278 5122
rect 28354 5070 28366 5122
rect 28418 5070 28430 5122
rect 29250 5070 29262 5122
rect 29314 5070 29326 5122
rect 22878 5058 22930 5070
rect 27918 5058 27970 5070
rect 29486 5058 29538 5070
rect 30158 5122 30210 5134
rect 30158 5058 30210 5070
rect 30830 5122 30882 5134
rect 30830 5058 30882 5070
rect 31278 5122 31330 5134
rect 31278 5058 31330 5070
rect 32398 5122 32450 5134
rect 37438 5122 37490 5134
rect 49310 5122 49362 5134
rect 50430 5122 50482 5134
rect 32610 5070 32622 5122
rect 32674 5070 32686 5122
rect 36418 5070 36430 5122
rect 36482 5070 36494 5122
rect 37090 5070 37102 5122
rect 37154 5070 37166 5122
rect 37538 5070 37550 5122
rect 37602 5070 37614 5122
rect 38882 5070 38894 5122
rect 38946 5070 38958 5122
rect 42018 5070 42030 5122
rect 42082 5070 42094 5122
rect 42466 5070 42478 5122
rect 42530 5070 42542 5122
rect 44818 5070 44830 5122
rect 44882 5070 44894 5122
rect 46834 5070 46846 5122
rect 46898 5070 46910 5122
rect 49858 5070 49870 5122
rect 49922 5070 49934 5122
rect 32398 5058 32450 5070
rect 37438 5058 37490 5070
rect 49310 5058 49362 5070
rect 50430 5058 50482 5070
rect 51774 5122 51826 5134
rect 51774 5058 51826 5070
rect 52782 5122 52834 5134
rect 75630 5122 75682 5134
rect 77198 5122 77250 5134
rect 54226 5070 54238 5122
rect 54290 5070 54302 5122
rect 57138 5070 57150 5122
rect 57202 5070 57214 5122
rect 60498 5070 60510 5122
rect 60562 5070 60574 5122
rect 63522 5070 63534 5122
rect 63586 5070 63598 5122
rect 68338 5070 68350 5122
rect 68402 5070 68414 5122
rect 71362 5070 71374 5122
rect 71426 5070 71438 5122
rect 76290 5070 76302 5122
rect 76354 5070 76366 5122
rect 77746 5070 77758 5122
rect 77810 5070 77822 5122
rect 52782 5058 52834 5070
rect 75630 5058 75682 5070
rect 77198 5058 77250 5070
rect 6750 5010 6802 5022
rect 2034 4958 2046 5010
rect 2098 4958 2110 5010
rect 6750 4946 6802 4958
rect 9214 5010 9266 5022
rect 9214 4946 9266 4958
rect 9886 5010 9938 5022
rect 9886 4946 9938 4958
rect 10670 5010 10722 5022
rect 10670 4946 10722 4958
rect 12574 5010 12626 5022
rect 12574 4946 12626 4958
rect 13694 5010 13746 5022
rect 13694 4946 13746 4958
rect 18174 5010 18226 5022
rect 18174 4946 18226 4958
rect 18510 5010 18562 5022
rect 18510 4946 18562 4958
rect 20414 5010 20466 5022
rect 20414 4946 20466 4958
rect 22542 5010 22594 5022
rect 22542 4946 22594 4958
rect 27582 5010 27634 5022
rect 27582 4946 27634 4958
rect 28590 5010 28642 5022
rect 28590 4946 28642 4958
rect 30718 5010 30770 5022
rect 35870 5010 35922 5022
rect 32722 4958 32734 5010
rect 32786 4958 32798 5010
rect 30718 4946 30770 4958
rect 35870 4946 35922 4958
rect 38334 5010 38386 5022
rect 40014 5010 40066 5022
rect 43598 5010 43650 5022
rect 38994 4958 39006 5010
rect 39058 4958 39070 5010
rect 39666 4958 39678 5010
rect 39730 4958 39742 5010
rect 40562 4958 40574 5010
rect 40626 4958 40638 5010
rect 38334 4946 38386 4958
rect 40014 4946 40066 4958
rect 43598 4946 43650 4958
rect 45390 5010 45442 5022
rect 45390 4946 45442 4958
rect 47406 5010 47458 5022
rect 47406 4946 47458 4958
rect 48974 5010 49026 5022
rect 48974 4946 49026 4958
rect 49646 5010 49698 5022
rect 77522 4958 77534 5010
rect 77586 4958 77598 5010
rect 49646 4946 49698 4958
rect 5182 4898 5234 4910
rect 5182 4834 5234 4846
rect 8654 4898 8706 4910
rect 8654 4834 8706 4846
rect 10110 4898 10162 4910
rect 10110 4834 10162 4846
rect 11790 4898 11842 4910
rect 11790 4834 11842 4846
rect 12350 4898 12402 4910
rect 12350 4834 12402 4846
rect 20862 4898 20914 4910
rect 20862 4834 20914 4846
rect 21870 4898 21922 4910
rect 21870 4834 21922 4846
rect 27022 4898 27074 4910
rect 27022 4834 27074 4846
rect 30046 4898 30098 4910
rect 30046 4834 30098 4846
rect 33966 4898 34018 4910
rect 33966 4834 34018 4846
rect 42926 4898 42978 4910
rect 42926 4834 42978 4846
rect 53342 4898 53394 4910
rect 53342 4834 53394 4846
rect 61518 4898 61570 4910
rect 61518 4834 61570 4846
rect 67454 4898 67506 4910
rect 67454 4834 67506 4846
rect 72270 4898 72322 4910
rect 75170 4846 75182 4898
rect 75234 4846 75246 4898
rect 72270 4834 72322 4846
rect 1344 4730 78624 4764
rect 1344 4678 19838 4730
rect 19890 4678 19942 4730
rect 19994 4678 20046 4730
rect 20098 4678 50558 4730
rect 50610 4678 50662 4730
rect 50714 4678 50766 4730
rect 50818 4678 78624 4730
rect 1344 4644 78624 4678
rect 6190 4562 6242 4574
rect 6190 4498 6242 4510
rect 7534 4562 7586 4574
rect 7534 4498 7586 4510
rect 8206 4562 8258 4574
rect 8206 4498 8258 4510
rect 8990 4562 9042 4574
rect 8990 4498 9042 4510
rect 9998 4562 10050 4574
rect 9998 4498 10050 4510
rect 15374 4562 15426 4574
rect 15374 4498 15426 4510
rect 15822 4562 15874 4574
rect 15822 4498 15874 4510
rect 16718 4562 16770 4574
rect 16718 4498 16770 4510
rect 17838 4562 17890 4574
rect 17838 4498 17890 4510
rect 18622 4562 18674 4574
rect 18622 4498 18674 4510
rect 19294 4562 19346 4574
rect 19294 4498 19346 4510
rect 22654 4562 22706 4574
rect 40910 4562 40962 4574
rect 55918 4562 55970 4574
rect 40226 4510 40238 4562
rect 40290 4510 40302 4562
rect 43810 4510 43822 4562
rect 43874 4510 43886 4562
rect 48738 4510 48750 4562
rect 48802 4510 48814 4562
rect 22654 4498 22706 4510
rect 40910 4498 40962 4510
rect 55918 4498 55970 4510
rect 62526 4562 62578 4574
rect 62526 4498 62578 4510
rect 63198 4562 63250 4574
rect 63198 4498 63250 4510
rect 63534 4562 63586 4574
rect 63534 4498 63586 4510
rect 71038 4562 71090 4574
rect 71038 4498 71090 4510
rect 78206 4562 78258 4574
rect 78206 4498 78258 4510
rect 5182 4450 5234 4462
rect 5182 4386 5234 4398
rect 5854 4450 5906 4462
rect 5854 4386 5906 4398
rect 6974 4450 7026 4462
rect 6974 4386 7026 4398
rect 7646 4450 7698 4462
rect 7646 4386 7698 4398
rect 8318 4450 8370 4462
rect 8318 4386 8370 4398
rect 10334 4450 10386 4462
rect 10334 4386 10386 4398
rect 10670 4450 10722 4462
rect 14814 4450 14866 4462
rect 11778 4398 11790 4450
rect 11842 4398 11854 4450
rect 10670 4386 10722 4398
rect 14814 4386 14866 4398
rect 15486 4450 15538 4462
rect 15486 4386 15538 4398
rect 16158 4450 16210 4462
rect 16158 4386 16210 4398
rect 18286 4450 18338 4462
rect 18286 4386 18338 4398
rect 19630 4450 19682 4462
rect 19630 4386 19682 4398
rect 19966 4450 20018 4462
rect 19966 4386 20018 4398
rect 21310 4450 21362 4462
rect 21310 4386 21362 4398
rect 21758 4450 21810 4462
rect 21758 4386 21810 4398
rect 21982 4450 22034 4462
rect 21982 4386 22034 4398
rect 23326 4450 23378 4462
rect 23326 4386 23378 4398
rect 23662 4450 23714 4462
rect 23662 4386 23714 4398
rect 23998 4450 24050 4462
rect 23998 4386 24050 4398
rect 24334 4450 24386 4462
rect 24334 4386 24386 4398
rect 24670 4450 24722 4462
rect 24670 4386 24722 4398
rect 29262 4450 29314 4462
rect 29262 4386 29314 4398
rect 31278 4450 31330 4462
rect 37102 4450 37154 4462
rect 34066 4398 34078 4450
rect 34130 4398 34142 4450
rect 31278 4386 31330 4398
rect 37102 4386 37154 4398
rect 39118 4450 39170 4462
rect 39118 4386 39170 4398
rect 41022 4450 41074 4462
rect 41022 4386 41074 4398
rect 42814 4450 42866 4462
rect 42814 4386 42866 4398
rect 45390 4450 45442 4462
rect 46386 4398 46398 4450
rect 46450 4398 46462 4450
rect 46610 4398 46622 4450
rect 46674 4398 46686 4450
rect 45390 4386 45442 4398
rect 38670 4338 38722 4350
rect 6738 4286 6750 4338
rect 6802 4286 6814 4338
rect 7298 4286 7310 4338
rect 7362 4286 7374 4338
rect 7970 4286 7982 4338
rect 8034 4286 8046 4338
rect 8754 4286 8766 4338
rect 8818 4286 8830 4338
rect 9762 4286 9774 4338
rect 9826 4286 9838 4338
rect 10994 4286 11006 4338
rect 11058 4286 11070 4338
rect 14578 4286 14590 4338
rect 14642 4286 14654 4338
rect 15138 4286 15150 4338
rect 15202 4286 15214 4338
rect 16482 4286 16494 4338
rect 16546 4286 16558 4338
rect 17602 4286 17614 4338
rect 17666 4286 17678 4338
rect 19058 4286 19070 4338
rect 19122 4286 19134 4338
rect 20290 4286 20302 4338
rect 20354 4286 20366 4338
rect 20962 4286 20974 4338
rect 21026 4286 21038 4338
rect 22418 4286 22430 4338
rect 22482 4286 22494 4338
rect 22978 4286 22990 4338
rect 23042 4286 23054 4338
rect 25218 4286 25230 4338
rect 25282 4286 25294 4338
rect 28690 4286 28702 4338
rect 28754 4286 28766 4338
rect 30706 4286 30718 4338
rect 30770 4286 30782 4338
rect 33394 4286 33406 4338
rect 33458 4286 33470 4338
rect 38098 4286 38110 4338
rect 38162 4286 38174 4338
rect 38670 4274 38722 4286
rect 41918 4338 41970 4350
rect 49086 4338 49138 4350
rect 42242 4286 42254 4338
rect 42306 4286 42318 4338
rect 44258 4286 44270 4338
rect 44322 4286 44334 4338
rect 47282 4286 47294 4338
rect 47346 4286 47358 4338
rect 49522 4286 49534 4338
rect 49586 4286 49598 4338
rect 52882 4286 52894 4338
rect 52946 4286 52958 4338
rect 56578 4286 56590 4338
rect 56642 4286 56654 4338
rect 61618 4286 61630 4338
rect 61682 4286 61694 4338
rect 64530 4286 64542 4338
rect 64594 4286 64606 4338
rect 67330 4286 67342 4338
rect 67394 4286 67406 4338
rect 72258 4286 72270 4338
rect 72322 4286 72334 4338
rect 75394 4286 75406 4338
rect 75458 4286 75470 4338
rect 41918 4274 41970 4286
rect 49086 4274 49138 4286
rect 2158 4226 2210 4238
rect 2158 4162 2210 4174
rect 4734 4226 4786 4238
rect 4734 4162 4786 4174
rect 5630 4226 5682 4238
rect 5630 4162 5682 4174
rect 13918 4226 13970 4238
rect 23214 4226 23266 4238
rect 52558 4226 52610 4238
rect 70478 4226 70530 4238
rect 21074 4174 21086 4226
rect 21138 4174 21150 4226
rect 21634 4174 21646 4226
rect 21698 4174 21710 4226
rect 26002 4174 26014 4226
rect 26066 4174 26078 4226
rect 28130 4174 28142 4226
rect 28194 4174 28206 4226
rect 31826 4174 31838 4226
rect 31890 4174 31902 4226
rect 36194 4174 36206 4226
rect 36258 4174 36270 4226
rect 41458 4174 41470 4226
rect 41522 4174 41534 4226
rect 65538 4174 65550 4226
rect 65602 4174 65614 4226
rect 13918 4162 13970 4174
rect 23214 4162 23266 4174
rect 52558 4162 52610 4174
rect 70478 4162 70530 4174
rect 71710 4226 71762 4238
rect 71710 4162 71762 4174
rect 16830 4114 16882 4126
rect 16830 4050 16882 4062
rect 17950 4114 18002 4126
rect 17950 4050 18002 4062
rect 20302 4114 20354 4126
rect 20302 4050 20354 4062
rect 20638 4114 20690 4126
rect 20638 4050 20690 4062
rect 50542 4114 50594 4126
rect 50542 4050 50594 4062
rect 53902 4114 53954 4126
rect 53902 4050 53954 4062
rect 57598 4114 57650 4126
rect 57598 4050 57650 4062
rect 59726 4114 59778 4126
rect 59726 4050 59778 4062
rect 68350 4114 68402 4126
rect 68350 4050 68402 4062
rect 73278 4114 73330 4126
rect 73278 4050 73330 4062
rect 76190 4114 76242 4126
rect 76190 4050 76242 4062
rect 1344 3946 78624 3980
rect 1344 3894 4478 3946
rect 4530 3894 4582 3946
rect 4634 3894 4686 3946
rect 4738 3894 35198 3946
rect 35250 3894 35302 3946
rect 35354 3894 35406 3946
rect 35458 3894 65918 3946
rect 65970 3894 66022 3946
rect 66074 3894 66126 3946
rect 66178 3894 78624 3946
rect 1344 3860 78624 3894
rect 11566 3778 11618 3790
rect 11566 3714 11618 3726
rect 13694 3778 13746 3790
rect 13694 3714 13746 3726
rect 23326 3778 23378 3790
rect 23326 3714 23378 3726
rect 39118 3778 39170 3790
rect 39118 3714 39170 3726
rect 47630 3778 47682 3790
rect 47630 3714 47682 3726
rect 67454 3778 67506 3790
rect 67454 3714 67506 3726
rect 75070 3778 75122 3790
rect 75070 3714 75122 3726
rect 11118 3666 11170 3678
rect 47406 3666 47458 3678
rect 54238 3666 54290 3678
rect 23090 3614 23102 3666
rect 23154 3614 23166 3666
rect 32498 3614 32510 3666
rect 32562 3614 32574 3666
rect 42802 3614 42814 3666
rect 42866 3614 42878 3666
rect 45714 3614 45726 3666
rect 45778 3614 45790 3666
rect 47954 3614 47966 3666
rect 48018 3614 48030 3666
rect 11118 3602 11170 3614
rect 47406 3602 47458 3614
rect 54238 3602 54290 3614
rect 56030 3666 56082 3678
rect 56030 3602 56082 3614
rect 58046 3666 58098 3678
rect 58046 3602 58098 3614
rect 59054 3666 59106 3678
rect 65662 3666 65714 3678
rect 63858 3614 63870 3666
rect 63922 3614 63934 3666
rect 59054 3602 59106 3614
rect 65662 3602 65714 3614
rect 69806 3666 69858 3678
rect 69806 3602 69858 3614
rect 71262 3666 71314 3678
rect 71262 3602 71314 3614
rect 73614 3666 73666 3678
rect 73614 3602 73666 3614
rect 5742 3554 5794 3566
rect 4722 3502 4734 3554
rect 4786 3502 4798 3554
rect 5742 3490 5794 3502
rect 6414 3554 6466 3566
rect 8430 3554 8482 3566
rect 7186 3502 7198 3554
rect 7250 3502 7262 3554
rect 7858 3502 7870 3554
rect 7922 3502 7934 3554
rect 6414 3490 6466 3502
rect 8430 3490 8482 3502
rect 9550 3554 9602 3566
rect 9550 3490 9602 3502
rect 10222 3554 10274 3566
rect 13582 3554 13634 3566
rect 14702 3554 14754 3566
rect 10882 3502 10894 3554
rect 10946 3502 10958 3554
rect 11554 3502 11566 3554
rect 11618 3502 11630 3554
rect 13346 3502 13358 3554
rect 13410 3502 13422 3554
rect 14130 3502 14142 3554
rect 14194 3502 14206 3554
rect 10222 3490 10274 3502
rect 13582 3490 13634 3502
rect 14702 3490 14754 3502
rect 15374 3554 15426 3566
rect 17166 3554 17218 3566
rect 16146 3502 16158 3554
rect 16210 3502 16222 3554
rect 15374 3490 15426 3502
rect 17166 3490 17218 3502
rect 17838 3554 17890 3566
rect 19854 3554 19906 3566
rect 18610 3502 18622 3554
rect 18674 3502 18686 3554
rect 19282 3502 19294 3554
rect 19346 3502 19358 3554
rect 17838 3490 17890 3502
rect 19854 3490 19906 3502
rect 20974 3554 21026 3566
rect 22318 3554 22370 3566
rect 23662 3554 23714 3566
rect 21746 3502 21758 3554
rect 21810 3502 21822 3554
rect 22978 3502 22990 3554
rect 23042 3502 23054 3554
rect 20974 3490 21026 3502
rect 22318 3490 22370 3502
rect 23662 3490 23714 3502
rect 24782 3554 24834 3566
rect 24782 3490 24834 3502
rect 25342 3554 25394 3566
rect 25342 3490 25394 3502
rect 26126 3554 26178 3566
rect 61854 3554 61906 3566
rect 76974 3554 77026 3566
rect 27570 3502 27582 3554
rect 27634 3502 27646 3554
rect 30706 3502 30718 3554
rect 30770 3502 30782 3554
rect 31378 3502 31390 3554
rect 31442 3502 31454 3554
rect 33954 3502 33966 3554
rect 34018 3502 34030 3554
rect 35074 3502 35086 3554
rect 35138 3502 35150 3554
rect 36866 3502 36878 3554
rect 36930 3502 36942 3554
rect 39218 3502 39230 3554
rect 39282 3502 39294 3554
rect 41346 3502 41358 3554
rect 41410 3502 41422 3554
rect 43026 3502 43038 3554
rect 43090 3502 43102 3554
rect 43698 3502 43710 3554
rect 43762 3502 43774 3554
rect 45266 3502 45278 3554
rect 45330 3502 45342 3554
rect 48514 3502 48526 3554
rect 48578 3502 48590 3554
rect 49186 3502 49198 3554
rect 49250 3502 49262 3554
rect 49858 3502 49870 3554
rect 49922 3502 49934 3554
rect 50530 3502 50542 3554
rect 50594 3502 50606 3554
rect 51650 3502 51662 3554
rect 51714 3502 51726 3554
rect 52322 3502 52334 3554
rect 52386 3502 52398 3554
rect 52994 3502 53006 3554
rect 53058 3502 53070 3554
rect 53666 3502 53678 3554
rect 53730 3502 53742 3554
rect 55458 3502 55470 3554
rect 55522 3502 55534 3554
rect 60946 3502 60958 3554
rect 61010 3502 61022 3554
rect 63074 3502 63086 3554
rect 63138 3502 63150 3554
rect 66434 3502 66446 3554
rect 66498 3502 66510 3554
rect 70242 3502 70254 3554
rect 70306 3502 70318 3554
rect 74050 3502 74062 3554
rect 74114 3502 74126 3554
rect 26126 3490 26178 3502
rect 61854 3490 61906 3502
rect 76974 3490 77026 3502
rect 77870 3554 77922 3566
rect 77870 3490 77922 3502
rect 1710 3442 1762 3454
rect 2382 3442 2434 3454
rect 3166 3442 3218 3454
rect 2034 3390 2046 3442
rect 2098 3390 2110 3442
rect 2706 3390 2718 3442
rect 2770 3390 2782 3442
rect 1710 3378 1762 3390
rect 2382 3378 2434 3390
rect 3166 3378 3218 3390
rect 3726 3442 3778 3454
rect 3726 3378 3778 3390
rect 3950 3442 4002 3454
rect 3950 3378 4002 3390
rect 4286 3442 4338 3454
rect 4286 3378 4338 3390
rect 4958 3442 5010 3454
rect 4958 3378 5010 3390
rect 6078 3442 6130 3454
rect 6078 3378 6130 3390
rect 6750 3442 6802 3454
rect 6750 3378 6802 3390
rect 7422 3442 7474 3454
rect 7422 3378 7474 3390
rect 8094 3442 8146 3454
rect 8094 3378 8146 3390
rect 9886 3442 9938 3454
rect 9886 3378 9938 3390
rect 10558 3442 10610 3454
rect 10558 3378 10610 3390
rect 11230 3442 11282 3454
rect 11230 3378 11282 3390
rect 11902 3442 11954 3454
rect 11902 3378 11954 3390
rect 12238 3442 12290 3454
rect 12238 3378 12290 3390
rect 12574 3442 12626 3454
rect 12574 3378 12626 3390
rect 15038 3442 15090 3454
rect 15038 3378 15090 3390
rect 15710 3442 15762 3454
rect 15710 3378 15762 3390
rect 16382 3442 16434 3454
rect 16382 3378 16434 3390
rect 17502 3442 17554 3454
rect 17502 3378 17554 3390
rect 18174 3442 18226 3454
rect 18174 3378 18226 3390
rect 19518 3442 19570 3454
rect 19518 3378 19570 3390
rect 20190 3442 20242 3454
rect 20190 3378 20242 3390
rect 21310 3442 21362 3454
rect 21310 3378 21362 3390
rect 21982 3442 22034 3454
rect 21982 3378 22034 3390
rect 23998 3442 24050 3454
rect 23998 3378 24050 3390
rect 26462 3442 26514 3454
rect 26462 3378 26514 3390
rect 26798 3442 26850 3454
rect 26798 3378 26850 3390
rect 27134 3442 27186 3454
rect 27134 3378 27186 3390
rect 28590 3442 28642 3454
rect 28590 3378 28642 3390
rect 29262 3442 29314 3454
rect 29262 3378 29314 3390
rect 29598 3442 29650 3454
rect 29598 3378 29650 3390
rect 29934 3442 29986 3454
rect 29934 3378 29986 3390
rect 30270 3442 30322 3454
rect 30270 3378 30322 3390
rect 30942 3442 30994 3454
rect 30942 3378 30994 3390
rect 32174 3442 32226 3454
rect 48302 3442 48354 3454
rect 33618 3390 33630 3442
rect 33682 3390 33694 3442
rect 35298 3390 35310 3442
rect 35362 3390 35374 3442
rect 36642 3390 36654 3442
rect 36706 3390 36718 3442
rect 37650 3390 37662 3442
rect 37714 3390 37726 3442
rect 41458 3390 41470 3442
rect 41522 3390 41534 3442
rect 42466 3390 42478 3442
rect 42530 3390 42542 3442
rect 44370 3390 44382 3442
rect 44434 3390 44446 3442
rect 45154 3390 45166 3442
rect 45218 3390 45230 3442
rect 32174 3378 32226 3390
rect 48302 3378 48354 3390
rect 48974 3442 49026 3454
rect 48974 3378 49026 3390
rect 49646 3442 49698 3454
rect 49646 3378 49698 3390
rect 50318 3442 50370 3454
rect 50318 3378 50370 3390
rect 51214 3442 51266 3454
rect 77310 3442 77362 3454
rect 52098 3390 52110 3442
rect 52162 3390 52174 3442
rect 52770 3390 52782 3442
rect 52834 3390 52846 3442
rect 53442 3390 53454 3442
rect 53506 3390 53518 3442
rect 78194 3390 78206 3442
rect 78258 3390 78270 3442
rect 51214 3378 51266 3390
rect 77310 3378 77362 3390
rect 8766 3330 8818 3342
rect 8766 3266 8818 3278
rect 14366 3330 14418 3342
rect 14366 3266 14418 3278
rect 18846 3330 18898 3342
rect 25902 3330 25954 3342
rect 22642 3278 22654 3330
rect 22706 3278 22718 3330
rect 18846 3266 18898 3278
rect 25902 3266 25954 3278
rect 27806 3330 27858 3342
rect 27806 3266 27858 3278
rect 28926 3330 28978 3342
rect 28926 3266 28978 3278
rect 31614 3330 31666 3342
rect 31614 3266 31666 3278
rect 1344 3162 78624 3196
rect 1344 3110 19838 3162
rect 19890 3110 19942 3162
rect 19994 3110 20046 3162
rect 20098 3110 50558 3162
rect 50610 3110 50662 3162
rect 50714 3110 50766 3162
rect 50818 3110 78624 3162
rect 1344 3076 78624 3110
rect 7186 2942 7198 2994
rect 7250 2991 7262 2994
rect 9650 2991 9662 2994
rect 7250 2945 9662 2991
rect 7250 2942 7262 2945
rect 9650 2942 9662 2945
rect 9714 2942 9726 2994
rect 12226 2942 12238 2994
rect 12290 2991 12302 2994
rect 16370 2991 16382 2994
rect 12290 2945 16382 2991
rect 12290 2942 12302 2945
rect 16370 2942 16382 2945
rect 16434 2942 16446 2994
rect 29138 1374 29150 1426
rect 29202 1423 29214 1426
rect 29698 1423 29710 1426
rect 29202 1377 29710 1423
rect 29202 1374 29214 1377
rect 29698 1374 29710 1377
rect 29762 1374 29774 1426
<< via1 >>
rect 69022 77198 69074 77250
rect 70030 77198 70082 77250
rect 70254 77198 70306 77250
rect 42814 77086 42866 77138
rect 43598 77086 43650 77138
rect 50878 77086 50930 77138
rect 51774 77086 51826 77138
rect 52110 77086 52162 77138
rect 64318 77086 64370 77138
rect 65326 77086 65378 77138
rect 66334 77086 66386 77138
rect 67118 77086 67170 77138
rect 71038 77086 71090 77138
rect 72270 77086 72322 77138
rect 75182 77086 75234 77138
rect 75630 77086 75682 77138
rect 76414 77086 76466 77138
rect 37214 76974 37266 77026
rect 38110 76974 38162 77026
rect 43710 76974 43762 77026
rect 43934 76974 43986 77026
rect 44494 76974 44546 77026
rect 45502 76974 45554 77026
rect 46734 76974 46786 77026
rect 47518 76974 47570 77026
rect 48302 76974 48354 77026
rect 48862 76974 48914 77026
rect 50094 76974 50146 77026
rect 51550 76974 51602 77026
rect 53006 76974 53058 77026
rect 62302 76974 62354 77026
rect 63310 76974 63362 77026
rect 63646 76974 63698 77026
rect 64654 76974 64706 77026
rect 65662 76974 65714 77026
rect 66446 76974 66498 77026
rect 67678 76974 67730 77026
rect 68462 76974 68514 77026
rect 69022 76974 69074 77026
rect 70142 76974 70194 77026
rect 74398 76974 74450 77026
rect 74958 76974 75010 77026
rect 75742 76974 75794 77026
rect 19838 76806 19890 76858
rect 19942 76806 19994 76858
rect 20046 76806 20098 76858
rect 50558 76806 50610 76858
rect 50662 76806 50714 76858
rect 50766 76806 50818 76858
rect 4622 76638 4674 76690
rect 15374 76638 15426 76690
rect 21086 76638 21138 76690
rect 24894 76638 24946 76690
rect 25566 76638 25618 76690
rect 26238 76638 26290 76690
rect 26910 76638 26962 76690
rect 27582 76638 27634 76690
rect 28366 76638 28418 76690
rect 28926 76638 28978 76690
rect 29598 76638 29650 76690
rect 30270 76638 30322 76690
rect 30942 76638 30994 76690
rect 31502 76638 31554 76690
rect 32286 76638 32338 76690
rect 36878 76638 36930 76690
rect 38334 76638 38386 76690
rect 39230 76638 39282 76690
rect 40126 76638 40178 76690
rect 41022 76638 41074 76690
rect 42030 76638 42082 76690
rect 42366 76638 42418 76690
rect 43598 76638 43650 76690
rect 44494 76638 44546 76690
rect 48302 76638 48354 76690
rect 49198 76638 49250 76690
rect 50094 76638 50146 76690
rect 51214 76638 51266 76690
rect 52110 76638 52162 76690
rect 53006 76638 53058 76690
rect 53902 76638 53954 76690
rect 55134 76638 55186 76690
rect 59838 76638 59890 76690
rect 63310 76638 63362 76690
rect 63982 76638 64034 76690
rect 64654 76638 64706 76690
rect 65326 76638 65378 76690
rect 66446 76638 66498 76690
rect 67118 76638 67170 76690
rect 67790 76638 67842 76690
rect 68462 76638 68514 76690
rect 69358 76638 69410 76690
rect 70254 76638 70306 76690
rect 72270 76638 72322 76690
rect 76078 76638 76130 76690
rect 77310 76638 77362 76690
rect 4958 76526 5010 76578
rect 5518 76526 5570 76578
rect 19294 76526 19346 76578
rect 36206 76526 36258 76578
rect 45950 76526 46002 76578
rect 61742 76526 61794 76578
rect 62638 76526 62690 76578
rect 63646 76526 63698 76578
rect 64318 76526 64370 76578
rect 64990 76526 65042 76578
rect 65662 76526 65714 76578
rect 66782 76526 66834 76578
rect 67454 76526 67506 76578
rect 68126 76526 68178 76578
rect 69694 76526 69746 76578
rect 70590 76526 70642 76578
rect 70926 76526 70978 76578
rect 71262 76526 71314 76578
rect 71598 76526 71650 76578
rect 71934 76526 71986 76578
rect 72606 76526 72658 76578
rect 72942 76526 72994 76578
rect 74062 76526 74114 76578
rect 74734 76526 74786 76578
rect 75070 76526 75122 76578
rect 75406 76526 75458 76578
rect 75742 76526 75794 76578
rect 76414 76526 76466 76578
rect 78206 76526 78258 76578
rect 4286 76414 4338 76466
rect 5742 76414 5794 76466
rect 12462 76414 12514 76466
rect 16382 76414 16434 76466
rect 18062 76414 18114 76466
rect 23774 76414 23826 76466
rect 35086 76414 35138 76466
rect 36430 76414 36482 76466
rect 46734 76414 46786 76466
rect 47854 76414 47906 76466
rect 58270 76414 58322 76466
rect 58830 76414 58882 76466
rect 62078 76414 62130 76466
rect 62862 76414 62914 76466
rect 73166 76414 73218 76466
rect 74286 76414 74338 76466
rect 77870 76414 77922 76466
rect 13358 76302 13410 76354
rect 17166 76302 17218 76354
rect 21646 76302 21698 76354
rect 33406 76302 33458 76354
rect 37438 76302 37490 76354
rect 37886 76302 37938 76354
rect 38782 76302 38834 76354
rect 40686 76302 40738 76354
rect 41582 76302 41634 76354
rect 42926 76302 42978 76354
rect 44046 76302 44098 76354
rect 44942 76302 44994 76354
rect 45502 76302 45554 76354
rect 46286 76302 46338 76354
rect 47406 76302 47458 76354
rect 48862 76302 48914 76354
rect 49646 76302 49698 76354
rect 50542 76302 50594 76354
rect 51662 76302 51714 76354
rect 52558 76302 52610 76354
rect 53454 76302 53506 76354
rect 54462 76302 54514 76354
rect 55918 76302 55970 76354
rect 69022 76302 69074 76354
rect 76750 76302 76802 76354
rect 1934 76190 1986 76242
rect 11566 76190 11618 76242
rect 4478 76022 4530 76074
rect 4582 76022 4634 76074
rect 4686 76022 4738 76074
rect 35198 76022 35250 76074
rect 35302 76022 35354 76074
rect 35406 76022 35458 76074
rect 65918 76022 65970 76074
rect 66022 76022 66074 76074
rect 66126 76022 66178 76074
rect 11902 75854 11954 75906
rect 16830 75854 16882 75906
rect 21982 75854 22034 75906
rect 45838 75854 45890 75906
rect 46510 75854 46562 75906
rect 56702 75854 56754 75906
rect 63310 75854 63362 75906
rect 63758 75854 63810 75906
rect 1934 75742 1986 75794
rect 18622 75742 18674 75794
rect 32734 75742 32786 75794
rect 35198 75742 35250 75794
rect 37214 75742 37266 75794
rect 39454 75742 39506 75794
rect 41470 75742 41522 75794
rect 42478 75742 42530 75794
rect 43374 75742 43426 75794
rect 43934 75742 43986 75794
rect 44382 75742 44434 75794
rect 46062 75742 46114 75794
rect 46622 75742 46674 75794
rect 48078 75742 48130 75794
rect 48526 75742 48578 75794
rect 49086 75742 49138 75794
rect 49534 75742 49586 75794
rect 50766 75742 50818 75794
rect 51214 75742 51266 75794
rect 51774 75742 51826 75794
rect 52222 75742 52274 75794
rect 63758 75742 63810 75794
rect 64206 75742 64258 75794
rect 64990 75742 65042 75794
rect 65998 75742 66050 75794
rect 66446 75742 66498 75794
rect 67006 75742 67058 75794
rect 67566 75742 67618 75794
rect 68462 75742 68514 75794
rect 69134 75742 69186 75794
rect 70030 75742 70082 75794
rect 70702 75742 70754 75794
rect 71374 75742 71426 75794
rect 71934 75742 71986 75794
rect 72382 75742 72434 75794
rect 73390 75742 73442 75794
rect 73950 75742 74002 75794
rect 74510 75742 74562 75794
rect 75070 75742 75122 75794
rect 77758 75742 77810 75794
rect 4286 75630 4338 75682
rect 4958 75630 5010 75682
rect 12574 75630 12626 75682
rect 13582 75630 13634 75682
rect 14702 75630 14754 75682
rect 17838 75630 17890 75682
rect 20302 75630 20354 75682
rect 23886 75630 23938 75682
rect 24782 75630 24834 75682
rect 25230 75630 25282 75682
rect 32958 75630 33010 75682
rect 33518 75630 33570 75682
rect 33966 75630 34018 75682
rect 34414 75630 34466 75682
rect 34750 75630 34802 75682
rect 35646 75630 35698 75682
rect 36206 75630 36258 75682
rect 37438 75630 37490 75682
rect 37998 75630 38050 75682
rect 38334 75630 38386 75682
rect 38894 75630 38946 75682
rect 40910 75630 40962 75682
rect 41694 75630 41746 75682
rect 45054 75630 45106 75682
rect 47070 75630 47122 75682
rect 47630 75630 47682 75682
rect 49758 75630 49810 75682
rect 50318 75630 50370 75682
rect 52670 75630 52722 75682
rect 53230 75630 53282 75682
rect 53790 75630 53842 75682
rect 54350 75630 54402 75682
rect 54686 75630 54738 75682
rect 55246 75630 55298 75682
rect 55694 75630 55746 75682
rect 56142 75630 56194 75682
rect 59054 75630 59106 75682
rect 61742 75630 61794 75682
rect 63310 75630 63362 75682
rect 65214 75630 65266 75682
rect 72606 75630 72658 75682
rect 75406 75630 75458 75682
rect 76190 75630 76242 75682
rect 76862 75630 76914 75682
rect 4622 75518 4674 75570
rect 24222 75518 24274 75570
rect 45614 75518 45666 75570
rect 61182 75518 61234 75570
rect 62078 75518 62130 75570
rect 75630 75518 75682 75570
rect 76526 75518 76578 75570
rect 77198 75518 77250 75570
rect 78206 75518 78258 75570
rect 14254 75406 14306 75458
rect 42030 75406 42082 75458
rect 59390 75406 59442 75458
rect 59726 75406 59778 75458
rect 60510 75406 60562 75458
rect 60846 75406 60898 75458
rect 62414 75406 62466 75458
rect 62862 75406 62914 75458
rect 65550 75406 65602 75458
rect 72942 75406 72994 75458
rect 19838 75238 19890 75290
rect 19942 75238 19994 75290
rect 20046 75238 20098 75290
rect 50558 75238 50610 75290
rect 50662 75238 50714 75290
rect 50766 75238 50818 75290
rect 4622 75070 4674 75122
rect 12910 75070 12962 75122
rect 23102 75070 23154 75122
rect 23550 75070 23602 75122
rect 34638 75070 34690 75122
rect 35534 75070 35586 75122
rect 35982 75070 36034 75122
rect 36766 75070 36818 75122
rect 37662 75070 37714 75122
rect 46846 75070 46898 75122
rect 52782 75070 52834 75122
rect 53566 75070 53618 75122
rect 54462 75070 54514 75122
rect 55358 75070 55410 75122
rect 57598 75070 57650 75122
rect 61294 75070 61346 75122
rect 61742 75070 61794 75122
rect 62190 75070 62242 75122
rect 64654 75070 64706 75122
rect 74062 75070 74114 75122
rect 74510 75070 74562 75122
rect 74958 75070 75010 75122
rect 76862 75070 76914 75122
rect 78206 75070 78258 75122
rect 15262 74958 15314 75010
rect 75406 74958 75458 75010
rect 75630 74958 75682 75010
rect 75966 74958 76018 75010
rect 4174 74846 4226 74898
rect 4846 74846 4898 74898
rect 13470 74846 13522 74898
rect 16494 74846 16546 74898
rect 22766 74846 22818 74898
rect 60398 74846 60450 74898
rect 60846 74846 60898 74898
rect 77310 74846 77362 74898
rect 2158 74734 2210 74786
rect 17950 74734 18002 74786
rect 18286 74734 18338 74786
rect 19406 74734 19458 74786
rect 19854 74734 19906 74786
rect 20414 74734 20466 74786
rect 35086 74734 35138 74786
rect 38222 74734 38274 74786
rect 38782 74734 38834 74786
rect 58046 74734 58098 74786
rect 76414 74734 76466 74786
rect 77758 74734 77810 74786
rect 37438 74622 37490 74674
rect 38222 74622 38274 74674
rect 4478 74454 4530 74506
rect 4582 74454 4634 74506
rect 4686 74454 4738 74506
rect 35198 74454 35250 74506
rect 35302 74454 35354 74506
rect 35406 74454 35458 74506
rect 65918 74454 65970 74506
rect 66022 74454 66074 74506
rect 66126 74454 66178 74506
rect 15934 74286 15986 74338
rect 19182 74286 19234 74338
rect 76078 74286 76130 74338
rect 76414 74286 76466 74338
rect 1934 74174 1986 74226
rect 11230 74174 11282 74226
rect 58494 74174 58546 74226
rect 59166 74174 59218 74226
rect 59502 74174 59554 74226
rect 75742 74174 75794 74226
rect 76414 74174 76466 74226
rect 4286 74062 4338 74114
rect 4846 74062 4898 74114
rect 12686 74062 12738 74114
rect 17614 74062 17666 74114
rect 18174 74062 18226 74114
rect 75294 74062 75346 74114
rect 76974 74062 77026 74114
rect 77534 74062 77586 74114
rect 78094 74062 78146 74114
rect 4622 73950 4674 74002
rect 14030 73950 14082 74002
rect 14366 73950 14418 74002
rect 22990 73950 23042 74002
rect 77870 73950 77922 74002
rect 19838 73670 19890 73722
rect 19942 73670 19994 73722
rect 20046 73670 20098 73722
rect 50558 73670 50610 73722
rect 50662 73670 50714 73722
rect 50766 73670 50818 73722
rect 76190 73502 76242 73554
rect 76638 73502 76690 73554
rect 77198 73502 77250 73554
rect 77646 73502 77698 73554
rect 78206 73502 78258 73554
rect 4622 73390 4674 73442
rect 12126 73390 12178 73442
rect 77870 73390 77922 73442
rect 4286 73278 4338 73330
rect 4846 73278 4898 73330
rect 13918 73278 13970 73330
rect 16382 73278 16434 73330
rect 14590 73166 14642 73218
rect 18062 73166 18114 73218
rect 1934 73054 1986 73106
rect 4478 72886 4530 72938
rect 4582 72886 4634 72938
rect 4686 72886 4738 72938
rect 35198 72886 35250 72938
rect 35302 72886 35354 72938
rect 35406 72886 35458 72938
rect 65918 72886 65970 72938
rect 66022 72886 66074 72938
rect 66126 72886 66178 72938
rect 1934 72606 1986 72658
rect 77198 72606 77250 72658
rect 3838 72494 3890 72546
rect 77646 72382 77698 72434
rect 78206 72382 78258 72434
rect 14142 72270 14194 72322
rect 77870 72270 77922 72322
rect 19838 72102 19890 72154
rect 19942 72102 19994 72154
rect 20046 72102 20098 72154
rect 50558 72102 50610 72154
rect 50662 72102 50714 72154
rect 50766 72102 50818 72154
rect 3166 71934 3218 71986
rect 3502 71934 3554 71986
rect 4174 71934 4226 71986
rect 2494 71822 2546 71874
rect 3838 71822 3890 71874
rect 4510 71822 4562 71874
rect 77870 71822 77922 71874
rect 2158 71710 2210 71762
rect 2942 71710 2994 71762
rect 78206 71710 78258 71762
rect 1934 71598 1986 71650
rect 77646 71598 77698 71650
rect 4478 71318 4530 71370
rect 4582 71318 4634 71370
rect 4686 71318 4738 71370
rect 35198 71318 35250 71370
rect 35302 71318 35354 71370
rect 35406 71318 35458 71370
rect 65918 71318 65970 71370
rect 66022 71318 66074 71370
rect 66126 71318 66178 71370
rect 1934 71038 1986 71090
rect 3950 70926 4002 70978
rect 77646 70926 77698 70978
rect 77422 70702 77474 70754
rect 78206 70702 78258 70754
rect 19838 70534 19890 70586
rect 19942 70534 19994 70586
rect 20046 70534 20098 70586
rect 50558 70534 50610 70586
rect 50662 70534 50714 70586
rect 50766 70534 50818 70586
rect 3838 70142 3890 70194
rect 1934 69918 1986 69970
rect 4478 69750 4530 69802
rect 4582 69750 4634 69802
rect 4686 69750 4738 69802
rect 35198 69750 35250 69802
rect 35302 69750 35354 69802
rect 35406 69750 35458 69802
rect 65918 69750 65970 69802
rect 66022 69750 66074 69802
rect 66126 69750 66178 69802
rect 2942 69358 2994 69410
rect 2382 69246 2434 69298
rect 2718 69246 2770 69298
rect 2046 69134 2098 69186
rect 77646 69134 77698 69186
rect 77870 69134 77922 69186
rect 78206 69134 78258 69186
rect 19838 68966 19890 69018
rect 19942 68966 19994 69018
rect 20046 68966 20098 69018
rect 50558 68966 50610 69018
rect 50662 68966 50714 69018
rect 50766 68966 50818 69018
rect 2046 68574 2098 68626
rect 77422 68574 77474 68626
rect 78206 68574 78258 68626
rect 77646 68462 77698 68514
rect 2718 68350 2770 68402
rect 4478 68182 4530 68234
rect 4582 68182 4634 68234
rect 4686 68182 4738 68234
rect 35198 68182 35250 68234
rect 35302 68182 35354 68234
rect 35406 68182 35458 68234
rect 65918 68182 65970 68234
rect 66022 68182 66074 68234
rect 66126 68182 66178 68234
rect 1934 67902 1986 67954
rect 3838 67790 3890 67842
rect 19838 67398 19890 67450
rect 19942 67398 19994 67450
rect 20046 67398 20098 67450
rect 50558 67398 50610 67450
rect 50662 67398 50714 67450
rect 50766 67398 50818 67450
rect 3390 67230 3442 67282
rect 2046 67118 2098 67170
rect 2382 67118 2434 67170
rect 3054 67118 3106 67170
rect 77870 67118 77922 67170
rect 2718 67006 2770 67058
rect 3614 67006 3666 67058
rect 78206 67006 78258 67058
rect 77646 66894 77698 66946
rect 4478 66614 4530 66666
rect 4582 66614 4634 66666
rect 4686 66614 4738 66666
rect 35198 66614 35250 66666
rect 35302 66614 35354 66666
rect 35406 66614 35458 66666
rect 65918 66614 65970 66666
rect 66022 66614 66074 66666
rect 66126 66614 66178 66666
rect 2046 66222 2098 66274
rect 2718 65998 2770 66050
rect 77646 65998 77698 66050
rect 77870 65998 77922 66050
rect 78206 65998 78258 66050
rect 19838 65830 19890 65882
rect 19942 65830 19994 65882
rect 20046 65830 20098 65882
rect 50558 65830 50610 65882
rect 50662 65830 50714 65882
rect 50766 65830 50818 65882
rect 4286 65438 4338 65490
rect 1934 65214 1986 65266
rect 4478 65046 4530 65098
rect 4582 65046 4634 65098
rect 4686 65046 4738 65098
rect 35198 65046 35250 65098
rect 35302 65046 35354 65098
rect 35406 65046 35458 65098
rect 65918 65046 65970 65098
rect 66022 65046 66074 65098
rect 66126 65046 66178 65098
rect 1934 64766 1986 64818
rect 3838 64654 3890 64706
rect 77646 64654 77698 64706
rect 4622 64542 4674 64594
rect 4958 64542 5010 64594
rect 77422 64542 77474 64594
rect 78206 64542 78258 64594
rect 19838 64262 19890 64314
rect 19942 64262 19994 64314
rect 20046 64262 20098 64314
rect 50558 64262 50610 64314
rect 50662 64262 50714 64314
rect 50766 64262 50818 64314
rect 3838 64094 3890 64146
rect 2494 63982 2546 64034
rect 3166 63982 3218 64034
rect 2270 63870 2322 63922
rect 2942 63870 2994 63922
rect 3614 63870 3666 63922
rect 77422 63870 77474 63922
rect 77646 63870 77698 63922
rect 78206 63870 78258 63922
rect 4478 63478 4530 63530
rect 4582 63478 4634 63530
rect 4686 63478 4738 63530
rect 35198 63478 35250 63530
rect 35302 63478 35354 63530
rect 35406 63478 35458 63530
rect 65918 63478 65970 63530
rect 66022 63478 66074 63530
rect 66126 63478 66178 63530
rect 1934 63198 1986 63250
rect 3838 63086 3890 63138
rect 78206 62974 78258 63026
rect 77646 62862 77698 62914
rect 77870 62862 77922 62914
rect 19838 62694 19890 62746
rect 19942 62694 19994 62746
rect 20046 62694 20098 62746
rect 50558 62694 50610 62746
rect 50662 62694 50714 62746
rect 50766 62694 50818 62746
rect 3838 62302 3890 62354
rect 1934 62078 1986 62130
rect 4478 61910 4530 61962
rect 4582 61910 4634 61962
rect 4686 61910 4738 61962
rect 35198 61910 35250 61962
rect 35302 61910 35354 61962
rect 35406 61910 35458 61962
rect 65918 61910 65970 61962
rect 66022 61910 66074 61962
rect 66126 61910 66178 61962
rect 2270 61518 2322 61570
rect 3614 61518 3666 61570
rect 77646 61518 77698 61570
rect 2718 61406 2770 61458
rect 3054 61406 3106 61458
rect 3390 61406 3442 61458
rect 2046 61294 2098 61346
rect 4286 61294 4338 61346
rect 77422 61294 77474 61346
rect 78206 61294 78258 61346
rect 19838 61126 19890 61178
rect 19942 61126 19994 61178
rect 20046 61126 20098 61178
rect 50558 61126 50610 61178
rect 50662 61126 50714 61178
rect 50766 61126 50818 61178
rect 77870 60846 77922 60898
rect 2046 60734 2098 60786
rect 77646 60734 77698 60786
rect 78206 60734 78258 60786
rect 2718 60510 2770 60562
rect 4478 60342 4530 60394
rect 4582 60342 4634 60394
rect 4686 60342 4738 60394
rect 35198 60342 35250 60394
rect 35302 60342 35354 60394
rect 35406 60342 35458 60394
rect 65918 60342 65970 60394
rect 66022 60342 66074 60394
rect 66126 60342 66178 60394
rect 1934 60062 1986 60114
rect 3838 59950 3890 60002
rect 19838 59558 19890 59610
rect 19942 59558 19994 59610
rect 20046 59558 20098 59610
rect 50558 59558 50610 59610
rect 50662 59558 50714 59610
rect 50766 59558 50818 59610
rect 2718 59390 2770 59442
rect 2046 59278 2098 59330
rect 2382 59166 2434 59218
rect 2942 59166 2994 59218
rect 3502 59166 3554 59218
rect 78206 59166 78258 59218
rect 77422 59054 77474 59106
rect 77646 59054 77698 59106
rect 4478 58774 4530 58826
rect 4582 58774 4634 58826
rect 4686 58774 4738 58826
rect 35198 58774 35250 58826
rect 35302 58774 35354 58826
rect 35406 58774 35458 58826
rect 65918 58774 65970 58826
rect 66022 58774 66074 58826
rect 66126 58774 66178 58826
rect 2046 58382 2098 58434
rect 2718 58158 2770 58210
rect 77646 58158 77698 58210
rect 77870 58158 77922 58210
rect 78206 58158 78258 58210
rect 19838 57990 19890 58042
rect 19942 57990 19994 58042
rect 20046 57990 20098 58042
rect 50558 57990 50610 58042
rect 50662 57990 50714 58042
rect 50766 57990 50818 58042
rect 4286 57598 4338 57650
rect 1934 57374 1986 57426
rect 4478 57206 4530 57258
rect 4582 57206 4634 57258
rect 4686 57206 4738 57258
rect 35198 57206 35250 57258
rect 35302 57206 35354 57258
rect 35406 57206 35458 57258
rect 65918 57206 65970 57258
rect 66022 57206 66074 57258
rect 66126 57206 66178 57258
rect 1934 56926 1986 56978
rect 3838 56814 3890 56866
rect 4846 56814 4898 56866
rect 4622 56702 4674 56754
rect 77646 56702 77698 56754
rect 78206 56702 78258 56754
rect 77870 56590 77922 56642
rect 19838 56422 19890 56474
rect 19942 56422 19994 56474
rect 20046 56422 20098 56474
rect 50558 56422 50610 56474
rect 50662 56422 50714 56474
rect 50766 56422 50818 56474
rect 2718 56254 2770 56306
rect 3726 56254 3778 56306
rect 2046 56142 2098 56194
rect 2382 56142 2434 56194
rect 3390 56142 3442 56194
rect 77870 56142 77922 56194
rect 2942 56030 2994 56082
rect 78206 56030 78258 56082
rect 77646 55918 77698 55970
rect 4478 55638 4530 55690
rect 4582 55638 4634 55690
rect 4686 55638 4738 55690
rect 35198 55638 35250 55690
rect 35302 55638 35354 55690
rect 35406 55638 35458 55690
rect 65918 55638 65970 55690
rect 66022 55638 66074 55690
rect 66126 55638 66178 55690
rect 2046 55246 2098 55298
rect 78206 55134 78258 55186
rect 2718 55022 2770 55074
rect 77646 55022 77698 55074
rect 77870 55022 77922 55074
rect 19838 54854 19890 54906
rect 19942 54854 19994 54906
rect 20046 54854 20098 54906
rect 50558 54854 50610 54906
rect 50662 54854 50714 54906
rect 50766 54854 50818 54906
rect 3838 54462 3890 54514
rect 1934 54238 1986 54290
rect 4478 54070 4530 54122
rect 4582 54070 4634 54122
rect 4686 54070 4738 54122
rect 35198 54070 35250 54122
rect 35302 54070 35354 54122
rect 35406 54070 35458 54122
rect 65918 54070 65970 54122
rect 66022 54070 66074 54122
rect 66126 54070 66178 54122
rect 2942 53678 2994 53730
rect 2158 53566 2210 53618
rect 3166 53566 3218 53618
rect 3502 53566 3554 53618
rect 3838 53566 3890 53618
rect 77870 53566 77922 53618
rect 78206 53566 78258 53618
rect 1934 53454 1986 53506
rect 2494 53454 2546 53506
rect 77646 53454 77698 53506
rect 19838 53286 19890 53338
rect 19942 53286 19994 53338
rect 20046 53286 20098 53338
rect 50558 53286 50610 53338
rect 50662 53286 50714 53338
rect 50766 53286 50818 53338
rect 77870 53006 77922 53058
rect 3950 52894 4002 52946
rect 78206 52894 78258 52946
rect 77646 52782 77698 52834
rect 1934 52670 1986 52722
rect 4478 52502 4530 52554
rect 4582 52502 4634 52554
rect 4686 52502 4738 52554
rect 35198 52502 35250 52554
rect 35302 52502 35354 52554
rect 35406 52502 35458 52554
rect 65918 52502 65970 52554
rect 66022 52502 66074 52554
rect 66126 52502 66178 52554
rect 1934 52222 1986 52274
rect 3838 52110 3890 52162
rect 19838 51718 19890 51770
rect 19942 51718 19994 51770
rect 20046 51718 20098 51770
rect 50558 51718 50610 51770
rect 50662 51718 50714 51770
rect 50766 51718 50818 51770
rect 2494 51550 2546 51602
rect 3502 51550 3554 51602
rect 2830 51438 2882 51490
rect 3838 51438 3890 51490
rect 77870 51438 77922 51490
rect 2270 51326 2322 51378
rect 3166 51326 3218 51378
rect 78206 51326 78258 51378
rect 77646 51214 77698 51266
rect 4478 50934 4530 50986
rect 4582 50934 4634 50986
rect 4686 50934 4738 50986
rect 35198 50934 35250 50986
rect 35302 50934 35354 50986
rect 35406 50934 35458 50986
rect 65918 50934 65970 50986
rect 66022 50934 66074 50986
rect 66126 50934 66178 50986
rect 1934 50654 1986 50706
rect 3838 50542 3890 50594
rect 77646 50430 77698 50482
rect 78206 50430 78258 50482
rect 77870 50318 77922 50370
rect 19838 50150 19890 50202
rect 19942 50150 19994 50202
rect 20046 50150 20098 50202
rect 50558 50150 50610 50202
rect 50662 50150 50714 50202
rect 50766 50150 50818 50202
rect 3838 49758 3890 49810
rect 1934 49534 1986 49586
rect 4478 49366 4530 49418
rect 4582 49366 4634 49418
rect 4686 49366 4738 49418
rect 35198 49366 35250 49418
rect 35302 49366 35354 49418
rect 35406 49366 35458 49418
rect 65918 49366 65970 49418
rect 66022 49366 66074 49418
rect 66126 49366 66178 49418
rect 1934 49086 1986 49138
rect 3838 48974 3890 49026
rect 77646 48862 77698 48914
rect 78206 48862 78258 48914
rect 77870 48750 77922 48802
rect 19838 48582 19890 48634
rect 19942 48582 19994 48634
rect 20046 48582 20098 48634
rect 50558 48582 50610 48634
rect 50662 48582 50714 48634
rect 50766 48582 50818 48634
rect 2718 48414 2770 48466
rect 3390 48414 3442 48466
rect 2046 48302 2098 48354
rect 77870 48302 77922 48354
rect 2382 48190 2434 48242
rect 2942 48190 2994 48242
rect 3614 48190 3666 48242
rect 78206 48190 78258 48242
rect 77646 48078 77698 48130
rect 4478 47798 4530 47850
rect 4582 47798 4634 47850
rect 4686 47798 4738 47850
rect 35198 47798 35250 47850
rect 35302 47798 35354 47850
rect 35406 47798 35458 47850
rect 65918 47798 65970 47850
rect 66022 47798 66074 47850
rect 66126 47798 66178 47850
rect 2046 47406 2098 47458
rect 77646 47294 77698 47346
rect 78206 47294 78258 47346
rect 2718 47182 2770 47234
rect 77870 47182 77922 47234
rect 19838 47014 19890 47066
rect 19942 47014 19994 47066
rect 20046 47014 20098 47066
rect 50558 47014 50610 47066
rect 50662 47014 50714 47066
rect 50766 47014 50818 47066
rect 3838 46622 3890 46674
rect 1934 46398 1986 46450
rect 4478 46230 4530 46282
rect 4582 46230 4634 46282
rect 4686 46230 4738 46282
rect 35198 46230 35250 46282
rect 35302 46230 35354 46282
rect 35406 46230 35458 46282
rect 65918 46230 65970 46282
rect 66022 46230 66074 46282
rect 66126 46230 66178 46282
rect 2382 45838 2434 45890
rect 2830 45838 2882 45890
rect 3614 45838 3666 45890
rect 3054 45726 3106 45778
rect 3390 45726 3442 45778
rect 4286 45726 4338 45778
rect 78206 45726 78258 45778
rect 2046 45614 2098 45666
rect 77646 45614 77698 45666
rect 77870 45614 77922 45666
rect 19838 45446 19890 45498
rect 19942 45446 19994 45498
rect 20046 45446 20098 45498
rect 50558 45446 50610 45498
rect 50662 45446 50714 45498
rect 50766 45446 50818 45498
rect 77870 45166 77922 45218
rect 2046 45054 2098 45106
rect 78206 45054 78258 45106
rect 77646 44942 77698 44994
rect 2718 44830 2770 44882
rect 4478 44662 4530 44714
rect 4582 44662 4634 44714
rect 4686 44662 4738 44714
rect 35198 44662 35250 44714
rect 35302 44662 35354 44714
rect 35406 44662 35458 44714
rect 65918 44662 65970 44714
rect 66022 44662 66074 44714
rect 66126 44662 66178 44714
rect 2046 44270 2098 44322
rect 2718 44046 2770 44098
rect 77982 44046 78034 44098
rect 19838 43878 19890 43930
rect 19942 43878 19994 43930
rect 20046 43878 20098 43930
rect 50558 43878 50610 43930
rect 50662 43878 50714 43930
rect 50766 43878 50818 43930
rect 2046 43710 2098 43762
rect 2718 43598 2770 43650
rect 77870 43598 77922 43650
rect 2270 43486 2322 43538
rect 2942 43486 2994 43538
rect 77086 43486 77138 43538
rect 78206 43486 78258 43538
rect 77646 43374 77698 43426
rect 4478 43094 4530 43146
rect 4582 43094 4634 43146
rect 4686 43094 4738 43146
rect 35198 43094 35250 43146
rect 35302 43094 35354 43146
rect 35406 43094 35458 43146
rect 65918 43094 65970 43146
rect 66022 43094 66074 43146
rect 66126 43094 66178 43146
rect 1934 42814 1986 42866
rect 55806 42814 55858 42866
rect 56702 42814 56754 42866
rect 57598 42814 57650 42866
rect 58494 42814 58546 42866
rect 62414 42814 62466 42866
rect 75294 42814 75346 42866
rect 76526 42814 76578 42866
rect 3838 42702 3890 42754
rect 57150 42702 57202 42754
rect 58046 42702 58098 42754
rect 76750 42702 76802 42754
rect 77086 42702 77138 42754
rect 77422 42590 77474 42642
rect 77758 42590 77810 42642
rect 55246 42478 55298 42530
rect 56142 42478 56194 42530
rect 77086 42478 77138 42530
rect 78094 42478 78146 42530
rect 19838 42310 19890 42362
rect 19942 42310 19994 42362
rect 20046 42310 20098 42362
rect 50558 42310 50610 42362
rect 50662 42310 50714 42362
rect 50766 42310 50818 42362
rect 55022 42142 55074 42194
rect 57150 42142 57202 42194
rect 58046 42142 58098 42194
rect 62862 42030 62914 42082
rect 75294 42030 75346 42082
rect 3838 41918 3890 41970
rect 4734 41918 4786 41970
rect 61630 41918 61682 41970
rect 62750 41918 62802 41970
rect 63310 41918 63362 41970
rect 64542 41918 64594 41970
rect 73950 41918 74002 41970
rect 74958 41918 75010 41970
rect 75630 41918 75682 41970
rect 55582 41806 55634 41858
rect 56142 41806 56194 41858
rect 56590 41806 56642 41858
rect 57486 41806 57538 41858
rect 62190 41806 62242 41858
rect 63086 41806 63138 41858
rect 63646 41806 63698 41858
rect 70590 41806 70642 41858
rect 71038 41806 71090 41858
rect 74734 41806 74786 41858
rect 77982 41806 78034 41858
rect 1934 41694 1986 41746
rect 55358 41694 55410 41746
rect 55806 41694 55858 41746
rect 56030 41694 56082 41746
rect 56814 41694 56866 41746
rect 57710 41694 57762 41746
rect 4478 41526 4530 41578
rect 4582 41526 4634 41578
rect 4686 41526 4738 41578
rect 35198 41526 35250 41578
rect 35302 41526 35354 41578
rect 35406 41526 35458 41578
rect 65918 41526 65970 41578
rect 66022 41526 66074 41578
rect 66126 41526 66178 41578
rect 55470 41358 55522 41410
rect 55806 41358 55858 41410
rect 71374 41358 71426 41410
rect 74622 41358 74674 41410
rect 75518 41358 75570 41410
rect 1934 41246 1986 41298
rect 4734 41246 4786 41298
rect 57150 41246 57202 41298
rect 61518 41246 61570 41298
rect 65326 41246 65378 41298
rect 70814 41246 70866 41298
rect 71486 41246 71538 41298
rect 71934 41246 71986 41298
rect 72046 41246 72098 41298
rect 75182 41246 75234 41298
rect 78094 41246 78146 41298
rect 4062 41134 4114 41186
rect 55246 41134 55298 41186
rect 60510 41134 60562 41186
rect 61854 41134 61906 41186
rect 62190 41134 62242 41186
rect 62414 41134 62466 41186
rect 62974 41134 63026 41186
rect 63310 41134 63362 41186
rect 64430 41134 64482 41186
rect 64878 41134 64930 41186
rect 65662 41134 65714 41186
rect 66782 41134 66834 41186
rect 71710 41134 71762 41186
rect 73502 41134 73554 41186
rect 74062 41134 74114 41186
rect 74286 41134 74338 41186
rect 74958 41134 75010 41186
rect 76414 41134 76466 41186
rect 76750 41134 76802 41186
rect 77422 41134 77474 41186
rect 58382 41022 58434 41074
rect 58718 41022 58770 41074
rect 61070 41022 61122 41074
rect 63422 41022 63474 41074
rect 65774 41022 65826 41074
rect 69582 41022 69634 41074
rect 73166 41022 73218 41074
rect 73726 41022 73778 41074
rect 76190 41022 76242 41074
rect 77086 41022 77138 41074
rect 77646 41022 77698 41074
rect 54910 40910 54962 40962
rect 56254 40910 56306 40962
rect 62078 40910 62130 40962
rect 62974 40910 63026 40962
rect 66670 40910 66722 40962
rect 69022 40910 69074 40962
rect 69246 40910 69298 40962
rect 70030 40910 70082 40962
rect 70366 40910 70418 40962
rect 73390 40910 73442 40962
rect 76638 40910 76690 40962
rect 77198 40910 77250 40962
rect 19838 40742 19890 40794
rect 19942 40742 19994 40794
rect 20046 40742 20098 40794
rect 50558 40742 50610 40794
rect 50662 40742 50714 40794
rect 50766 40742 50818 40794
rect 2270 40574 2322 40626
rect 63534 40574 63586 40626
rect 67454 40574 67506 40626
rect 68350 40574 68402 40626
rect 69582 40574 69634 40626
rect 70254 40574 70306 40626
rect 74622 40574 74674 40626
rect 4062 40462 4114 40514
rect 4510 40462 4562 40514
rect 59838 40462 59890 40514
rect 61518 40462 61570 40514
rect 62526 40462 62578 40514
rect 65102 40462 65154 40514
rect 66334 40462 66386 40514
rect 67902 40462 67954 40514
rect 75294 40462 75346 40514
rect 76526 40462 76578 40514
rect 1710 40350 1762 40402
rect 2606 40350 2658 40402
rect 3166 40350 3218 40402
rect 3502 40350 3554 40402
rect 4958 40350 5010 40402
rect 5406 40350 5458 40402
rect 60062 40350 60114 40402
rect 60734 40350 60786 40402
rect 61070 40350 61122 40402
rect 62190 40350 62242 40402
rect 63086 40350 63138 40402
rect 63422 40350 63474 40402
rect 64430 40350 64482 40402
rect 65550 40350 65602 40402
rect 65886 40350 65938 40402
rect 66782 40350 66834 40402
rect 68574 40350 68626 40402
rect 69134 40350 69186 40402
rect 73166 40350 73218 40402
rect 73614 40350 73666 40402
rect 74286 40350 74338 40402
rect 75070 40350 75122 40402
rect 78206 40350 78258 40402
rect 60174 40238 60226 40290
rect 61406 40238 61458 40290
rect 64878 40238 64930 40290
rect 66446 40238 66498 40290
rect 70702 40238 70754 40290
rect 73390 40238 73442 40290
rect 72942 40126 72994 40178
rect 4478 39958 4530 40010
rect 4582 39958 4634 40010
rect 4686 39958 4738 40010
rect 35198 39958 35250 40010
rect 35302 39958 35354 40010
rect 35406 39958 35458 40010
rect 65918 39958 65970 40010
rect 66022 39958 66074 40010
rect 66126 39958 66178 40010
rect 1934 39678 1986 39730
rect 62302 39678 62354 39730
rect 62638 39678 62690 39730
rect 63198 39678 63250 39730
rect 66222 39678 66274 39730
rect 67118 39678 67170 39730
rect 69022 39678 69074 39730
rect 71374 39678 71426 39730
rect 71822 39678 71874 39730
rect 73166 39678 73218 39730
rect 74622 39678 74674 39730
rect 76750 39678 76802 39730
rect 77982 39678 78034 39730
rect 3838 39566 3890 39618
rect 4734 39566 4786 39618
rect 60734 39566 60786 39618
rect 61070 39566 61122 39618
rect 65662 39566 65714 39618
rect 66110 39566 66162 39618
rect 68574 39566 68626 39618
rect 69582 39566 69634 39618
rect 70254 39566 70306 39618
rect 70702 39566 70754 39618
rect 72830 39566 72882 39618
rect 72942 39566 72994 39618
rect 74958 39566 75010 39618
rect 75406 39566 75458 39618
rect 75630 39566 75682 39618
rect 76526 39566 76578 39618
rect 77310 39566 77362 39618
rect 61182 39454 61234 39506
rect 63982 39454 64034 39506
rect 66558 39454 66610 39506
rect 69246 39454 69298 39506
rect 70926 39454 70978 39506
rect 73278 39454 73330 39506
rect 73838 39454 73890 39506
rect 74174 39454 74226 39506
rect 76190 39454 76242 39506
rect 77870 39454 77922 39506
rect 78094 39454 78146 39506
rect 60622 39342 60674 39394
rect 63646 39342 63698 39394
rect 64318 39342 64370 39394
rect 67566 39342 67618 39394
rect 70478 39342 70530 39394
rect 72382 39342 72434 39394
rect 75294 39342 75346 39394
rect 19838 39174 19890 39226
rect 19942 39174 19994 39226
rect 20046 39174 20098 39226
rect 50558 39174 50610 39226
rect 50662 39174 50714 39226
rect 50766 39174 50818 39226
rect 41134 39006 41186 39058
rect 42926 39006 42978 39058
rect 43262 39006 43314 39058
rect 60958 39006 61010 39058
rect 63310 39006 63362 39058
rect 72830 39006 72882 39058
rect 75966 39006 76018 39058
rect 78206 39006 78258 39058
rect 41246 38894 41298 38946
rect 42254 38894 42306 38946
rect 42702 38894 42754 38946
rect 67006 38894 67058 38946
rect 67678 38894 67730 38946
rect 69918 38894 69970 38946
rect 71374 38894 71426 38946
rect 72494 38894 72546 38946
rect 73166 38894 73218 38946
rect 73502 38894 73554 38946
rect 74510 38894 74562 38946
rect 75406 38894 75458 38946
rect 76526 38894 76578 38946
rect 77534 38894 77586 38946
rect 2046 38782 2098 38834
rect 40910 38782 40962 38834
rect 41694 38782 41746 38834
rect 42590 38782 42642 38834
rect 43710 38782 43762 38834
rect 63534 38782 63586 38834
rect 65214 38782 65266 38834
rect 65774 38782 65826 38834
rect 66110 38782 66162 38834
rect 67230 38782 67282 38834
rect 68126 38782 68178 38834
rect 68574 38782 68626 38834
rect 69022 38782 69074 38834
rect 69582 38782 69634 38834
rect 70366 38782 70418 38834
rect 70702 38782 70754 38834
rect 70926 38782 70978 38834
rect 71598 38782 71650 38834
rect 74174 38782 74226 38834
rect 74734 38782 74786 38834
rect 75070 38782 75122 38834
rect 76302 38782 76354 38834
rect 76974 38782 77026 38834
rect 77086 38782 77138 38834
rect 77646 38782 77698 38834
rect 3390 38670 3442 38722
rect 41582 38670 41634 38722
rect 62974 38670 63026 38722
rect 66558 38670 66610 38722
rect 67678 38670 67730 38722
rect 69470 38670 69522 38722
rect 70590 38670 70642 38722
rect 74958 38670 75010 38722
rect 76750 38670 76802 38722
rect 77310 38670 77362 38722
rect 4478 38390 4530 38442
rect 4582 38390 4634 38442
rect 4686 38390 4738 38442
rect 35198 38390 35250 38442
rect 35302 38390 35354 38442
rect 35406 38390 35458 38442
rect 65918 38390 65970 38442
rect 66022 38390 66074 38442
rect 66126 38390 66178 38442
rect 72718 38222 72770 38274
rect 73278 38222 73330 38274
rect 77310 38222 77362 38274
rect 2046 38110 2098 38162
rect 2942 38110 2994 38162
rect 41470 38110 41522 38162
rect 67342 38110 67394 38162
rect 69918 38110 69970 38162
rect 72158 38110 72210 38162
rect 72606 38110 72658 38162
rect 75742 38110 75794 38162
rect 76414 38110 76466 38162
rect 77982 38110 78034 38162
rect 2494 37998 2546 38050
rect 66110 37998 66162 38050
rect 66558 37998 66610 38050
rect 68350 37998 68402 38050
rect 69358 37998 69410 38050
rect 70254 37998 70306 38050
rect 70590 37998 70642 38050
rect 70814 37998 70866 38050
rect 71150 37998 71202 38050
rect 71374 37998 71426 38050
rect 73054 37998 73106 38050
rect 74510 37998 74562 38050
rect 74846 37998 74898 38050
rect 75070 37998 75122 38050
rect 77198 37998 77250 38050
rect 77534 37998 77586 38050
rect 69246 37886 69298 37938
rect 71710 37886 71762 37938
rect 73838 37886 73890 37938
rect 74174 37886 74226 37938
rect 76190 37886 76242 37938
rect 67790 37774 67842 37826
rect 68574 37774 68626 37826
rect 70366 37774 70418 37826
rect 71598 37774 71650 37826
rect 73502 37774 73554 37826
rect 74622 37774 74674 37826
rect 76414 37774 76466 37826
rect 19838 37606 19890 37658
rect 19942 37606 19994 37658
rect 20046 37606 20098 37658
rect 50558 37606 50610 37658
rect 50662 37606 50714 37658
rect 50766 37606 50818 37658
rect 68462 37438 68514 37490
rect 69470 37438 69522 37490
rect 69806 37438 69858 37490
rect 70814 37438 70866 37490
rect 71150 37438 71202 37490
rect 71486 37438 71538 37490
rect 76414 37438 76466 37490
rect 2046 37326 2098 37378
rect 72270 37326 72322 37378
rect 72830 37326 72882 37378
rect 73726 37326 73778 37378
rect 74062 37326 74114 37378
rect 75630 37326 75682 37378
rect 76190 37326 76242 37378
rect 1710 37214 1762 37266
rect 68686 37214 68738 37266
rect 69134 37214 69186 37266
rect 70030 37214 70082 37266
rect 70590 37214 70642 37266
rect 72494 37214 72546 37266
rect 73054 37214 73106 37266
rect 73390 37214 73442 37266
rect 74286 37214 74338 37266
rect 74622 37214 74674 37266
rect 75070 37214 75122 37266
rect 75406 37214 75458 37266
rect 76078 37214 76130 37266
rect 76526 37214 76578 37266
rect 77310 37214 77362 37266
rect 77870 37214 77922 37266
rect 2494 37102 2546 37154
rect 68126 37102 68178 37154
rect 72382 37102 72434 37154
rect 73278 37102 73330 37154
rect 74510 37102 74562 37154
rect 75182 37102 75234 37154
rect 77422 37102 77474 37154
rect 77534 36990 77586 37042
rect 4478 36822 4530 36874
rect 4582 36822 4634 36874
rect 4686 36822 4738 36874
rect 35198 36822 35250 36874
rect 35302 36822 35354 36874
rect 35406 36822 35458 36874
rect 65918 36822 65970 36874
rect 66022 36822 66074 36874
rect 66126 36822 66178 36874
rect 76302 36654 76354 36706
rect 68798 36542 68850 36594
rect 71262 36542 71314 36594
rect 71710 36542 71762 36594
rect 72606 36542 72658 36594
rect 73838 36542 73890 36594
rect 74398 36542 74450 36594
rect 75518 36542 75570 36594
rect 77086 36542 77138 36594
rect 69694 36430 69746 36482
rect 72158 36430 72210 36482
rect 72830 36430 72882 36482
rect 73166 36430 73218 36482
rect 73390 36430 73442 36482
rect 74734 36430 74786 36482
rect 75294 36430 75346 36482
rect 76526 36430 76578 36482
rect 76862 36430 76914 36482
rect 1710 36318 1762 36370
rect 45054 36318 45106 36370
rect 45614 36318 45666 36370
rect 74958 36318 75010 36370
rect 75630 36318 75682 36370
rect 77870 36318 77922 36370
rect 78206 36318 78258 36370
rect 2046 36206 2098 36258
rect 2494 36206 2546 36258
rect 45166 36206 45218 36258
rect 73054 36206 73106 36258
rect 19838 36038 19890 36090
rect 19942 36038 19994 36090
rect 20046 36038 20098 36090
rect 50558 36038 50610 36090
rect 50662 36038 50714 36090
rect 50766 36038 50818 36090
rect 44718 35870 44770 35922
rect 56814 35870 56866 35922
rect 71374 35870 71426 35922
rect 72606 35870 72658 35922
rect 74286 35870 74338 35922
rect 77310 35870 77362 35922
rect 77982 35870 78034 35922
rect 45054 35758 45106 35810
rect 54238 35758 54290 35810
rect 55358 35758 55410 35810
rect 72942 35758 72994 35810
rect 74174 35758 74226 35810
rect 75182 35758 75234 35810
rect 76302 35758 76354 35810
rect 76974 35758 77026 35810
rect 77534 35758 77586 35810
rect 78094 35758 78146 35810
rect 45726 35646 45778 35698
rect 45950 35646 46002 35698
rect 46174 35646 46226 35698
rect 46398 35646 46450 35698
rect 54014 35646 54066 35698
rect 55022 35646 55074 35698
rect 72270 35646 72322 35698
rect 73166 35646 73218 35698
rect 74062 35646 74114 35698
rect 74622 35646 74674 35698
rect 74734 35646 74786 35698
rect 75406 35646 75458 35698
rect 76078 35646 76130 35698
rect 76750 35646 76802 35698
rect 77310 35646 77362 35698
rect 54686 35534 54738 35586
rect 55694 35534 55746 35586
rect 71710 35534 71762 35586
rect 74958 35534 75010 35586
rect 76526 35534 76578 35586
rect 45166 35422 45218 35474
rect 77870 35422 77922 35474
rect 4478 35254 4530 35306
rect 4582 35254 4634 35306
rect 4686 35254 4738 35306
rect 35198 35254 35250 35306
rect 35302 35254 35354 35306
rect 35406 35254 35458 35306
rect 65918 35254 65970 35306
rect 66022 35254 66074 35306
rect 66126 35254 66178 35306
rect 55022 34974 55074 35026
rect 55358 34974 55410 35026
rect 72606 34974 72658 35026
rect 76302 34974 76354 35026
rect 77198 34974 77250 35026
rect 45726 34862 45778 34914
rect 46174 34862 46226 34914
rect 46622 34862 46674 34914
rect 46846 34862 46898 34914
rect 46958 34862 47010 34914
rect 47182 34862 47234 34914
rect 53902 34862 53954 34914
rect 72830 34862 72882 34914
rect 73278 34862 73330 34914
rect 73950 34862 74002 34914
rect 74846 34862 74898 34914
rect 75406 34862 75458 34914
rect 76190 34862 76242 34914
rect 76862 34862 76914 34914
rect 77870 34862 77922 34914
rect 1710 34750 1762 34802
rect 2494 34750 2546 34802
rect 45166 34750 45218 34802
rect 45278 34750 45330 34802
rect 46398 34750 46450 34802
rect 53790 34750 53842 34802
rect 73502 34750 73554 34802
rect 75630 34750 75682 34802
rect 78206 34750 78258 34802
rect 2046 34638 2098 34690
rect 44382 34638 44434 34690
rect 46062 34638 46114 34690
rect 54014 34638 54066 34690
rect 71822 34638 71874 34690
rect 72158 34638 72210 34690
rect 73054 34638 73106 34690
rect 74174 34638 74226 34690
rect 74622 34638 74674 34690
rect 19838 34470 19890 34522
rect 19942 34470 19994 34522
rect 20046 34470 20098 34522
rect 50558 34470 50610 34522
rect 50662 34470 50714 34522
rect 50766 34470 50818 34522
rect 78206 34302 78258 34354
rect 2046 34190 2098 34242
rect 46286 34190 46338 34242
rect 71150 34190 71202 34242
rect 71486 34190 71538 34242
rect 72606 34190 72658 34242
rect 73166 34190 73218 34242
rect 73502 34190 73554 34242
rect 74622 34190 74674 34242
rect 75294 34190 75346 34242
rect 75966 34190 76018 34242
rect 77534 34190 77586 34242
rect 1710 34078 1762 34130
rect 45838 34078 45890 34130
rect 46510 34078 46562 34130
rect 71710 34078 71762 34130
rect 72158 34078 72210 34130
rect 72718 34078 72770 34130
rect 73726 34078 73778 34130
rect 74286 34078 74338 34130
rect 75070 34078 75122 34130
rect 75742 34078 75794 34130
rect 76302 34078 76354 34130
rect 76526 34078 76578 34130
rect 76862 34078 76914 34130
rect 77086 34078 77138 34130
rect 77646 34078 77698 34130
rect 2494 33966 2546 34018
rect 46062 33966 46114 34018
rect 70926 33966 70978 34018
rect 71262 33966 71314 34018
rect 72382 33966 72434 34018
rect 73278 33966 73330 34018
rect 76414 33966 76466 34018
rect 77310 33966 77362 34018
rect 4478 33686 4530 33738
rect 4582 33686 4634 33738
rect 4686 33686 4738 33738
rect 35198 33686 35250 33738
rect 35302 33686 35354 33738
rect 35406 33686 35458 33738
rect 65918 33686 65970 33738
rect 66022 33686 66074 33738
rect 66126 33686 66178 33738
rect 45278 33518 45330 33570
rect 71486 33518 71538 33570
rect 72046 33518 72098 33570
rect 73950 33518 74002 33570
rect 53118 33406 53170 33458
rect 54126 33406 54178 33458
rect 71150 33406 71202 33458
rect 72046 33406 72098 33458
rect 73838 33406 73890 33458
rect 74398 33406 74450 33458
rect 74846 33406 74898 33458
rect 78318 33406 78370 33458
rect 46846 33294 46898 33346
rect 53006 33294 53058 33346
rect 72718 33294 72770 33346
rect 74510 33294 74562 33346
rect 75294 33294 75346 33346
rect 76862 33294 76914 33346
rect 77086 33294 77138 33346
rect 77758 33294 77810 33346
rect 45166 33182 45218 33234
rect 45726 33182 45778 33234
rect 46398 33182 46450 33234
rect 47070 33182 47122 33234
rect 53342 33182 53394 33234
rect 76526 33182 76578 33234
rect 77422 33182 77474 33234
rect 1710 33070 1762 33122
rect 2046 33070 2098 33122
rect 2494 33070 2546 33122
rect 46062 33070 46114 33122
rect 71598 33070 71650 33122
rect 72942 33070 72994 33122
rect 73726 33070 73778 33122
rect 76638 33070 76690 33122
rect 19838 32902 19890 32954
rect 19942 32902 19994 32954
rect 20046 32902 20098 32954
rect 50558 32902 50610 32954
rect 50662 32902 50714 32954
rect 50766 32902 50818 32954
rect 70926 32734 70978 32786
rect 74174 32734 74226 32786
rect 77758 32734 77810 32786
rect 45502 32622 45554 32674
rect 45838 32622 45890 32674
rect 46174 32622 46226 32674
rect 71710 32622 71762 32674
rect 72382 32622 72434 32674
rect 72718 32622 72770 32674
rect 76750 32622 76802 32674
rect 77534 32622 77586 32674
rect 71038 32510 71090 32562
rect 71374 32510 71426 32562
rect 73726 32510 73778 32562
rect 74398 32510 74450 32562
rect 74958 32510 75010 32562
rect 75518 32510 75570 32562
rect 76414 32510 76466 32562
rect 77310 32510 77362 32562
rect 71262 32398 71314 32450
rect 73502 32398 73554 32450
rect 74286 32398 74338 32450
rect 75406 32398 75458 32450
rect 77870 32398 77922 32450
rect 74846 32286 74898 32338
rect 4478 32118 4530 32170
rect 4582 32118 4634 32170
rect 4686 32118 4738 32170
rect 35198 32118 35250 32170
rect 35302 32118 35354 32170
rect 35406 32118 35458 32170
rect 65918 32118 65970 32170
rect 66022 32118 66074 32170
rect 66126 32118 66178 32170
rect 77534 31950 77586 32002
rect 52782 31838 52834 31890
rect 75294 31838 75346 31890
rect 75742 31838 75794 31890
rect 77646 31838 77698 31890
rect 44942 31726 44994 31778
rect 45950 31726 46002 31778
rect 46174 31726 46226 31778
rect 51102 31726 51154 31778
rect 70926 31726 70978 31778
rect 71710 31726 71762 31778
rect 72270 31726 72322 31778
rect 72606 31726 72658 31778
rect 73054 31726 73106 31778
rect 73726 31726 73778 31778
rect 74062 31726 74114 31778
rect 76526 31726 76578 31778
rect 76862 31726 76914 31778
rect 77870 31726 77922 31778
rect 1710 31614 1762 31666
rect 45054 31614 45106 31666
rect 46398 31614 46450 31666
rect 46622 31614 46674 31666
rect 51438 31614 51490 31666
rect 71262 31614 71314 31666
rect 71486 31614 71538 31666
rect 72158 31614 72210 31666
rect 73278 31614 73330 31666
rect 74622 31614 74674 31666
rect 77086 31614 77138 31666
rect 2046 31502 2098 31554
rect 2494 31502 2546 31554
rect 45502 31502 45554 31554
rect 51662 31502 51714 31554
rect 71150 31502 71202 31554
rect 72046 31502 72098 31554
rect 72830 31502 72882 31554
rect 74510 31502 74562 31554
rect 74734 31502 74786 31554
rect 76638 31502 76690 31554
rect 19838 31334 19890 31386
rect 19942 31334 19994 31386
rect 20046 31334 20098 31386
rect 50558 31334 50610 31386
rect 50662 31334 50714 31386
rect 50766 31334 50818 31386
rect 44270 31166 44322 31218
rect 52334 31166 52386 31218
rect 52782 31166 52834 31218
rect 71822 31166 71874 31218
rect 72718 31166 72770 31218
rect 73502 31166 73554 31218
rect 75854 31166 75906 31218
rect 2046 31054 2098 31106
rect 44606 31054 44658 31106
rect 45726 31054 45778 31106
rect 46398 31054 46450 31106
rect 46622 31054 46674 31106
rect 47294 31054 47346 31106
rect 50318 31054 50370 31106
rect 51438 31054 51490 31106
rect 70926 31054 70978 31106
rect 74510 31054 74562 31106
rect 75182 31054 75234 31106
rect 75518 31054 75570 31106
rect 76190 31054 76242 31106
rect 77422 31054 77474 31106
rect 1710 30942 1762 30994
rect 44718 30942 44770 30994
rect 45502 30942 45554 30994
rect 45950 30942 46002 30994
rect 46174 30942 46226 30994
rect 46958 30942 47010 30994
rect 47406 30942 47458 30994
rect 50542 30942 50594 30994
rect 51102 30942 51154 30994
rect 73838 30942 73890 30994
rect 74174 30942 74226 30994
rect 74846 30942 74898 30994
rect 76526 30942 76578 30994
rect 76638 30942 76690 30994
rect 76974 30942 77026 30994
rect 77646 30942 77698 30994
rect 2494 30830 2546 30882
rect 47070 30830 47122 30882
rect 50766 30830 50818 30882
rect 71374 30830 71426 30882
rect 76302 30830 76354 30882
rect 77198 30830 77250 30882
rect 78206 30830 78258 30882
rect 51214 30718 51266 30770
rect 71262 30718 71314 30770
rect 71822 30718 71874 30770
rect 4478 30550 4530 30602
rect 4582 30550 4634 30602
rect 4686 30550 4738 30602
rect 35198 30550 35250 30602
rect 35302 30550 35354 30602
rect 35406 30550 35458 30602
rect 65918 30550 65970 30602
rect 66022 30550 66074 30602
rect 66126 30550 66178 30602
rect 45502 30382 45554 30434
rect 45838 30382 45890 30434
rect 77534 30382 77586 30434
rect 74062 30270 74114 30322
rect 77646 30270 77698 30322
rect 44942 30158 44994 30210
rect 46174 30158 46226 30210
rect 46398 30158 46450 30210
rect 46622 30158 46674 30210
rect 47070 30158 47122 30210
rect 50654 30158 50706 30210
rect 51774 30158 51826 30210
rect 71822 30158 71874 30210
rect 73278 30158 73330 30210
rect 73950 30158 74002 30210
rect 74958 30158 75010 30210
rect 75182 30158 75234 30210
rect 76638 30158 76690 30210
rect 76750 30158 76802 30210
rect 77870 30158 77922 30210
rect 44830 30046 44882 30098
rect 46062 30046 46114 30098
rect 47294 30046 47346 30098
rect 50766 30046 50818 30098
rect 51326 30046 51378 30098
rect 71598 30046 71650 30098
rect 72494 30046 72546 30098
rect 72718 30046 72770 30098
rect 73054 30046 73106 30098
rect 76302 30046 76354 30098
rect 45390 29934 45442 29986
rect 72830 29934 72882 29986
rect 76414 29934 76466 29986
rect 19838 29766 19890 29818
rect 19942 29766 19994 29818
rect 20046 29766 20098 29818
rect 50558 29766 50610 29818
rect 50662 29766 50714 29818
rect 50766 29766 50818 29818
rect 45166 29598 45218 29650
rect 72382 29598 72434 29650
rect 72606 29598 72658 29650
rect 73278 29598 73330 29650
rect 73502 29598 73554 29650
rect 77870 29598 77922 29650
rect 2046 29486 2098 29538
rect 44830 29486 44882 29538
rect 45054 29486 45106 29538
rect 71710 29486 71762 29538
rect 74398 29486 74450 29538
rect 74958 29486 75010 29538
rect 75518 29486 75570 29538
rect 76078 29486 76130 29538
rect 78206 29486 78258 29538
rect 1710 29374 1762 29426
rect 71038 29374 71090 29426
rect 71374 29374 71426 29426
rect 72830 29374 72882 29426
rect 73726 29374 73778 29426
rect 74622 29374 74674 29426
rect 76414 29374 76466 29426
rect 76638 29374 76690 29426
rect 77534 29374 77586 29426
rect 2494 29262 2546 29314
rect 72718 29262 72770 29314
rect 73614 29262 73666 29314
rect 75406 29262 75458 29314
rect 76190 29262 76242 29314
rect 77422 29262 77474 29314
rect 75742 29150 75794 29202
rect 77198 29150 77250 29202
rect 4478 28982 4530 29034
rect 4582 28982 4634 29034
rect 4686 28982 4738 29034
rect 35198 28982 35250 29034
rect 35302 28982 35354 29034
rect 35406 28982 35458 29034
rect 65918 28982 65970 29034
rect 66022 28982 66074 29034
rect 66126 28982 66178 29034
rect 77198 28814 77250 28866
rect 37550 28702 37602 28754
rect 40910 28702 40962 28754
rect 71262 28702 71314 28754
rect 71710 28702 71762 28754
rect 72158 28702 72210 28754
rect 73390 28702 73442 28754
rect 73726 28702 73778 28754
rect 77310 28702 77362 28754
rect 1710 28590 1762 28642
rect 2494 28590 2546 28642
rect 37886 28590 37938 28642
rect 38334 28590 38386 28642
rect 72382 28590 72434 28642
rect 74286 28590 74338 28642
rect 75406 28590 75458 28642
rect 75630 28590 75682 28642
rect 76526 28590 76578 28642
rect 76638 28590 76690 28642
rect 77534 28590 77586 28642
rect 78206 28590 78258 28642
rect 2046 28478 2098 28530
rect 38782 28478 38834 28530
rect 72718 28478 72770 28530
rect 75070 28478 75122 28530
rect 75182 28478 75234 28530
rect 76190 28478 76242 28530
rect 77870 28478 77922 28530
rect 37998 28366 38050 28418
rect 74510 28366 74562 28418
rect 76302 28366 76354 28418
rect 19838 28198 19890 28250
rect 19942 28198 19994 28250
rect 20046 28198 20098 28250
rect 50558 28198 50610 28250
rect 50662 28198 50714 28250
rect 50766 28198 50818 28250
rect 34750 28030 34802 28082
rect 37102 28030 37154 28082
rect 37662 28030 37714 28082
rect 39902 28030 39954 28082
rect 40350 28030 40402 28082
rect 42478 28030 42530 28082
rect 44606 28030 44658 28082
rect 70702 28030 70754 28082
rect 71822 28030 71874 28082
rect 75966 28030 76018 28082
rect 76750 28030 76802 28082
rect 77870 28030 77922 28082
rect 35086 27918 35138 27970
rect 38782 27918 38834 27970
rect 41918 27918 41970 27970
rect 44942 27918 44994 27970
rect 72718 27918 72770 27970
rect 72942 27918 72994 27970
rect 73278 27918 73330 27970
rect 74174 27918 74226 27970
rect 74958 27918 75010 27970
rect 75854 27918 75906 27970
rect 76190 27918 76242 27970
rect 76414 27918 76466 27970
rect 78206 27918 78258 27970
rect 35310 27806 35362 27858
rect 36206 27806 36258 27858
rect 36654 27806 36706 27858
rect 37886 27806 37938 27858
rect 39006 27806 39058 27858
rect 39454 27806 39506 27858
rect 41022 27806 41074 27858
rect 41470 27806 41522 27858
rect 70254 27806 70306 27858
rect 70926 27806 70978 27858
rect 73502 27806 73554 27858
rect 73726 27806 73778 27858
rect 74286 27806 74338 27858
rect 74734 27806 74786 27858
rect 75294 27806 75346 27858
rect 77086 27806 77138 27858
rect 77646 27806 77698 27858
rect 35534 27694 35586 27746
rect 38558 27694 38610 27746
rect 41358 27694 41410 27746
rect 70814 27694 70866 27746
rect 73054 27694 73106 27746
rect 73950 27694 74002 27746
rect 75182 27694 75234 27746
rect 45054 27582 45106 27634
rect 4478 27414 4530 27466
rect 4582 27414 4634 27466
rect 4686 27414 4738 27466
rect 35198 27414 35250 27466
rect 35302 27414 35354 27466
rect 35406 27414 35458 27466
rect 65918 27414 65970 27466
rect 66022 27414 66074 27466
rect 66126 27414 66178 27466
rect 76190 27246 76242 27298
rect 76862 27246 76914 27298
rect 43822 27134 43874 27186
rect 44830 27134 44882 27186
rect 45390 27134 45442 27186
rect 46398 27134 46450 27186
rect 50318 27134 50370 27186
rect 50766 27134 50818 27186
rect 71934 27134 71986 27186
rect 75406 27134 75458 27186
rect 76974 27134 77026 27186
rect 34078 27022 34130 27074
rect 34750 27022 34802 27074
rect 35758 27022 35810 27074
rect 36206 27022 36258 27074
rect 36990 27022 37042 27074
rect 37438 27022 37490 27074
rect 38110 27022 38162 27074
rect 38670 27022 38722 27074
rect 39790 27022 39842 27074
rect 40686 27022 40738 27074
rect 41022 27022 41074 27074
rect 42142 27022 42194 27074
rect 43038 27022 43090 27074
rect 46174 27022 46226 27074
rect 47070 27022 47122 27074
rect 47294 27022 47346 27074
rect 49086 27022 49138 27074
rect 49646 27022 49698 27074
rect 70590 27022 70642 27074
rect 71038 27022 71090 27074
rect 72382 27022 72434 27074
rect 73390 27022 73442 27074
rect 73502 27022 73554 27074
rect 75294 27022 75346 27074
rect 77198 27022 77250 27074
rect 1710 26910 1762 26962
rect 2046 26910 2098 26962
rect 2494 26910 2546 26962
rect 34974 26910 35026 26962
rect 35646 26910 35698 26962
rect 38782 26910 38834 26962
rect 40574 26910 40626 26962
rect 41694 26910 41746 26962
rect 44942 26910 44994 26962
rect 46622 26910 46674 26962
rect 46846 26910 46898 26962
rect 47518 26910 47570 26962
rect 47742 26910 47794 26962
rect 49758 26910 49810 26962
rect 73054 26910 73106 26962
rect 74286 26910 74338 26962
rect 74622 26910 74674 26962
rect 75630 26910 75682 26962
rect 76526 26910 76578 26962
rect 77534 26910 77586 26962
rect 77870 26910 77922 26962
rect 33966 26798 34018 26850
rect 36206 26798 36258 26850
rect 38334 26798 38386 26850
rect 39790 26798 39842 26850
rect 41134 26798 41186 26850
rect 42478 26798 42530 26850
rect 44382 26798 44434 26850
rect 49198 26798 49250 26850
rect 49422 26798 49474 26850
rect 49982 26798 50034 26850
rect 71150 26798 71202 26850
rect 71262 26798 71314 26850
rect 72830 26798 72882 26850
rect 73166 26798 73218 26850
rect 76302 26798 76354 26850
rect 19838 26630 19890 26682
rect 19942 26630 19994 26682
rect 20046 26630 20098 26682
rect 50558 26630 50610 26682
rect 50662 26630 50714 26682
rect 50766 26630 50818 26682
rect 35198 26462 35250 26514
rect 42590 26462 42642 26514
rect 44046 26462 44098 26514
rect 44606 26462 44658 26514
rect 47518 26462 47570 26514
rect 50094 26462 50146 26514
rect 50542 26462 50594 26514
rect 70926 26462 70978 26514
rect 76974 26462 77026 26514
rect 77198 26462 77250 26514
rect 77870 26462 77922 26514
rect 2046 26350 2098 26402
rect 35870 26350 35922 26402
rect 38782 26350 38834 26402
rect 41694 26350 41746 26402
rect 43038 26350 43090 26402
rect 44942 26350 44994 26402
rect 46062 26350 46114 26402
rect 46734 26350 46786 26402
rect 47630 26350 47682 26402
rect 48862 26350 48914 26402
rect 49310 26350 49362 26402
rect 49422 26350 49474 26402
rect 75630 26350 75682 26402
rect 76302 26350 76354 26402
rect 77534 26350 77586 26402
rect 1710 26238 1762 26290
rect 35982 26238 36034 26290
rect 36318 26238 36370 26290
rect 37326 26238 37378 26290
rect 37774 26238 37826 26290
rect 38110 26238 38162 26290
rect 39230 26238 39282 26290
rect 40350 26238 40402 26290
rect 41022 26238 41074 26290
rect 41806 26238 41858 26290
rect 43598 26238 43650 26290
rect 44158 26238 44210 26290
rect 45054 26238 45106 26290
rect 45838 26238 45890 26290
rect 46286 26238 46338 26290
rect 46510 26238 46562 26290
rect 46846 26238 46898 26290
rect 47182 26238 47234 26290
rect 47742 26238 47794 26290
rect 48750 26238 48802 26290
rect 71150 26238 71202 26290
rect 71374 26238 71426 26290
rect 72382 26238 72434 26290
rect 73502 26238 73554 26290
rect 74286 26238 74338 26290
rect 74846 26238 74898 26290
rect 75406 26238 75458 26290
rect 75966 26238 76018 26290
rect 78206 26238 78258 26290
rect 2494 26126 2546 26178
rect 35758 26126 35810 26178
rect 38558 26126 38610 26178
rect 39902 26126 39954 26178
rect 41470 26126 41522 26178
rect 48862 26014 48914 26066
rect 70814 26126 70866 26178
rect 71262 26126 71314 26178
rect 72942 26126 72994 26178
rect 73278 26126 73330 26178
rect 49422 26014 49474 26066
rect 70590 26014 70642 26066
rect 74062 26014 74114 26066
rect 4478 25846 4530 25898
rect 4582 25846 4634 25898
rect 4686 25846 4738 25898
rect 35198 25846 35250 25898
rect 35302 25846 35354 25898
rect 35406 25846 35458 25898
rect 65918 25846 65970 25898
rect 66022 25846 66074 25898
rect 66126 25846 66178 25898
rect 47070 25678 47122 25730
rect 72718 25678 72770 25730
rect 74398 25678 74450 25730
rect 77758 25678 77810 25730
rect 78094 25678 78146 25730
rect 35870 25566 35922 25618
rect 37774 25566 37826 25618
rect 44046 25566 44098 25618
rect 46958 25566 47010 25618
rect 47518 25566 47570 25618
rect 47966 25566 48018 25618
rect 63310 25566 63362 25618
rect 71038 25566 71090 25618
rect 37326 25454 37378 25506
rect 38110 25454 38162 25506
rect 38334 25454 38386 25506
rect 40350 25454 40402 25506
rect 42478 25454 42530 25506
rect 43374 25454 43426 25506
rect 44830 25454 44882 25506
rect 45726 25454 45778 25506
rect 62862 25454 62914 25506
rect 63198 25454 63250 25506
rect 70814 25454 70866 25506
rect 71822 25454 71874 25506
rect 72158 25454 72210 25506
rect 72494 25454 72546 25506
rect 73278 25454 73330 25506
rect 73838 25454 73890 25506
rect 74174 25454 74226 25506
rect 74958 25454 75010 25506
rect 75518 25454 75570 25506
rect 76750 25454 76802 25506
rect 77422 25454 77474 25506
rect 2046 25342 2098 25394
rect 23998 25342 24050 25394
rect 27134 25342 27186 25394
rect 36430 25342 36482 25394
rect 40462 25342 40514 25394
rect 42142 25342 42194 25394
rect 42590 25342 42642 25394
rect 44942 25342 44994 25394
rect 46286 25342 46338 25394
rect 46622 25342 46674 25394
rect 70702 25342 70754 25394
rect 76414 25342 76466 25394
rect 77086 25342 77138 25394
rect 1710 25230 1762 25282
rect 2494 25230 2546 25282
rect 23662 25230 23714 25282
rect 24110 25230 24162 25282
rect 24334 25230 24386 25282
rect 27022 25230 27074 25282
rect 35534 25230 35586 25282
rect 40014 25230 40066 25282
rect 41806 25230 41858 25282
rect 43486 25230 43538 25282
rect 45838 25230 45890 25282
rect 63422 25230 63474 25282
rect 77982 25230 78034 25282
rect 19838 25062 19890 25114
rect 19942 25062 19994 25114
rect 20046 25062 20098 25114
rect 50558 25062 50610 25114
rect 50662 25062 50714 25114
rect 50766 25062 50818 25114
rect 25342 24894 25394 24946
rect 34974 24894 35026 24946
rect 35310 24894 35362 24946
rect 37438 24894 37490 24946
rect 39454 24894 39506 24946
rect 40350 24894 40402 24946
rect 44382 24894 44434 24946
rect 45950 24894 46002 24946
rect 48190 24894 48242 24946
rect 63198 24894 63250 24946
rect 63982 24894 64034 24946
rect 71710 24894 71762 24946
rect 74174 24894 74226 24946
rect 74958 24894 75010 24946
rect 75406 24894 75458 24946
rect 76190 24894 76242 24946
rect 77646 24894 77698 24946
rect 35758 24782 35810 24834
rect 41694 24782 41746 24834
rect 44942 24782 44994 24834
rect 46622 24782 46674 24834
rect 46958 24782 47010 24834
rect 47294 24782 47346 24834
rect 76078 24782 76130 24834
rect 77086 24782 77138 24834
rect 77534 24782 77586 24834
rect 77758 24782 77810 24834
rect 17502 24670 17554 24722
rect 20638 24670 20690 24722
rect 25566 24670 25618 24722
rect 25790 24670 25842 24722
rect 27246 24670 27298 24722
rect 30382 24670 30434 24722
rect 30494 24670 30546 24722
rect 35086 24670 35138 24722
rect 35422 24670 35474 24722
rect 35982 24670 36034 24722
rect 37550 24670 37602 24722
rect 37886 24670 37938 24722
rect 39342 24670 39394 24722
rect 40126 24670 40178 24722
rect 40910 24670 40962 24722
rect 44158 24670 44210 24722
rect 45278 24670 45330 24722
rect 45614 24670 45666 24722
rect 46398 24670 46450 24722
rect 48862 24670 48914 24722
rect 62750 24670 62802 24722
rect 63422 24670 63474 24722
rect 72158 24670 72210 24722
rect 73054 24670 73106 24722
rect 73502 24670 73554 24722
rect 74622 24670 74674 24722
rect 75630 24670 75682 24722
rect 18174 24558 18226 24610
rect 20302 24558 20354 24610
rect 21422 24558 21474 24610
rect 23550 24558 23602 24610
rect 23886 24558 23938 24610
rect 24222 24558 24274 24610
rect 25678 24558 25730 24610
rect 27918 24558 27970 24610
rect 30046 24558 30098 24610
rect 43822 24558 43874 24610
rect 47854 24558 47906 24610
rect 63310 24558 63362 24610
rect 71374 24558 71426 24610
rect 77198 24558 77250 24610
rect 39454 24446 39506 24498
rect 72382 24446 72434 24498
rect 75294 24446 75346 24498
rect 76302 24446 76354 24498
rect 76862 24446 76914 24498
rect 4478 24278 4530 24330
rect 4582 24278 4634 24330
rect 4686 24278 4738 24330
rect 35198 24278 35250 24330
rect 35302 24278 35354 24330
rect 35406 24278 35458 24330
rect 65918 24278 65970 24330
rect 66022 24278 66074 24330
rect 66126 24278 66178 24330
rect 35982 24110 36034 24162
rect 75294 24110 75346 24162
rect 76190 24110 76242 24162
rect 76526 24110 76578 24162
rect 17166 23998 17218 24050
rect 17614 23998 17666 24050
rect 19742 23998 19794 24050
rect 20078 23998 20130 24050
rect 21758 23998 21810 24050
rect 23326 23998 23378 24050
rect 25006 23998 25058 24050
rect 27134 23998 27186 24050
rect 28030 23998 28082 24050
rect 42366 23998 42418 24050
rect 43262 23998 43314 24050
rect 44158 23998 44210 24050
rect 48302 23998 48354 24050
rect 74286 23998 74338 24050
rect 17726 23886 17778 23938
rect 18174 23886 18226 23938
rect 18286 23886 18338 23938
rect 18622 23886 18674 23938
rect 20750 23886 20802 23938
rect 21198 23886 21250 23938
rect 23662 23886 23714 23938
rect 23998 23886 24050 23938
rect 24334 23886 24386 23938
rect 27470 23886 27522 23938
rect 34750 23886 34802 23938
rect 35870 23886 35922 23938
rect 38222 23886 38274 23938
rect 39454 23886 39506 23938
rect 40350 23886 40402 23938
rect 41806 23886 41858 23938
rect 42702 23886 42754 23938
rect 46062 23886 46114 23938
rect 46510 23886 46562 23938
rect 46734 23886 46786 23938
rect 72270 23886 72322 23938
rect 73278 23886 73330 23938
rect 73614 23886 73666 23938
rect 75406 23886 75458 23938
rect 1710 23774 1762 23826
rect 2046 23774 2098 23826
rect 18510 23774 18562 23826
rect 20414 23774 20466 23826
rect 27918 23774 27970 23826
rect 35646 23774 35698 23826
rect 37102 23774 37154 23826
rect 37214 23774 37266 23826
rect 37662 23774 37714 23826
rect 37774 23774 37826 23826
rect 40462 23774 40514 23826
rect 43598 23774 43650 23826
rect 43710 23774 43762 23826
rect 44830 23774 44882 23826
rect 45390 23774 45442 23826
rect 47070 23774 47122 23826
rect 47182 23774 47234 23826
rect 47630 23774 47682 23826
rect 47742 23774 47794 23826
rect 48750 23774 48802 23826
rect 73726 23774 73778 23826
rect 74622 23774 74674 23826
rect 74958 23774 75010 23826
rect 76862 23774 76914 23826
rect 77198 23774 77250 23826
rect 77870 23774 77922 23826
rect 78206 23774 78258 23826
rect 2494 23662 2546 23714
rect 17502 23662 17554 23714
rect 19406 23662 19458 23714
rect 20526 23662 20578 23714
rect 21646 23662 21698 23714
rect 21870 23662 21922 23714
rect 22318 23662 22370 23714
rect 23774 23662 23826 23714
rect 28142 23662 28194 23714
rect 34302 23662 34354 23714
rect 35086 23662 35138 23714
rect 35982 23662 36034 23714
rect 37438 23662 37490 23714
rect 37998 23662 38050 23714
rect 39342 23662 39394 23714
rect 43934 23662 43986 23714
rect 44270 23662 44322 23714
rect 44942 23662 44994 23714
rect 45166 23662 45218 23714
rect 45502 23662 45554 23714
rect 46398 23662 46450 23714
rect 47406 23662 47458 23714
rect 47966 23662 48018 23714
rect 49310 23662 49362 23714
rect 49646 23662 49698 23714
rect 72158 23662 72210 23714
rect 75518 23662 75570 23714
rect 76414 23662 76466 23714
rect 19838 23494 19890 23546
rect 19942 23494 19994 23546
rect 20046 23494 20098 23546
rect 50558 23494 50610 23546
rect 50662 23494 50714 23546
rect 50766 23494 50818 23546
rect 18398 23326 18450 23378
rect 24222 23326 24274 23378
rect 25790 23326 25842 23378
rect 27582 23326 27634 23378
rect 33742 23326 33794 23378
rect 34526 23326 34578 23378
rect 35086 23326 35138 23378
rect 36654 23326 36706 23378
rect 43374 23326 43426 23378
rect 45726 23326 45778 23378
rect 47182 23326 47234 23378
rect 51102 23326 51154 23378
rect 71710 23326 71762 23378
rect 74398 23326 74450 23378
rect 2046 23214 2098 23266
rect 17502 23214 17554 23266
rect 17614 23214 17666 23266
rect 19518 23214 19570 23266
rect 19630 23214 19682 23266
rect 23886 23214 23938 23266
rect 23998 23214 24050 23266
rect 35870 23214 35922 23266
rect 41246 23214 41298 23266
rect 41694 23214 41746 23266
rect 42814 23214 42866 23266
rect 44494 23214 44546 23266
rect 46510 23214 46562 23266
rect 47518 23214 47570 23266
rect 47966 23214 48018 23266
rect 76862 23214 76914 23266
rect 77086 23214 77138 23266
rect 77534 23214 77586 23266
rect 77758 23214 77810 23266
rect 1710 23102 1762 23154
rect 19854 23102 19906 23154
rect 20302 23102 20354 23154
rect 25118 23102 25170 23154
rect 25566 23102 25618 23154
rect 26910 23102 26962 23154
rect 27358 23102 27410 23154
rect 27918 23102 27970 23154
rect 34190 23102 34242 23154
rect 34302 23102 34354 23154
rect 34638 23102 34690 23154
rect 35198 23102 35250 23154
rect 35758 23102 35810 23154
rect 37326 23102 37378 23154
rect 37662 23102 37714 23154
rect 39790 23102 39842 23154
rect 40910 23102 40962 23154
rect 41582 23102 41634 23154
rect 42366 23102 42418 23154
rect 44158 23102 44210 23154
rect 45614 23102 45666 23154
rect 47854 23102 47906 23154
rect 48190 23102 48242 23154
rect 48862 23102 48914 23154
rect 72158 23102 72210 23154
rect 72942 23102 72994 23154
rect 73502 23102 73554 23154
rect 74510 23102 74562 23154
rect 74846 23102 74898 23154
rect 75966 23102 76018 23154
rect 76190 23102 76242 23154
rect 2494 22990 2546 23042
rect 16830 22990 16882 23042
rect 19182 22990 19234 23042
rect 21086 22990 21138 23042
rect 23214 22990 23266 23042
rect 24558 22990 24610 23042
rect 25678 22990 25730 23042
rect 27470 22990 27522 23042
rect 28702 22990 28754 23042
rect 30830 22990 30882 23042
rect 39454 22990 39506 23042
rect 40350 22990 40402 23042
rect 42254 22990 42306 23042
rect 49198 22990 49250 23042
rect 49310 22990 49362 23042
rect 17502 22878 17554 22930
rect 35086 22878 35138 22930
rect 41694 22878 41746 22930
rect 48750 22878 48802 22930
rect 49870 22990 49922 23042
rect 50206 22990 50258 23042
rect 74846 22990 74898 23042
rect 77198 22990 77250 23042
rect 77870 22990 77922 23042
rect 50206 22878 50258 22930
rect 72382 22878 72434 22930
rect 75070 22878 75122 22930
rect 76414 22878 76466 22930
rect 76638 22878 76690 22930
rect 4478 22710 4530 22762
rect 4582 22710 4634 22762
rect 4686 22710 4738 22762
rect 35198 22710 35250 22762
rect 35302 22710 35354 22762
rect 35406 22710 35458 22762
rect 65918 22710 65970 22762
rect 66022 22710 66074 22762
rect 66126 22710 66178 22762
rect 50542 22542 50594 22594
rect 51102 22542 51154 22594
rect 51326 22542 51378 22594
rect 51774 22542 51826 22594
rect 74174 22542 74226 22594
rect 77534 22542 77586 22594
rect 77870 22542 77922 22594
rect 19406 22430 19458 22482
rect 20414 22430 20466 22482
rect 21758 22430 21810 22482
rect 23102 22430 23154 22482
rect 25118 22430 25170 22482
rect 27246 22430 27298 22482
rect 37326 22430 37378 22482
rect 42030 22430 42082 22482
rect 43374 22430 43426 22482
rect 44830 22430 44882 22482
rect 48638 22430 48690 22482
rect 50430 22430 50482 22482
rect 51774 22430 51826 22482
rect 53790 22430 53842 22482
rect 54238 22430 54290 22482
rect 71710 22430 71762 22482
rect 72158 22430 72210 22482
rect 72494 22430 72546 22482
rect 75070 22430 75122 22482
rect 76526 22430 76578 22482
rect 16606 22318 16658 22370
rect 19966 22318 20018 22370
rect 21198 22318 21250 22370
rect 23550 22318 23602 22370
rect 24334 22318 24386 22370
rect 27582 22318 27634 22370
rect 30830 22318 30882 22370
rect 30942 22318 30994 22370
rect 34302 22318 34354 22370
rect 35310 22318 35362 22370
rect 37774 22318 37826 22370
rect 39006 22318 39058 22370
rect 41358 22318 41410 22370
rect 42478 22318 42530 22370
rect 43822 22318 43874 22370
rect 45390 22318 45442 22370
rect 46062 22318 46114 22370
rect 46510 22318 46562 22370
rect 46734 22318 46786 22370
rect 47406 22318 47458 22370
rect 47518 22318 47570 22370
rect 49422 22318 49474 22370
rect 49982 22318 50034 22370
rect 52782 22318 52834 22370
rect 53342 22318 53394 22370
rect 72270 22318 72322 22370
rect 73278 22318 73330 22370
rect 73614 22318 73666 22370
rect 73950 22318 74002 22370
rect 74958 22318 75010 22370
rect 17278 22206 17330 22258
rect 19742 22206 19794 22258
rect 20750 22206 20802 22258
rect 23774 22206 23826 22258
rect 33518 22206 33570 22258
rect 35758 22206 35810 22258
rect 39454 22206 39506 22258
rect 41246 22206 41298 22258
rect 44942 22206 44994 22258
rect 47070 22206 47122 22258
rect 47966 22206 48018 22258
rect 48078 22206 48130 22258
rect 76750 22206 76802 22258
rect 21646 22094 21698 22146
rect 21870 22094 21922 22146
rect 22990 22094 23042 22146
rect 27694 22094 27746 22146
rect 34302 22094 34354 22146
rect 40574 22094 40626 22146
rect 44270 22094 44322 22146
rect 45614 22094 45666 22146
rect 46398 22094 46450 22146
rect 47294 22094 47346 22146
rect 48302 22094 48354 22146
rect 49086 22094 49138 22146
rect 50878 22094 50930 22146
rect 51438 22094 51490 22146
rect 77086 22094 77138 22146
rect 77758 22094 77810 22146
rect 19838 21926 19890 21978
rect 19942 21926 19994 21978
rect 20046 21926 20098 21978
rect 50558 21926 50610 21978
rect 50662 21926 50714 21978
rect 50766 21926 50818 21978
rect 2046 21758 2098 21810
rect 17502 21758 17554 21810
rect 17838 21758 17890 21810
rect 24222 21758 24274 21810
rect 26238 21758 26290 21810
rect 35422 21758 35474 21810
rect 36206 21758 36258 21810
rect 38222 21758 38274 21810
rect 41246 21758 41298 21810
rect 47742 21758 47794 21810
rect 48862 21758 48914 21810
rect 55022 21758 55074 21810
rect 56030 21758 56082 21810
rect 70030 21758 70082 21810
rect 74622 21758 74674 21810
rect 75854 21758 75906 21810
rect 77310 21758 77362 21810
rect 77870 21758 77922 21810
rect 22318 21646 22370 21698
rect 23886 21646 23938 21698
rect 23998 21646 24050 21698
rect 25678 21646 25730 21698
rect 37438 21646 37490 21698
rect 39454 21646 39506 21698
rect 42478 21646 42530 21698
rect 44046 21646 44098 21698
rect 46174 21646 46226 21698
rect 49870 21646 49922 21698
rect 50878 21646 50930 21698
rect 51774 21646 51826 21698
rect 54462 21646 54514 21698
rect 55582 21646 55634 21698
rect 72270 21646 72322 21698
rect 75182 21646 75234 21698
rect 76638 21646 76690 21698
rect 77198 21646 77250 21698
rect 78206 21646 78258 21698
rect 1710 21534 1762 21586
rect 17726 21534 17778 21586
rect 17950 21534 18002 21586
rect 19182 21534 19234 21586
rect 22542 21534 22594 21586
rect 26462 21534 26514 21586
rect 35086 21534 35138 21586
rect 35534 21534 35586 21586
rect 35758 21534 35810 21586
rect 35982 21534 36034 21586
rect 36430 21534 36482 21586
rect 36542 21534 36594 21586
rect 37550 21534 37602 21586
rect 39230 21534 39282 21586
rect 44942 21534 44994 21586
rect 45838 21534 45890 21586
rect 47406 21534 47458 21586
rect 47630 21534 47682 21586
rect 47966 21534 48018 21586
rect 48750 21534 48802 21586
rect 49422 21534 49474 21586
rect 50206 21534 50258 21586
rect 51326 21534 51378 21586
rect 52222 21534 52274 21586
rect 52782 21534 52834 21586
rect 53118 21534 53170 21586
rect 54350 21534 54402 21586
rect 54910 21534 54962 21586
rect 70254 21534 70306 21586
rect 71374 21534 71426 21586
rect 71598 21534 71650 21586
rect 72606 21534 72658 21586
rect 73278 21534 73330 21586
rect 74062 21534 74114 21586
rect 74846 21534 74898 21586
rect 75518 21534 75570 21586
rect 76862 21534 76914 21586
rect 77534 21534 77586 21586
rect 2494 21422 2546 21474
rect 18398 21422 18450 21474
rect 19854 21422 19906 21474
rect 21982 21422 22034 21474
rect 23550 21422 23602 21474
rect 33294 21422 33346 21474
rect 33630 21422 33682 21474
rect 34526 21422 34578 21474
rect 34862 21422 34914 21474
rect 43262 21422 43314 21474
rect 46622 21422 46674 21474
rect 50878 21422 50930 21474
rect 52334 21422 52386 21474
rect 53678 21422 53730 21474
rect 70590 21422 70642 21474
rect 73054 21422 73106 21474
rect 76526 21422 76578 21474
rect 42030 21310 42082 21362
rect 4478 21142 4530 21194
rect 4582 21142 4634 21194
rect 4686 21142 4738 21194
rect 35198 21142 35250 21194
rect 35302 21142 35354 21194
rect 35406 21142 35458 21194
rect 65918 21142 65970 21194
rect 66022 21142 66074 21194
rect 66126 21142 66178 21194
rect 75294 20974 75346 21026
rect 77086 20974 77138 21026
rect 77422 20974 77474 21026
rect 21758 20862 21810 20914
rect 25006 20862 25058 20914
rect 30158 20862 30210 20914
rect 33630 20862 33682 20914
rect 34414 20862 34466 20914
rect 35310 20862 35362 20914
rect 38110 20862 38162 20914
rect 46174 20862 46226 20914
rect 47070 20862 47122 20914
rect 51326 20862 51378 20914
rect 57150 20862 57202 20914
rect 70926 20862 70978 20914
rect 71262 20862 71314 20914
rect 72158 20862 72210 20914
rect 72942 20862 72994 20914
rect 73838 20862 73890 20914
rect 74734 20862 74786 20914
rect 77534 20862 77586 20914
rect 78318 20862 78370 20914
rect 18622 20750 18674 20802
rect 22094 20750 22146 20802
rect 25342 20750 25394 20802
rect 26014 20750 26066 20802
rect 27246 20750 27298 20802
rect 29038 20750 29090 20802
rect 29486 20750 29538 20802
rect 30830 20750 30882 20802
rect 34190 20750 34242 20802
rect 34862 20750 34914 20802
rect 35758 20750 35810 20802
rect 36430 20750 36482 20802
rect 37886 20750 37938 20802
rect 39342 20750 39394 20802
rect 41246 20750 41298 20802
rect 42926 20750 42978 20802
rect 43262 20750 43314 20802
rect 44830 20750 44882 20802
rect 45278 20750 45330 20802
rect 45726 20750 45778 20802
rect 46622 20750 46674 20802
rect 47182 20750 47234 20802
rect 48302 20750 48354 20802
rect 49422 20750 49474 20802
rect 49758 20750 49810 20802
rect 50430 20750 50482 20802
rect 51662 20750 51714 20802
rect 52782 20750 52834 20802
rect 53230 20750 53282 20802
rect 54126 20750 54178 20802
rect 54686 20750 54738 20802
rect 55582 20750 55634 20802
rect 56142 20750 56194 20802
rect 71038 20750 71090 20802
rect 72046 20750 72098 20802
rect 72718 20750 72770 20802
rect 73502 20750 73554 20802
rect 76750 20750 76802 20802
rect 77758 20750 77810 20802
rect 2046 20638 2098 20690
rect 18958 20638 19010 20690
rect 19070 20638 19122 20690
rect 22878 20638 22930 20690
rect 25678 20638 25730 20690
rect 26350 20638 26402 20690
rect 30382 20638 30434 20690
rect 31502 20638 31554 20690
rect 34638 20638 34690 20690
rect 35198 20638 35250 20690
rect 35534 20638 35586 20690
rect 36094 20638 36146 20690
rect 36990 20638 37042 20690
rect 38334 20638 38386 20690
rect 38558 20638 38610 20690
rect 39006 20638 39058 20690
rect 40014 20638 40066 20690
rect 40350 20638 40402 20690
rect 41134 20638 41186 20690
rect 47742 20638 47794 20690
rect 48638 20638 48690 20690
rect 50654 20638 50706 20690
rect 53454 20638 53506 20690
rect 55246 20638 55298 20690
rect 56254 20638 56306 20690
rect 75630 20638 75682 20690
rect 1710 20526 1762 20578
rect 2494 20526 2546 20578
rect 19294 20526 19346 20578
rect 20638 20526 20690 20578
rect 21646 20526 21698 20578
rect 26126 20526 26178 20578
rect 26574 20526 26626 20578
rect 26910 20526 26962 20578
rect 27358 20526 27410 20578
rect 27582 20526 27634 20578
rect 27918 20526 27970 20578
rect 29598 20526 29650 20578
rect 29710 20526 29762 20578
rect 37326 20526 37378 20578
rect 39678 20526 39730 20578
rect 40686 20526 40738 20578
rect 43038 20526 43090 20578
rect 49198 20526 49250 20578
rect 49870 20526 49922 20578
rect 52894 20526 52946 20578
rect 54238 20526 54290 20578
rect 55694 20526 55746 20578
rect 75406 20526 75458 20578
rect 76302 20526 76354 20578
rect 76974 20526 77026 20578
rect 19838 20358 19890 20410
rect 19942 20358 19994 20410
rect 20046 20358 20098 20410
rect 50558 20358 50610 20410
rect 50662 20358 50714 20410
rect 50766 20358 50818 20410
rect 18734 20190 18786 20242
rect 31502 20190 31554 20242
rect 33966 20190 34018 20242
rect 34414 20190 34466 20242
rect 39678 20190 39730 20242
rect 42814 20190 42866 20242
rect 46510 20190 46562 20242
rect 48078 20190 48130 20242
rect 52894 20190 52946 20242
rect 54350 20190 54402 20242
rect 72606 20190 72658 20242
rect 74622 20190 74674 20242
rect 18398 20078 18450 20130
rect 25230 20078 25282 20130
rect 26238 20078 26290 20130
rect 26350 20078 26402 20130
rect 26910 20078 26962 20130
rect 28478 20078 28530 20130
rect 31390 20078 31442 20130
rect 33518 20078 33570 20130
rect 34862 20078 34914 20130
rect 35534 20078 35586 20130
rect 36318 20078 36370 20130
rect 38782 20078 38834 20130
rect 41358 20078 41410 20130
rect 42926 20078 42978 20130
rect 44494 20078 44546 20130
rect 46958 20078 47010 20130
rect 49422 20078 49474 20130
rect 52110 20078 52162 20130
rect 53454 20078 53506 20130
rect 55246 20078 55298 20130
rect 56702 20078 56754 20130
rect 75182 20078 75234 20130
rect 76190 20078 76242 20130
rect 76302 20078 76354 20130
rect 76750 20078 76802 20130
rect 77086 20078 77138 20130
rect 77870 20078 77922 20130
rect 24670 19966 24722 20018
rect 26574 19966 26626 20018
rect 27806 19966 27858 20018
rect 30942 19966 30994 20018
rect 31614 19966 31666 20018
rect 35422 19966 35474 20018
rect 36206 19966 36258 20018
rect 37662 19966 37714 20018
rect 37998 19966 38050 20018
rect 39342 19966 39394 20018
rect 39678 19966 39730 20018
rect 39902 19966 39954 20018
rect 41134 19966 41186 20018
rect 43038 19966 43090 20018
rect 44718 19966 44770 20018
rect 46622 19966 46674 20018
rect 48862 19966 48914 20018
rect 50094 19966 50146 20018
rect 51102 19966 51154 20018
rect 51438 19966 51490 20018
rect 52782 19966 52834 20018
rect 53342 19966 53394 20018
rect 54462 19966 54514 20018
rect 54798 19966 54850 20018
rect 55806 19966 55858 20018
rect 76078 19966 76130 20018
rect 78094 19966 78146 20018
rect 19630 19854 19682 19906
rect 25566 19854 25618 19906
rect 27470 19854 27522 19906
rect 30606 19854 30658 19906
rect 32174 19854 32226 19906
rect 32622 19854 32674 19906
rect 33406 19854 33458 19906
rect 33854 19854 33906 19906
rect 34302 19854 34354 19906
rect 34750 19854 34802 19906
rect 48190 19854 48242 19906
rect 77646 19854 77698 19906
rect 4478 19574 4530 19626
rect 4582 19574 4634 19626
rect 4686 19574 4738 19626
rect 35198 19574 35250 19626
rect 35302 19574 35354 19626
rect 35406 19574 35458 19626
rect 65918 19574 65970 19626
rect 66022 19574 66074 19626
rect 66126 19574 66178 19626
rect 76750 19406 76802 19458
rect 77422 19406 77474 19458
rect 18846 19294 18898 19346
rect 20302 19294 20354 19346
rect 21758 19294 21810 19346
rect 22766 19294 22818 19346
rect 24446 19294 24498 19346
rect 35534 19294 35586 19346
rect 36430 19294 36482 19346
rect 38110 19294 38162 19346
rect 43934 19294 43986 19346
rect 48526 19294 48578 19346
rect 51774 19294 51826 19346
rect 78318 19294 78370 19346
rect 19742 19182 19794 19234
rect 20414 19182 20466 19234
rect 22318 19182 22370 19234
rect 22654 19182 22706 19234
rect 26350 19182 26402 19234
rect 26686 19182 26738 19234
rect 27022 19182 27074 19234
rect 27694 19182 27746 19234
rect 34414 19182 34466 19234
rect 35646 19182 35698 19234
rect 35870 19182 35922 19234
rect 38334 19182 38386 19234
rect 38558 19182 38610 19234
rect 38782 19182 38834 19234
rect 39230 19182 39282 19234
rect 39342 19182 39394 19234
rect 40798 19182 40850 19234
rect 42254 19182 42306 19234
rect 43374 19182 43426 19234
rect 44830 19182 44882 19234
rect 45390 19182 45442 19234
rect 47070 19182 47122 19234
rect 49870 19182 49922 19234
rect 50990 19182 51042 19234
rect 52670 19182 52722 19234
rect 53230 19182 53282 19234
rect 53902 19182 53954 19234
rect 55470 19182 55522 19234
rect 56142 19182 56194 19234
rect 76862 19182 76914 19234
rect 77758 19182 77810 19234
rect 1710 19070 1762 19122
rect 2046 19070 2098 19122
rect 2494 19070 2546 19122
rect 19182 19070 19234 19122
rect 19294 19070 19346 19122
rect 21982 19070 22034 19122
rect 22878 19070 22930 19122
rect 23550 19070 23602 19122
rect 23886 19070 23938 19122
rect 24782 19070 24834 19122
rect 25118 19070 25170 19122
rect 25454 19070 25506 19122
rect 25790 19070 25842 19122
rect 29150 19070 29202 19122
rect 29486 19070 29538 19122
rect 30270 19070 30322 19122
rect 35422 19070 35474 19122
rect 37662 19070 37714 19122
rect 37998 19070 38050 19122
rect 40126 19070 40178 19122
rect 40462 19070 40514 19122
rect 41246 19070 41298 19122
rect 42926 19070 42978 19122
rect 46958 19070 47010 19122
rect 49310 19070 49362 19122
rect 51102 19070 51154 19122
rect 54126 19070 54178 19122
rect 57374 19070 57426 19122
rect 19518 18958 19570 19010
rect 20190 18958 20242 19010
rect 23102 18958 23154 19010
rect 26462 18958 26514 19010
rect 27470 18958 27522 19010
rect 27582 18958 27634 19010
rect 28142 18958 28194 19010
rect 28590 18958 28642 19010
rect 37326 18958 37378 19010
rect 39118 18958 39170 19010
rect 39790 18958 39842 19010
rect 40574 18958 40626 19010
rect 46846 18958 46898 19010
rect 55358 18958 55410 19010
rect 76526 18958 76578 19010
rect 76974 18958 77026 19010
rect 77534 18958 77586 19010
rect 19838 18790 19890 18842
rect 19942 18790 19994 18842
rect 20046 18790 20098 18842
rect 50558 18790 50610 18842
rect 50662 18790 50714 18842
rect 50766 18790 50818 18842
rect 17614 18622 17666 18674
rect 18062 18622 18114 18674
rect 40014 18622 40066 18674
rect 41694 18622 41746 18674
rect 46958 18622 47010 18674
rect 49870 18622 49922 18674
rect 54014 18622 54066 18674
rect 77534 18622 77586 18674
rect 77870 18622 77922 18674
rect 2046 18510 2098 18562
rect 18174 18510 18226 18562
rect 27134 18510 27186 18562
rect 40910 18510 40962 18562
rect 41582 18510 41634 18562
rect 42142 18510 42194 18562
rect 44046 18510 44098 18562
rect 47518 18510 47570 18562
rect 48862 18510 48914 18562
rect 51102 18510 51154 18562
rect 53454 18510 53506 18562
rect 55694 18510 55746 18562
rect 1710 18398 1762 18450
rect 18622 18398 18674 18450
rect 21870 18398 21922 18450
rect 26462 18398 26514 18450
rect 29710 18398 29762 18450
rect 34414 18398 34466 18450
rect 40238 18398 40290 18450
rect 41134 18398 41186 18450
rect 41918 18398 41970 18450
rect 42478 18398 42530 18450
rect 43934 18398 43986 18450
rect 44830 18398 44882 18450
rect 45278 18398 45330 18450
rect 46846 18398 46898 18450
rect 47406 18398 47458 18450
rect 48974 18398 49026 18450
rect 51326 18398 51378 18450
rect 53678 18398 53730 18450
rect 55134 18398 55186 18450
rect 57150 18398 57202 18450
rect 77310 18398 77362 18450
rect 78206 18398 78258 18450
rect 2494 18286 2546 18338
rect 19294 18286 19346 18338
rect 21422 18286 21474 18338
rect 22542 18286 22594 18338
rect 24670 18286 24722 18338
rect 25342 18286 25394 18338
rect 25678 18286 25730 18338
rect 29262 18286 29314 18338
rect 30382 18286 30434 18338
rect 32510 18286 32562 18338
rect 33182 18286 33234 18338
rect 33518 18286 33570 18338
rect 33742 18286 33794 18338
rect 38446 18286 38498 18338
rect 52446 18286 52498 18338
rect 56702 18286 56754 18338
rect 76974 18286 77026 18338
rect 18062 18174 18114 18226
rect 43710 18174 43762 18226
rect 4478 18006 4530 18058
rect 4582 18006 4634 18058
rect 4686 18006 4738 18058
rect 35198 18006 35250 18058
rect 35302 18006 35354 18058
rect 35406 18006 35458 18058
rect 65918 18006 65970 18058
rect 66022 18006 66074 18058
rect 66126 18006 66178 18058
rect 33854 17838 33906 17890
rect 37998 17838 38050 17890
rect 20638 17726 20690 17778
rect 21422 17726 21474 17778
rect 22430 17726 22482 17778
rect 28590 17726 28642 17778
rect 33406 17726 33458 17778
rect 33742 17726 33794 17778
rect 34750 17726 34802 17778
rect 35310 17726 35362 17778
rect 46062 17726 46114 17778
rect 50206 17726 50258 17778
rect 50766 17726 50818 17778
rect 52110 17726 52162 17778
rect 19070 17614 19122 17666
rect 19406 17614 19458 17666
rect 20190 17614 20242 17666
rect 20526 17614 20578 17666
rect 20750 17614 20802 17666
rect 21982 17614 22034 17666
rect 22318 17614 22370 17666
rect 28142 17614 28194 17666
rect 30718 17614 30770 17666
rect 31166 17614 31218 17666
rect 31390 17614 31442 17666
rect 35086 17614 35138 17666
rect 35534 17614 35586 17666
rect 35758 17614 35810 17666
rect 36430 17614 36482 17666
rect 37886 17614 37938 17666
rect 39006 17614 39058 17666
rect 39790 17614 39842 17666
rect 40574 17614 40626 17666
rect 41694 17614 41746 17666
rect 42926 17614 42978 17666
rect 43150 17614 43202 17666
rect 45278 17614 45330 17666
rect 45950 17614 46002 17666
rect 47294 17614 47346 17666
rect 48750 17614 48802 17666
rect 50990 17614 51042 17666
rect 51662 17614 51714 17666
rect 53230 17614 53282 17666
rect 54798 17614 54850 17666
rect 55694 17614 55746 17666
rect 56590 17614 56642 17666
rect 56814 17614 56866 17666
rect 58718 17614 58770 17666
rect 1710 17502 1762 17554
rect 18734 17502 18786 17554
rect 22542 17502 22594 17554
rect 25118 17502 25170 17554
rect 31278 17502 31330 17554
rect 34190 17502 34242 17554
rect 34302 17502 34354 17554
rect 34638 17502 34690 17554
rect 36990 17502 37042 17554
rect 37326 17502 37378 17554
rect 37550 17502 37602 17554
rect 38446 17502 38498 17554
rect 38782 17502 38834 17554
rect 39342 17502 39394 17554
rect 39678 17502 39730 17554
rect 40238 17502 40290 17554
rect 41470 17502 41522 17554
rect 46174 17502 46226 17554
rect 46958 17502 47010 17554
rect 48862 17502 48914 17554
rect 50878 17502 50930 17554
rect 53454 17502 53506 17554
rect 58830 17502 58882 17554
rect 70814 17502 70866 17554
rect 77646 17502 77698 17554
rect 77870 17502 77922 17554
rect 78206 17502 78258 17554
rect 2046 17390 2098 17442
rect 2494 17390 2546 17442
rect 19182 17390 19234 17442
rect 29262 17390 29314 17442
rect 32734 17390 32786 17442
rect 36094 17390 36146 17442
rect 37214 17390 37266 17442
rect 38558 17390 38610 17442
rect 39566 17390 39618 17442
rect 40350 17390 40402 17442
rect 43038 17390 43090 17442
rect 48414 17390 48466 17442
rect 55022 17390 55074 17442
rect 58382 17390 58434 17442
rect 70254 17390 70306 17442
rect 70478 17390 70530 17442
rect 19838 17222 19890 17274
rect 19942 17222 19994 17274
rect 20046 17222 20098 17274
rect 50558 17222 50610 17274
rect 50662 17222 50714 17274
rect 50766 17222 50818 17274
rect 22766 17054 22818 17106
rect 33406 17054 33458 17106
rect 35422 17054 35474 17106
rect 35982 17054 36034 17106
rect 37774 17054 37826 17106
rect 38670 17054 38722 17106
rect 39454 17054 39506 17106
rect 40462 17054 40514 17106
rect 41694 17054 41746 17106
rect 42030 17054 42082 17106
rect 42254 17054 42306 17106
rect 43934 17054 43986 17106
rect 50430 17054 50482 17106
rect 53454 17054 53506 17106
rect 56814 17054 56866 17106
rect 57150 17054 57202 17106
rect 77870 17054 77922 17106
rect 32286 16942 32338 16994
rect 36094 16942 36146 16994
rect 36990 16942 37042 16994
rect 37326 16942 37378 16994
rect 38782 16942 38834 16994
rect 39678 16942 39730 16994
rect 41134 16942 41186 16994
rect 41358 16942 41410 16994
rect 41470 16942 41522 16994
rect 42590 16942 42642 16994
rect 45278 16942 45330 16994
rect 47518 16942 47570 16994
rect 49086 16942 49138 16994
rect 51102 16942 51154 16994
rect 52334 16942 52386 16994
rect 54574 16942 54626 16994
rect 25342 16830 25394 16882
rect 28702 16830 28754 16882
rect 29486 16830 29538 16882
rect 33854 16830 33906 16882
rect 34302 16830 34354 16882
rect 35646 16830 35698 16882
rect 36206 16830 36258 16882
rect 37662 16830 37714 16882
rect 38222 16830 38274 16882
rect 39230 16830 39282 16882
rect 39790 16830 39842 16882
rect 41918 16830 41970 16882
rect 42702 16830 42754 16882
rect 46398 16830 46450 16882
rect 46734 16830 46786 16882
rect 47294 16830 47346 16882
rect 49310 16830 49362 16882
rect 51438 16830 51490 16882
rect 52558 16830 52610 16882
rect 54686 16830 54738 16882
rect 56030 16830 56082 16882
rect 77646 16830 77698 16882
rect 78206 16830 78258 16882
rect 26126 16718 26178 16770
rect 28254 16718 28306 16770
rect 31614 16718 31666 16770
rect 31950 16718 32002 16770
rect 47742 16718 47794 16770
rect 38334 16606 38386 16658
rect 4478 16438 4530 16490
rect 4582 16438 4634 16490
rect 4686 16438 4738 16490
rect 35198 16438 35250 16490
rect 35302 16438 35354 16490
rect 35406 16438 35458 16490
rect 65918 16438 65970 16490
rect 66022 16438 66074 16490
rect 66126 16438 66178 16490
rect 37438 16270 37490 16322
rect 37998 16270 38050 16322
rect 38334 16270 38386 16322
rect 25566 16158 25618 16210
rect 26686 16158 26738 16210
rect 28142 16158 28194 16210
rect 32062 16158 32114 16210
rect 35310 16158 35362 16210
rect 35646 16158 35698 16210
rect 36542 16158 36594 16210
rect 37326 16158 37378 16210
rect 37886 16158 37938 16210
rect 38334 16158 38386 16210
rect 38782 16158 38834 16210
rect 40686 16158 40738 16210
rect 41134 16158 41186 16210
rect 41582 16158 41634 16210
rect 43934 16158 43986 16210
rect 45054 16158 45106 16210
rect 45502 16158 45554 16210
rect 45838 16158 45890 16210
rect 51102 16158 51154 16210
rect 52110 16158 52162 16210
rect 26574 16046 26626 16098
rect 28254 16046 28306 16098
rect 28702 16046 28754 16098
rect 29150 16046 29202 16098
rect 32510 16046 32562 16098
rect 39230 16046 39282 16098
rect 39678 16046 39730 16098
rect 39790 16046 39842 16098
rect 43374 16046 43426 16098
rect 43710 16046 43762 16098
rect 46174 16046 46226 16098
rect 47854 16046 47906 16098
rect 48974 16046 49026 16098
rect 52670 16046 52722 16098
rect 53678 16046 53730 16098
rect 54574 16046 54626 16098
rect 54798 16046 54850 16098
rect 1710 15934 1762 15986
rect 2046 15934 2098 15986
rect 29934 15934 29986 15986
rect 33182 15934 33234 15986
rect 35982 15934 36034 15986
rect 41918 15934 41970 15986
rect 42478 15934 42530 15986
rect 43486 15934 43538 15986
rect 47182 15934 47234 15986
rect 49422 15934 49474 15986
rect 77870 15934 77922 15986
rect 78206 15934 78258 15986
rect 2494 15822 2546 15874
rect 26014 15822 26066 15874
rect 26350 15822 26402 15874
rect 26798 15822 26850 15874
rect 27246 15822 27298 15874
rect 27470 15822 27522 15874
rect 27582 15822 27634 15874
rect 27694 15822 27746 15874
rect 28030 15822 28082 15874
rect 39566 15822 39618 15874
rect 41806 15822 41858 15874
rect 42814 15822 42866 15874
rect 44046 15822 44098 15874
rect 46510 15822 46562 15874
rect 47966 15822 48018 15874
rect 50430 15822 50482 15874
rect 51662 15822 51714 15874
rect 53790 15822 53842 15874
rect 77646 15822 77698 15874
rect 19838 15654 19890 15706
rect 19942 15654 19994 15706
rect 20046 15654 20098 15706
rect 50558 15654 50610 15706
rect 50662 15654 50714 15706
rect 50766 15654 50818 15706
rect 33406 15486 33458 15538
rect 33518 15486 33570 15538
rect 38558 15486 38610 15538
rect 41134 15486 41186 15538
rect 41582 15486 41634 15538
rect 46174 15486 46226 15538
rect 46622 15486 46674 15538
rect 47182 15486 47234 15538
rect 47966 15486 48018 15538
rect 53454 15486 53506 15538
rect 2046 15374 2098 15426
rect 27918 15374 27970 15426
rect 31614 15374 31666 15426
rect 31950 15374 32002 15426
rect 39230 15374 39282 15426
rect 48750 15374 48802 15426
rect 50654 15374 50706 15426
rect 52782 15374 52834 15426
rect 54574 15374 54626 15426
rect 1710 15262 1762 15314
rect 31054 15262 31106 15314
rect 32958 15262 33010 15314
rect 33630 15262 33682 15314
rect 35086 15262 35138 15314
rect 39454 15262 39506 15314
rect 39902 15262 39954 15314
rect 40126 15262 40178 15314
rect 42142 15262 42194 15314
rect 45390 15262 45442 15314
rect 45502 15262 45554 15314
rect 49758 15262 49810 15314
rect 50878 15262 50930 15314
rect 52558 15262 52610 15314
rect 54462 15262 54514 15314
rect 2494 15150 2546 15202
rect 35870 15150 35922 15202
rect 37998 15150 38050 15202
rect 38446 15150 38498 15202
rect 38894 15150 38946 15202
rect 40014 15150 40066 15202
rect 42926 15150 42978 15202
rect 45054 15150 45106 15202
rect 51662 15150 51714 15202
rect 4478 14870 4530 14922
rect 4582 14870 4634 14922
rect 4686 14870 4738 14922
rect 35198 14870 35250 14922
rect 35302 14870 35354 14922
rect 35406 14870 35458 14922
rect 65918 14870 65970 14922
rect 66022 14870 66074 14922
rect 66126 14870 66178 14922
rect 30830 14702 30882 14754
rect 31502 14702 31554 14754
rect 52110 14702 52162 14754
rect 25678 14590 25730 14642
rect 27806 14590 27858 14642
rect 28478 14590 28530 14642
rect 29598 14590 29650 14642
rect 30830 14590 30882 14642
rect 34638 14590 34690 14642
rect 35198 14590 35250 14642
rect 35870 14590 35922 14642
rect 37214 14590 37266 14642
rect 38334 14590 38386 14642
rect 38670 14590 38722 14642
rect 39790 14590 39842 14642
rect 41918 14590 41970 14642
rect 42814 14590 42866 14642
rect 43374 14590 43426 14642
rect 43934 14590 43986 14642
rect 44270 14590 44322 14642
rect 46286 14590 46338 14642
rect 51102 14590 51154 14642
rect 53118 14590 53170 14642
rect 19966 14478 20018 14530
rect 24894 14478 24946 14530
rect 28254 14478 28306 14530
rect 29038 14478 29090 14530
rect 29486 14478 29538 14530
rect 29710 14478 29762 14530
rect 31838 14478 31890 14530
rect 35758 14478 35810 14530
rect 39006 14478 39058 14530
rect 42702 14478 42754 14530
rect 46510 14478 46562 14530
rect 47742 14478 47794 14530
rect 48750 14478 48802 14530
rect 51326 14478 51378 14530
rect 52670 14478 52722 14530
rect 19854 14366 19906 14418
rect 30046 14366 30098 14418
rect 32510 14366 32562 14418
rect 43262 14366 43314 14418
rect 48974 14366 49026 14418
rect 77870 14366 77922 14418
rect 78206 14366 78258 14418
rect 20078 14254 20130 14306
rect 20302 14254 20354 14306
rect 21422 14254 21474 14306
rect 30382 14254 30434 14306
rect 31278 14254 31330 14306
rect 35534 14254 35586 14306
rect 35982 14254 36034 14306
rect 42478 14254 42530 14306
rect 42926 14254 42978 14306
rect 48190 14254 48242 14306
rect 77646 14254 77698 14306
rect 19838 14086 19890 14138
rect 19942 14086 19994 14138
rect 20046 14086 20098 14138
rect 50558 14086 50610 14138
rect 50662 14086 50714 14138
rect 50766 14086 50818 14138
rect 2046 13918 2098 13970
rect 19182 13918 19234 13970
rect 22878 13918 22930 13970
rect 26238 13918 26290 13970
rect 27246 13918 27298 13970
rect 28814 13918 28866 13970
rect 29598 13918 29650 13970
rect 30942 13918 30994 13970
rect 33406 13918 33458 13970
rect 33518 13918 33570 13970
rect 33630 13918 33682 13970
rect 34078 13918 34130 13970
rect 35310 13918 35362 13970
rect 38558 13918 38610 13970
rect 39118 13918 39170 13970
rect 39342 13918 39394 13970
rect 41246 13918 41298 13970
rect 41470 13918 41522 13970
rect 45390 13918 45442 13970
rect 48078 13918 48130 13970
rect 48862 13918 48914 13970
rect 52670 13918 52722 13970
rect 55134 13918 55186 13970
rect 77870 13918 77922 13970
rect 18622 13806 18674 13858
rect 26462 13806 26514 13858
rect 26574 13806 26626 13858
rect 27022 13806 27074 13858
rect 28030 13806 28082 13858
rect 28478 13806 28530 13858
rect 28590 13806 28642 13858
rect 29038 13806 29090 13858
rect 29822 13806 29874 13858
rect 29934 13806 29986 13858
rect 31166 13806 31218 13858
rect 31726 13806 31778 13858
rect 32286 13806 32338 13858
rect 34638 13806 34690 13858
rect 34974 13806 35026 13858
rect 37774 13806 37826 13858
rect 38222 13806 38274 13858
rect 38334 13806 38386 13858
rect 38782 13806 38834 13858
rect 39566 13806 39618 13858
rect 54238 13806 54290 13858
rect 1710 13694 1762 13746
rect 18958 13694 19010 13746
rect 19518 13694 19570 13746
rect 19854 13694 19906 13746
rect 26910 13694 26962 13746
rect 27806 13694 27858 13746
rect 29374 13694 29426 13746
rect 31278 13694 31330 13746
rect 31614 13694 31666 13746
rect 31950 13694 32002 13746
rect 32174 13694 32226 13746
rect 32958 13694 33010 13746
rect 35646 13694 35698 13746
rect 37662 13694 37714 13746
rect 37998 13694 38050 13746
rect 39678 13694 39730 13746
rect 40798 13694 40850 13746
rect 42142 13694 42194 13746
rect 45278 13694 45330 13746
rect 52222 13694 52274 13746
rect 52894 13694 52946 13746
rect 53902 13694 53954 13746
rect 78206 13694 78258 13746
rect 2494 13582 2546 13634
rect 19070 13582 19122 13634
rect 20638 13582 20690 13634
rect 41358 13582 41410 13634
rect 42814 13582 42866 13634
rect 44942 13582 44994 13634
rect 46622 13582 46674 13634
rect 77646 13582 77698 13634
rect 32286 13470 32338 13522
rect 4478 13302 4530 13354
rect 4582 13302 4634 13354
rect 4686 13302 4738 13354
rect 35198 13302 35250 13354
rect 35302 13302 35354 13354
rect 35406 13302 35458 13354
rect 65918 13302 65970 13354
rect 66022 13302 66074 13354
rect 66126 13302 66178 13354
rect 20078 13134 20130 13186
rect 20414 13134 20466 13186
rect 12462 13022 12514 13074
rect 19518 13022 19570 13074
rect 25454 13022 25506 13074
rect 36430 13022 36482 13074
rect 37774 13022 37826 13074
rect 40238 13022 40290 13074
rect 42366 13022 42418 13074
rect 43150 13022 43202 13074
rect 74510 13022 74562 13074
rect 74734 13022 74786 13074
rect 74958 13022 75010 13074
rect 76302 13022 76354 13074
rect 16606 12910 16658 12962
rect 22542 12910 22594 12962
rect 28366 12910 28418 12962
rect 31614 12910 31666 12962
rect 32174 12910 32226 12962
rect 33630 12910 33682 12962
rect 38446 12910 38498 12962
rect 39566 12910 39618 12962
rect 42590 12910 42642 12962
rect 43038 12910 43090 12962
rect 43262 12910 43314 12962
rect 1710 12798 1762 12850
rect 2046 12798 2098 12850
rect 17390 12798 17442 12850
rect 23326 12798 23378 12850
rect 29486 12798 29538 12850
rect 31838 12798 31890 12850
rect 34302 12798 34354 12850
rect 37438 12798 37490 12850
rect 2494 12686 2546 12738
rect 20302 12686 20354 12738
rect 28590 12686 28642 12738
rect 29822 12686 29874 12738
rect 32286 12686 32338 12738
rect 32510 12686 32562 12738
rect 37102 12686 37154 12738
rect 37886 12686 37938 12738
rect 38782 12686 38834 12738
rect 75294 12686 75346 12738
rect 19838 12518 19890 12570
rect 19942 12518 19994 12570
rect 20046 12518 20098 12570
rect 50558 12518 50610 12570
rect 50662 12518 50714 12570
rect 50766 12518 50818 12570
rect 11902 12350 11954 12402
rect 15598 12350 15650 12402
rect 17390 12350 17442 12402
rect 18510 12350 18562 12402
rect 25454 12350 25506 12402
rect 35086 12350 35138 12402
rect 35198 12350 35250 12402
rect 35310 12350 35362 12402
rect 35758 12350 35810 12402
rect 41246 12350 41298 12402
rect 41582 12350 41634 12402
rect 17614 12238 17666 12290
rect 17838 12238 17890 12290
rect 18062 12238 18114 12290
rect 25678 12238 25730 12290
rect 26462 12238 26514 12290
rect 35646 12238 35698 12290
rect 36206 12238 36258 12290
rect 40910 12238 40962 12290
rect 41022 12238 41074 12290
rect 77534 12238 77586 12290
rect 9550 12126 9602 12178
rect 11678 12126 11730 12178
rect 12350 12126 12402 12178
rect 12686 12126 12738 12178
rect 21870 12126 21922 12178
rect 25230 12126 25282 12178
rect 29710 12126 29762 12178
rect 34638 12126 34690 12178
rect 37550 12126 37602 12178
rect 77758 12126 77810 12178
rect 9774 12014 9826 12066
rect 9886 12014 9938 12066
rect 11790 12014 11842 12066
rect 13358 12014 13410 12066
rect 17726 12014 17778 12066
rect 22542 12014 22594 12066
rect 24670 12014 24722 12066
rect 25342 12014 25394 12066
rect 26462 12014 26514 12066
rect 30382 12014 30434 12066
rect 32510 12014 32562 12066
rect 37214 12014 37266 12066
rect 38222 12014 38274 12066
rect 40350 12014 40402 12066
rect 26238 11902 26290 11954
rect 4478 11734 4530 11786
rect 4582 11734 4634 11786
rect 4686 11734 4738 11786
rect 35198 11734 35250 11786
rect 35302 11734 35354 11786
rect 35406 11734 35458 11786
rect 65918 11734 65970 11786
rect 66022 11734 66074 11786
rect 66126 11734 66178 11786
rect 37774 11566 37826 11618
rect 9774 11454 9826 11506
rect 11902 11454 11954 11506
rect 14478 11454 14530 11506
rect 18286 11454 18338 11506
rect 20750 11454 20802 11506
rect 22542 11454 22594 11506
rect 23214 11454 23266 11506
rect 26462 11454 26514 11506
rect 28590 11454 28642 11506
rect 30158 11454 30210 11506
rect 32398 11454 32450 11506
rect 32622 11454 32674 11506
rect 36430 11454 36482 11506
rect 76526 11454 76578 11506
rect 9102 11342 9154 11394
rect 13694 11342 13746 11394
rect 15374 11342 15426 11394
rect 19406 11342 19458 11394
rect 19854 11342 19906 11394
rect 19966 11342 20018 11394
rect 20414 11342 20466 11394
rect 22318 11342 22370 11394
rect 22990 11342 23042 11394
rect 25006 11342 25058 11394
rect 25454 11342 25506 11394
rect 25790 11342 25842 11394
rect 31950 11342 32002 11394
rect 32398 11342 32450 11394
rect 32622 11342 32674 11394
rect 32958 11342 33010 11394
rect 33630 11342 33682 11394
rect 37102 11342 37154 11394
rect 38670 11342 38722 11394
rect 78206 11342 78258 11394
rect 1710 11230 1762 11282
rect 2494 11230 2546 11282
rect 16046 11230 16098 11282
rect 22654 11230 22706 11282
rect 23326 11230 23378 11282
rect 24894 11230 24946 11282
rect 30382 11230 30434 11282
rect 31838 11230 31890 11282
rect 34302 11230 34354 11282
rect 37662 11230 37714 11282
rect 41358 11230 41410 11282
rect 44830 11230 44882 11282
rect 77198 11230 77250 11282
rect 77534 11230 77586 11282
rect 77870 11230 77922 11282
rect 2046 11118 2098 11170
rect 13470 11118 13522 11170
rect 13582 11118 13634 11170
rect 13918 11118 13970 11170
rect 19182 11118 19234 11170
rect 19294 11118 19346 11170
rect 19742 11118 19794 11170
rect 24782 11118 24834 11170
rect 30158 11118 30210 11170
rect 31726 11118 31778 11170
rect 33070 11118 33122 11170
rect 33182 11118 33234 11170
rect 37326 11118 37378 11170
rect 38334 11118 38386 11170
rect 44942 11118 44994 11170
rect 76974 11118 77026 11170
rect 19838 10950 19890 11002
rect 19942 10950 19994 11002
rect 20046 10950 20098 11002
rect 50558 10950 50610 11002
rect 50662 10950 50714 11002
rect 50766 10950 50818 11002
rect 2046 10782 2098 10834
rect 13246 10782 13298 10834
rect 17950 10782 18002 10834
rect 21646 10782 21698 10834
rect 25230 10782 25282 10834
rect 26462 10782 26514 10834
rect 26574 10782 26626 10834
rect 32510 10782 32562 10834
rect 39342 10782 39394 10834
rect 39454 10782 39506 10834
rect 39566 10782 39618 10834
rect 40238 10782 40290 10834
rect 13134 10670 13186 10722
rect 13358 10670 13410 10722
rect 19406 10670 19458 10722
rect 25678 10670 25730 10722
rect 40350 10670 40402 10722
rect 1710 10558 1762 10610
rect 9550 10558 9602 10610
rect 17726 10558 17778 10610
rect 17838 10558 17890 10610
rect 18398 10558 18450 10610
rect 18734 10558 18786 10610
rect 22654 10558 22706 10610
rect 25454 10558 25506 10610
rect 26014 10558 26066 10610
rect 26686 10558 26738 10610
rect 28478 10558 28530 10610
rect 36990 10558 37042 10610
rect 38894 10558 38946 10610
rect 41358 10558 41410 10610
rect 78206 10558 78258 10610
rect 2494 10446 2546 10498
rect 10334 10446 10386 10498
rect 12462 10446 12514 10498
rect 14142 10446 14194 10498
rect 14478 10446 14530 10498
rect 15150 10446 15202 10498
rect 15598 10446 15650 10498
rect 16046 10446 16098 10498
rect 22878 10446 22930 10498
rect 22990 10446 23042 10498
rect 25342 10446 25394 10498
rect 25790 10446 25842 10498
rect 26014 10446 26066 10498
rect 29150 10446 29202 10498
rect 31278 10446 31330 10498
rect 34078 10446 34130 10498
rect 41022 10446 41074 10498
rect 42142 10446 42194 10498
rect 44270 10446 44322 10498
rect 76526 10446 76578 10498
rect 4478 10166 4530 10218
rect 4582 10166 4634 10218
rect 4686 10166 4738 10218
rect 35198 10166 35250 10218
rect 35302 10166 35354 10218
rect 35406 10166 35458 10218
rect 65918 10166 65970 10218
rect 66022 10166 66074 10218
rect 66126 10166 66178 10218
rect 29150 9998 29202 10050
rect 33966 9998 34018 10050
rect 35758 9998 35810 10050
rect 37438 9998 37490 10050
rect 9438 9886 9490 9938
rect 12462 9886 12514 9938
rect 12686 9886 12738 9938
rect 15374 9886 15426 9938
rect 27806 9886 27858 9938
rect 34190 9886 34242 9938
rect 34974 9886 35026 9938
rect 40350 9886 40402 9938
rect 41022 9886 41074 9938
rect 44270 9886 44322 9938
rect 44942 9886 44994 9938
rect 11790 9774 11842 9826
rect 12014 9774 12066 9826
rect 12350 9774 12402 9826
rect 12798 9774 12850 9826
rect 20302 9774 20354 9826
rect 20862 9774 20914 9826
rect 22766 9774 22818 9826
rect 32398 9774 32450 9826
rect 33070 9774 33122 9826
rect 33294 9774 33346 9826
rect 35870 9774 35922 9826
rect 36206 9774 36258 9826
rect 37326 9774 37378 9826
rect 38110 9774 38162 9826
rect 38670 9774 38722 9826
rect 39230 9774 39282 9826
rect 39454 9774 39506 9826
rect 39790 9774 39842 9826
rect 41358 9774 41410 9826
rect 1710 9662 1762 9714
rect 2046 9662 2098 9714
rect 9550 9662 9602 9714
rect 11902 9662 11954 9714
rect 13470 9662 13522 9714
rect 14702 9662 14754 9714
rect 23662 9662 23714 9714
rect 26910 9662 26962 9714
rect 29486 9662 29538 9714
rect 32622 9662 32674 9714
rect 33182 9662 33234 9714
rect 33518 9662 33570 9714
rect 34638 9662 34690 9714
rect 36542 9662 36594 9714
rect 40686 9662 40738 9714
rect 42142 9662 42194 9714
rect 45278 9662 45330 9714
rect 77646 9662 77698 9714
rect 78206 9662 78258 9714
rect 2494 9550 2546 9602
rect 9326 9550 9378 9602
rect 13806 9550 13858 9602
rect 14478 9550 14530 9602
rect 14590 9550 14642 9602
rect 27246 9550 27298 9602
rect 28590 9550 28642 9602
rect 29262 9550 29314 9602
rect 29934 9550 29986 9602
rect 30382 9550 30434 9602
rect 31838 9550 31890 9602
rect 32174 9550 32226 9602
rect 32286 9550 32338 9602
rect 34190 9550 34242 9602
rect 34862 9550 34914 9602
rect 35758 9550 35810 9602
rect 36318 9550 36370 9602
rect 37438 9550 37490 9602
rect 37886 9550 37938 9602
rect 38782 9550 38834 9602
rect 38894 9550 38946 9602
rect 39678 9550 39730 9602
rect 75294 9550 75346 9602
rect 75742 9550 75794 9602
rect 76302 9550 76354 9602
rect 76974 9550 77026 9602
rect 77870 9550 77922 9602
rect 19838 9382 19890 9434
rect 19942 9382 19994 9434
rect 20046 9382 20098 9434
rect 50558 9382 50610 9434
rect 50662 9382 50714 9434
rect 50766 9382 50818 9434
rect 12574 9214 12626 9266
rect 13022 9214 13074 9266
rect 13358 9214 13410 9266
rect 16718 9214 16770 9266
rect 17614 9214 17666 9266
rect 18510 9214 18562 9266
rect 18622 9214 18674 9266
rect 18846 9214 18898 9266
rect 22318 9214 22370 9266
rect 24670 9214 24722 9266
rect 25230 9214 25282 9266
rect 25566 9214 25618 9266
rect 33518 9214 33570 9266
rect 43374 9214 43426 9266
rect 43486 9214 43538 9266
rect 43598 9214 43650 9266
rect 43934 9214 43986 9266
rect 44046 9214 44098 9266
rect 44158 9214 44210 9266
rect 44382 9214 44434 9266
rect 45614 9214 45666 9266
rect 46062 9214 46114 9266
rect 14478 9102 14530 9154
rect 17726 9102 17778 9154
rect 34974 9102 35026 9154
rect 38222 9102 38274 9154
rect 42702 9102 42754 9154
rect 44942 9102 44994 9154
rect 45054 9102 45106 9154
rect 9662 8990 9714 9042
rect 13694 8990 13746 9042
rect 17390 8990 17442 9042
rect 18398 8990 18450 9042
rect 19406 8990 19458 9042
rect 25902 8990 25954 9042
rect 29598 8990 29650 9042
rect 33182 8990 33234 9042
rect 34190 8990 34242 9042
rect 37438 8990 37490 9042
rect 41022 8990 41074 9042
rect 41134 8990 41186 9042
rect 41246 8990 41298 9042
rect 41470 8990 41522 9042
rect 41918 8990 41970 9042
rect 42142 8990 42194 9042
rect 42926 8990 42978 9042
rect 75294 8990 75346 9042
rect 77758 8990 77810 9042
rect 10334 8878 10386 8930
rect 20078 8878 20130 8930
rect 22990 8878 23042 8930
rect 23550 8878 23602 8930
rect 24334 8878 24386 8930
rect 26686 8878 26738 8930
rect 28814 8878 28866 8930
rect 30270 8878 30322 8930
rect 32398 8878 32450 8930
rect 37102 8878 37154 8930
rect 40350 8878 40402 8930
rect 44942 8766 44994 8818
rect 73390 8766 73442 8818
rect 75854 8766 75906 8818
rect 4478 8598 4530 8650
rect 4582 8598 4634 8650
rect 4686 8598 4738 8650
rect 35198 8598 35250 8650
rect 35302 8598 35354 8650
rect 35406 8598 35458 8650
rect 65918 8598 65970 8650
rect 66022 8598 66074 8650
rect 66126 8598 66178 8650
rect 28142 8430 28194 8482
rect 9326 8318 9378 8370
rect 17838 8318 17890 8370
rect 19966 8318 20018 8370
rect 22878 8318 22930 8370
rect 25006 8318 25058 8370
rect 26910 8318 26962 8370
rect 27358 8318 27410 8370
rect 27470 8318 27522 8370
rect 30158 8318 30210 8370
rect 30270 8318 30322 8370
rect 31166 8318 31218 8370
rect 34638 8318 34690 8370
rect 36430 8318 36482 8370
rect 38782 8318 38834 8370
rect 40126 8318 40178 8370
rect 42590 8318 42642 8370
rect 45278 8318 45330 8370
rect 74286 8318 74338 8370
rect 11006 8206 11058 8258
rect 11790 8206 11842 8258
rect 12014 8206 12066 8258
rect 12350 8206 12402 8258
rect 14926 8206 14978 8258
rect 18622 8206 18674 8258
rect 19854 8206 19906 8258
rect 20078 8206 20130 8258
rect 20526 8206 20578 8258
rect 22094 8206 22146 8258
rect 25566 8206 25618 8258
rect 25790 8206 25842 8258
rect 26238 8206 26290 8258
rect 26798 8206 26850 8258
rect 29934 8206 29986 8258
rect 32174 8206 32226 8258
rect 32958 8206 33010 8258
rect 33854 8206 33906 8258
rect 34750 8206 34802 8258
rect 38894 8206 38946 8258
rect 40686 8206 40738 8258
rect 40798 8206 40850 8258
rect 41806 8206 41858 8258
rect 43038 8206 43090 8258
rect 43598 8206 43650 8258
rect 75518 8206 75570 8258
rect 76862 8206 76914 8258
rect 78094 8206 78146 8258
rect 1710 8094 1762 8146
rect 2046 8094 2098 8146
rect 9438 8094 9490 8146
rect 11902 8094 11954 8146
rect 13022 8094 13074 8146
rect 14254 8094 14306 8146
rect 14590 8094 14642 8146
rect 15710 8094 15762 8146
rect 18846 8094 18898 8146
rect 21310 8094 21362 8146
rect 26574 8094 26626 8146
rect 28142 8094 28194 8146
rect 28254 8094 28306 8146
rect 31950 8094 32002 8146
rect 34302 8094 34354 8146
rect 35422 8094 35474 8146
rect 36094 8094 36146 8146
rect 37102 8094 37154 8146
rect 37774 8094 37826 8146
rect 39230 8094 39282 8146
rect 41134 8094 41186 8146
rect 42926 8094 42978 8146
rect 44270 8094 44322 8146
rect 77198 8094 77250 8146
rect 77534 8094 77586 8146
rect 77870 8094 77922 8146
rect 2494 7982 2546 8034
rect 9214 7982 9266 8034
rect 10670 7982 10722 8034
rect 11454 7982 11506 8034
rect 14030 7982 14082 8034
rect 18398 7982 18450 8034
rect 18510 7982 18562 8034
rect 19630 7982 19682 8034
rect 21646 7982 21698 8034
rect 25678 7982 25730 8034
rect 27022 7982 27074 8034
rect 27582 7982 27634 8034
rect 29710 7982 29762 8034
rect 30830 7982 30882 8034
rect 31726 7982 31778 8034
rect 33294 7982 33346 8034
rect 34526 7982 34578 8034
rect 34974 7982 35026 8034
rect 35758 7982 35810 8034
rect 36318 7982 36370 8034
rect 37438 7982 37490 8034
rect 38110 7982 38162 8034
rect 44158 7982 44210 8034
rect 44830 7982 44882 8034
rect 45950 7982 46002 8034
rect 46286 7982 46338 8034
rect 76302 7982 76354 8034
rect 19838 7814 19890 7866
rect 19942 7814 19994 7866
rect 20046 7814 20098 7866
rect 50558 7814 50610 7866
rect 50662 7814 50714 7866
rect 50766 7814 50818 7866
rect 2046 7646 2098 7698
rect 15710 7646 15762 7698
rect 16494 7646 16546 7698
rect 16942 7646 16994 7698
rect 17950 7646 18002 7698
rect 18398 7646 18450 7698
rect 19406 7646 19458 7698
rect 20302 7646 20354 7698
rect 20638 7646 20690 7698
rect 21422 7646 21474 7698
rect 25342 7646 25394 7698
rect 26350 7646 26402 7698
rect 26574 7646 26626 7698
rect 28142 7646 28194 7698
rect 29038 7646 29090 7698
rect 33406 7646 33458 7698
rect 38222 7646 38274 7698
rect 42926 7646 42978 7698
rect 66670 7646 66722 7698
rect 15822 7534 15874 7586
rect 19742 7534 19794 7586
rect 19966 7534 20018 7586
rect 26910 7534 26962 7586
rect 27694 7534 27746 7586
rect 30270 7534 30322 7586
rect 31278 7534 31330 7586
rect 32062 7534 32114 7586
rect 32286 7534 32338 7586
rect 34078 7534 34130 7586
rect 38782 7534 38834 7586
rect 39342 7534 39394 7586
rect 41246 7534 41298 7586
rect 43038 7534 43090 7586
rect 44494 7534 44546 7586
rect 46062 7534 46114 7586
rect 71710 7534 71762 7586
rect 1710 7422 1762 7474
rect 10558 7422 10610 7474
rect 14030 7422 14082 7474
rect 14254 7422 14306 7474
rect 14702 7422 14754 7474
rect 15486 7422 15538 7474
rect 18174 7422 18226 7474
rect 18846 7422 18898 7474
rect 21198 7422 21250 7474
rect 21870 7422 21922 7474
rect 27806 7422 27858 7474
rect 29598 7422 29650 7474
rect 29934 7422 29986 7474
rect 30942 7422 30994 7474
rect 33070 7422 33122 7474
rect 33742 7422 33794 7474
rect 34526 7422 34578 7474
rect 35310 7422 35362 7474
rect 40238 7422 40290 7474
rect 41582 7422 41634 7474
rect 41918 7422 41970 7474
rect 43934 7422 43986 7474
rect 46286 7422 46338 7474
rect 46846 7422 46898 7474
rect 67006 7422 67058 7474
rect 72382 7422 72434 7474
rect 75294 7422 75346 7474
rect 2494 7310 2546 7362
rect 9886 7310 9938 7362
rect 10334 7310 10386 7362
rect 11342 7310 11394 7362
rect 13470 7310 13522 7362
rect 14142 7310 14194 7362
rect 15262 7310 15314 7362
rect 18286 7310 18338 7362
rect 19630 7310 19682 7362
rect 22542 7310 22594 7362
rect 24670 7310 24722 7362
rect 25790 7310 25842 7362
rect 28478 7310 28530 7362
rect 28702 7310 28754 7362
rect 29374 7310 29426 7362
rect 31838 7310 31890 7362
rect 32398 7310 32450 7362
rect 37438 7310 37490 7362
rect 39902 7310 39954 7362
rect 41470 7310 41522 7362
rect 47518 7310 47570 7362
rect 48078 7310 48130 7362
rect 60174 7310 60226 7362
rect 68574 7310 68626 7362
rect 73950 7310 74002 7362
rect 27694 7198 27746 7250
rect 38558 7198 38610 7250
rect 76302 7198 76354 7250
rect 4478 7030 4530 7082
rect 4582 7030 4634 7082
rect 4686 7030 4738 7082
rect 35198 7030 35250 7082
rect 35302 7030 35354 7082
rect 35406 7030 35458 7082
rect 65918 7030 65970 7082
rect 66022 7030 66074 7082
rect 66126 7030 66178 7082
rect 9438 6862 9490 6914
rect 11230 6862 11282 6914
rect 8318 6750 8370 6802
rect 8430 6750 8482 6802
rect 8990 6750 9042 6802
rect 9102 6750 9154 6802
rect 9774 6750 9826 6802
rect 11118 6750 11170 6802
rect 19294 6750 19346 6802
rect 20750 6750 20802 6802
rect 23886 6750 23938 6802
rect 26126 6750 26178 6802
rect 33294 6750 33346 6802
rect 40126 6750 40178 6802
rect 42254 6750 42306 6802
rect 10334 6638 10386 6690
rect 10894 6638 10946 6690
rect 13806 6638 13858 6690
rect 15038 6638 15090 6690
rect 16382 6638 16434 6690
rect 17166 6638 17218 6690
rect 20078 6638 20130 6690
rect 22430 6638 22482 6690
rect 26014 6638 26066 6690
rect 26238 6638 26290 6690
rect 26686 6638 26738 6690
rect 27246 6638 27298 6690
rect 28366 6638 28418 6690
rect 28590 6638 28642 6690
rect 29822 6638 29874 6690
rect 30494 6638 30546 6690
rect 34414 6638 34466 6690
rect 34638 6638 34690 6690
rect 34862 6638 34914 6690
rect 35870 6638 35922 6690
rect 37326 6638 37378 6690
rect 37998 6638 38050 6690
rect 40462 6638 40514 6690
rect 44270 6638 44322 6690
rect 46510 6638 46562 6690
rect 47070 6638 47122 6690
rect 50206 6638 50258 6690
rect 51102 6638 51154 6690
rect 51550 6638 51602 6690
rect 59502 6638 59554 6690
rect 60062 6638 60114 6690
rect 60510 6638 60562 6690
rect 63422 6638 63474 6690
rect 67902 6638 67954 6690
rect 68350 6638 68402 6690
rect 71262 6638 71314 6690
rect 74510 6638 74562 6690
rect 74734 6638 74786 6690
rect 76190 6638 76242 6690
rect 76414 6638 76466 6690
rect 10110 6526 10162 6578
rect 16158 6526 16210 6578
rect 19854 6526 19906 6578
rect 23214 6526 23266 6578
rect 23326 6526 23378 6578
rect 23438 6526 23490 6578
rect 23774 6526 23826 6578
rect 25342 6526 25394 6578
rect 25678 6526 25730 6578
rect 28030 6526 28082 6578
rect 29262 6526 29314 6578
rect 29374 6526 29426 6578
rect 31166 6526 31218 6578
rect 33742 6526 33794 6578
rect 33966 6526 34018 6578
rect 35086 6526 35138 6578
rect 36094 6526 36146 6578
rect 41582 6526 41634 6578
rect 44158 6526 44210 6578
rect 46062 6526 46114 6578
rect 48638 6526 48690 6578
rect 50766 6526 50818 6578
rect 77198 6526 77250 6578
rect 77534 6526 77586 6578
rect 77870 6526 77922 6578
rect 78206 6526 78258 6578
rect 7422 6414 7474 6466
rect 7870 6414 7922 6466
rect 8206 6414 8258 6466
rect 8878 6414 8930 6466
rect 9550 6414 9602 6466
rect 12126 6414 12178 6466
rect 12574 6414 12626 6466
rect 13022 6414 13074 6466
rect 13470 6414 13522 6466
rect 14478 6414 14530 6466
rect 14702 6414 14754 6466
rect 15710 6414 15762 6466
rect 21534 6414 21586 6466
rect 21982 6414 22034 6466
rect 22206 6414 22258 6466
rect 23998 6414 24050 6466
rect 24670 6414 24722 6466
rect 25118 6414 25170 6466
rect 26910 6414 26962 6466
rect 27806 6414 27858 6466
rect 29038 6414 29090 6466
rect 30046 6414 30098 6466
rect 33854 6414 33906 6466
rect 34750 6414 34802 6466
rect 36430 6414 36482 6466
rect 46622 6414 46674 6466
rect 49086 6414 49138 6466
rect 52110 6414 52162 6466
rect 56814 6414 56866 6466
rect 61518 6414 61570 6466
rect 64430 6414 64482 6466
rect 67342 6414 67394 6466
rect 69358 6414 69410 6466
rect 72270 6414 72322 6466
rect 75070 6414 75122 6466
rect 75518 6414 75570 6466
rect 76750 6414 76802 6466
rect 19838 6246 19890 6298
rect 19942 6246 19994 6298
rect 20046 6246 20098 6298
rect 50558 6246 50610 6298
rect 50662 6246 50714 6298
rect 50766 6246 50818 6298
rect 2046 6078 2098 6130
rect 14254 6078 14306 6130
rect 15598 6078 15650 6130
rect 18062 6078 18114 6130
rect 18846 6078 18898 6130
rect 19854 6078 19906 6130
rect 20190 6078 20242 6130
rect 8990 5966 9042 6018
rect 13582 5966 13634 6018
rect 13918 5966 13970 6018
rect 14702 5966 14754 6018
rect 17502 5966 17554 6018
rect 17838 5966 17890 6018
rect 22094 6078 22146 6130
rect 22654 6078 22706 6130
rect 23550 6078 23602 6130
rect 24782 6078 24834 6130
rect 25902 6078 25954 6130
rect 26350 6078 26402 6130
rect 26798 6078 26850 6130
rect 27582 6078 27634 6130
rect 28030 6078 28082 6130
rect 22206 5966 22258 6018
rect 22766 5966 22818 6018
rect 23886 5966 23938 6018
rect 24110 5966 24162 6018
rect 27470 5966 27522 6018
rect 28926 5966 28978 6018
rect 29038 6022 29090 6074
rect 29262 6078 29314 6130
rect 29822 6078 29874 6130
rect 31390 6078 31442 6130
rect 33182 6078 33234 6130
rect 33294 6078 33346 6130
rect 35198 6078 35250 6130
rect 44942 6078 44994 6130
rect 56030 6078 56082 6130
rect 63198 6078 63250 6130
rect 63870 6078 63922 6130
rect 78318 6078 78370 6130
rect 29486 5966 29538 6018
rect 30494 5966 30546 6018
rect 31838 5966 31890 6018
rect 32062 5966 32114 6018
rect 34750 5966 34802 6018
rect 35646 5966 35698 6018
rect 37662 5966 37714 6018
rect 39342 5966 39394 6018
rect 40126 5966 40178 6018
rect 42590 5966 42642 6018
rect 45614 5966 45666 6018
rect 47742 5966 47794 6018
rect 1710 5854 1762 5906
rect 8654 5854 8706 5906
rect 9886 5854 9938 5906
rect 10222 5854 10274 5906
rect 14478 5854 14530 5906
rect 15374 5854 15426 5906
rect 17726 5854 17778 5906
rect 21198 5854 21250 5906
rect 21534 5854 21586 5906
rect 21870 5854 21922 5906
rect 22542 5854 22594 5906
rect 25678 5854 25730 5906
rect 26574 5854 26626 5906
rect 28366 5854 28418 5906
rect 28590 5854 28642 5906
rect 30158 5854 30210 5906
rect 30830 5854 30882 5906
rect 31054 5854 31106 5906
rect 32622 5854 32674 5906
rect 33070 5854 33122 5906
rect 33742 5854 33794 5906
rect 34414 5854 34466 5906
rect 35086 5854 35138 5906
rect 37102 5854 37154 5906
rect 39230 5854 39282 5906
rect 42478 5854 42530 5906
rect 44494 5854 44546 5906
rect 46958 5854 47010 5906
rect 47966 5854 48018 5906
rect 48750 5854 48802 5906
rect 49198 5854 49250 5906
rect 56926 5854 56978 5906
rect 59838 5854 59890 5906
rect 64430 5854 64482 5906
rect 67342 5854 67394 5906
rect 71038 5854 71090 5906
rect 72270 5854 72322 5906
rect 75182 5854 75234 5906
rect 2494 5742 2546 5794
rect 6190 5742 6242 5794
rect 6638 5742 6690 5794
rect 7086 5742 7138 5794
rect 7534 5742 7586 5794
rect 7982 5742 8034 5794
rect 8430 5742 8482 5794
rect 8766 5742 8818 5794
rect 10894 5742 10946 5794
rect 13022 5742 13074 5794
rect 14366 5742 14418 5794
rect 16494 5742 16546 5794
rect 16942 5742 16994 5794
rect 17390 5742 17442 5794
rect 18398 5742 18450 5794
rect 19294 5742 19346 5794
rect 20974 5742 21026 5794
rect 21310 5742 21362 5794
rect 23998 5742 24050 5794
rect 25454 5742 25506 5794
rect 26462 5742 26514 5794
rect 30270 5742 30322 5794
rect 34190 5742 34242 5794
rect 34526 5742 34578 5794
rect 40462 5742 40514 5794
rect 41022 5742 41074 5794
rect 41470 5742 41522 5794
rect 42254 5742 42306 5794
rect 46734 5742 46786 5794
rect 49758 5742 49810 5794
rect 50206 5742 50258 5794
rect 50990 5742 51042 5794
rect 51438 5742 51490 5794
rect 52558 5742 52610 5794
rect 65550 5742 65602 5794
rect 68910 5742 68962 5794
rect 70478 5742 70530 5794
rect 71710 5742 71762 5794
rect 7422 5630 7474 5682
rect 8094 5630 8146 5682
rect 15710 5630 15762 5682
rect 26014 5630 26066 5682
rect 27694 5630 27746 5682
rect 31726 5630 31778 5682
rect 47294 5630 47346 5682
rect 57934 5630 57986 5682
rect 60846 5630 60898 5682
rect 73278 5630 73330 5682
rect 76190 5630 76242 5682
rect 4478 5462 4530 5514
rect 4582 5462 4634 5514
rect 4686 5462 4738 5514
rect 35198 5462 35250 5514
rect 35302 5462 35354 5514
rect 35406 5462 35458 5514
rect 65918 5462 65970 5514
rect 66022 5462 66074 5514
rect 66126 5462 66178 5514
rect 7198 5294 7250 5346
rect 7870 5294 7922 5346
rect 21758 5294 21810 5346
rect 22094 5294 22146 5346
rect 27246 5294 27298 5346
rect 29598 5294 29650 5346
rect 30270 5294 30322 5346
rect 30942 5294 30994 5346
rect 37102 5294 37154 5346
rect 37438 5294 37490 5346
rect 50318 5294 50370 5346
rect 50990 5294 51042 5346
rect 51998 5294 52050 5346
rect 67342 5294 67394 5346
rect 67566 5294 67618 5346
rect 74846 5294 74898 5346
rect 7422 5182 7474 5234
rect 7870 5182 7922 5234
rect 8318 5182 8370 5234
rect 10222 5182 10274 5234
rect 10782 5182 10834 5234
rect 10894 5182 10946 5234
rect 13582 5182 13634 5234
rect 15150 5182 15202 5234
rect 17278 5182 17330 5234
rect 17950 5182 18002 5234
rect 18622 5182 18674 5234
rect 19966 5182 20018 5234
rect 21534 5182 21586 5234
rect 23998 5182 24050 5234
rect 26126 5182 26178 5234
rect 26686 5182 26738 5234
rect 27134 5182 27186 5234
rect 31838 5182 31890 5234
rect 46958 5182 47010 5234
rect 50878 5182 50930 5234
rect 51326 5182 51378 5234
rect 54014 5182 54066 5234
rect 55246 5182 55298 5234
rect 58158 5182 58210 5234
rect 64430 5182 64482 5234
rect 66446 5182 66498 5234
rect 67118 5182 67170 5234
rect 69358 5182 69410 5234
rect 74398 5182 74450 5234
rect 74622 5182 74674 5234
rect 76638 5182 76690 5234
rect 1710 5070 1762 5122
rect 2494 5070 2546 5122
rect 6190 5070 6242 5122
rect 6526 5070 6578 5122
rect 8766 5070 8818 5122
rect 8878 5070 8930 5122
rect 9550 5070 9602 5122
rect 11566 5070 11618 5122
rect 11902 5070 11954 5122
rect 12462 5070 12514 5122
rect 13022 5070 13074 5122
rect 13470 5070 13522 5122
rect 14142 5070 14194 5122
rect 14366 5070 14418 5122
rect 17838 5070 17890 5122
rect 18846 5070 18898 5122
rect 19518 5070 19570 5122
rect 22878 5070 22930 5122
rect 23214 5070 23266 5122
rect 27918 5070 27970 5122
rect 28366 5070 28418 5122
rect 29262 5070 29314 5122
rect 29486 5070 29538 5122
rect 30158 5070 30210 5122
rect 30830 5070 30882 5122
rect 31278 5070 31330 5122
rect 32398 5070 32450 5122
rect 32622 5070 32674 5122
rect 36430 5070 36482 5122
rect 37102 5070 37154 5122
rect 37438 5070 37490 5122
rect 37550 5070 37602 5122
rect 38894 5070 38946 5122
rect 42030 5070 42082 5122
rect 42478 5070 42530 5122
rect 44830 5070 44882 5122
rect 46846 5070 46898 5122
rect 49310 5070 49362 5122
rect 49870 5070 49922 5122
rect 50430 5070 50482 5122
rect 51774 5070 51826 5122
rect 52782 5070 52834 5122
rect 54238 5070 54290 5122
rect 57150 5070 57202 5122
rect 60510 5070 60562 5122
rect 63534 5070 63586 5122
rect 68350 5070 68402 5122
rect 71374 5070 71426 5122
rect 75630 5070 75682 5122
rect 76302 5070 76354 5122
rect 77198 5070 77250 5122
rect 77758 5070 77810 5122
rect 2046 4958 2098 5010
rect 6750 4958 6802 5010
rect 9214 4958 9266 5010
rect 9886 4958 9938 5010
rect 10670 4958 10722 5010
rect 12574 4958 12626 5010
rect 13694 4958 13746 5010
rect 18174 4958 18226 5010
rect 18510 4958 18562 5010
rect 20414 4958 20466 5010
rect 22542 4958 22594 5010
rect 27582 4958 27634 5010
rect 28590 4958 28642 5010
rect 30718 4958 30770 5010
rect 32734 4958 32786 5010
rect 35870 4958 35922 5010
rect 38334 4958 38386 5010
rect 39006 4958 39058 5010
rect 39678 4958 39730 5010
rect 40014 4958 40066 5010
rect 40574 4958 40626 5010
rect 43598 4958 43650 5010
rect 45390 4958 45442 5010
rect 47406 4958 47458 5010
rect 48974 4958 49026 5010
rect 49646 4958 49698 5010
rect 77534 4958 77586 5010
rect 5182 4846 5234 4898
rect 8654 4846 8706 4898
rect 10110 4846 10162 4898
rect 11790 4846 11842 4898
rect 12350 4846 12402 4898
rect 20862 4846 20914 4898
rect 21870 4846 21922 4898
rect 27022 4846 27074 4898
rect 30046 4846 30098 4898
rect 33966 4846 34018 4898
rect 42926 4846 42978 4898
rect 53342 4846 53394 4898
rect 61518 4846 61570 4898
rect 67454 4846 67506 4898
rect 72270 4846 72322 4898
rect 75182 4846 75234 4898
rect 19838 4678 19890 4730
rect 19942 4678 19994 4730
rect 20046 4678 20098 4730
rect 50558 4678 50610 4730
rect 50662 4678 50714 4730
rect 50766 4678 50818 4730
rect 6190 4510 6242 4562
rect 7534 4510 7586 4562
rect 8206 4510 8258 4562
rect 8990 4510 9042 4562
rect 9998 4510 10050 4562
rect 15374 4510 15426 4562
rect 15822 4510 15874 4562
rect 16718 4510 16770 4562
rect 17838 4510 17890 4562
rect 18622 4510 18674 4562
rect 19294 4510 19346 4562
rect 22654 4510 22706 4562
rect 40238 4510 40290 4562
rect 40910 4510 40962 4562
rect 43822 4510 43874 4562
rect 48750 4510 48802 4562
rect 55918 4510 55970 4562
rect 62526 4510 62578 4562
rect 63198 4510 63250 4562
rect 63534 4510 63586 4562
rect 71038 4510 71090 4562
rect 78206 4510 78258 4562
rect 5182 4398 5234 4450
rect 5854 4398 5906 4450
rect 6974 4398 7026 4450
rect 7646 4398 7698 4450
rect 8318 4398 8370 4450
rect 10334 4398 10386 4450
rect 10670 4398 10722 4450
rect 11790 4398 11842 4450
rect 14814 4398 14866 4450
rect 15486 4398 15538 4450
rect 16158 4398 16210 4450
rect 18286 4398 18338 4450
rect 19630 4398 19682 4450
rect 19966 4398 20018 4450
rect 21310 4398 21362 4450
rect 21758 4398 21810 4450
rect 21982 4398 22034 4450
rect 23326 4398 23378 4450
rect 23662 4398 23714 4450
rect 23998 4398 24050 4450
rect 24334 4398 24386 4450
rect 24670 4398 24722 4450
rect 29262 4398 29314 4450
rect 31278 4398 31330 4450
rect 34078 4398 34130 4450
rect 37102 4398 37154 4450
rect 39118 4398 39170 4450
rect 41022 4398 41074 4450
rect 42814 4398 42866 4450
rect 45390 4398 45442 4450
rect 46398 4398 46450 4450
rect 46622 4398 46674 4450
rect 6750 4286 6802 4338
rect 7310 4286 7362 4338
rect 7982 4286 8034 4338
rect 8766 4286 8818 4338
rect 9774 4286 9826 4338
rect 11006 4286 11058 4338
rect 14590 4286 14642 4338
rect 15150 4286 15202 4338
rect 16494 4286 16546 4338
rect 17614 4286 17666 4338
rect 19070 4286 19122 4338
rect 20302 4286 20354 4338
rect 20974 4286 21026 4338
rect 22430 4286 22482 4338
rect 22990 4286 23042 4338
rect 25230 4286 25282 4338
rect 28702 4286 28754 4338
rect 30718 4286 30770 4338
rect 33406 4286 33458 4338
rect 38110 4286 38162 4338
rect 38670 4286 38722 4338
rect 41918 4286 41970 4338
rect 42254 4286 42306 4338
rect 44270 4286 44322 4338
rect 47294 4286 47346 4338
rect 49086 4286 49138 4338
rect 49534 4286 49586 4338
rect 52894 4286 52946 4338
rect 56590 4286 56642 4338
rect 61630 4286 61682 4338
rect 64542 4286 64594 4338
rect 67342 4286 67394 4338
rect 72270 4286 72322 4338
rect 75406 4286 75458 4338
rect 2158 4174 2210 4226
rect 4734 4174 4786 4226
rect 5630 4174 5682 4226
rect 13918 4174 13970 4226
rect 21086 4174 21138 4226
rect 21646 4174 21698 4226
rect 23214 4174 23266 4226
rect 26014 4174 26066 4226
rect 28142 4174 28194 4226
rect 31838 4174 31890 4226
rect 36206 4174 36258 4226
rect 41470 4174 41522 4226
rect 52558 4174 52610 4226
rect 65550 4174 65602 4226
rect 70478 4174 70530 4226
rect 71710 4174 71762 4226
rect 16830 4062 16882 4114
rect 17950 4062 18002 4114
rect 20302 4062 20354 4114
rect 20638 4062 20690 4114
rect 50542 4062 50594 4114
rect 53902 4062 53954 4114
rect 57598 4062 57650 4114
rect 59726 4062 59778 4114
rect 68350 4062 68402 4114
rect 73278 4062 73330 4114
rect 76190 4062 76242 4114
rect 4478 3894 4530 3946
rect 4582 3894 4634 3946
rect 4686 3894 4738 3946
rect 35198 3894 35250 3946
rect 35302 3894 35354 3946
rect 35406 3894 35458 3946
rect 65918 3894 65970 3946
rect 66022 3894 66074 3946
rect 66126 3894 66178 3946
rect 11566 3726 11618 3778
rect 13694 3726 13746 3778
rect 23326 3726 23378 3778
rect 39118 3726 39170 3778
rect 47630 3726 47682 3778
rect 67454 3726 67506 3778
rect 75070 3726 75122 3778
rect 11118 3614 11170 3666
rect 23102 3614 23154 3666
rect 32510 3614 32562 3666
rect 42814 3614 42866 3666
rect 45726 3614 45778 3666
rect 47406 3614 47458 3666
rect 47966 3614 48018 3666
rect 54238 3614 54290 3666
rect 56030 3614 56082 3666
rect 58046 3614 58098 3666
rect 59054 3614 59106 3666
rect 63870 3614 63922 3666
rect 65662 3614 65714 3666
rect 69806 3614 69858 3666
rect 71262 3614 71314 3666
rect 73614 3614 73666 3666
rect 4734 3502 4786 3554
rect 5742 3502 5794 3554
rect 6414 3502 6466 3554
rect 7198 3502 7250 3554
rect 7870 3502 7922 3554
rect 8430 3502 8482 3554
rect 9550 3502 9602 3554
rect 10222 3502 10274 3554
rect 10894 3502 10946 3554
rect 11566 3502 11618 3554
rect 13358 3502 13410 3554
rect 13582 3502 13634 3554
rect 14142 3502 14194 3554
rect 14702 3502 14754 3554
rect 15374 3502 15426 3554
rect 16158 3502 16210 3554
rect 17166 3502 17218 3554
rect 17838 3502 17890 3554
rect 18622 3502 18674 3554
rect 19294 3502 19346 3554
rect 19854 3502 19906 3554
rect 20974 3502 21026 3554
rect 21758 3502 21810 3554
rect 22318 3502 22370 3554
rect 22990 3502 23042 3554
rect 23662 3502 23714 3554
rect 24782 3502 24834 3554
rect 25342 3502 25394 3554
rect 26126 3502 26178 3554
rect 27582 3502 27634 3554
rect 30718 3502 30770 3554
rect 31390 3502 31442 3554
rect 33966 3502 34018 3554
rect 35086 3502 35138 3554
rect 36878 3502 36930 3554
rect 39230 3502 39282 3554
rect 41358 3502 41410 3554
rect 43038 3502 43090 3554
rect 43710 3502 43762 3554
rect 45278 3502 45330 3554
rect 48526 3502 48578 3554
rect 49198 3502 49250 3554
rect 49870 3502 49922 3554
rect 50542 3502 50594 3554
rect 51662 3502 51714 3554
rect 52334 3502 52386 3554
rect 53006 3502 53058 3554
rect 53678 3502 53730 3554
rect 55470 3502 55522 3554
rect 60958 3502 61010 3554
rect 61854 3502 61906 3554
rect 63086 3502 63138 3554
rect 66446 3502 66498 3554
rect 70254 3502 70306 3554
rect 74062 3502 74114 3554
rect 76974 3502 77026 3554
rect 77870 3502 77922 3554
rect 1710 3390 1762 3442
rect 2046 3390 2098 3442
rect 2382 3390 2434 3442
rect 2718 3390 2770 3442
rect 3166 3390 3218 3442
rect 3726 3390 3778 3442
rect 3950 3390 4002 3442
rect 4286 3390 4338 3442
rect 4958 3390 5010 3442
rect 6078 3390 6130 3442
rect 6750 3390 6802 3442
rect 7422 3390 7474 3442
rect 8094 3390 8146 3442
rect 9886 3390 9938 3442
rect 10558 3390 10610 3442
rect 11230 3390 11282 3442
rect 11902 3390 11954 3442
rect 12238 3390 12290 3442
rect 12574 3390 12626 3442
rect 15038 3390 15090 3442
rect 15710 3390 15762 3442
rect 16382 3390 16434 3442
rect 17502 3390 17554 3442
rect 18174 3390 18226 3442
rect 19518 3390 19570 3442
rect 20190 3390 20242 3442
rect 21310 3390 21362 3442
rect 21982 3390 22034 3442
rect 23998 3390 24050 3442
rect 26462 3390 26514 3442
rect 26798 3390 26850 3442
rect 27134 3390 27186 3442
rect 28590 3390 28642 3442
rect 29262 3390 29314 3442
rect 29598 3390 29650 3442
rect 29934 3390 29986 3442
rect 30270 3390 30322 3442
rect 30942 3390 30994 3442
rect 32174 3390 32226 3442
rect 33630 3390 33682 3442
rect 35310 3390 35362 3442
rect 36654 3390 36706 3442
rect 37662 3390 37714 3442
rect 41470 3390 41522 3442
rect 42478 3390 42530 3442
rect 44382 3390 44434 3442
rect 45166 3390 45218 3442
rect 48302 3390 48354 3442
rect 48974 3390 49026 3442
rect 49646 3390 49698 3442
rect 50318 3390 50370 3442
rect 51214 3390 51266 3442
rect 52110 3390 52162 3442
rect 52782 3390 52834 3442
rect 53454 3390 53506 3442
rect 77310 3390 77362 3442
rect 78206 3390 78258 3442
rect 8766 3278 8818 3330
rect 14366 3278 14418 3330
rect 18846 3278 18898 3330
rect 22654 3278 22706 3330
rect 25902 3278 25954 3330
rect 27806 3278 27858 3330
rect 28926 3278 28978 3330
rect 31614 3278 31666 3330
rect 19838 3110 19890 3162
rect 19942 3110 19994 3162
rect 20046 3110 20098 3162
rect 50558 3110 50610 3162
rect 50662 3110 50714 3162
rect 50766 3110 50818 3162
rect 7198 2942 7250 2994
rect 9662 2942 9714 2994
rect 12238 2942 12290 2994
rect 16382 2942 16434 2994
rect 29150 1374 29202 1426
rect 29710 1374 29762 1426
<< metal2 >>
rect 448 79200 560 80000
rect 1120 79200 1232 80000
rect 1792 79200 1904 80000
rect 2464 79200 2576 80000
rect 3136 79200 3248 80000
rect 3808 79200 3920 80000
rect 4480 79200 4592 80000
rect 5152 79200 5264 80000
rect 5824 79200 5936 80000
rect 6496 79200 6608 80000
rect 7168 79200 7280 80000
rect 7840 79200 7952 80000
rect 8512 79200 8624 80000
rect 9184 79200 9296 80000
rect 9856 79200 9968 80000
rect 10528 79200 10640 80000
rect 11200 79200 11312 80000
rect 11872 79200 11984 80000
rect 12544 79200 12656 80000
rect 13216 79200 13328 80000
rect 13888 79200 14000 80000
rect 14560 79200 14672 80000
rect 15232 79200 15344 80000
rect 15904 79200 16016 80000
rect 16576 79200 16688 80000
rect 17248 79200 17360 80000
rect 17920 79200 18032 80000
rect 18592 79200 18704 80000
rect 19264 79200 19376 80000
rect 19936 79200 20048 80000
rect 20608 79200 20720 80000
rect 21280 79200 21392 80000
rect 21952 79200 22064 80000
rect 22624 79200 22736 80000
rect 23296 79200 23408 80000
rect 23968 79200 24080 80000
rect 24640 79200 24752 80000
rect 25312 79200 25424 80000
rect 25984 79200 26096 80000
rect 26656 79200 26768 80000
rect 27328 79200 27440 80000
rect 28000 79200 28112 80000
rect 28672 79200 28784 80000
rect 29344 79200 29456 80000
rect 30016 79200 30128 80000
rect 30688 79200 30800 80000
rect 31360 79200 31472 80000
rect 32032 79200 32144 80000
rect 32704 79200 32816 80000
rect 33376 79200 33488 80000
rect 34048 79200 34160 80000
rect 34720 79200 34832 80000
rect 35392 79200 35504 80000
rect 36064 79200 36176 80000
rect 36736 79200 36848 80000
rect 37408 79200 37520 80000
rect 38080 79200 38192 80000
rect 38752 79200 38864 80000
rect 39424 79200 39536 80000
rect 40096 79200 40208 80000
rect 40768 79200 40880 80000
rect 41440 79200 41552 80000
rect 42112 79200 42224 80000
rect 42784 79200 42896 80000
rect 43456 79200 43568 80000
rect 44128 79200 44240 80000
rect 44800 79200 44912 80000
rect 45472 79200 45584 80000
rect 46144 79200 46256 80000
rect 46816 79200 46928 80000
rect 47488 79200 47600 80000
rect 48160 79200 48272 80000
rect 48832 79200 48944 80000
rect 49504 79200 49616 80000
rect 50176 79200 50288 80000
rect 50848 79200 50960 80000
rect 51520 79200 51632 80000
rect 52192 79200 52304 80000
rect 52864 79200 52976 80000
rect 53536 79200 53648 80000
rect 54208 79200 54320 80000
rect 54880 79200 54992 80000
rect 55552 79200 55664 80000
rect 56224 79200 56336 80000
rect 56896 79200 57008 80000
rect 57568 79200 57680 80000
rect 58240 79200 58352 80000
rect 58912 79200 59024 80000
rect 59584 79200 59696 80000
rect 60256 79200 60368 80000
rect 60928 79200 61040 80000
rect 61600 79200 61712 80000
rect 62272 79200 62384 80000
rect 62944 79200 63056 80000
rect 63616 79200 63728 80000
rect 64288 79200 64400 80000
rect 64960 79200 65072 80000
rect 65632 79200 65744 80000
rect 66304 79200 66416 80000
rect 66976 79200 67088 80000
rect 67648 79200 67760 80000
rect 68320 79200 68432 80000
rect 68992 79200 69104 80000
rect 69664 79200 69776 80000
rect 70336 79200 70448 80000
rect 71008 79200 71120 80000
rect 71680 79200 71792 80000
rect 72352 79200 72464 80000
rect 73024 79200 73136 80000
rect 73696 79200 73808 80000
rect 74368 79200 74480 80000
rect 75040 79200 75152 80000
rect 75712 79200 75824 80000
rect 76384 79200 76496 80000
rect 77056 79200 77168 80000
rect 77728 79200 77840 80000
rect 78400 79200 78512 80000
rect 79072 79200 79184 80000
rect 2156 77364 2212 77374
rect 1932 76244 1988 76254
rect 1932 76150 1988 76188
rect 1932 75794 1988 75806
rect 1932 75742 1934 75794
rect 1986 75742 1988 75794
rect 1932 75348 1988 75742
rect 1932 75282 1988 75292
rect 2156 74786 2212 77308
rect 4620 76692 4676 76702
rect 4172 76690 4676 76692
rect 4172 76638 4622 76690
rect 4674 76638 4676 76690
rect 4172 76636 4676 76638
rect 4172 74898 4228 76636
rect 4620 76626 4676 76636
rect 4956 76580 5012 76590
rect 5516 76580 5572 76590
rect 4956 76578 5572 76580
rect 4956 76526 4958 76578
rect 5010 76526 5518 76578
rect 5570 76526 5572 76578
rect 4956 76524 5572 76526
rect 4284 76466 4340 76478
rect 4284 76414 4286 76466
rect 4338 76414 4340 76466
rect 4284 75908 4340 76414
rect 4476 76076 4740 76086
rect 4532 76020 4580 76076
rect 4636 76020 4684 76076
rect 4476 76010 4740 76020
rect 4284 75852 4676 75908
rect 4284 75684 4340 75694
rect 4284 75682 4564 75684
rect 4284 75630 4286 75682
rect 4338 75630 4564 75682
rect 4284 75628 4564 75630
rect 4284 75618 4340 75628
rect 4508 75124 4564 75628
rect 4620 75570 4676 75852
rect 4956 75682 5012 76524
rect 5516 76514 5572 76524
rect 4956 75630 4958 75682
rect 5010 75630 5012 75682
rect 4956 75618 5012 75630
rect 5740 76466 5796 76478
rect 5740 76414 5742 76466
rect 5794 76414 5796 76466
rect 4620 75518 4622 75570
rect 4674 75518 4676 75570
rect 4620 75506 4676 75518
rect 4620 75124 4676 75134
rect 4508 75122 4676 75124
rect 4508 75070 4622 75122
rect 4674 75070 4676 75122
rect 4508 75068 4676 75070
rect 4620 75058 4676 75068
rect 4172 74846 4174 74898
rect 4226 74846 4228 74898
rect 4172 74834 4228 74846
rect 4844 74898 4900 74910
rect 4844 74846 4846 74898
rect 4898 74846 4900 74898
rect 2156 74734 2158 74786
rect 2210 74734 2212 74786
rect 2156 74722 2212 74734
rect 4476 74508 4740 74518
rect 4532 74452 4580 74508
rect 4636 74452 4684 74508
rect 4476 74442 4740 74452
rect 1932 74228 1988 74238
rect 1932 74134 1988 74172
rect 4284 74116 4340 74126
rect 4284 74114 4676 74116
rect 4284 74062 4286 74114
rect 4338 74062 4676 74114
rect 4284 74060 4676 74062
rect 4284 74050 4340 74060
rect 4620 74002 4676 74060
rect 4620 73950 4622 74002
rect 4674 73950 4676 74002
rect 4620 73938 4676 73950
rect 4844 74114 4900 74846
rect 4844 74062 4846 74114
rect 4898 74062 4900 74114
rect 4620 73444 4676 73454
rect 4284 73442 4676 73444
rect 4284 73390 4622 73442
rect 4674 73390 4676 73442
rect 4284 73388 4676 73390
rect 4284 73330 4340 73388
rect 4620 73378 4676 73388
rect 4284 73278 4286 73330
rect 4338 73278 4340 73330
rect 4284 73266 4340 73278
rect 4844 73330 4900 74062
rect 4844 73278 4846 73330
rect 4898 73278 4900 73330
rect 1932 73108 1988 73118
rect 1932 73014 1988 73052
rect 4476 72940 4740 72950
rect 4532 72884 4580 72940
rect 4636 72884 4684 72940
rect 4476 72874 4740 72884
rect 1932 72658 1988 72670
rect 1932 72606 1934 72658
rect 1986 72606 1988 72658
rect 1932 71988 1988 72606
rect 3836 72548 3892 72558
rect 3500 72546 3892 72548
rect 3500 72494 3838 72546
rect 3890 72494 3892 72546
rect 3500 72492 3892 72494
rect 1932 71922 1988 71932
rect 3164 71988 3220 71998
rect 3164 71894 3220 71932
rect 3500 71986 3556 72492
rect 3836 72482 3892 72492
rect 4844 72212 4900 73278
rect 3500 71934 3502 71986
rect 3554 71934 3556 71986
rect 3500 71922 3556 71934
rect 3836 72156 4900 72212
rect 2492 71876 2548 71886
rect 2492 71782 2548 71820
rect 2940 71876 2996 71886
rect 2156 71762 2212 71774
rect 2156 71710 2158 71762
rect 2210 71710 2212 71762
rect 1932 71652 1988 71662
rect 2156 71652 2212 71710
rect 1820 71650 2212 71652
rect 1820 71598 1934 71650
rect 1986 71598 2212 71650
rect 1820 71596 2212 71598
rect 2940 71762 2996 71820
rect 3836 71874 3892 72156
rect 3836 71822 3838 71874
rect 3890 71822 3892 71874
rect 3836 71810 3892 71822
rect 3948 71988 4004 71998
rect 2940 71710 2942 71762
rect 2994 71710 2996 71762
rect 1820 43708 1876 71596
rect 1932 71586 1988 71596
rect 1932 71090 1988 71102
rect 1932 71038 1934 71090
rect 1986 71038 1988 71090
rect 1932 70644 1988 71038
rect 1932 70578 1988 70588
rect 2716 70196 2772 70206
rect 1932 69970 1988 69982
rect 1932 69918 1934 69970
rect 1986 69918 1988 69970
rect 1932 69524 1988 69918
rect 1932 69458 1988 69468
rect 2380 69298 2436 69310
rect 2380 69246 2382 69298
rect 2434 69246 2436 69298
rect 2044 69186 2100 69198
rect 2044 69134 2046 69186
rect 2098 69134 2100 69186
rect 2044 68626 2100 69134
rect 2044 68574 2046 68626
rect 2098 68574 2100 68626
rect 2044 68562 2100 68574
rect 1932 67954 1988 67966
rect 1932 67902 1934 67954
rect 1986 67902 1988 67954
rect 1932 67284 1988 67902
rect 1932 67218 1988 67228
rect 2044 67170 2100 67182
rect 2044 67118 2046 67170
rect 2098 67118 2100 67170
rect 2044 66274 2100 67118
rect 2380 67172 2436 69246
rect 2716 69298 2772 70140
rect 2940 69410 2996 71710
rect 3948 70978 4004 71932
rect 4172 71986 4228 72156
rect 4172 71934 4174 71986
rect 4226 71934 4228 71986
rect 4172 71922 4228 71934
rect 4508 71876 4564 71886
rect 4508 71782 4564 71820
rect 5740 71876 5796 76414
rect 11228 74226 11284 79200
rect 11564 76242 11620 76254
rect 11564 76190 11566 76242
rect 11618 76190 11620 76242
rect 11564 75572 11620 76190
rect 11900 76244 11956 79200
rect 12460 76466 12516 76478
rect 12460 76414 12462 76466
rect 12514 76414 12516 76466
rect 12460 76356 12516 76414
rect 12460 76290 12516 76300
rect 11900 76188 12068 76244
rect 11900 75908 11956 75918
rect 11900 75814 11956 75852
rect 11564 75506 11620 75516
rect 11228 74174 11230 74226
rect 11282 74174 11284 74226
rect 11228 74162 11284 74174
rect 11676 74900 11732 74910
rect 5740 71810 5796 71820
rect 4476 71372 4740 71382
rect 4532 71316 4580 71372
rect 4636 71316 4684 71372
rect 4476 71306 4740 71316
rect 3948 70926 3950 70978
rect 4002 70926 4004 70978
rect 3948 70914 4004 70926
rect 3836 70196 3892 70206
rect 3836 70102 3892 70140
rect 4476 69804 4740 69814
rect 4532 69748 4580 69804
rect 4636 69748 4684 69804
rect 4476 69738 4740 69748
rect 2940 69358 2942 69410
rect 2994 69358 2996 69410
rect 2940 69346 2996 69358
rect 2716 69246 2718 69298
rect 2770 69246 2772 69298
rect 2716 69234 2772 69246
rect 2716 68404 2772 68414
rect 2716 68310 2772 68348
rect 4476 68236 4740 68246
rect 4532 68180 4580 68236
rect 4636 68180 4684 68236
rect 4476 68170 4740 68180
rect 3836 67844 3892 67854
rect 3388 67842 3892 67844
rect 3388 67790 3838 67842
rect 3890 67790 3892 67842
rect 3388 67788 3892 67790
rect 3388 67282 3444 67788
rect 3836 67778 3892 67788
rect 3388 67230 3390 67282
rect 3442 67230 3444 67282
rect 3388 67218 3444 67230
rect 2380 67078 2436 67116
rect 3052 67172 3108 67182
rect 2716 67060 2772 67070
rect 2044 66222 2046 66274
rect 2098 66222 2100 66274
rect 2044 66210 2100 66222
rect 2492 67058 2772 67060
rect 2492 67006 2718 67058
rect 2770 67006 2772 67058
rect 2492 67004 2772 67006
rect 3052 67060 3108 67116
rect 3612 67060 3668 67070
rect 3052 67058 3668 67060
rect 3052 67006 3614 67058
rect 3666 67006 3668 67058
rect 3052 67004 3668 67006
rect 1932 65268 1988 65278
rect 1932 65174 1988 65212
rect 1932 64818 1988 64830
rect 1932 64766 1934 64818
rect 1986 64766 1988 64818
rect 1932 63924 1988 64766
rect 2492 64260 2548 67004
rect 2716 66994 2772 67004
rect 3612 66994 3668 67004
rect 4476 66668 4740 66678
rect 4532 66612 4580 66668
rect 4636 66612 4684 66668
rect 4476 66602 4740 66612
rect 2716 66052 2772 66062
rect 2716 65958 2772 65996
rect 4284 65490 4340 65502
rect 4284 65438 4286 65490
rect 4338 65438 4340 65490
rect 4284 64932 4340 65438
rect 4476 65100 4740 65110
rect 4532 65044 4580 65100
rect 4636 65044 4684 65100
rect 4476 65034 4740 65044
rect 4284 64876 4676 64932
rect 3836 64706 3892 64718
rect 3836 64654 3838 64706
rect 3890 64654 3892 64706
rect 1932 63858 1988 63868
rect 2268 64204 2548 64260
rect 3612 64596 3668 64606
rect 2268 63922 2324 64204
rect 2268 63870 2270 63922
rect 2322 63870 2324 63922
rect 1932 63250 1988 63262
rect 1932 63198 1934 63250
rect 1986 63198 1988 63250
rect 1932 62804 1988 63198
rect 1932 62738 1988 62748
rect 1932 62130 1988 62142
rect 1932 62078 1934 62130
rect 1986 62078 1988 62130
rect 1932 61684 1988 62078
rect 1932 61618 1988 61628
rect 2268 61572 2324 63870
rect 2492 64034 2548 64046
rect 2492 63982 2494 64034
rect 2546 63982 2548 64034
rect 2492 63924 2548 63982
rect 3164 64034 3220 64046
rect 3164 63982 3166 64034
rect 3218 63982 3220 64034
rect 2492 63858 2548 63868
rect 2940 63924 2996 63934
rect 2940 61572 2996 63868
rect 3164 63140 3220 63982
rect 3612 63924 3668 64540
rect 3836 64146 3892 64654
rect 4620 64594 4676 64876
rect 4620 64542 4622 64594
rect 4674 64542 4676 64594
rect 4620 64530 4676 64542
rect 4956 64596 5012 64606
rect 4956 64502 5012 64540
rect 3836 64094 3838 64146
rect 3890 64094 3892 64146
rect 3836 64082 3892 64094
rect 3612 63830 3668 63868
rect 4476 63532 4740 63542
rect 4532 63476 4580 63532
rect 4636 63476 4684 63532
rect 4476 63466 4740 63476
rect 3836 63140 3892 63150
rect 3164 63138 3892 63140
rect 3164 63086 3838 63138
rect 3890 63086 3892 63138
rect 3164 63084 3892 63086
rect 3836 63074 3892 63084
rect 3836 62356 3892 62366
rect 2268 61570 2772 61572
rect 2268 61518 2270 61570
rect 2322 61518 2772 61570
rect 2268 61516 2772 61518
rect 2268 61506 2324 61516
rect 2716 61458 2772 61516
rect 2940 61506 2996 61516
rect 3388 62354 3892 62356
rect 3388 62302 3838 62354
rect 3890 62302 3892 62354
rect 3388 62300 3892 62302
rect 2716 61406 2718 61458
rect 2770 61406 2772 61458
rect 2716 61394 2772 61406
rect 3052 61458 3108 61470
rect 3052 61406 3054 61458
rect 3106 61406 3108 61458
rect 2044 61346 2100 61358
rect 2044 61294 2046 61346
rect 2098 61294 2100 61346
rect 2044 60786 2100 61294
rect 3052 61348 3108 61406
rect 3388 61458 3444 62300
rect 3836 62290 3892 62300
rect 4476 61964 4740 61974
rect 4532 61908 4580 61964
rect 4636 61908 4684 61964
rect 4476 61898 4740 61908
rect 3612 61572 3668 61582
rect 3612 61478 3668 61516
rect 3388 61406 3390 61458
rect 3442 61406 3444 61458
rect 3388 61394 3444 61406
rect 3052 61282 3108 61292
rect 4172 61348 4228 61358
rect 4284 61348 4340 61358
rect 4228 61346 4340 61348
rect 4228 61294 4286 61346
rect 4338 61294 4340 61346
rect 4228 61292 4340 61294
rect 2044 60734 2046 60786
rect 2098 60734 2100 60786
rect 2044 60722 2100 60734
rect 2716 60564 2772 60574
rect 2716 60470 2772 60508
rect 1932 60114 1988 60126
rect 1932 60062 1934 60114
rect 1986 60062 1988 60114
rect 1932 59444 1988 60062
rect 1932 59378 1988 59388
rect 2716 60004 2772 60014
rect 2716 59442 2772 59948
rect 3836 60004 3892 60014
rect 3836 59910 3892 59948
rect 2716 59390 2718 59442
rect 2770 59390 2772 59442
rect 2716 59378 2772 59390
rect 2044 59330 2100 59342
rect 2044 59278 2046 59330
rect 2098 59278 2100 59330
rect 2044 58434 2100 59278
rect 2044 58382 2046 58434
rect 2098 58382 2100 58434
rect 2044 58370 2100 58382
rect 2156 59220 2212 59230
rect 1932 57428 1988 57438
rect 1932 57334 1988 57372
rect 1932 56978 1988 56990
rect 1932 56926 1934 56978
rect 1986 56926 1988 56978
rect 1932 56084 1988 56926
rect 1932 56018 1988 56028
rect 2044 56194 2100 56206
rect 2044 56142 2046 56194
rect 2098 56142 2100 56194
rect 2044 55298 2100 56142
rect 2044 55246 2046 55298
rect 2098 55246 2100 55298
rect 2044 55234 2100 55246
rect 1932 54290 1988 54302
rect 1932 54238 1934 54290
rect 1986 54238 1988 54290
rect 1932 53844 1988 54238
rect 1932 53778 1988 53788
rect 2156 53618 2212 59164
rect 2380 59218 2436 59230
rect 2380 59166 2382 59218
rect 2434 59166 2436 59218
rect 2380 56308 2436 59166
rect 2940 59220 2996 59230
rect 2940 59126 2996 59164
rect 3500 59220 3556 59230
rect 3500 59126 3556 59164
rect 2716 58212 2772 58222
rect 2716 58118 2772 58156
rect 3836 56868 3892 56878
rect 3724 56866 3892 56868
rect 3724 56814 3838 56866
rect 3890 56814 3892 56866
rect 3724 56812 3892 56814
rect 2716 56308 2772 56318
rect 2380 56306 2772 56308
rect 2380 56254 2718 56306
rect 2770 56254 2772 56306
rect 2380 56252 2772 56254
rect 2380 56194 2436 56252
rect 2380 56142 2382 56194
rect 2434 56142 2436 56194
rect 2380 56130 2436 56142
rect 2716 56196 2772 56252
rect 3724 56306 3780 56812
rect 3836 56802 3892 56812
rect 3724 56254 3726 56306
rect 3778 56254 3780 56306
rect 3724 56242 3780 56254
rect 2716 56130 2772 56140
rect 3388 56196 3444 56206
rect 3388 56102 3444 56140
rect 2940 56082 2996 56094
rect 2940 56030 2942 56082
rect 2994 56030 2996 56082
rect 2716 55076 2772 55086
rect 2716 54982 2772 55020
rect 2156 53566 2158 53618
rect 2210 53566 2212 53618
rect 1932 53508 1988 53518
rect 2156 53508 2212 53566
rect 2940 53730 2996 56030
rect 4172 55468 4228 61292
rect 4284 61282 4340 61292
rect 4476 60396 4740 60406
rect 4532 60340 4580 60396
rect 4636 60340 4684 60396
rect 4476 60330 4740 60340
rect 4476 58828 4740 58838
rect 4532 58772 4580 58828
rect 4636 58772 4684 58828
rect 4476 58762 4740 58772
rect 4284 57650 4340 57662
rect 4284 57598 4286 57650
rect 4338 57598 4340 57650
rect 4284 56756 4340 57598
rect 4476 57260 4740 57270
rect 4532 57204 4580 57260
rect 4636 57204 4684 57260
rect 4476 57194 4740 57204
rect 4844 56866 4900 56878
rect 4844 56814 4846 56866
rect 4898 56814 4900 56866
rect 4620 56756 4676 56766
rect 4284 56754 4676 56756
rect 4284 56702 4622 56754
rect 4674 56702 4676 56754
rect 4284 56700 4676 56702
rect 4620 56690 4676 56700
rect 4844 56196 4900 56814
rect 4844 56130 4900 56140
rect 4476 55692 4740 55702
rect 4532 55636 4580 55692
rect 4636 55636 4684 55692
rect 4476 55626 4740 55636
rect 4060 55412 4228 55468
rect 3836 54516 3892 54526
rect 2940 53678 2942 53730
rect 2994 53678 2996 53730
rect 1932 53506 2212 53508
rect 1932 53454 1934 53506
rect 1986 53454 2212 53506
rect 1932 53452 2212 53454
rect 1932 53442 1988 53452
rect 1932 52724 1988 52734
rect 1932 52630 1988 52668
rect 1932 52274 1988 52286
rect 1932 52222 1934 52274
rect 1986 52222 1988 52274
rect 1932 51604 1988 52222
rect 1932 51538 1988 51548
rect 1932 50708 1988 50718
rect 1932 50614 1988 50652
rect 1932 49588 1988 49598
rect 1932 49494 1988 49532
rect 1932 49138 1988 49150
rect 1932 49086 1934 49138
rect 1986 49086 1988 49138
rect 1932 48244 1988 49086
rect 1932 48178 1988 48188
rect 2044 48354 2100 48366
rect 2044 48302 2046 48354
rect 2098 48302 2100 48354
rect 2044 47458 2100 48302
rect 2044 47406 2046 47458
rect 2098 47406 2100 47458
rect 2044 47394 2100 47406
rect 1932 46450 1988 46462
rect 1932 46398 1934 46450
rect 1986 46398 1988 46450
rect 1932 46004 1988 46398
rect 1932 45938 1988 45948
rect 2044 45666 2100 45678
rect 2044 45614 2046 45666
rect 2098 45614 2100 45666
rect 2044 45106 2100 45614
rect 2044 45054 2046 45106
rect 2098 45054 2100 45106
rect 2044 45042 2100 45054
rect 1708 43652 1876 43708
rect 2044 44322 2100 44334
rect 2044 44270 2046 44322
rect 2098 44270 2100 44322
rect 2044 43762 2100 44270
rect 2044 43710 2046 43762
rect 2098 43710 2100 43762
rect 2044 43698 2100 43710
rect 2156 43708 2212 53452
rect 2492 53508 2548 53518
rect 2492 53414 2548 53452
rect 2940 53508 2996 53678
rect 3500 54514 3892 54516
rect 3500 54462 3838 54514
rect 3890 54462 3892 54514
rect 3500 54460 3892 54462
rect 3164 53620 3220 53630
rect 3164 53526 3220 53564
rect 3500 53618 3556 54460
rect 3836 54450 3892 54460
rect 3500 53566 3502 53618
rect 3554 53566 3556 53618
rect 3500 53554 3556 53566
rect 3836 53618 3892 53630
rect 3836 53566 3838 53618
rect 3890 53566 3892 53618
rect 2940 53442 2996 53452
rect 3836 53508 3892 53566
rect 3836 52724 3892 53452
rect 3948 53620 4004 53630
rect 3948 52946 4004 53564
rect 3948 52894 3950 52946
rect 4002 52894 4004 52946
rect 3948 52882 4004 52894
rect 3836 52668 4004 52724
rect 3836 52164 3892 52174
rect 3500 52162 3892 52164
rect 3500 52110 3838 52162
rect 3890 52110 3892 52162
rect 3500 52108 3892 52110
rect 2492 51660 2996 51716
rect 2492 51602 2548 51660
rect 2492 51550 2494 51602
rect 2546 51550 2548 51602
rect 2492 51538 2548 51550
rect 2828 51490 2884 51502
rect 2828 51438 2830 51490
rect 2882 51438 2884 51490
rect 2268 51378 2324 51390
rect 2268 51326 2270 51378
rect 2322 51326 2324 51378
rect 2268 45108 2324 51326
rect 2828 50596 2884 51438
rect 2940 51380 2996 51660
rect 3500 51602 3556 52108
rect 3836 52098 3892 52108
rect 3500 51550 3502 51602
rect 3554 51550 3556 51602
rect 3500 51538 3556 51550
rect 3836 51492 3892 51502
rect 3948 51492 4004 52668
rect 3836 51490 4004 51492
rect 3836 51438 3838 51490
rect 3890 51438 4004 51490
rect 3836 51436 4004 51438
rect 3836 51426 3892 51436
rect 3164 51380 3220 51390
rect 2940 51378 3220 51380
rect 2940 51326 3166 51378
rect 3218 51326 3220 51378
rect 2940 51324 3220 51326
rect 2828 50530 2884 50540
rect 3164 49588 3220 51324
rect 3836 50596 3892 50606
rect 3836 50502 3892 50540
rect 3836 49812 3892 49822
rect 3164 49522 3220 49532
rect 3388 49810 3892 49812
rect 3388 49758 3838 49810
rect 3890 49758 3892 49810
rect 3388 49756 3892 49758
rect 2716 49028 2772 49038
rect 2716 48466 2772 48972
rect 2716 48414 2718 48466
rect 2770 48414 2772 48466
rect 2716 48402 2772 48414
rect 3388 48466 3444 49756
rect 3836 49746 3892 49756
rect 3388 48414 3390 48466
rect 3442 48414 3444 48466
rect 3388 48402 3444 48414
rect 3612 49588 3668 49598
rect 2380 48244 2436 48254
rect 2940 48244 2996 48254
rect 2380 48242 2996 48244
rect 2380 48190 2382 48242
rect 2434 48190 2942 48242
rect 2994 48190 2996 48242
rect 2380 48188 2996 48190
rect 2380 45892 2436 48188
rect 2940 48178 2996 48188
rect 3612 48242 3668 49532
rect 3836 49028 3892 49038
rect 3836 48934 3892 48972
rect 3612 48190 3614 48242
rect 3666 48190 3668 48242
rect 3612 48178 3668 48190
rect 2716 47236 2772 47246
rect 2716 47142 2772 47180
rect 3836 46676 3892 46686
rect 3388 46674 3892 46676
rect 3388 46622 3838 46674
rect 3890 46622 3892 46674
rect 3388 46620 3892 46622
rect 2380 45798 2436 45836
rect 2828 45890 2884 45902
rect 2828 45838 2830 45890
rect 2882 45838 2884 45890
rect 2828 45780 2884 45838
rect 2828 45714 2884 45724
rect 3052 45892 3108 45902
rect 3052 45778 3108 45836
rect 3052 45726 3054 45778
rect 3106 45726 3108 45778
rect 3052 45714 3108 45726
rect 3276 45780 3332 45790
rect 2268 45052 2996 45108
rect 2716 44884 2772 44894
rect 2716 44790 2772 44828
rect 2716 44100 2772 44110
rect 2716 44006 2772 44044
rect 2156 43652 2660 43708
rect 1708 41972 1764 43652
rect 2268 43540 2324 43550
rect 2044 43484 2268 43540
rect 1932 42868 1988 42878
rect 1932 42774 1988 42812
rect 1708 40402 1764 41916
rect 1932 41748 1988 41758
rect 1932 41654 1988 41692
rect 1708 40350 1710 40402
rect 1762 40350 1764 40402
rect 1708 40338 1764 40350
rect 1932 41298 1988 41310
rect 1932 41246 1934 41298
rect 1986 41246 1988 41298
rect 1932 40404 1988 41246
rect 1932 40338 1988 40348
rect 1932 39730 1988 39742
rect 1932 39678 1934 39730
rect 1986 39678 1988 39730
rect 1932 39284 1988 39678
rect 1932 39218 1988 39228
rect 2044 38834 2100 43484
rect 2268 43446 2324 43484
rect 2268 40628 2324 40638
rect 2268 40534 2324 40572
rect 2604 40402 2660 43652
rect 2716 43650 2772 43662
rect 2716 43598 2718 43650
rect 2770 43598 2772 43650
rect 2716 42756 2772 43598
rect 2828 43540 2884 43550
rect 2940 43540 2996 45052
rect 2884 43538 2996 43540
rect 2884 43486 2942 43538
rect 2994 43486 2996 43538
rect 2884 43484 2996 43486
rect 2828 43474 2884 43484
rect 2940 43446 2996 43484
rect 2716 42690 2772 42700
rect 2604 40350 2606 40402
rect 2658 40350 2660 40402
rect 2604 39620 2660 40350
rect 3164 40404 3220 40414
rect 3164 40310 3220 40348
rect 2604 39554 2660 39564
rect 2044 38782 2046 38834
rect 2098 38782 2100 38834
rect 2044 38162 2100 38782
rect 2940 38724 2996 38734
rect 2940 38164 2996 38668
rect 3276 38724 3332 45724
rect 3388 45778 3444 46620
rect 3836 46610 3892 46620
rect 3612 45892 3668 45902
rect 3612 45798 3668 45836
rect 3388 45726 3390 45778
rect 3442 45726 3444 45778
rect 3388 45714 3444 45726
rect 3836 42756 3892 42766
rect 3836 42662 3892 42700
rect 3836 41972 3892 41982
rect 3836 41878 3892 41916
rect 4060 41300 4116 55412
rect 4476 54124 4740 54134
rect 4532 54068 4580 54124
rect 4636 54068 4684 54124
rect 4476 54058 4740 54068
rect 4476 52556 4740 52566
rect 4532 52500 4580 52556
rect 4636 52500 4684 52556
rect 4476 52490 4740 52500
rect 4476 50988 4740 50998
rect 4532 50932 4580 50988
rect 4636 50932 4684 50988
rect 4476 50922 4740 50932
rect 4476 49420 4740 49430
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4476 49354 4740 49364
rect 4476 47852 4740 47862
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4476 47786 4740 47796
rect 4476 46284 4740 46294
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4476 46218 4740 46228
rect 4284 45780 4340 45790
rect 4284 45686 4340 45724
rect 4476 44716 4740 44726
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4476 44650 4740 44660
rect 4476 43148 4740 43158
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4476 43082 4740 43092
rect 4732 41972 4788 41982
rect 4732 41878 4788 41916
rect 4476 41580 4740 41590
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4476 41514 4740 41524
rect 4732 41300 4788 41310
rect 4060 41298 4788 41300
rect 4060 41246 4734 41298
rect 4786 41246 4788 41298
rect 4060 41244 4788 41246
rect 4060 41188 4116 41244
rect 4732 41234 4788 41244
rect 3500 41186 4116 41188
rect 3500 41134 4062 41186
rect 4114 41134 4116 41186
rect 3500 41132 4116 41134
rect 3500 40402 3556 41132
rect 4060 41122 4116 41132
rect 5404 40628 5460 40638
rect 4060 40516 4116 40526
rect 4060 40422 4116 40460
rect 4508 40516 4564 40526
rect 4508 40422 4564 40460
rect 5180 40516 5236 40526
rect 3500 40350 3502 40402
rect 3554 40350 3556 40402
rect 3500 40338 3556 40350
rect 4956 40404 5012 40414
rect 4956 40310 5012 40348
rect 4476 40012 4740 40022
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4476 39946 4740 39956
rect 3836 39620 3892 39630
rect 3836 39526 3892 39564
rect 4732 39620 4788 39630
rect 4732 39526 4788 39564
rect 5180 39396 5236 40460
rect 5180 39330 5236 39340
rect 5404 40402 5460 40572
rect 5404 40350 5406 40402
rect 5458 40350 5460 40402
rect 3276 38658 3332 38668
rect 3388 38722 3444 38734
rect 3388 38670 3390 38722
rect 3442 38670 3444 38722
rect 2044 38110 2046 38162
rect 2098 38110 2100 38162
rect 2044 38098 2100 38110
rect 2492 38162 2996 38164
rect 2492 38110 2942 38162
rect 2994 38110 2996 38162
rect 2492 38108 2996 38110
rect 2492 38050 2548 38108
rect 2940 38098 2996 38108
rect 3388 38164 3444 38670
rect 4476 38444 4740 38454
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4476 38378 4740 38388
rect 3388 38098 3444 38108
rect 2492 37998 2494 38050
rect 2546 37998 2548 38050
rect 2492 37986 2548 37998
rect 2044 37380 2100 37390
rect 2044 37286 2100 37324
rect 1708 37266 1764 37278
rect 1708 37214 1710 37266
rect 1762 37214 1764 37266
rect 1708 37044 1764 37214
rect 1708 36978 1764 36988
rect 2492 37154 2548 37166
rect 2492 37102 2494 37154
rect 2546 37102 2548 37154
rect 2492 37044 2548 37102
rect 2492 36978 2548 36988
rect 4476 36876 4740 36886
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4476 36810 4740 36820
rect 1708 36370 1764 36382
rect 1708 36318 1710 36370
rect 1762 36318 1764 36370
rect 1708 35924 1764 36318
rect 2044 36260 2100 36270
rect 2044 36166 2100 36204
rect 2492 36258 2548 36270
rect 2492 36206 2494 36258
rect 2546 36206 2548 36258
rect 1708 35858 1764 35868
rect 2492 35924 2548 36206
rect 2492 35858 2548 35868
rect 4476 35308 4740 35318
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4476 35242 4740 35252
rect 1708 34804 1764 34814
rect 1708 34710 1764 34748
rect 2492 34804 2548 34814
rect 2492 34710 2548 34748
rect 2044 34692 2100 34702
rect 2044 34598 2100 34636
rect 2044 34242 2100 34254
rect 2044 34190 2046 34242
rect 2098 34190 2100 34242
rect 1708 34130 1764 34142
rect 1708 34078 1710 34130
rect 1762 34078 1764 34130
rect 1708 33684 1764 34078
rect 1708 33618 1764 33628
rect 2044 33348 2100 34190
rect 2492 34018 2548 34030
rect 2492 33966 2494 34018
rect 2546 33966 2548 34018
rect 2492 33684 2548 33966
rect 4476 33740 4740 33750
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4476 33674 4740 33684
rect 2492 33618 2548 33628
rect 2044 33282 2100 33292
rect 1708 33122 1764 33134
rect 1708 33070 1710 33122
rect 1762 33070 1764 33122
rect 1708 32564 1764 33070
rect 2044 33124 2100 33134
rect 2044 33030 2100 33068
rect 2492 33122 2548 33134
rect 2492 33070 2494 33122
rect 2546 33070 2548 33122
rect 1708 32498 1764 32508
rect 2492 32564 2548 33070
rect 2492 32498 2548 32508
rect 4476 32172 4740 32182
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4476 32106 4740 32116
rect 1708 31666 1764 31678
rect 1708 31614 1710 31666
rect 1762 31614 1764 31666
rect 1708 31444 1764 31614
rect 2044 31556 2100 31566
rect 2044 31462 2100 31500
rect 2492 31554 2548 31566
rect 2492 31502 2494 31554
rect 2546 31502 2548 31554
rect 1708 31378 1764 31388
rect 2492 31444 2548 31502
rect 2492 31378 2548 31388
rect 2044 31108 2100 31118
rect 2044 31014 2100 31052
rect 1708 30994 1764 31006
rect 1708 30942 1710 30994
rect 1762 30942 1764 30994
rect 1708 30884 1764 30942
rect 1708 30324 1764 30828
rect 2492 30884 2548 30894
rect 2492 30790 2548 30828
rect 4476 30604 4740 30614
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4476 30538 4740 30548
rect 1708 30258 1764 30268
rect 2044 29540 2100 29550
rect 2044 29446 2100 29484
rect 1708 29426 1764 29438
rect 1708 29374 1710 29426
rect 1762 29374 1764 29426
rect 1708 29204 1764 29374
rect 1708 29138 1764 29148
rect 2492 29314 2548 29326
rect 2492 29262 2494 29314
rect 2546 29262 2548 29314
rect 2492 29204 2548 29262
rect 2492 29138 2548 29148
rect 4476 29036 4740 29046
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4476 28970 4740 28980
rect 1708 28642 1764 28654
rect 1708 28590 1710 28642
rect 1762 28590 1764 28642
rect 1708 28084 1764 28590
rect 2044 28644 2100 28654
rect 2044 28530 2100 28588
rect 2044 28478 2046 28530
rect 2098 28478 2100 28530
rect 2044 28466 2100 28478
rect 2492 28642 2548 28654
rect 2492 28590 2494 28642
rect 2546 28590 2548 28642
rect 1708 28018 1764 28028
rect 2492 28084 2548 28590
rect 2492 28018 2548 28028
rect 5404 27748 5460 40350
rect 5404 27682 5460 27692
rect 2044 27636 2100 27646
rect 1708 26964 1764 26974
rect 1708 26870 1764 26908
rect 2044 26962 2100 27580
rect 4476 27468 4740 27478
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4476 27402 4740 27412
rect 2044 26910 2046 26962
rect 2098 26910 2100 26962
rect 2044 26898 2100 26910
rect 2492 26964 2548 26974
rect 2492 26870 2548 26908
rect 2156 26516 2212 26526
rect 2044 26404 2100 26414
rect 2044 26310 2100 26348
rect 1708 26290 1764 26302
rect 1708 26238 1710 26290
rect 1762 26238 1764 26290
rect 1708 25844 1764 26238
rect 1708 25778 1764 25788
rect 2044 25396 2100 25406
rect 2156 25396 2212 26460
rect 2492 26178 2548 26190
rect 2492 26126 2494 26178
rect 2546 26126 2548 26178
rect 2492 25844 2548 26126
rect 4476 25900 4740 25910
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4476 25834 4740 25844
rect 2492 25778 2548 25788
rect 2044 25394 2212 25396
rect 2044 25342 2046 25394
rect 2098 25342 2212 25394
rect 2044 25340 2212 25342
rect 2044 25330 2100 25340
rect 1708 25282 1764 25294
rect 1708 25230 1710 25282
rect 1762 25230 1764 25282
rect 1708 24724 1764 25230
rect 1708 24658 1764 24668
rect 2492 25282 2548 25294
rect 2492 25230 2494 25282
rect 2546 25230 2548 25282
rect 2492 24724 2548 25230
rect 2492 24658 2548 24668
rect 4476 24332 4740 24342
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4476 24266 4740 24276
rect 2044 24052 2100 24062
rect 1708 23826 1764 23838
rect 1708 23774 1710 23826
rect 1762 23774 1764 23826
rect 1708 23604 1764 23774
rect 2044 23826 2100 23996
rect 2044 23774 2046 23826
rect 2098 23774 2100 23826
rect 2044 23762 2100 23774
rect 1708 23538 1764 23548
rect 2492 23714 2548 23726
rect 2492 23662 2494 23714
rect 2546 23662 2548 23714
rect 2492 23604 2548 23662
rect 2492 23538 2548 23548
rect 11564 23604 11620 23614
rect 2156 23492 2212 23502
rect 2044 23266 2100 23278
rect 2044 23214 2046 23266
rect 2098 23214 2100 23266
rect 1708 23154 1764 23166
rect 1708 23102 1710 23154
rect 1762 23102 1764 23154
rect 1708 23044 1764 23102
rect 1708 22484 1764 22988
rect 2044 22932 2100 23214
rect 2044 22866 2100 22876
rect 2156 22596 2212 23436
rect 2492 23044 2548 23054
rect 2492 22950 2548 22988
rect 4476 22764 4740 22774
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4476 22698 4740 22708
rect 1708 22418 1764 22428
rect 2044 22540 2212 22596
rect 2044 21810 2100 22540
rect 2044 21758 2046 21810
rect 2098 21758 2100 21810
rect 2044 21746 2100 21758
rect 2156 21812 2212 21822
rect 1708 21586 1764 21598
rect 1708 21534 1710 21586
rect 1762 21534 1764 21586
rect 1708 21364 1764 21534
rect 1708 21298 1764 21308
rect 2044 20692 2100 20702
rect 2156 20692 2212 21756
rect 2492 21474 2548 21486
rect 2492 21422 2494 21474
rect 2546 21422 2548 21474
rect 2492 21364 2548 21422
rect 2492 21298 2548 21308
rect 4476 21196 4740 21206
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4476 21130 4740 21140
rect 2044 20690 2212 20692
rect 2044 20638 2046 20690
rect 2098 20638 2212 20690
rect 2044 20636 2212 20638
rect 2044 20626 2100 20636
rect 1708 20578 1764 20590
rect 1708 20526 1710 20578
rect 1762 20526 1764 20578
rect 1708 20244 1764 20526
rect 2492 20578 2548 20590
rect 2492 20526 2494 20578
rect 2546 20526 2548 20578
rect 1708 20178 1764 20188
rect 2044 20356 2100 20366
rect 1708 19124 1764 19134
rect 1708 19030 1764 19068
rect 2044 19122 2100 20300
rect 2492 20244 2548 20526
rect 2492 20178 2548 20188
rect 7532 19796 7588 19806
rect 4476 19628 4740 19638
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4476 19562 4740 19572
rect 2044 19070 2046 19122
rect 2098 19070 2100 19122
rect 2044 19058 2100 19070
rect 2492 19124 2548 19134
rect 2492 19030 2548 19068
rect 2044 18562 2100 18574
rect 2044 18510 2046 18562
rect 2098 18510 2100 18562
rect 1708 18450 1764 18462
rect 1708 18398 1710 18450
rect 1762 18398 1764 18450
rect 1708 18004 1764 18398
rect 1708 17938 1764 17948
rect 2044 17892 2100 18510
rect 2492 18338 2548 18350
rect 2492 18286 2494 18338
rect 2546 18286 2548 18338
rect 2492 18004 2548 18286
rect 4476 18060 4740 18070
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4476 17994 4740 18004
rect 2492 17938 2548 17948
rect 2044 17826 2100 17836
rect 1708 17554 1764 17566
rect 1708 17502 1710 17554
rect 1762 17502 1764 17554
rect 1708 17444 1764 17502
rect 1708 16884 1764 17388
rect 2044 17442 2100 17454
rect 2044 17390 2046 17442
rect 2098 17390 2100 17442
rect 2044 17108 2100 17390
rect 2492 17444 2548 17454
rect 2492 17350 2548 17388
rect 2044 17042 2100 17052
rect 1708 16818 1764 16828
rect 4476 16492 4740 16502
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4476 16426 4740 16436
rect 2044 16324 2100 16334
rect 1932 16100 1988 16110
rect 1708 15986 1764 15998
rect 1708 15934 1710 15986
rect 1762 15934 1764 15986
rect 1708 15764 1764 15934
rect 1708 15698 1764 15708
rect 1708 15314 1764 15326
rect 1708 15262 1710 15314
rect 1762 15262 1764 15314
rect 1708 14644 1764 15262
rect 1708 14578 1764 14588
rect 1708 13746 1764 13758
rect 1708 13694 1710 13746
rect 1762 13694 1764 13746
rect 1708 13524 1764 13694
rect 1708 13458 1764 13468
rect 1708 12850 1764 12862
rect 1708 12798 1710 12850
rect 1762 12798 1764 12850
rect 1708 12404 1764 12798
rect 1708 12338 1764 12348
rect 1708 11284 1764 11294
rect 1708 11190 1764 11228
rect 1708 10610 1764 10622
rect 1708 10558 1710 10610
rect 1762 10558 1764 10610
rect 1708 10164 1764 10558
rect 1708 10098 1764 10108
rect 1708 9714 1764 9726
rect 1708 9662 1710 9714
rect 1762 9662 1764 9714
rect 1708 9604 1764 9662
rect 1708 9044 1764 9548
rect 1708 8978 1764 8988
rect 1708 8146 1764 8158
rect 1708 8094 1710 8146
rect 1762 8094 1764 8146
rect 1708 7924 1764 8094
rect 1708 7858 1764 7868
rect 1708 7474 1764 7486
rect 1708 7422 1710 7474
rect 1762 7422 1764 7474
rect 1708 7364 1764 7422
rect 1708 6804 1764 7308
rect 1708 6738 1764 6748
rect 1932 6132 1988 16044
rect 2044 15986 2100 16268
rect 2044 15934 2046 15986
rect 2098 15934 2100 15986
rect 2044 15922 2100 15934
rect 5964 15988 6020 15998
rect 2492 15874 2548 15886
rect 2492 15822 2494 15874
rect 2546 15822 2548 15874
rect 2492 15764 2548 15822
rect 2492 15698 2548 15708
rect 2044 15428 2100 15438
rect 2044 15334 2100 15372
rect 2492 15202 2548 15214
rect 2492 15150 2494 15202
rect 2546 15150 2548 15202
rect 2156 14756 2212 14766
rect 2044 13972 2100 13982
rect 2044 13878 2100 13916
rect 2044 12852 2100 12862
rect 2156 12852 2212 14700
rect 2492 14644 2548 15150
rect 4476 14924 4740 14934
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4476 14858 4740 14868
rect 2492 14578 2548 14588
rect 2492 13634 2548 13646
rect 2492 13582 2494 13634
rect 2546 13582 2548 13634
rect 2492 13524 2548 13582
rect 2492 13458 2548 13468
rect 4476 13356 4740 13366
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4476 13290 4740 13300
rect 2044 12850 2212 12852
rect 2044 12798 2046 12850
rect 2098 12798 2212 12850
rect 2044 12796 2212 12798
rect 2044 12786 2100 12796
rect 2492 12738 2548 12750
rect 2492 12686 2494 12738
rect 2546 12686 2548 12738
rect 2492 12404 2548 12686
rect 2492 12338 2548 12348
rect 2156 12292 2212 12302
rect 2044 11172 2100 11182
rect 2044 11078 2100 11116
rect 2044 10836 2100 10846
rect 2156 10836 2212 12236
rect 4476 11788 4740 11798
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4476 11722 4740 11732
rect 2492 11284 2548 11294
rect 2492 11190 2548 11228
rect 2044 10834 2212 10836
rect 2044 10782 2046 10834
rect 2098 10782 2212 10834
rect 2044 10780 2212 10782
rect 2380 10948 2436 10958
rect 2044 10770 2100 10780
rect 2044 10052 2100 10062
rect 2044 9714 2100 9996
rect 2044 9662 2046 9714
rect 2098 9662 2100 9714
rect 2044 9650 2100 9662
rect 2380 8428 2436 10892
rect 2492 10498 2548 10510
rect 2492 10446 2494 10498
rect 2546 10446 2548 10498
rect 2492 10164 2548 10446
rect 4476 10220 4740 10230
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4476 10154 4740 10164
rect 2492 10098 2548 10108
rect 2492 9604 2548 9614
rect 2492 9510 2548 9548
rect 4476 8652 4740 8662
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4476 8586 4740 8596
rect 2044 8372 2436 8428
rect 2044 8146 2100 8372
rect 2044 8094 2046 8146
rect 2098 8094 2100 8146
rect 2044 8082 2100 8094
rect 2492 8034 2548 8046
rect 2492 7982 2494 8034
rect 2546 7982 2548 8034
rect 2492 7924 2548 7982
rect 2492 7858 2548 7868
rect 2044 7700 2100 7710
rect 2044 7606 2100 7644
rect 2492 7364 2548 7374
rect 2492 7270 2548 7308
rect 4476 7084 4740 7094
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4476 7018 4740 7028
rect 2716 6804 2772 6814
rect 2044 6132 2100 6142
rect 1932 6130 2100 6132
rect 1932 6078 2046 6130
rect 2098 6078 2100 6130
rect 1932 6076 2100 6078
rect 2044 6066 2100 6076
rect 1708 5906 1764 5918
rect 1708 5854 1710 5906
rect 1762 5854 1764 5906
rect 1708 5684 1764 5854
rect 1708 5618 1764 5628
rect 2044 5796 2100 5806
rect 1708 5122 1764 5134
rect 1708 5070 1710 5122
rect 1762 5070 1764 5122
rect 1708 4564 1764 5070
rect 2044 5010 2100 5740
rect 2492 5794 2548 5806
rect 2492 5742 2494 5794
rect 2546 5742 2548 5794
rect 2492 5684 2548 5742
rect 2492 5618 2548 5628
rect 2044 4958 2046 5010
rect 2098 4958 2100 5010
rect 2044 4946 2100 4958
rect 2492 5122 2548 5134
rect 2492 5070 2494 5122
rect 2546 5070 2548 5122
rect 1708 4498 1764 4508
rect 2044 4788 2100 4798
rect 1708 3444 1764 3454
rect 1708 3350 1764 3388
rect 2044 3442 2100 4732
rect 2492 4564 2548 5070
rect 2492 4498 2548 4508
rect 2044 3390 2046 3442
rect 2098 3390 2100 3442
rect 2044 3378 2100 3390
rect 2156 4226 2212 4238
rect 2156 4174 2158 4226
rect 2210 4174 2212 4226
rect 2156 3444 2212 4174
rect 2380 3444 2436 3454
rect 2156 3442 2436 3444
rect 2156 3390 2382 3442
rect 2434 3390 2436 3442
rect 2156 3388 2436 3390
rect 2380 2324 2436 3388
rect 2716 3442 2772 6748
rect 4284 5684 4340 5694
rect 2716 3390 2718 3442
rect 2770 3390 2772 3442
rect 2716 3378 2772 3390
rect 3164 3444 3220 3454
rect 3164 3350 3220 3388
rect 3724 3444 3780 3454
rect 3948 3444 4004 3454
rect 3724 3442 4004 3444
rect 3724 3390 3726 3442
rect 3778 3390 3950 3442
rect 4002 3390 4004 3442
rect 3724 3388 4004 3390
rect 4284 3442 4340 5628
rect 4476 5516 4740 5526
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4476 5450 4740 5460
rect 4956 5348 5012 5358
rect 4732 4228 4788 4238
rect 4732 4226 4900 4228
rect 4732 4174 4734 4226
rect 4786 4174 4900 4226
rect 4732 4172 4900 4174
rect 4732 4162 4788 4172
rect 4476 3948 4740 3958
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4476 3882 4740 3892
rect 4284 3390 4286 3442
rect 4338 3390 4340 3442
rect 3724 3378 3780 3388
rect 3948 3332 4116 3388
rect 4284 3378 4340 3390
rect 4732 3556 4788 3566
rect 4844 3556 4900 4172
rect 4732 3554 4900 3556
rect 4732 3502 4734 3554
rect 4786 3502 4900 3554
rect 4732 3500 4900 3502
rect 4732 3444 4788 3500
rect 4732 3378 4788 3388
rect 4956 3442 5012 5292
rect 5180 4900 5236 4910
rect 5180 4806 5236 4844
rect 5964 4788 6020 15932
rect 6972 14532 7028 14542
rect 6636 13076 6692 13086
rect 6636 7700 6692 13020
rect 6636 7634 6692 7644
rect 6300 6468 6356 6478
rect 6188 5796 6244 5806
rect 5964 4722 6020 4732
rect 6076 5794 6244 5796
rect 6076 5742 6190 5794
rect 6242 5742 6244 5794
rect 6076 5740 6244 5742
rect 6076 4564 6132 5740
rect 6188 5730 6244 5740
rect 6188 5122 6244 5134
rect 6188 5070 6190 5122
rect 6242 5070 6244 5122
rect 6188 4788 6244 5070
rect 6188 4722 6244 4732
rect 5964 4508 6132 4564
rect 6188 4564 6244 4574
rect 6300 4564 6356 6412
rect 6748 5908 6804 5918
rect 6636 5794 6692 5806
rect 6636 5742 6638 5794
rect 6690 5742 6692 5794
rect 6524 5124 6580 5134
rect 6636 5124 6692 5742
rect 6524 5122 6692 5124
rect 6524 5070 6526 5122
rect 6578 5070 6692 5122
rect 6524 5068 6692 5070
rect 6188 4562 6356 4564
rect 6188 4510 6190 4562
rect 6242 4510 6356 4562
rect 6188 4508 6356 4510
rect 6412 4900 6468 4910
rect 5180 4452 5236 4462
rect 5852 4452 5908 4462
rect 5180 4450 5908 4452
rect 5180 4398 5182 4450
rect 5234 4398 5854 4450
rect 5906 4398 5908 4450
rect 5180 4396 5908 4398
rect 5180 4386 5236 4396
rect 5628 4226 5684 4238
rect 5628 4174 5630 4226
rect 5682 4174 5684 4226
rect 5628 3892 5684 4174
rect 5628 3826 5684 3836
rect 5740 3668 5796 3678
rect 5740 3554 5796 3612
rect 5740 3502 5742 3554
rect 5794 3502 5796 3554
rect 5740 3490 5796 3502
rect 4956 3390 4958 3442
rect 5010 3390 5012 3442
rect 4956 3378 5012 3390
rect 2380 2258 2436 2268
rect 4060 756 4116 3332
rect 5852 2884 5908 4396
rect 5964 3668 6020 4508
rect 6188 4498 6244 4508
rect 5964 3602 6020 3612
rect 6076 4340 6132 4350
rect 6076 3442 6132 4284
rect 6412 3780 6468 4844
rect 6412 3554 6468 3724
rect 6412 3502 6414 3554
rect 6466 3502 6468 3554
rect 6412 3490 6468 3502
rect 6076 3390 6078 3442
rect 6130 3390 6132 3442
rect 6076 3378 6132 3390
rect 6300 3444 6356 3454
rect 5628 2828 5908 2884
rect 4732 924 5012 980
rect 4732 756 4788 924
rect 4956 800 5012 924
rect 5628 800 5684 2828
rect 6300 800 6356 3388
rect 6524 3388 6580 5068
rect 6748 5010 6804 5852
rect 6972 5796 7028 14476
rect 7420 6916 7476 6926
rect 7308 6860 7420 6916
rect 6972 5730 7028 5740
rect 7084 5794 7140 5806
rect 7084 5742 7086 5794
rect 7138 5742 7140 5794
rect 6748 4958 6750 5010
rect 6802 4958 6804 5010
rect 6748 4946 6804 4958
rect 6860 4900 6916 4910
rect 6748 4338 6804 4350
rect 6748 4286 6750 4338
rect 6802 4286 6804 4338
rect 6748 3892 6804 4286
rect 6748 3826 6804 3836
rect 6748 3444 6804 3454
rect 6860 3444 6916 4844
rect 7084 4676 7140 5742
rect 7196 5796 7252 5806
rect 7196 5346 7252 5740
rect 7196 5294 7198 5346
rect 7250 5294 7252 5346
rect 7196 5282 7252 5294
rect 7084 4610 7140 4620
rect 7308 4564 7364 6860
rect 7420 6850 7476 6860
rect 7532 6804 7588 19740
rect 9996 18004 10052 18014
rect 9548 12180 9604 12190
rect 8988 12178 9604 12180
rect 8988 12126 9550 12178
rect 9602 12126 9604 12178
rect 8988 12124 9604 12126
rect 7532 6738 7588 6748
rect 8316 9604 8372 9614
rect 8316 6802 8372 9548
rect 8876 8484 8932 8494
rect 8764 8428 8876 8484
rect 8316 6750 8318 6802
rect 8370 6750 8372 6802
rect 8316 6738 8372 6750
rect 8428 6804 8484 6814
rect 8428 6710 8484 6748
rect 7420 6466 7476 6478
rect 7420 6414 7422 6466
rect 7474 6414 7476 6466
rect 7420 5682 7476 6414
rect 7868 6466 7924 6478
rect 7868 6414 7870 6466
rect 7922 6414 7924 6466
rect 7532 5796 7588 5806
rect 7532 5794 7812 5796
rect 7532 5742 7534 5794
rect 7586 5742 7812 5794
rect 7532 5740 7812 5742
rect 7532 5730 7588 5740
rect 7420 5630 7422 5682
rect 7474 5630 7476 5682
rect 7420 5618 7476 5630
rect 7420 5460 7476 5470
rect 7420 5234 7476 5404
rect 7420 5182 7422 5234
rect 7474 5182 7476 5234
rect 7420 5170 7476 5182
rect 7532 4564 7588 4574
rect 7308 4562 7588 4564
rect 7308 4510 7534 4562
rect 7586 4510 7588 4562
rect 7308 4508 7588 4510
rect 7532 4498 7588 4508
rect 6972 4452 7028 4462
rect 7644 4452 7700 4462
rect 6972 4450 7364 4452
rect 6972 4398 6974 4450
rect 7026 4398 7364 4450
rect 6972 4396 7364 4398
rect 6972 4386 7028 4396
rect 7308 4338 7364 4396
rect 7644 4358 7700 4396
rect 7308 4286 7310 4338
rect 7362 4286 7364 4338
rect 7308 4274 7364 4286
rect 7420 4116 7476 4126
rect 6748 3442 6916 3444
rect 6748 3390 6750 3442
rect 6802 3390 6916 3442
rect 6748 3388 6916 3390
rect 7196 3556 7252 3566
rect 6524 3332 6692 3388
rect 6748 3378 6804 3388
rect 6636 3220 6692 3332
rect 6636 3164 7028 3220
rect 6972 800 7028 3164
rect 7196 2994 7252 3500
rect 7420 3442 7476 4060
rect 7420 3390 7422 3442
rect 7474 3390 7476 3442
rect 7420 3378 7476 3390
rect 7644 3892 7700 3902
rect 7756 3892 7812 5740
rect 7868 5572 7924 6414
rect 8204 6468 8260 6478
rect 8204 6374 8260 6412
rect 8316 6132 8372 6142
rect 7868 5506 7924 5516
rect 7980 5794 8036 5806
rect 7980 5742 7982 5794
rect 8034 5742 8036 5794
rect 7868 5346 7924 5358
rect 7868 5294 7870 5346
rect 7922 5294 7924 5346
rect 7868 5234 7924 5294
rect 7868 5182 7870 5234
rect 7922 5182 7924 5234
rect 7868 5170 7924 5182
rect 7980 4564 8036 5742
rect 7980 4498 8036 4508
rect 8092 5682 8148 5694
rect 8092 5630 8094 5682
rect 8146 5630 8148 5682
rect 7980 4340 8036 4350
rect 7980 4246 8036 4284
rect 8092 4228 8148 5630
rect 8204 5236 8260 5246
rect 8204 4562 8260 5180
rect 8316 5234 8372 6076
rect 8652 5908 8708 5946
rect 8652 5842 8708 5852
rect 8316 5182 8318 5234
rect 8370 5182 8372 5234
rect 8316 5170 8372 5182
rect 8428 5794 8484 5806
rect 8428 5742 8430 5794
rect 8482 5742 8484 5794
rect 8428 5012 8484 5742
rect 8764 5794 8820 8428
rect 8876 8418 8932 8428
rect 8988 6802 9044 12124
rect 9548 12114 9604 12124
rect 9772 12066 9828 12078
rect 9772 12014 9774 12066
rect 9826 12014 9828 12066
rect 9772 11506 9828 12014
rect 9884 12068 9940 12078
rect 9884 11974 9940 12012
rect 9772 11454 9774 11506
rect 9826 11454 9828 11506
rect 9772 11442 9828 11454
rect 9100 11396 9156 11406
rect 9100 11394 9604 11396
rect 9100 11342 9102 11394
rect 9154 11342 9604 11394
rect 9100 11340 9604 11342
rect 9100 11330 9156 11340
rect 9548 10612 9604 11340
rect 9996 10948 10052 17948
rect 9996 10882 10052 10892
rect 10108 14644 10164 14654
rect 9548 10610 9716 10612
rect 9548 10558 9550 10610
rect 9602 10558 9716 10610
rect 9548 10556 9716 10558
rect 9548 10546 9604 10556
rect 9436 10500 9492 10510
rect 9436 9938 9492 10444
rect 9436 9886 9438 9938
rect 9490 9886 9492 9938
rect 9436 9874 9492 9886
rect 9548 9716 9604 9726
rect 9548 9622 9604 9660
rect 9324 9604 9380 9614
rect 9324 9510 9380 9548
rect 9660 9042 9716 10556
rect 10108 10052 10164 14588
rect 11564 11172 11620 23548
rect 11676 21700 11732 74844
rect 12012 73444 12068 76188
rect 12572 75908 12628 79200
rect 13244 76132 13300 79200
rect 13356 76356 13412 76366
rect 13356 76262 13412 76300
rect 12572 75842 12628 75852
rect 12908 76076 13300 76132
rect 12572 75684 12628 75694
rect 12124 73444 12180 73454
rect 12012 73442 12180 73444
rect 12012 73390 12126 73442
rect 12178 73390 12180 73442
rect 12012 73388 12180 73390
rect 12124 73378 12180 73388
rect 12572 72772 12628 75628
rect 12908 75122 12964 76076
rect 13580 75684 13636 75694
rect 13580 75590 13636 75628
rect 13916 75572 13972 79200
rect 13916 75506 13972 75516
rect 14140 76356 14196 76366
rect 12908 75070 12910 75122
rect 12962 75070 12964 75122
rect 12908 75058 12964 75070
rect 13468 74900 13524 74910
rect 13468 74806 13524 74844
rect 14140 74676 14196 76300
rect 14252 75458 14308 75470
rect 14252 75406 14254 75458
rect 14306 75406 14308 75458
rect 14252 74900 14308 75406
rect 14252 74834 14308 74844
rect 14140 74620 14308 74676
rect 12460 72716 12628 72772
rect 12684 74114 12740 74126
rect 12684 74062 12686 74114
rect 12738 74062 12740 74114
rect 12684 74004 12740 74062
rect 12460 24500 12516 72716
rect 12684 55468 12740 73948
rect 14028 74002 14084 74014
rect 14028 73950 14030 74002
rect 14082 73950 14084 74002
rect 13916 73330 13972 73342
rect 13916 73278 13918 73330
rect 13970 73278 13972 73330
rect 13916 72324 13972 73278
rect 14028 73332 14084 73950
rect 14028 73266 14084 73276
rect 14140 72324 14196 72334
rect 13916 72322 14196 72324
rect 13916 72270 14142 72322
rect 14194 72270 14196 72322
rect 13916 72268 14196 72270
rect 14140 55468 14196 72268
rect 12460 23548 12516 24444
rect 11676 21634 11732 21644
rect 12348 23492 12516 23548
rect 12572 55412 12740 55468
rect 13468 55412 14196 55468
rect 12572 23548 12628 55412
rect 13468 25284 13524 55412
rect 13468 23604 13524 25228
rect 14252 24836 14308 74620
rect 14364 74004 14420 74014
rect 14364 73910 14420 73948
rect 14588 73218 14644 79200
rect 14700 75684 14756 75694
rect 14700 75590 14756 75628
rect 15260 75010 15316 79200
rect 15372 76692 15428 76702
rect 15372 76598 15428 76636
rect 15260 74958 15262 75010
rect 15314 74958 15316 75010
rect 15260 74946 15316 74958
rect 15932 74338 15988 79200
rect 16604 76692 16660 79200
rect 16604 76626 16660 76636
rect 16380 76466 16436 76478
rect 16380 76414 16382 76466
rect 16434 76414 16436 76466
rect 16380 76356 16436 76414
rect 16380 76290 16436 76300
rect 17164 76356 17220 76366
rect 17164 76262 17220 76300
rect 16828 75908 16884 75918
rect 17276 75908 17332 79200
rect 16828 75906 17332 75908
rect 16828 75854 16830 75906
rect 16882 75854 17332 75906
rect 16828 75852 17332 75854
rect 16828 75842 16884 75852
rect 15932 74286 15934 74338
rect 15986 74286 15988 74338
rect 15932 74274 15988 74286
rect 16492 75684 16548 75694
rect 16492 74898 16548 75628
rect 17836 75682 17892 75694
rect 17836 75630 17838 75682
rect 17890 75630 17892 75682
rect 17836 75012 17892 75630
rect 17948 75572 18004 79200
rect 18060 76468 18116 76478
rect 18060 76374 18116 76412
rect 18620 75794 18676 79200
rect 19292 76578 19348 79200
rect 19964 77028 20020 79200
rect 19964 76972 20244 77028
rect 19836 76860 20100 76870
rect 19892 76804 19940 76860
rect 19996 76804 20044 76860
rect 19836 76794 20100 76804
rect 20188 76692 20244 76972
rect 19292 76526 19294 76578
rect 19346 76526 19348 76578
rect 19292 76514 19348 76526
rect 20076 76636 20244 76692
rect 18620 75742 18622 75794
rect 18674 75742 18676 75794
rect 18620 75730 18676 75742
rect 19404 76468 19460 76478
rect 17948 75506 18004 75516
rect 19180 75572 19236 75582
rect 17836 74956 18116 75012
rect 16492 74846 16494 74898
rect 16546 74846 16548 74898
rect 14588 73166 14590 73218
rect 14642 73166 14644 73218
rect 14588 73154 14644 73166
rect 16268 73332 16324 73342
rect 16380 73332 16436 73342
rect 16324 73330 16436 73332
rect 16324 73278 16382 73330
rect 16434 73278 16436 73330
rect 16324 73276 16436 73278
rect 14252 24770 14308 24780
rect 14812 24836 14868 24846
rect 12572 23492 12852 23548
rect 13468 23538 13524 23548
rect 13804 23604 13860 23614
rect 12348 15092 12404 23492
rect 12796 23156 12852 23492
rect 12348 15036 12516 15092
rect 12460 13076 12516 15036
rect 11900 13074 12516 13076
rect 11900 13022 12462 13074
rect 12514 13022 12516 13074
rect 11900 13020 12516 13022
rect 11900 12402 11956 13020
rect 12460 13010 12516 13020
rect 12796 12964 12852 23100
rect 13804 15148 13860 23548
rect 14028 18564 14084 18574
rect 14028 15148 14084 18508
rect 13804 15092 13972 15148
rect 14028 15092 14420 15148
rect 11900 12350 11902 12402
rect 11954 12350 11956 12402
rect 11564 11106 11620 11116
rect 11676 12178 11732 12190
rect 11676 12126 11678 12178
rect 11730 12126 11732 12178
rect 10332 10500 10388 10510
rect 10332 10406 10388 10444
rect 11676 10164 11732 12126
rect 11788 12068 11844 12078
rect 11788 11974 11844 12012
rect 11900 11506 11956 12350
rect 12572 12908 12852 12964
rect 11900 11454 11902 11506
rect 11954 11454 11956 11506
rect 11900 11442 11956 11454
rect 12348 12178 12404 12190
rect 12348 12126 12350 12178
rect 12402 12126 12404 12178
rect 12012 11172 12068 11182
rect 11788 10164 11844 10174
rect 11676 10108 11788 10164
rect 10108 9986 10164 9996
rect 11788 9826 11844 10108
rect 11788 9774 11790 9826
rect 11842 9774 11844 9826
rect 9660 8990 9662 9042
rect 9714 8990 9716 9042
rect 9324 8932 9380 8942
rect 9324 8370 9380 8876
rect 9324 8318 9326 8370
rect 9378 8318 9380 8370
rect 9324 8306 9380 8318
rect 9436 8148 9492 8158
rect 9436 8054 9492 8092
rect 9212 8036 9268 8046
rect 9212 8034 9380 8036
rect 9212 7982 9214 8034
rect 9266 7982 9380 8034
rect 9212 7980 9380 7982
rect 9212 7970 9268 7980
rect 9324 6916 9380 7980
rect 9660 7812 9716 8990
rect 11116 9604 11172 9614
rect 10332 8932 10388 8942
rect 10332 8838 10388 8876
rect 11004 8260 11060 8270
rect 11004 8166 11060 8204
rect 10668 8034 10724 8046
rect 10668 7982 10670 8034
rect 10722 7982 10724 8034
rect 9660 7746 9716 7756
rect 10556 7812 10612 7822
rect 10556 7474 10612 7756
rect 10556 7422 10558 7474
rect 10610 7422 10612 7474
rect 9884 7362 9940 7374
rect 9884 7310 9886 7362
rect 9938 7310 9940 7362
rect 9436 6916 9492 6926
rect 9324 6914 9492 6916
rect 9324 6862 9438 6914
rect 9490 6862 9492 6914
rect 9324 6860 9492 6862
rect 9884 6916 9940 7310
rect 10332 7364 10388 7374
rect 10332 7362 10500 7364
rect 10332 7310 10334 7362
rect 10386 7310 10500 7362
rect 10332 7308 10500 7310
rect 10332 7298 10388 7308
rect 9884 6860 10276 6916
rect 9436 6850 9492 6860
rect 8988 6750 8990 6802
rect 9042 6750 9044 6802
rect 8988 6738 9044 6750
rect 9100 6804 9156 6814
rect 8764 5742 8766 5794
rect 8818 5742 8820 5794
rect 8764 5730 8820 5742
rect 8876 6466 8932 6478
rect 8876 6414 8878 6466
rect 8930 6414 8932 6466
rect 8876 5348 8932 6414
rect 8988 6020 9044 6030
rect 9100 6020 9156 6748
rect 9772 6804 9828 6814
rect 9828 6748 10052 6804
rect 9772 6710 9828 6748
rect 9884 6580 9940 6590
rect 9996 6580 10052 6748
rect 10220 6692 10276 6860
rect 10332 6692 10388 6702
rect 10220 6690 10388 6692
rect 10220 6638 10334 6690
rect 10386 6638 10388 6690
rect 10220 6636 10388 6638
rect 10108 6580 10164 6590
rect 9996 6578 10164 6580
rect 9996 6526 10110 6578
rect 10162 6526 10164 6578
rect 9996 6524 10164 6526
rect 8988 6018 9156 6020
rect 8988 5966 8990 6018
rect 9042 5966 9156 6018
rect 8988 5964 9156 5966
rect 9548 6466 9604 6478
rect 9548 6414 9550 6466
rect 9602 6414 9604 6466
rect 8988 5954 9044 5964
rect 9548 5684 9604 6414
rect 9884 6132 9940 6524
rect 10108 6514 10164 6524
rect 10332 6132 10388 6636
rect 10444 6244 10500 7308
rect 10444 6178 10500 6188
rect 9884 6076 10052 6132
rect 9884 5908 9940 5918
rect 9884 5814 9940 5852
rect 9548 5618 9604 5628
rect 9436 5572 9492 5582
rect 8876 5282 8932 5292
rect 9324 5460 9380 5470
rect 8764 5124 8820 5134
rect 8764 5030 8820 5068
rect 8876 5122 8932 5134
rect 8876 5070 8878 5122
rect 8930 5070 8932 5122
rect 8428 4946 8484 4956
rect 8876 5012 8932 5070
rect 9212 5012 9268 5022
rect 8876 4956 9212 5012
rect 8652 4900 8708 4910
rect 8652 4806 8708 4844
rect 8876 4676 8932 4956
rect 9212 4918 9268 4956
rect 9324 4788 9380 5404
rect 8204 4510 8206 4562
rect 8258 4510 8260 4562
rect 8204 4498 8260 4510
rect 8316 4620 8932 4676
rect 8988 4732 9380 4788
rect 8316 4452 8372 4620
rect 8988 4562 9044 4732
rect 8988 4510 8990 4562
rect 9042 4510 9044 4562
rect 8988 4498 9044 4510
rect 9436 4564 9492 5516
rect 9548 5348 9604 5358
rect 9548 5122 9604 5292
rect 9548 5070 9550 5122
rect 9602 5070 9604 5122
rect 9548 5058 9604 5070
rect 9884 5012 9940 5022
rect 9884 4918 9940 4956
rect 8316 4358 8372 4396
rect 8764 4452 8820 4462
rect 8764 4338 8820 4396
rect 8764 4286 8766 4338
rect 8818 4286 8820 4338
rect 8092 4172 8484 4228
rect 7868 3892 7924 3902
rect 7756 3836 7868 3892
rect 7196 2942 7198 2994
rect 7250 2942 7252 2994
rect 7196 2930 7252 2942
rect 7644 800 7700 3836
rect 7868 3554 7924 3836
rect 7868 3502 7870 3554
rect 7922 3502 7924 3554
rect 7868 3490 7924 3502
rect 8316 3668 8372 3678
rect 8092 3444 8148 3482
rect 8092 3378 8148 3388
rect 8316 800 8372 3612
rect 8428 3668 8484 4172
rect 8764 4004 8820 4286
rect 8764 3938 8820 3948
rect 8988 3780 9044 3790
rect 8540 3668 8596 3678
rect 8428 3612 8540 3668
rect 8428 3554 8484 3612
rect 8540 3602 8596 3612
rect 8428 3502 8430 3554
rect 8482 3502 8484 3554
rect 8428 3490 8484 3502
rect 8764 3330 8820 3342
rect 8764 3278 8766 3330
rect 8818 3278 8820 3330
rect 8764 3220 8820 3278
rect 8764 3154 8820 3164
rect 8988 800 9044 3724
rect 9436 3556 9492 4508
rect 9772 4788 9828 4798
rect 9772 4452 9828 4732
rect 9996 4562 10052 6076
rect 10108 6076 10388 6132
rect 10108 5348 10164 6076
rect 10556 6020 10612 7422
rect 10220 5964 10612 6020
rect 10220 5906 10276 5964
rect 10220 5854 10222 5906
rect 10274 5854 10276 5906
rect 10220 5842 10276 5854
rect 10108 5282 10164 5292
rect 10220 5234 10276 5246
rect 10220 5182 10222 5234
rect 10274 5182 10276 5234
rect 9996 4510 9998 4562
rect 10050 4510 10052 4562
rect 9996 4498 10052 4510
rect 10108 4898 10164 4910
rect 10108 4846 10110 4898
rect 10162 4846 10164 4898
rect 9772 4338 9828 4396
rect 9772 4286 9774 4338
rect 9826 4286 9828 4338
rect 9772 4274 9828 4286
rect 9884 4340 9940 4350
rect 9548 3556 9604 3566
rect 9436 3554 9604 3556
rect 9436 3502 9550 3554
rect 9602 3502 9604 3554
rect 9436 3500 9604 3502
rect 9548 3490 9604 3500
rect 9884 3442 9940 4284
rect 10108 4116 10164 4846
rect 10220 4228 10276 5182
rect 10332 4900 10388 4910
rect 10332 4450 10388 4844
rect 10556 4788 10612 5964
rect 10668 6020 10724 7982
rect 11116 7476 11172 9548
rect 11788 8258 11844 9774
rect 12012 9826 12068 11116
rect 12012 9774 12014 9826
rect 12066 9774 12068 9826
rect 12012 9762 12068 9774
rect 12348 9828 12404 12126
rect 12460 11172 12516 11182
rect 12460 10498 12516 11116
rect 12460 10446 12462 10498
rect 12514 10446 12516 10498
rect 12460 9938 12516 10446
rect 12460 9886 12462 9938
rect 12514 9886 12516 9938
rect 12460 9874 12516 9886
rect 11900 9716 11956 9726
rect 11900 9622 11956 9660
rect 11788 8206 11790 8258
rect 11842 8206 11844 8258
rect 11788 8194 11844 8206
rect 12012 8260 12068 8270
rect 12012 8166 12068 8204
rect 12348 8258 12404 9772
rect 12348 8206 12350 8258
rect 12402 8206 12404 8258
rect 12348 8194 12404 8206
rect 12572 9266 12628 12908
rect 12684 12178 12740 12190
rect 12684 12126 12686 12178
rect 12738 12126 12740 12178
rect 12684 11844 12740 12126
rect 13356 12068 13412 12078
rect 12684 11778 12740 11788
rect 13244 12066 13412 12068
rect 13244 12014 13358 12066
rect 13410 12014 13412 12066
rect 13244 12012 13412 12014
rect 13020 11172 13076 11182
rect 13020 10164 13076 11116
rect 13244 10834 13300 12012
rect 13356 12002 13412 12012
rect 13692 11508 13748 11518
rect 13692 11394 13748 11452
rect 13692 11342 13694 11394
rect 13746 11342 13748 11394
rect 13692 11330 13748 11342
rect 13916 11396 13972 15092
rect 13916 11340 14308 11396
rect 13468 11172 13524 11182
rect 13468 11078 13524 11116
rect 13580 11170 13636 11182
rect 13580 11118 13582 11170
rect 13634 11118 13636 11170
rect 13244 10782 13246 10834
rect 13298 10782 13300 10834
rect 13244 10770 13300 10782
rect 12684 9940 12740 9950
rect 12684 9938 12852 9940
rect 12684 9886 12686 9938
rect 12738 9886 12852 9938
rect 12684 9884 12852 9886
rect 12684 9874 12740 9884
rect 12796 9826 12852 9884
rect 12796 9774 12798 9826
rect 12850 9774 12852 9826
rect 12796 9762 12852 9774
rect 12572 9214 12574 9266
rect 12626 9214 12628 9266
rect 12572 8260 12628 9214
rect 13020 9266 13076 10108
rect 13020 9214 13022 9266
rect 13074 9214 13076 9266
rect 13020 9202 13076 9214
rect 13132 10722 13188 10734
rect 13132 10670 13134 10722
rect 13186 10670 13188 10722
rect 13132 8484 13188 10670
rect 13356 10724 13412 10734
rect 13580 10724 13636 11118
rect 13356 10722 13636 10724
rect 13356 10670 13358 10722
rect 13410 10670 13636 10722
rect 13356 10668 13636 10670
rect 13916 11170 13972 11182
rect 13916 11118 13918 11170
rect 13970 11118 13972 11170
rect 13356 10658 13412 10668
rect 13804 10500 13860 10510
rect 13580 10444 13804 10500
rect 13356 10164 13412 10174
rect 13356 9266 13412 10108
rect 13468 9828 13524 9838
rect 13468 9714 13524 9772
rect 13468 9662 13470 9714
rect 13522 9662 13524 9714
rect 13468 9650 13524 9662
rect 13356 9214 13358 9266
rect 13410 9214 13412 9266
rect 13356 9202 13412 9214
rect 13132 8418 13188 8428
rect 12572 8194 12628 8204
rect 11900 8148 11956 8158
rect 11900 8054 11956 8092
rect 13020 8148 13076 8158
rect 13020 8054 13076 8092
rect 11004 7420 11172 7476
rect 11452 8034 11508 8046
rect 11452 7982 11454 8034
rect 11506 7982 11508 8034
rect 11452 7476 11508 7982
rect 10892 6916 10948 6926
rect 10892 6690 10948 6860
rect 10892 6638 10894 6690
rect 10946 6638 10948 6690
rect 10892 6626 10948 6638
rect 11004 6020 11060 7420
rect 11452 7410 11508 7420
rect 13468 7476 13524 7486
rect 11340 7364 11396 7374
rect 11676 7364 11732 7374
rect 11116 7362 11396 7364
rect 11116 7310 11342 7362
rect 11394 7310 11396 7362
rect 11116 7308 11396 7310
rect 11116 6802 11172 7308
rect 11340 7298 11396 7308
rect 11564 7308 11676 7364
rect 11228 6916 11284 6926
rect 11228 6822 11284 6860
rect 11116 6750 11118 6802
rect 11170 6750 11172 6802
rect 11116 6738 11172 6750
rect 11228 6020 11284 6030
rect 11004 5964 11172 6020
rect 10668 5954 10724 5964
rect 10892 5796 10948 5806
rect 10780 5794 10948 5796
rect 10780 5742 10894 5794
rect 10946 5742 10948 5794
rect 10780 5740 10948 5742
rect 10668 5236 10724 5246
rect 10668 5010 10724 5180
rect 10780 5234 10836 5740
rect 10892 5730 10948 5740
rect 10780 5182 10782 5234
rect 10834 5182 10836 5234
rect 10780 5170 10836 5182
rect 10892 5236 10948 5246
rect 10892 5142 10948 5180
rect 10668 4958 10670 5010
rect 10722 4958 10724 5010
rect 10668 4946 10724 4958
rect 10556 4732 11060 4788
rect 10332 4398 10334 4450
rect 10386 4398 10388 4450
rect 10332 4386 10388 4398
rect 10668 4452 10724 4462
rect 10668 4450 10948 4452
rect 10668 4398 10670 4450
rect 10722 4398 10948 4450
rect 10668 4396 10948 4398
rect 10668 4386 10724 4396
rect 10220 4162 10276 4172
rect 10108 4050 10164 4060
rect 10892 4116 10948 4396
rect 11004 4338 11060 4732
rect 11004 4286 11006 4338
rect 11058 4286 11060 4338
rect 11004 4274 11060 4286
rect 10892 4050 10948 4060
rect 10332 4004 10388 4014
rect 10220 3780 10276 3790
rect 10220 3554 10276 3724
rect 10220 3502 10222 3554
rect 10274 3502 10276 3554
rect 10220 3490 10276 3502
rect 9884 3390 9886 3442
rect 9938 3390 9940 3442
rect 9884 3378 9940 3390
rect 9660 2994 9716 3006
rect 9660 2942 9662 2994
rect 9714 2942 9716 2994
rect 9660 800 9716 2942
rect 10332 800 10388 3948
rect 10780 4004 10836 4014
rect 10780 3780 10836 3948
rect 10780 3714 10836 3724
rect 11004 3780 11060 3790
rect 10556 3668 10612 3678
rect 10556 3442 10612 3612
rect 10556 3390 10558 3442
rect 10610 3390 10612 3442
rect 10556 3378 10612 3390
rect 10892 3554 10948 3566
rect 10892 3502 10894 3554
rect 10946 3502 10948 3554
rect 10892 3444 10948 3502
rect 10892 3378 10948 3388
rect 11004 800 11060 3724
rect 11116 3666 11172 5964
rect 11228 4004 11284 5964
rect 11228 3938 11284 3948
rect 11340 5348 11396 5358
rect 11564 5348 11620 7308
rect 11676 7298 11732 7308
rect 13468 7362 13524 7420
rect 13468 7310 13470 7362
rect 13522 7310 13524 7362
rect 13468 7298 13524 7310
rect 13244 6692 13300 6702
rect 12124 6468 12180 6478
rect 12124 6374 12180 6412
rect 12572 6466 12628 6478
rect 12572 6414 12574 6466
rect 12626 6414 12628 6466
rect 11116 3614 11118 3666
rect 11170 3614 11172 3666
rect 11116 3602 11172 3614
rect 11228 3444 11284 3482
rect 11228 3378 11284 3388
rect 11340 2436 11396 5292
rect 11452 5292 11620 5348
rect 12236 6244 12292 6254
rect 11452 4900 11508 5292
rect 11564 5124 11620 5134
rect 11564 5030 11620 5068
rect 11900 5124 11956 5134
rect 11900 5030 11956 5068
rect 11676 4900 11732 4910
rect 11452 4844 11620 4900
rect 11452 4116 11508 4126
rect 11452 3556 11508 4060
rect 11564 3778 11620 4844
rect 11564 3726 11566 3778
rect 11618 3726 11620 3778
rect 11564 3714 11620 3726
rect 11564 3556 11620 3566
rect 11452 3554 11620 3556
rect 11452 3502 11566 3554
rect 11618 3502 11620 3554
rect 11452 3500 11620 3502
rect 11564 3490 11620 3500
rect 11340 2370 11396 2380
rect 11676 800 11732 4844
rect 11788 4898 11844 4910
rect 11788 4846 11790 4898
rect 11842 4846 11844 4898
rect 11788 4450 11844 4846
rect 11788 4398 11790 4450
rect 11842 4398 11844 4450
rect 11788 4386 11844 4398
rect 11900 3444 11956 3482
rect 11900 3332 11956 3388
rect 11900 3266 11956 3276
rect 12236 3442 12292 6188
rect 12460 5796 12516 5806
rect 12460 5460 12516 5740
rect 12572 5684 12628 6414
rect 13020 6468 13076 6478
rect 13020 6466 13188 6468
rect 13020 6414 13022 6466
rect 13074 6414 13188 6466
rect 13020 6412 13188 6414
rect 13020 6402 13076 6412
rect 13020 6020 13076 6030
rect 12572 5618 12628 5628
rect 12908 5964 13020 6020
rect 12460 5404 12628 5460
rect 12460 5124 12516 5134
rect 12460 5030 12516 5068
rect 12572 5012 12628 5404
rect 12572 4918 12628 4956
rect 12348 4900 12404 4910
rect 12348 4806 12404 4844
rect 12572 4004 12628 4014
rect 12236 3390 12238 3442
rect 12290 3390 12292 3442
rect 12236 2994 12292 3390
rect 12236 2942 12238 2994
rect 12290 2942 12292 2994
rect 12236 2930 12292 2942
rect 12348 3556 12404 3566
rect 12348 800 12404 3500
rect 12572 3442 12628 3948
rect 12572 3390 12574 3442
rect 12626 3390 12628 3442
rect 12572 3378 12628 3390
rect 12908 3388 12964 5964
rect 13020 5954 13076 5964
rect 13020 5794 13076 5806
rect 13020 5742 13022 5794
rect 13074 5742 13076 5794
rect 13020 5572 13076 5742
rect 13132 5796 13188 6412
rect 13132 5730 13188 5740
rect 13244 6132 13300 6636
rect 13244 5572 13300 6076
rect 13020 5516 13300 5572
rect 13244 5348 13300 5516
rect 13244 5282 13300 5292
rect 13468 6468 13524 6478
rect 13020 5124 13076 5134
rect 13020 5030 13076 5068
rect 13468 5122 13524 6412
rect 13580 6020 13636 10444
rect 13804 10434 13860 10444
rect 13804 9940 13860 9950
rect 13804 9602 13860 9884
rect 13916 9828 13972 11118
rect 14140 10498 14196 10510
rect 14140 10446 14142 10498
rect 14194 10446 14196 10498
rect 13916 9762 13972 9772
rect 14028 10164 14084 10174
rect 13804 9550 13806 9602
rect 13858 9550 13860 9602
rect 13580 5926 13636 5964
rect 13692 9042 13748 9054
rect 13692 8990 13694 9042
rect 13746 8990 13748 9042
rect 13692 7812 13748 8990
rect 13804 8932 13860 9550
rect 13804 8866 13860 8876
rect 14028 8596 14084 10108
rect 14140 9940 14196 10446
rect 14140 9874 14196 9884
rect 13692 5572 13748 7756
rect 13804 8540 14084 8596
rect 13804 6690 13860 8540
rect 14252 8372 14308 11340
rect 13804 6638 13806 6690
rect 13858 6638 13860 6690
rect 13804 6626 13860 6638
rect 13916 8316 14308 8372
rect 13916 6692 13972 8316
rect 14252 8148 14308 8158
rect 14252 8054 14308 8092
rect 14028 8036 14084 8046
rect 14028 8034 14196 8036
rect 14028 7982 14030 8034
rect 14082 7982 14196 8034
rect 14028 7980 14196 7982
rect 14028 7970 14084 7980
rect 14140 7700 14196 7980
rect 14364 7924 14420 15092
rect 14476 11508 14532 11518
rect 14476 11414 14532 11452
rect 14476 10500 14532 10510
rect 14476 10406 14532 10444
rect 14700 9716 14756 9726
rect 14700 9622 14756 9660
rect 14476 9604 14532 9614
rect 14476 9510 14532 9548
rect 14588 9602 14644 9614
rect 14588 9550 14590 9602
rect 14642 9550 14644 9602
rect 14476 9156 14532 9166
rect 14588 9156 14644 9550
rect 14476 9154 14644 9156
rect 14476 9102 14478 9154
rect 14530 9102 14644 9154
rect 14476 9100 14644 9102
rect 14476 9090 14532 9100
rect 14588 8932 14644 8942
rect 14588 8146 14644 8876
rect 14588 8094 14590 8146
rect 14642 8094 14644 8146
rect 14588 8082 14644 8094
rect 14364 7858 14420 7868
rect 14140 7644 14420 7700
rect 13916 6626 13972 6636
rect 14028 7474 14084 7486
rect 14028 7422 14030 7474
rect 14082 7422 14084 7474
rect 14028 6468 14084 7422
rect 14252 7476 14308 7486
rect 14252 7382 14308 7420
rect 14140 7362 14196 7374
rect 14140 7310 14142 7362
rect 14194 7310 14196 7362
rect 14140 6916 14196 7310
rect 14140 6850 14196 6860
rect 14028 6132 14084 6412
rect 14252 6132 14308 6142
rect 14028 6130 14308 6132
rect 14028 6078 14254 6130
rect 14306 6078 14308 6130
rect 14028 6076 14308 6078
rect 14364 6132 14420 7644
rect 14700 7474 14756 7486
rect 14700 7422 14702 7474
rect 14754 7422 14756 7474
rect 14476 6468 14532 6478
rect 14476 6374 14532 6412
rect 14700 6468 14756 7422
rect 14812 7476 14868 24780
rect 16268 23604 16324 73276
rect 16380 73266 16436 73276
rect 16492 55468 16548 74846
rect 17948 74786 18004 74798
rect 17948 74734 17950 74786
rect 18002 74734 18004 74786
rect 17612 74114 17668 74126
rect 17612 74062 17614 74114
rect 17666 74062 17668 74114
rect 17612 73220 17668 74062
rect 17948 74116 18004 74734
rect 18060 74788 18116 74956
rect 18284 74788 18340 74798
rect 18060 74786 18340 74788
rect 18060 74734 18286 74786
rect 18338 74734 18340 74786
rect 18060 74732 18340 74734
rect 18172 74116 18228 74126
rect 17948 74114 18228 74116
rect 17948 74062 18174 74114
rect 18226 74062 18228 74114
rect 17948 74060 18228 74062
rect 17612 73154 17668 73164
rect 17836 73444 17892 73454
rect 16380 55412 16548 55468
rect 16380 43708 16436 55412
rect 16380 43652 16772 43708
rect 16268 23538 16324 23548
rect 16604 24724 16660 24734
rect 16604 22370 16660 24668
rect 16604 22318 16606 22370
rect 16658 22318 16660 22370
rect 16604 22306 16660 22318
rect 16716 23044 16772 43652
rect 17836 29428 17892 73388
rect 18172 73444 18228 74060
rect 18284 74004 18340 74732
rect 18284 73938 18340 73948
rect 18844 74788 18900 74798
rect 18172 73378 18228 73388
rect 18060 73220 18116 73230
rect 18116 73164 18340 73220
rect 18060 73126 18116 73164
rect 18284 67844 18340 73164
rect 18060 67788 18340 67844
rect 18060 43708 18116 67788
rect 18060 43652 18452 43708
rect 18060 29428 18116 29438
rect 17836 29372 18060 29428
rect 18060 29362 18116 29372
rect 17164 24836 17220 24846
rect 17164 24050 17220 24780
rect 17500 24724 17556 24734
rect 17500 24630 17556 24668
rect 17164 23998 17166 24050
rect 17218 23998 17220 24050
rect 17164 23828 17220 23998
rect 17612 24612 17668 24622
rect 17612 24050 17668 24556
rect 18172 24612 18228 24622
rect 18172 24518 18228 24556
rect 18396 24612 18452 43652
rect 18396 24546 18452 24556
rect 17612 23998 17614 24050
rect 17666 23998 17668 24050
rect 17612 23986 17668 23998
rect 17724 24276 17780 24286
rect 17724 23938 17780 24220
rect 18396 24276 18452 24286
rect 18172 23996 18340 24052
rect 17724 23886 17726 23938
rect 17778 23886 17780 23938
rect 17724 23874 17780 23886
rect 18060 23940 18116 23950
rect 17164 23762 17220 23772
rect 17500 23716 17556 23726
rect 17276 23714 17556 23716
rect 17276 23662 17502 23714
rect 17554 23662 17556 23714
rect 17276 23660 17556 23662
rect 16828 23268 16884 23278
rect 16828 23044 16884 23212
rect 16716 23042 16884 23044
rect 16716 22990 16830 23042
rect 16882 22990 16884 23042
rect 16716 22988 16884 22990
rect 15596 21700 15652 21710
rect 15596 21476 15652 21644
rect 15596 12402 15652 21420
rect 16716 18564 16772 22988
rect 16828 22978 16884 22988
rect 17276 22484 17332 23660
rect 17500 23650 17556 23660
rect 17948 23716 18004 23726
rect 17612 23492 17668 23502
rect 17500 23268 17556 23278
rect 17500 23174 17556 23212
rect 17612 23266 17668 23436
rect 17612 23214 17614 23266
rect 17666 23214 17668 23266
rect 17612 23202 17668 23214
rect 17164 22428 17332 22484
rect 17500 22930 17556 22942
rect 17500 22878 17502 22930
rect 17554 22878 17556 22930
rect 17164 21588 17220 22428
rect 17276 22260 17332 22270
rect 17276 22258 17444 22260
rect 17276 22206 17278 22258
rect 17330 22206 17444 22258
rect 17276 22204 17444 22206
rect 17276 22194 17332 22204
rect 17164 21522 17220 21532
rect 17276 22036 17332 22046
rect 16716 18498 16772 18508
rect 15596 12350 15598 12402
rect 15650 12350 15652 12402
rect 15372 11844 15428 11854
rect 15372 11394 15428 11788
rect 15596 11508 15652 12350
rect 16604 12962 16660 12974
rect 16604 12910 16606 12962
rect 16658 12910 16660 12962
rect 16604 11844 16660 12910
rect 16604 11778 16660 11788
rect 15596 11442 15652 11452
rect 15372 11342 15374 11394
rect 15426 11342 15428 11394
rect 15148 10498 15204 10510
rect 15148 10446 15150 10498
rect 15202 10446 15204 10498
rect 14812 7410 14868 7420
rect 14924 8596 14980 8606
rect 14924 8258 14980 8540
rect 14924 8206 14926 8258
rect 14978 8206 14980 8258
rect 14924 7812 14980 8206
rect 14924 6692 14980 7756
rect 14924 6626 14980 6636
rect 15036 8148 15092 8158
rect 15036 6690 15092 8092
rect 15036 6638 15038 6690
rect 15090 6638 15092 6690
rect 15036 6626 15092 6638
rect 14700 6374 14756 6412
rect 15148 6132 15204 10446
rect 15372 9938 15428 11342
rect 16044 11284 16100 11294
rect 16044 11282 16212 11284
rect 16044 11230 16046 11282
rect 16098 11230 16212 11282
rect 16044 11228 16212 11230
rect 16044 11218 16100 11228
rect 15596 10500 15652 10510
rect 15596 10498 15988 10500
rect 15596 10446 15598 10498
rect 15650 10446 15988 10498
rect 15596 10444 15988 10446
rect 15596 10434 15652 10444
rect 15372 9886 15374 9938
rect 15426 9886 15428 9938
rect 15372 8596 15428 9886
rect 15372 8530 15428 8540
rect 15596 9044 15652 9054
rect 15484 7476 15540 7514
rect 15484 7410 15540 7420
rect 15260 7364 15316 7374
rect 15260 7270 15316 7308
rect 14364 6076 14644 6132
rect 15148 6076 15540 6132
rect 14252 6066 14308 6076
rect 13916 6020 13972 6030
rect 13916 5926 13972 5964
rect 14476 5908 14532 5918
rect 14476 5814 14532 5852
rect 14364 5796 14420 5806
rect 13692 5506 13748 5516
rect 13804 5794 14420 5796
rect 13804 5742 14366 5794
rect 14418 5742 14420 5794
rect 13804 5740 14420 5742
rect 13692 5348 13748 5358
rect 13580 5236 13636 5246
rect 13580 5142 13636 5180
rect 13468 5070 13470 5122
rect 13522 5070 13524 5122
rect 13468 4900 13524 5070
rect 13692 5010 13748 5292
rect 13692 4958 13694 5010
rect 13746 4958 13748 5010
rect 13692 4946 13748 4958
rect 13468 4834 13524 4844
rect 13468 4452 13524 4462
rect 13356 4228 13412 4238
rect 13356 3554 13412 4172
rect 13356 3502 13358 3554
rect 13410 3502 13412 3554
rect 13356 3490 13412 3502
rect 12908 3332 13076 3388
rect 13020 800 13076 3332
rect 13468 3108 13524 4396
rect 13692 3780 13748 3790
rect 13804 3780 13860 5740
rect 14364 5730 14420 5740
rect 14364 5572 14420 5582
rect 14028 5348 14084 5358
rect 13916 5236 13972 5246
rect 13916 5012 13972 5180
rect 13916 4226 13972 4956
rect 13916 4174 13918 4226
rect 13970 4174 13972 4226
rect 13916 4162 13972 4174
rect 13692 3778 13860 3780
rect 13692 3726 13694 3778
rect 13746 3726 13860 3778
rect 13692 3724 13860 3726
rect 13692 3714 13748 3724
rect 13580 3556 13636 3566
rect 14028 3556 14084 5292
rect 14140 5124 14196 5134
rect 14140 5030 14196 5068
rect 14364 5122 14420 5516
rect 14364 5070 14366 5122
rect 14418 5070 14420 5122
rect 14364 5058 14420 5070
rect 14588 4900 14644 6076
rect 14700 6018 14756 6030
rect 14700 5966 14702 6018
rect 14754 5966 14756 6018
rect 14700 5124 14756 5966
rect 14812 6020 14868 6030
rect 14812 5572 14868 5964
rect 15372 5908 15428 5918
rect 14812 5506 14868 5516
rect 15260 5906 15428 5908
rect 15260 5854 15374 5906
rect 15426 5854 15428 5906
rect 15260 5852 15428 5854
rect 15260 5460 15316 5852
rect 15372 5842 15428 5852
rect 15260 5394 15316 5404
rect 15372 5684 15428 5694
rect 15148 5348 15204 5358
rect 15148 5234 15204 5292
rect 15372 5236 15428 5628
rect 15148 5182 15150 5234
rect 15202 5182 15204 5234
rect 15148 5170 15204 5182
rect 15260 5180 15428 5236
rect 14700 5058 14756 5068
rect 14588 4844 14756 4900
rect 14252 4564 14308 4574
rect 13580 3554 14084 3556
rect 13580 3502 13582 3554
rect 13634 3502 14084 3554
rect 13580 3500 14084 3502
rect 14140 3556 14196 3566
rect 13580 3490 13636 3500
rect 14140 3462 14196 3500
rect 13468 3052 13748 3108
rect 13692 800 13748 3052
rect 14252 2100 14308 4508
rect 14588 4338 14644 4350
rect 14588 4286 14590 4338
rect 14642 4286 14644 4338
rect 14588 3780 14644 4286
rect 14588 3714 14644 3724
rect 14700 3554 14756 4844
rect 14812 4452 14868 4462
rect 14812 4358 14868 4396
rect 15148 4338 15204 4350
rect 15148 4286 15150 4338
rect 15202 4286 15204 4338
rect 14700 3502 14702 3554
rect 14754 3502 14756 3554
rect 14700 3444 14756 3502
rect 14700 3378 14756 3388
rect 14812 3892 14868 3902
rect 14812 3388 14868 3836
rect 15036 3892 15092 3902
rect 15036 3442 15092 3836
rect 15036 3390 15038 3442
rect 15090 3390 15092 3442
rect 14364 3330 14420 3342
rect 14812 3332 14980 3388
rect 15036 3378 15092 3390
rect 14364 3278 14366 3330
rect 14418 3278 14420 3330
rect 14364 2324 14420 3278
rect 14924 3220 14980 3332
rect 15148 3220 15204 4286
rect 15260 4340 15316 5180
rect 15372 5012 15428 5022
rect 15372 4562 15428 4956
rect 15484 4788 15540 6076
rect 15596 6130 15652 8988
rect 15708 8146 15764 8158
rect 15708 8094 15710 8146
rect 15762 8094 15764 8146
rect 15708 7698 15764 8094
rect 15708 7646 15710 7698
rect 15762 7646 15764 7698
rect 15708 7634 15764 7646
rect 15820 8036 15876 8046
rect 15820 7586 15876 7980
rect 15820 7534 15822 7586
rect 15874 7534 15876 7586
rect 15820 7522 15876 7534
rect 15708 6468 15764 6478
rect 15708 6374 15764 6412
rect 15596 6078 15598 6130
rect 15650 6078 15652 6130
rect 15596 6066 15652 6078
rect 15708 5684 15764 5694
rect 15708 5682 15876 5684
rect 15708 5630 15710 5682
rect 15762 5630 15876 5682
rect 15708 5628 15876 5630
rect 15708 5618 15764 5628
rect 15484 4722 15540 4732
rect 15820 4564 15876 5628
rect 15372 4510 15374 4562
rect 15426 4510 15428 4562
rect 15372 4498 15428 4510
rect 15484 4562 15876 4564
rect 15484 4510 15822 4562
rect 15874 4510 15876 4562
rect 15484 4508 15876 4510
rect 15484 4450 15540 4508
rect 15820 4498 15876 4508
rect 15484 4398 15486 4450
rect 15538 4398 15540 4450
rect 15260 4284 15428 4340
rect 15372 3556 15428 4284
rect 15372 3462 15428 3500
rect 15484 3332 15540 4398
rect 15932 4340 15988 10444
rect 16044 10498 16100 10510
rect 16044 10446 16046 10498
rect 16098 10446 16100 10498
rect 16044 8148 16100 10446
rect 16156 9268 16212 11228
rect 16156 9202 16212 9212
rect 16716 9380 16772 9390
rect 16716 9268 16772 9324
rect 16716 9266 16996 9268
rect 16716 9214 16718 9266
rect 16770 9214 16996 9266
rect 16716 9212 16996 9214
rect 16716 9202 16772 9212
rect 16380 8596 16436 8606
rect 16044 8082 16100 8092
rect 16268 8540 16380 8596
rect 16156 6580 16212 6590
rect 16156 6486 16212 6524
rect 16156 6132 16212 6142
rect 15484 3266 15540 3276
rect 15596 4284 15988 4340
rect 16044 6076 16156 6132
rect 15596 3780 15652 4284
rect 14924 3164 15092 3220
rect 14364 2258 14420 2268
rect 14252 2044 14420 2100
rect 14364 800 14420 2044
rect 15036 800 15092 3164
rect 15148 3154 15204 3164
rect 15596 1764 15652 3724
rect 15708 3444 15764 3454
rect 16044 3444 16100 6076
rect 16156 6066 16212 6076
rect 16156 4452 16212 4462
rect 16268 4452 16324 8540
rect 16380 8530 16436 8540
rect 16716 8484 16772 8494
rect 16492 8372 16548 8382
rect 16492 7698 16548 8316
rect 16492 7646 16494 7698
rect 16546 7646 16548 7698
rect 16492 7634 16548 7646
rect 16380 6692 16436 6702
rect 16380 6598 16436 6636
rect 16492 5794 16548 5806
rect 16492 5742 16494 5794
rect 16546 5742 16548 5794
rect 16492 4564 16548 5742
rect 16492 4498 16548 4508
rect 16716 4562 16772 8428
rect 16940 7698 16996 9212
rect 16940 7646 16942 7698
rect 16994 7646 16996 7698
rect 16940 7634 16996 7646
rect 17052 7364 17108 7374
rect 16716 4510 16718 4562
rect 16770 4510 16772 4562
rect 16716 4498 16772 4510
rect 16828 5796 16884 5806
rect 16156 4450 16324 4452
rect 16156 4398 16158 4450
rect 16210 4398 16324 4450
rect 16156 4396 16324 4398
rect 16156 3554 16212 4396
rect 16492 4340 16548 4350
rect 16492 4246 16548 4284
rect 16828 4340 16884 5740
rect 16828 4274 16884 4284
rect 16940 5794 16996 5806
rect 16940 5742 16942 5794
rect 16994 5742 16996 5794
rect 16156 3502 16158 3554
rect 16210 3502 16212 3554
rect 16156 3490 16212 3502
rect 16828 4116 16884 4126
rect 15708 3442 16100 3444
rect 15708 3390 15710 3442
rect 15762 3390 16100 3442
rect 15708 3388 16100 3390
rect 16380 3444 16436 3454
rect 16828 3444 16884 4060
rect 16940 3780 16996 5742
rect 17052 4788 17108 7308
rect 17164 6692 17220 6702
rect 17164 6598 17220 6636
rect 17052 4722 17108 4732
rect 17164 6356 17220 6366
rect 16940 3714 16996 3724
rect 17052 4228 17108 4238
rect 16380 3442 16884 3444
rect 16380 3390 16382 3442
rect 16434 3390 16884 3442
rect 16380 3388 16884 3390
rect 15708 3378 15764 3388
rect 16380 3378 16436 3388
rect 16380 2994 16436 3006
rect 16380 2942 16382 2994
rect 16434 2942 16436 2994
rect 15596 1708 15764 1764
rect 15708 800 15764 1708
rect 16380 800 16436 2942
rect 17052 800 17108 4172
rect 17164 4228 17220 6300
rect 17276 5908 17332 21980
rect 17388 21588 17444 22204
rect 17500 21810 17556 22878
rect 17948 22036 18004 23660
rect 17948 21970 18004 21980
rect 17836 21812 17892 21822
rect 17500 21758 17502 21810
rect 17554 21758 17556 21810
rect 17500 21746 17556 21758
rect 17612 21810 17892 21812
rect 17612 21758 17838 21810
rect 17890 21758 17892 21810
rect 17612 21756 17892 21758
rect 17612 21588 17668 21756
rect 17836 21746 17892 21756
rect 17388 21532 17668 21588
rect 17724 21586 17780 21598
rect 17724 21534 17726 21586
rect 17778 21534 17780 21586
rect 17724 21364 17780 21534
rect 17948 21588 18004 21598
rect 17948 21494 18004 21532
rect 17724 21298 17780 21308
rect 17612 18676 17668 18686
rect 18060 18676 18116 23884
rect 18172 23938 18228 23996
rect 18172 23886 18174 23938
rect 18226 23886 18228 23938
rect 18172 23874 18228 23886
rect 18284 23938 18340 23996
rect 18284 23886 18286 23938
rect 18338 23886 18340 23938
rect 18284 23874 18340 23886
rect 18396 23378 18452 24220
rect 18620 23938 18676 23950
rect 18620 23886 18622 23938
rect 18674 23886 18676 23938
rect 18508 23828 18564 23838
rect 18508 23734 18564 23772
rect 18620 23828 18676 23886
rect 18732 23828 18788 23838
rect 18620 23772 18732 23828
rect 18620 23492 18676 23772
rect 18732 23762 18788 23772
rect 18620 23426 18676 23436
rect 18396 23326 18398 23378
rect 18450 23326 18452 23378
rect 18396 23314 18452 23326
rect 18732 22148 18788 22158
rect 18396 21474 18452 21486
rect 18396 21422 18398 21474
rect 18450 21422 18452 21474
rect 18396 21364 18452 21422
rect 18396 21298 18452 21308
rect 18620 20804 18676 20814
rect 18508 20748 18620 20804
rect 18396 20132 18452 20142
rect 17612 18674 18116 18676
rect 17612 18622 17614 18674
rect 17666 18622 18062 18674
rect 18114 18622 18116 18674
rect 17612 18620 18116 18622
rect 17612 18610 17668 18620
rect 17948 15148 18004 18620
rect 18060 18610 18116 18620
rect 18172 18676 18228 18686
rect 18396 18676 18452 20076
rect 18228 18620 18452 18676
rect 18172 18562 18228 18620
rect 18172 18510 18174 18562
rect 18226 18510 18228 18562
rect 18172 18498 18228 18510
rect 18060 18228 18116 18238
rect 18060 18134 18116 18172
rect 17500 15092 18004 15148
rect 17388 12850 17444 12862
rect 17388 12798 17390 12850
rect 17442 12798 17444 12850
rect 17388 12402 17444 12798
rect 17388 12350 17390 12402
rect 17442 12350 17444 12402
rect 17388 12338 17444 12350
rect 17388 9044 17444 9054
rect 17388 8950 17444 8988
rect 17500 8932 17556 15092
rect 18060 13636 18116 13646
rect 17612 12290 17668 12302
rect 17612 12238 17614 12290
rect 17666 12238 17668 12290
rect 17612 12068 17668 12238
rect 17836 12290 17892 12302
rect 17836 12238 17838 12290
rect 17890 12238 17892 12290
rect 17724 12068 17780 12078
rect 17612 12066 17780 12068
rect 17612 12014 17726 12066
rect 17778 12014 17780 12066
rect 17612 12012 17780 12014
rect 17724 12002 17780 12012
rect 17836 10948 17892 12238
rect 18060 12290 18116 13580
rect 18060 12238 18062 12290
rect 18114 12238 18116 12290
rect 18060 12226 18116 12238
rect 18508 12402 18564 20748
rect 18620 20710 18676 20748
rect 18732 20242 18788 22092
rect 18732 20190 18734 20242
rect 18786 20190 18788 20242
rect 18732 20178 18788 20190
rect 18844 19348 18900 74732
rect 19180 74338 19236 75516
rect 19180 74286 19182 74338
rect 19234 74286 19236 74338
rect 19180 74274 19236 74286
rect 19404 74786 19460 76412
rect 20076 75572 20132 76636
rect 20636 75908 20692 79200
rect 21084 76692 21140 76702
rect 21084 76598 21140 76636
rect 20636 75842 20692 75852
rect 20748 76356 20804 76366
rect 21308 76356 21364 79200
rect 21980 76692 22036 79200
rect 22652 77252 22708 79200
rect 22652 77196 23156 77252
rect 21980 76626 22036 76636
rect 21644 76356 21700 76366
rect 21308 76354 21700 76356
rect 21308 76302 21646 76354
rect 21698 76302 21700 76354
rect 21308 76300 21700 76302
rect 20300 75682 20356 75694
rect 20300 75630 20302 75682
rect 20354 75630 20356 75682
rect 20076 75516 20244 75572
rect 19836 75292 20100 75302
rect 19892 75236 19940 75292
rect 19996 75236 20044 75292
rect 19836 75226 20100 75236
rect 19404 74734 19406 74786
rect 19458 74734 19460 74786
rect 19404 55468 19460 74734
rect 19852 74788 19908 74798
rect 19852 74694 19908 74732
rect 20188 74564 20244 75516
rect 20300 74788 20356 75630
rect 20300 74722 20356 74732
rect 20412 74786 20468 74798
rect 20412 74734 20414 74786
rect 20466 74734 20468 74786
rect 20412 74564 20468 74734
rect 20188 74508 20468 74564
rect 19836 73724 20100 73734
rect 19892 73668 19940 73724
rect 19996 73668 20044 73724
rect 19836 73658 20100 73668
rect 19836 72156 20100 72166
rect 19892 72100 19940 72156
rect 19996 72100 20044 72156
rect 19836 72090 20100 72100
rect 19836 70588 20100 70598
rect 19892 70532 19940 70588
rect 19996 70532 20044 70588
rect 19836 70522 20100 70532
rect 19836 69020 20100 69030
rect 19892 68964 19940 69020
rect 19996 68964 20044 69020
rect 19836 68954 20100 68964
rect 19836 67452 20100 67462
rect 19892 67396 19940 67452
rect 19996 67396 20044 67452
rect 19836 67386 20100 67396
rect 19836 65884 20100 65894
rect 19892 65828 19940 65884
rect 19996 65828 20044 65884
rect 19836 65818 20100 65828
rect 19836 64316 20100 64326
rect 19892 64260 19940 64316
rect 19996 64260 20044 64316
rect 19836 64250 20100 64260
rect 19836 62748 20100 62758
rect 19892 62692 19940 62748
rect 19996 62692 20044 62748
rect 19836 62682 20100 62692
rect 19836 61180 20100 61190
rect 19892 61124 19940 61180
rect 19996 61124 20044 61180
rect 19836 61114 20100 61124
rect 19836 59612 20100 59622
rect 19892 59556 19940 59612
rect 19996 59556 20044 59612
rect 19836 59546 20100 59556
rect 19836 58044 20100 58054
rect 19892 57988 19940 58044
rect 19996 57988 20044 58044
rect 19836 57978 20100 57988
rect 19836 56476 20100 56486
rect 19892 56420 19940 56476
rect 19996 56420 20044 56476
rect 19836 56410 20100 56420
rect 19292 55412 19460 55468
rect 19180 23044 19236 23054
rect 19180 22036 19236 22988
rect 19180 21970 19236 21980
rect 19292 21924 19348 55412
rect 19836 54908 20100 54918
rect 19892 54852 19940 54908
rect 19996 54852 20044 54908
rect 19836 54842 20100 54852
rect 19836 53340 20100 53350
rect 19892 53284 19940 53340
rect 19996 53284 20044 53340
rect 19836 53274 20100 53284
rect 19836 51772 20100 51782
rect 19892 51716 19940 51772
rect 19996 51716 20044 51772
rect 19836 51706 20100 51716
rect 19836 50204 20100 50214
rect 19892 50148 19940 50204
rect 19996 50148 20044 50204
rect 19836 50138 20100 50148
rect 19836 48636 20100 48646
rect 19892 48580 19940 48636
rect 19996 48580 20044 48636
rect 19836 48570 20100 48580
rect 19836 47068 20100 47078
rect 19892 47012 19940 47068
rect 19996 47012 20044 47068
rect 19836 47002 20100 47012
rect 19836 45500 20100 45510
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 19836 45434 20100 45444
rect 19836 43932 20100 43942
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 19836 43866 20100 43876
rect 19836 42364 20100 42374
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 19836 42298 20100 42308
rect 19836 40796 20100 40806
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 19836 40730 20100 40740
rect 19836 39228 20100 39238
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 19836 39162 20100 39172
rect 19836 37660 20100 37670
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 19836 37594 20100 37604
rect 19836 36092 20100 36102
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 19836 36026 20100 36036
rect 19836 34524 20100 34534
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 19836 34458 20100 34468
rect 19836 32956 20100 32966
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 19836 32890 20100 32900
rect 20748 31948 20804 76300
rect 21644 76290 21700 76300
rect 21980 75908 22036 75918
rect 21980 75814 22036 75852
rect 23100 75122 23156 77196
rect 23100 75070 23102 75122
rect 23154 75070 23156 75122
rect 23100 75058 23156 75070
rect 23324 75124 23380 79200
rect 23772 76466 23828 76478
rect 23772 76414 23774 76466
rect 23826 76414 23828 76466
rect 23772 75684 23828 76414
rect 23772 75618 23828 75628
rect 23884 75682 23940 75694
rect 23884 75630 23886 75682
rect 23938 75630 23940 75682
rect 23884 75348 23940 75630
rect 23996 75572 24052 79200
rect 24668 76692 24724 79200
rect 24892 76692 24948 76702
rect 24668 76690 24948 76692
rect 24668 76638 24894 76690
rect 24946 76638 24948 76690
rect 24668 76636 24948 76638
rect 25340 76692 25396 79200
rect 25564 76692 25620 76702
rect 25340 76690 25620 76692
rect 25340 76638 25566 76690
rect 25618 76638 25620 76690
rect 25340 76636 25620 76638
rect 26012 76692 26068 79200
rect 26236 76692 26292 76702
rect 26012 76690 26292 76692
rect 26012 76638 26238 76690
rect 26290 76638 26292 76690
rect 26012 76636 26292 76638
rect 26684 76692 26740 79200
rect 26908 76692 26964 76702
rect 26684 76690 26964 76692
rect 26684 76638 26910 76690
rect 26962 76638 26964 76690
rect 26684 76636 26964 76638
rect 27356 76692 27412 79200
rect 28028 77924 28084 79200
rect 28028 77868 28420 77924
rect 27580 76692 27636 76702
rect 27356 76690 27636 76692
rect 27356 76638 27582 76690
rect 27634 76638 27636 76690
rect 27356 76636 27636 76638
rect 24892 76626 24948 76636
rect 25564 76626 25620 76636
rect 26236 76626 26292 76636
rect 26908 76626 26964 76636
rect 27580 76626 27636 76636
rect 28364 76690 28420 77868
rect 28364 76638 28366 76690
rect 28418 76638 28420 76690
rect 28364 76626 28420 76638
rect 28700 76692 28756 79200
rect 28924 76692 28980 76702
rect 28700 76690 28980 76692
rect 28700 76638 28926 76690
rect 28978 76638 28980 76690
rect 28700 76636 28980 76638
rect 29372 76692 29428 79200
rect 29596 76692 29652 76702
rect 29372 76690 29652 76692
rect 29372 76638 29598 76690
rect 29650 76638 29652 76690
rect 29372 76636 29652 76638
rect 30044 76692 30100 79200
rect 30268 76692 30324 76702
rect 30044 76690 30324 76692
rect 30044 76638 30270 76690
rect 30322 76638 30324 76690
rect 30044 76636 30324 76638
rect 30716 76692 30772 79200
rect 30940 76692 30996 76702
rect 30716 76690 30996 76692
rect 30716 76638 30942 76690
rect 30994 76638 30996 76690
rect 30716 76636 30996 76638
rect 31388 76692 31444 79200
rect 31500 76692 31556 76702
rect 31388 76690 31556 76692
rect 31388 76638 31502 76690
rect 31554 76638 31556 76690
rect 31388 76636 31556 76638
rect 32060 76692 32116 79200
rect 32284 76692 32340 76702
rect 32060 76690 32340 76692
rect 32060 76638 32286 76690
rect 32338 76638 32340 76690
rect 32060 76636 32340 76638
rect 28924 76626 28980 76636
rect 29596 76626 29652 76636
rect 30268 76626 30324 76636
rect 30940 76626 30996 76636
rect 31500 76626 31556 76636
rect 32284 76626 32340 76636
rect 32732 75796 32788 79200
rect 33404 76354 33460 79200
rect 33404 76302 33406 76354
rect 33458 76302 33460 76354
rect 33404 76290 33460 76302
rect 34076 75908 34132 79200
rect 34076 75852 34692 75908
rect 33628 75796 33684 75806
rect 32732 75794 33012 75796
rect 32732 75742 32734 75794
rect 32786 75742 33012 75794
rect 32732 75740 33012 75742
rect 32732 75730 32788 75740
rect 24780 75682 24836 75694
rect 24780 75630 24782 75682
rect 24834 75630 24836 75682
rect 24220 75572 24276 75582
rect 23996 75570 24276 75572
rect 23996 75518 24222 75570
rect 24274 75518 24276 75570
rect 23996 75516 24276 75518
rect 24220 75506 24276 75516
rect 24780 75348 24836 75630
rect 25228 75684 25284 75694
rect 25228 75590 25284 75628
rect 25900 75684 25956 75694
rect 23884 75292 24836 75348
rect 23548 75124 23604 75134
rect 23324 75122 23604 75124
rect 23324 75070 23550 75122
rect 23602 75070 23604 75122
rect 23324 75068 23604 75070
rect 23548 75058 23604 75068
rect 22764 74898 22820 74910
rect 22764 74846 22766 74898
rect 22818 74846 22820 74898
rect 20412 31892 20804 31948
rect 20860 74004 20916 74014
rect 22764 74004 22820 74846
rect 22988 74004 23044 74014
rect 22764 74002 23044 74004
rect 22764 73950 22990 74002
rect 23042 73950 23044 74002
rect 22764 73948 23044 73950
rect 19836 31388 20100 31398
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 19836 31322 20100 31332
rect 19836 29820 20100 29830
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 19836 29754 20100 29764
rect 19836 28252 20100 28262
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 19836 28186 20100 28196
rect 19836 26684 20100 26694
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 19836 26618 20100 26628
rect 19836 25116 20100 25126
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 19836 25050 20100 25060
rect 20300 24612 20356 24622
rect 20076 24610 20356 24612
rect 20076 24558 20302 24610
rect 20354 24558 20356 24610
rect 20076 24556 20356 24558
rect 19740 24276 19796 24286
rect 19740 24050 19796 24220
rect 19740 23998 19742 24050
rect 19794 23998 19796 24050
rect 19740 23986 19796 23998
rect 20076 24050 20132 24556
rect 20300 24546 20356 24556
rect 20412 24052 20468 31892
rect 20076 23998 20078 24050
rect 20130 23998 20132 24050
rect 20076 23986 20132 23998
rect 20188 23996 20468 24052
rect 20636 24724 20692 24734
rect 19516 23828 19572 23838
rect 19404 23714 19460 23726
rect 19404 23662 19406 23714
rect 19458 23662 19460 23714
rect 19404 23604 19460 23662
rect 19404 23538 19460 23548
rect 19516 23266 19572 23772
rect 19836 23548 20100 23558
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 19836 23482 20100 23492
rect 19516 23214 19518 23266
rect 19570 23214 19572 23266
rect 19404 22484 19460 22494
rect 19404 22390 19460 22428
rect 19516 22260 19572 23214
rect 19628 23266 19684 23278
rect 19628 23214 19630 23266
rect 19682 23214 19684 23266
rect 19628 23044 19684 23214
rect 19628 22978 19684 22988
rect 19852 23154 19908 23166
rect 19852 23102 19854 23154
rect 19906 23102 19908 23154
rect 19852 22372 19908 23102
rect 19852 22306 19908 22316
rect 19964 22370 20020 22382
rect 19964 22318 19966 22370
rect 20018 22318 20020 22370
rect 19740 22260 19796 22270
rect 19516 22258 19796 22260
rect 19516 22206 19742 22258
rect 19794 22206 19796 22258
rect 19516 22204 19796 22206
rect 19740 22194 19796 22204
rect 19852 22148 19908 22158
rect 19964 22148 20020 22318
rect 19908 22092 20020 22148
rect 19852 22082 19908 22092
rect 19836 21980 20100 21990
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 19292 21868 19460 21924
rect 19836 21914 20100 21924
rect 19180 21586 19236 21598
rect 19180 21534 19182 21586
rect 19234 21534 19236 21586
rect 19068 20804 19124 20814
rect 18956 20690 19012 20702
rect 18956 20638 18958 20690
rect 19010 20638 19012 20690
rect 18956 20132 19012 20638
rect 19068 20690 19124 20748
rect 19068 20638 19070 20690
rect 19122 20638 19124 20690
rect 19068 20626 19124 20638
rect 18956 20066 19012 20076
rect 19068 20468 19124 20478
rect 19068 19460 19124 20412
rect 19180 19908 19236 21534
rect 19292 20578 19348 20590
rect 19292 20526 19294 20578
rect 19346 20526 19348 20578
rect 19292 20244 19348 20526
rect 19404 20468 19460 21868
rect 19852 21474 19908 21486
rect 19852 21422 19854 21474
rect 19906 21422 19908 21474
rect 19852 20580 19908 21422
rect 20188 20804 20244 23996
rect 20412 23828 20468 23838
rect 20412 23734 20468 23772
rect 20524 23716 20580 23726
rect 20524 23622 20580 23660
rect 20188 20738 20244 20748
rect 20300 23156 20356 23166
rect 20636 23156 20692 24668
rect 20748 23940 20804 23978
rect 20748 23874 20804 23884
rect 20300 23154 20692 23156
rect 20300 23102 20302 23154
rect 20354 23102 20692 23154
rect 20300 23100 20692 23102
rect 19852 20524 20244 20580
rect 19404 20402 19460 20412
rect 19836 20412 20100 20422
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 19836 20346 20100 20356
rect 19292 20188 19796 20244
rect 19180 19842 19236 19852
rect 19628 19908 19684 19918
rect 19404 19572 19460 19582
rect 19404 19460 19460 19516
rect 19068 19404 19460 19460
rect 18844 19346 19348 19348
rect 18844 19294 18846 19346
rect 18898 19294 19348 19346
rect 18844 19292 19348 19294
rect 18620 18564 18676 18574
rect 18620 18450 18676 18508
rect 18620 18398 18622 18450
rect 18674 18398 18676 18450
rect 18620 18386 18676 18398
rect 18732 17556 18788 17566
rect 18620 13860 18676 13870
rect 18620 13766 18676 13804
rect 18508 12350 18510 12402
rect 18562 12350 18564 12402
rect 18508 11788 18564 12350
rect 18284 11732 18564 11788
rect 18284 11508 18340 11732
rect 17836 10882 17892 10892
rect 17948 11506 18340 11508
rect 17948 11454 18286 11506
rect 18338 11454 18340 11506
rect 17948 11452 18340 11454
rect 17948 10834 18004 11452
rect 18284 11442 18340 11452
rect 18732 10836 18788 17500
rect 17948 10782 17950 10834
rect 18002 10782 18004 10834
rect 17948 10770 18004 10782
rect 18620 10780 18788 10836
rect 17724 10612 17780 10622
rect 17724 10518 17780 10556
rect 17836 10610 17892 10622
rect 17836 10558 17838 10610
rect 17890 10558 17892 10610
rect 17612 9268 17668 9278
rect 17612 9174 17668 9212
rect 17724 9156 17780 9166
rect 17836 9156 17892 10558
rect 17724 9154 17892 9156
rect 17724 9102 17726 9154
rect 17778 9102 17892 9154
rect 17724 9100 17892 9102
rect 18284 10612 18340 10622
rect 17724 9090 17780 9100
rect 18284 9044 18340 10556
rect 18396 10610 18452 10622
rect 18396 10558 18398 10610
rect 18450 10558 18452 10610
rect 18396 9268 18452 10558
rect 18396 9202 18452 9212
rect 18508 9716 18564 9726
rect 18508 9266 18564 9660
rect 18508 9214 18510 9266
rect 18562 9214 18564 9266
rect 18508 9202 18564 9214
rect 18620 9380 18676 10780
rect 18620 9266 18676 9324
rect 18620 9214 18622 9266
rect 18674 9214 18676 9266
rect 18620 9202 18676 9214
rect 18732 10610 18788 10622
rect 18732 10558 18734 10610
rect 18786 10558 18788 10610
rect 18396 9044 18452 9054
rect 18284 9042 18452 9044
rect 18284 8990 18398 9042
rect 18450 8990 18452 9042
rect 18284 8988 18452 8990
rect 17500 8876 17892 8932
rect 17836 8372 17892 8876
rect 17836 8278 17892 8316
rect 18396 8036 18452 8988
rect 18732 9044 18788 10558
rect 18844 9492 18900 19292
rect 19180 19122 19236 19134
rect 19180 19070 19182 19122
rect 19234 19070 19236 19122
rect 19180 18676 19236 19070
rect 19292 19122 19348 19292
rect 19292 19070 19294 19122
rect 19346 19070 19348 19122
rect 19292 19058 19348 19070
rect 19068 17668 19124 17678
rect 19180 17668 19236 18620
rect 19292 18340 19348 18350
rect 19292 18246 19348 18284
rect 19404 17892 19460 19404
rect 19516 19012 19572 19022
rect 19516 18918 19572 18956
rect 19628 18564 19684 19852
rect 19740 19234 19796 20188
rect 20188 19348 20244 20524
rect 20300 19908 20356 23100
rect 20412 22484 20468 22494
rect 20412 22390 20468 22428
rect 20748 22258 20804 22270
rect 20748 22206 20750 22258
rect 20802 22206 20804 22258
rect 20748 21364 20804 22206
rect 20748 21298 20804 21308
rect 20300 19842 20356 19852
rect 20636 20578 20692 20590
rect 20636 20526 20638 20578
rect 20690 20526 20692 20578
rect 20300 19348 20356 19358
rect 20188 19346 20356 19348
rect 20188 19294 20302 19346
rect 20354 19294 20356 19346
rect 20188 19292 20356 19294
rect 20300 19282 20356 19292
rect 19740 19182 19742 19234
rect 19794 19182 19796 19234
rect 19740 19170 19796 19182
rect 20412 19236 20468 19246
rect 20412 19142 20468 19180
rect 20188 19010 20244 19022
rect 20188 18958 20190 19010
rect 20242 18958 20244 19010
rect 19836 18844 20100 18854
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 19836 18778 20100 18788
rect 20188 18676 20244 18958
rect 20188 18610 20244 18620
rect 20524 18900 20580 18910
rect 19404 17836 19572 17892
rect 19068 17666 19236 17668
rect 19068 17614 19070 17666
rect 19122 17614 19236 17666
rect 19068 17612 19236 17614
rect 19404 17668 19460 17678
rect 19068 17602 19124 17612
rect 19404 17574 19460 17612
rect 19292 17556 19348 17566
rect 19180 17500 19292 17556
rect 19180 17442 19236 17500
rect 19292 17490 19348 17500
rect 19180 17390 19182 17442
rect 19234 17390 19236 17442
rect 19180 17378 19236 17390
rect 19516 15148 19572 17836
rect 19180 15092 19572 15148
rect 18956 14308 19012 14318
rect 18956 13746 19012 14252
rect 19180 13970 19236 15092
rect 19180 13918 19182 13970
rect 19234 13918 19236 13970
rect 19180 13860 19236 13918
rect 19236 13804 19460 13860
rect 19180 13794 19236 13804
rect 18956 13694 18958 13746
rect 19010 13694 19012 13746
rect 18956 11172 19012 13694
rect 19068 13636 19124 13646
rect 19068 13542 19124 13580
rect 19404 13076 19460 13804
rect 19516 13748 19572 13758
rect 19628 13748 19684 18508
rect 20188 17668 20244 17678
rect 20188 17574 20244 17612
rect 20524 17666 20580 18844
rect 20636 18676 20692 20526
rect 20636 18610 20692 18620
rect 20748 19236 20804 19246
rect 20636 18340 20692 18350
rect 20636 17778 20692 18284
rect 20636 17726 20638 17778
rect 20690 17726 20692 17778
rect 20636 17714 20692 17726
rect 20524 17614 20526 17666
rect 20578 17614 20580 17666
rect 20524 17602 20580 17614
rect 20748 17666 20804 19180
rect 20748 17614 20750 17666
rect 20802 17614 20804 17666
rect 20748 17602 20804 17614
rect 20860 17556 20916 73948
rect 22988 55468 23044 73948
rect 24780 55468 24836 75292
rect 22428 55412 23044 55468
rect 24444 55412 24836 55468
rect 22428 43708 22484 55412
rect 22428 43652 22708 43708
rect 21420 24612 21476 24622
rect 21420 24610 21812 24612
rect 21420 24558 21422 24610
rect 21474 24558 21812 24610
rect 21420 24556 21812 24558
rect 21420 24546 21476 24556
rect 21756 24050 21812 24556
rect 21756 23998 21758 24050
rect 21810 23998 21812 24050
rect 21756 23986 21812 23998
rect 21196 23940 21252 23950
rect 21196 23846 21252 23884
rect 21644 23716 21700 23726
rect 21644 23622 21700 23660
rect 21868 23714 21924 23726
rect 21868 23662 21870 23714
rect 21922 23662 21924 23714
rect 21084 23044 21140 23054
rect 21084 23042 21812 23044
rect 21084 22990 21086 23042
rect 21138 22990 21812 23042
rect 21084 22988 21812 22990
rect 21084 22978 21140 22988
rect 21756 22482 21812 22988
rect 21756 22430 21758 22482
rect 21810 22430 21812 22482
rect 21756 22418 21812 22430
rect 21196 22372 21252 22382
rect 21196 22278 21252 22316
rect 21644 22146 21700 22158
rect 21644 22094 21646 22146
rect 21698 22094 21700 22146
rect 21644 22036 21700 22094
rect 21644 21970 21700 21980
rect 21868 22146 21924 23662
rect 22316 23716 22372 23726
rect 22316 23622 22372 23660
rect 21868 22094 21870 22146
rect 21922 22094 21924 22146
rect 21868 21700 21924 22094
rect 21868 21634 21924 21644
rect 22092 21924 22148 21934
rect 21980 21476 22036 21486
rect 21756 21474 22036 21476
rect 21756 21422 21982 21474
rect 22034 21422 22036 21474
rect 21756 21420 22036 21422
rect 21756 20914 21812 21420
rect 21980 21410 22036 21420
rect 21756 20862 21758 20914
rect 21810 20862 21812 20914
rect 21756 20850 21812 20862
rect 22092 20804 22148 21868
rect 22316 21700 22372 21710
rect 22316 21606 22372 21644
rect 21868 20802 22148 20804
rect 21868 20750 22094 20802
rect 22146 20750 22148 20802
rect 21868 20748 22148 20750
rect 21644 20578 21700 20590
rect 21644 20526 21646 20578
rect 21698 20526 21700 20578
rect 21420 19124 21476 19134
rect 21420 18338 21476 19068
rect 21420 18286 21422 18338
rect 21474 18286 21476 18338
rect 21420 18274 21476 18286
rect 21532 18900 21588 18910
rect 21420 17780 21476 17790
rect 21532 17780 21588 18844
rect 21644 18676 21700 20526
rect 21756 19460 21812 19470
rect 21756 19346 21812 19404
rect 21756 19294 21758 19346
rect 21810 19294 21812 19346
rect 21756 19282 21812 19294
rect 21644 18610 21700 18620
rect 21420 17778 21588 17780
rect 21420 17726 21422 17778
rect 21474 17726 21588 17778
rect 21420 17724 21588 17726
rect 21868 18450 21924 20748
rect 22092 20738 22148 20748
rect 22540 21586 22596 21598
rect 22540 21534 22542 21586
rect 22594 21534 22596 21586
rect 22540 19348 22596 21534
rect 22652 20132 22708 43652
rect 23996 25394 24052 25406
rect 23996 25342 23998 25394
rect 24050 25342 24052 25394
rect 23660 25284 23716 25294
rect 23660 25190 23716 25228
rect 23548 24612 23604 24622
rect 23884 24612 23940 24622
rect 23548 24610 23940 24612
rect 23548 24558 23550 24610
rect 23602 24558 23886 24610
rect 23938 24558 23940 24610
rect 23548 24556 23940 24558
rect 23548 24546 23604 24556
rect 23884 24546 23940 24556
rect 23324 24500 23380 24510
rect 23324 24052 23380 24444
rect 23996 24164 24052 25342
rect 24108 25284 24164 25294
rect 24108 25190 24164 25228
rect 24332 25282 24388 25294
rect 24332 25230 24334 25282
rect 24386 25230 24388 25282
rect 24332 25060 24388 25230
rect 24332 24994 24388 25004
rect 23660 24108 24052 24164
rect 24220 24610 24276 24622
rect 24220 24558 24222 24610
rect 24274 24558 24276 24610
rect 23324 24050 23604 24052
rect 23324 23998 23326 24050
rect 23378 23998 23604 24050
rect 23324 23996 23604 23998
rect 23324 23986 23380 23996
rect 23548 23716 23604 23996
rect 23660 23938 23716 24108
rect 23660 23886 23662 23938
rect 23714 23886 23716 23938
rect 23660 23874 23716 23886
rect 23772 23716 23828 23726
rect 23548 23714 23828 23716
rect 23548 23662 23774 23714
rect 23826 23662 23828 23714
rect 23548 23660 23828 23662
rect 23772 23650 23828 23660
rect 23884 23268 23940 24108
rect 23996 23940 24052 23950
rect 23996 23846 24052 23884
rect 24220 23716 24276 24558
rect 24220 23650 24276 23660
rect 24332 23938 24388 23950
rect 24332 23886 24334 23938
rect 24386 23886 24388 23938
rect 24220 23380 24276 23390
rect 24108 23378 24276 23380
rect 24108 23326 24222 23378
rect 24274 23326 24276 23378
rect 24108 23324 24276 23326
rect 23772 23266 23940 23268
rect 23772 23214 23886 23266
rect 23938 23214 23940 23266
rect 23772 23212 23940 23214
rect 23212 23042 23268 23054
rect 23212 22990 23214 23042
rect 23266 22990 23268 23042
rect 23100 22484 23156 22494
rect 23212 22484 23268 22990
rect 23100 22482 23268 22484
rect 23100 22430 23102 22482
rect 23154 22430 23268 22482
rect 23100 22428 23268 22430
rect 23100 22418 23156 22428
rect 23548 22370 23604 22382
rect 23548 22318 23550 22370
rect 23602 22318 23604 22370
rect 22988 22146 23044 22158
rect 22988 22094 22990 22146
rect 23042 22094 23044 22146
rect 22988 22036 23044 22094
rect 23548 22148 23604 22318
rect 23772 22258 23828 23212
rect 23884 23202 23940 23212
rect 23996 23266 24052 23278
rect 23996 23214 23998 23266
rect 24050 23214 24052 23266
rect 23996 23156 24052 23214
rect 24108 23268 24164 23324
rect 24220 23314 24276 23324
rect 24108 23202 24164 23212
rect 23996 23090 24052 23100
rect 24220 23156 24276 23166
rect 23772 22206 23774 22258
rect 23826 22206 23828 22258
rect 23604 22092 23716 22148
rect 23548 22082 23604 22092
rect 22988 21970 23044 21980
rect 23548 21476 23604 21486
rect 23548 21382 23604 21420
rect 23660 20804 23716 22092
rect 23772 21700 23828 22206
rect 24220 21810 24276 23100
rect 24332 22370 24388 23886
rect 24332 22318 24334 22370
rect 24386 22318 24388 22370
rect 24332 21924 24388 22318
rect 24332 21858 24388 21868
rect 24220 21758 24222 21810
rect 24274 21758 24276 21810
rect 24220 21746 24276 21758
rect 23884 21700 23940 21710
rect 23772 21698 23940 21700
rect 23772 21646 23886 21698
rect 23938 21646 23940 21698
rect 23772 21644 23940 21646
rect 23884 21634 23940 21644
rect 23996 21698 24052 21710
rect 23996 21646 23998 21698
rect 24050 21646 24052 21698
rect 23996 21476 24052 21646
rect 24444 21700 24500 55412
rect 25900 26908 25956 75628
rect 30156 75684 30212 75694
rect 26908 40404 26964 40414
rect 26908 38948 26964 40348
rect 26908 38882 26964 38892
rect 26908 37380 26964 37390
rect 26908 36372 26964 37324
rect 26908 36306 26964 36316
rect 28476 33124 28532 33134
rect 28476 31668 28532 33068
rect 30156 31948 30212 75628
rect 32956 75682 33012 75740
rect 32956 75630 32958 75682
rect 33010 75630 33012 75682
rect 32956 75618 33012 75630
rect 33516 75684 33572 75694
rect 33516 75590 33572 75628
rect 33628 75460 33684 75740
rect 33964 75684 34020 75694
rect 34076 75684 34132 75852
rect 33964 75682 34132 75684
rect 33964 75630 33966 75682
rect 34018 75630 34132 75682
rect 33964 75628 34132 75630
rect 34412 75682 34468 75694
rect 34412 75630 34414 75682
rect 34466 75630 34468 75682
rect 33964 75618 34020 75628
rect 33516 75404 33684 75460
rect 28476 31602 28532 31612
rect 29932 31892 30212 31948
rect 31052 74788 31108 74798
rect 26908 31108 26964 31118
rect 26908 30100 26964 31052
rect 26908 30034 26964 30044
rect 25900 26852 26740 26908
rect 25228 25060 25284 25070
rect 25284 25004 25396 25060
rect 25228 24994 25284 25004
rect 25340 24946 25396 25004
rect 25340 24894 25342 24946
rect 25394 24894 25396 24946
rect 25340 24882 25396 24894
rect 25564 24724 25620 24734
rect 25564 24630 25620 24668
rect 25788 24722 25844 24734
rect 25788 24670 25790 24722
rect 25842 24670 25844 24722
rect 25004 24612 25060 24622
rect 25004 24050 25060 24556
rect 25676 24612 25732 24622
rect 25676 24518 25732 24556
rect 25004 23998 25006 24050
rect 25058 23998 25060 24050
rect 25004 23986 25060 23998
rect 25788 23380 25844 24670
rect 25788 23378 26068 23380
rect 25788 23326 25790 23378
rect 25842 23326 26068 23378
rect 25788 23324 26068 23326
rect 25788 23314 25844 23324
rect 26012 23268 26068 23324
rect 26068 23212 26292 23268
rect 26012 23202 26068 23212
rect 25116 23156 25172 23166
rect 25116 23062 25172 23100
rect 25564 23156 25620 23166
rect 25564 23062 25620 23100
rect 24556 23044 24612 23054
rect 24556 22950 24612 22988
rect 25676 23042 25732 23054
rect 25676 22990 25678 23042
rect 25730 22990 25732 23042
rect 25676 22708 25732 22990
rect 25116 22652 25732 22708
rect 25116 22482 25172 22652
rect 25116 22430 25118 22482
rect 25170 22430 25172 22482
rect 25116 22418 25172 22430
rect 26236 21810 26292 23212
rect 26236 21758 26238 21810
rect 26290 21758 26292 21810
rect 26236 21746 26292 21758
rect 25676 21700 25732 21710
rect 24444 21634 24500 21644
rect 25564 21644 25676 21700
rect 23996 21410 24052 21420
rect 25004 20916 25060 20926
rect 25004 20914 25284 20916
rect 25004 20862 25006 20914
rect 25058 20862 25284 20914
rect 25004 20860 25284 20862
rect 25004 20850 25060 20860
rect 23660 20738 23716 20748
rect 24780 20804 24836 20814
rect 22652 20066 22708 20076
rect 22876 20690 22932 20702
rect 22876 20638 22878 20690
rect 22930 20638 22932 20690
rect 21980 19236 22036 19246
rect 21980 19122 22036 19180
rect 22316 19236 22372 19246
rect 22540 19236 22596 19292
rect 22764 19348 22820 19358
rect 22876 19348 22932 20638
rect 23212 20132 23268 20142
rect 22764 19346 22932 19348
rect 22764 19294 22766 19346
rect 22818 19294 22932 19346
rect 22764 19292 22932 19294
rect 22988 19460 23044 19470
rect 22764 19282 22820 19292
rect 22316 19234 22596 19236
rect 22316 19182 22318 19234
rect 22370 19182 22596 19234
rect 22316 19180 22596 19182
rect 22652 19236 22708 19246
rect 22316 19170 22372 19180
rect 21980 19070 21982 19122
rect 22034 19070 22036 19122
rect 21980 19058 22036 19070
rect 21868 18398 21870 18450
rect 21922 18398 21924 18450
rect 21420 17714 21476 17724
rect 20860 17490 20916 17500
rect 21868 17556 21924 18398
rect 22540 18338 22596 18350
rect 22540 18286 22542 18338
rect 22594 18286 22596 18338
rect 21980 18228 22036 18238
rect 21980 17666 22036 18172
rect 21980 17614 21982 17666
rect 22034 17614 22036 17666
rect 21980 17602 22036 17614
rect 22316 18228 22372 18238
rect 22316 17666 22372 18172
rect 22428 17780 22484 17790
rect 22540 17780 22596 18286
rect 22428 17778 22596 17780
rect 22428 17726 22430 17778
rect 22482 17726 22596 17778
rect 22428 17724 22596 17726
rect 22428 17714 22484 17724
rect 22316 17614 22318 17666
rect 22370 17614 22372 17666
rect 21868 17490 21924 17500
rect 22316 17332 22372 17614
rect 22540 17556 22596 17566
rect 22652 17556 22708 19180
rect 22876 19124 22932 19134
rect 22988 19124 23044 19404
rect 22876 19122 23044 19124
rect 22876 19070 22878 19122
rect 22930 19070 23044 19122
rect 22876 19068 23044 19070
rect 22876 19058 22932 19068
rect 23100 19012 23156 19022
rect 23100 18918 23156 18956
rect 22540 17554 22708 17556
rect 22540 17502 22542 17554
rect 22594 17502 22708 17554
rect 22540 17500 22708 17502
rect 22540 17490 22596 17500
rect 19836 17276 20100 17286
rect 22316 17276 22820 17332
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 19836 17210 20100 17220
rect 22764 17106 22820 17276
rect 22764 17054 22766 17106
rect 22818 17054 22820 17106
rect 22764 17042 22820 17054
rect 19836 15708 20100 15718
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 19836 15642 20100 15652
rect 23212 15148 23268 20076
rect 24668 20018 24724 20030
rect 24668 19966 24670 20018
rect 24722 19966 24724 20018
rect 24668 19908 24724 19966
rect 24668 19842 24724 19852
rect 24444 19572 24500 19582
rect 24444 19346 24500 19516
rect 24444 19294 24446 19346
rect 24498 19294 24500 19346
rect 23548 19124 23604 19134
rect 23548 19030 23604 19068
rect 23884 19122 23940 19134
rect 23884 19070 23886 19122
rect 23938 19070 23940 19122
rect 23884 18900 23940 19070
rect 24444 19012 24500 19294
rect 24780 19122 24836 20748
rect 24780 19070 24782 19122
rect 24834 19070 24836 19122
rect 24780 19058 24836 19070
rect 24892 20580 24948 20590
rect 24444 18946 24500 18956
rect 23884 18834 23940 18844
rect 24668 18340 24724 18350
rect 24668 18246 24724 18284
rect 22876 15092 23268 15148
rect 21868 14868 21924 14878
rect 19964 14532 20020 14542
rect 19964 14530 20244 14532
rect 19964 14478 19966 14530
rect 20018 14478 20244 14530
rect 19964 14476 20244 14478
rect 19964 14466 20020 14476
rect 19852 14418 19908 14430
rect 19852 14366 19854 14418
rect 19906 14366 19908 14418
rect 19740 14308 19796 14318
rect 19852 14308 19908 14366
rect 19796 14252 19908 14308
rect 20076 14308 20132 14346
rect 19740 14242 19796 14252
rect 20076 14242 20132 14252
rect 19836 14140 20100 14150
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 19836 14074 20100 14084
rect 20188 13972 20244 14476
rect 20076 13916 20244 13972
rect 20300 14306 20356 14318
rect 20300 14254 20302 14306
rect 20354 14254 20356 14306
rect 19852 13748 19908 13758
rect 19628 13746 19908 13748
rect 19628 13694 19854 13746
rect 19906 13694 19908 13746
rect 19628 13692 19908 13694
rect 19516 13654 19572 13692
rect 19852 13682 19908 13692
rect 20076 13186 20132 13916
rect 20076 13134 20078 13186
rect 20130 13134 20132 13186
rect 20076 13122 20132 13134
rect 20300 13748 20356 14254
rect 21420 14308 21476 14318
rect 21420 14214 21476 14252
rect 19516 13076 19572 13086
rect 19404 13074 19572 13076
rect 19404 13022 19518 13074
rect 19570 13022 19572 13074
rect 19404 13020 19572 13022
rect 19516 13010 19572 13020
rect 20300 12964 20356 13692
rect 20636 13636 20692 13646
rect 20412 13634 20692 13636
rect 20412 13582 20638 13634
rect 20690 13582 20692 13634
rect 20412 13580 20692 13582
rect 20412 13186 20468 13580
rect 20636 13570 20692 13580
rect 20412 13134 20414 13186
rect 20466 13134 20468 13186
rect 20412 13122 20468 13134
rect 20300 12908 20468 12964
rect 20300 12740 20356 12750
rect 20188 12738 20356 12740
rect 20188 12686 20302 12738
rect 20354 12686 20356 12738
rect 20188 12684 20356 12686
rect 19836 12572 20100 12582
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 19836 12506 20100 12516
rect 19964 11508 20020 11518
rect 19404 11396 19460 11406
rect 19852 11396 19908 11406
rect 19404 11394 19908 11396
rect 19404 11342 19406 11394
rect 19458 11342 19854 11394
rect 19906 11342 19908 11394
rect 19404 11340 19908 11342
rect 19404 11330 19460 11340
rect 19852 11330 19908 11340
rect 19964 11394 20020 11452
rect 19964 11342 19966 11394
rect 20018 11342 20020 11394
rect 19964 11330 20020 11342
rect 18956 11106 19012 11116
rect 19180 11170 19236 11182
rect 19180 11118 19182 11170
rect 19234 11118 19236 11170
rect 18844 9436 19012 9492
rect 18732 8978 18788 8988
rect 18844 9268 18900 9278
rect 18732 8820 18788 8830
rect 18620 8372 18676 8382
rect 18620 8258 18676 8316
rect 18620 8206 18622 8258
rect 18674 8206 18676 8258
rect 18620 8194 18676 8206
rect 18284 8034 18452 8036
rect 18284 7982 18398 8034
rect 18450 7982 18452 8034
rect 18284 7980 18452 7982
rect 17948 7924 18004 7934
rect 18284 7924 18340 7980
rect 18396 7970 18452 7980
rect 18508 8036 18564 8046
rect 18732 8036 18788 8764
rect 18508 7942 18564 7980
rect 18620 7980 18788 8036
rect 18844 8146 18900 9212
rect 18844 8094 18846 8146
rect 18898 8094 18900 8146
rect 17836 7812 17892 7822
rect 17612 7588 17668 7598
rect 17276 5234 17332 5852
rect 17388 6020 17444 6030
rect 17388 5794 17444 5964
rect 17388 5742 17390 5794
rect 17442 5742 17444 5794
rect 17388 5730 17444 5742
rect 17500 6018 17556 6030
rect 17500 5966 17502 6018
rect 17554 5966 17556 6018
rect 17276 5182 17278 5234
rect 17330 5182 17332 5234
rect 17276 5170 17332 5182
rect 17388 5236 17444 5246
rect 17276 4228 17332 4238
rect 17164 4172 17276 4228
rect 17164 3554 17220 4172
rect 17276 4162 17332 4172
rect 17164 3502 17166 3554
rect 17218 3502 17220 3554
rect 17164 3490 17220 3502
rect 17388 3444 17444 5180
rect 17500 5124 17556 5966
rect 17612 5684 17668 7532
rect 17836 7476 17892 7756
rect 17948 7698 18004 7868
rect 17948 7646 17950 7698
rect 18002 7646 18004 7698
rect 17948 7634 18004 7646
rect 18172 7868 18340 7924
rect 17836 7420 18004 7476
rect 17836 6018 17892 6030
rect 17836 5966 17838 6018
rect 17890 5966 17892 6018
rect 17724 5908 17780 5918
rect 17836 5908 17892 5966
rect 17724 5906 17892 5908
rect 17724 5854 17726 5906
rect 17778 5854 17892 5906
rect 17724 5852 17892 5854
rect 17724 5842 17780 5852
rect 17612 5628 17780 5684
rect 17500 5058 17556 5068
rect 17724 4900 17780 5628
rect 17836 5572 17892 5582
rect 17836 5122 17892 5516
rect 17948 5234 18004 7420
rect 18172 7474 18228 7868
rect 18396 7812 18452 7822
rect 18396 7698 18452 7756
rect 18396 7646 18398 7698
rect 18450 7646 18452 7698
rect 18396 7634 18452 7646
rect 18172 7422 18174 7474
rect 18226 7422 18228 7474
rect 18172 6692 18228 7422
rect 18172 6626 18228 6636
rect 18284 7362 18340 7374
rect 18284 7310 18286 7362
rect 18338 7310 18340 7362
rect 18060 6132 18116 6142
rect 18284 6132 18340 7310
rect 18060 6130 18340 6132
rect 18060 6078 18062 6130
rect 18114 6078 18340 6130
rect 18060 6076 18340 6078
rect 18396 7252 18452 7262
rect 18060 6066 18116 6076
rect 18396 6020 18452 7196
rect 18172 5964 18452 6020
rect 18172 5236 18228 5964
rect 18396 5794 18452 5806
rect 18396 5742 18398 5794
rect 18450 5742 18452 5794
rect 18396 5348 18452 5742
rect 18396 5282 18452 5292
rect 17948 5182 17950 5234
rect 18002 5182 18004 5234
rect 17948 5170 18004 5182
rect 18060 5180 18228 5236
rect 18620 5234 18676 7980
rect 18844 7700 18900 8094
rect 18844 7474 18900 7644
rect 18844 7422 18846 7474
rect 18898 7422 18900 7474
rect 18844 7410 18900 7422
rect 18956 7812 19012 9436
rect 19180 8484 19236 11118
rect 19292 11170 19348 11182
rect 19740 11172 19796 11210
rect 19292 11118 19294 11170
rect 19346 11118 19348 11170
rect 19292 10724 19348 11118
rect 19628 11116 19740 11172
rect 19404 10724 19460 10734
rect 19292 10722 19460 10724
rect 19292 10670 19406 10722
rect 19458 10670 19460 10722
rect 19292 10668 19460 10670
rect 19404 10658 19460 10668
rect 19404 9044 19460 9054
rect 19404 8950 19460 8988
rect 19180 8418 19236 8428
rect 19516 8932 19572 8942
rect 19404 8260 19460 8270
rect 19012 7756 19348 7812
rect 18620 5182 18622 5234
rect 18674 5182 18676 5234
rect 17836 5070 17838 5122
rect 17890 5070 17892 5122
rect 17836 5058 17892 5070
rect 17948 5012 18004 5022
rect 17724 4844 17892 4900
rect 17836 4562 17892 4844
rect 17836 4510 17838 4562
rect 17890 4510 17892 4562
rect 17836 4498 17892 4510
rect 17612 4340 17668 4350
rect 17500 4338 17668 4340
rect 17500 4286 17614 4338
rect 17666 4286 17668 4338
rect 17500 4284 17668 4286
rect 17500 3668 17556 4284
rect 17612 4274 17668 4284
rect 17836 4340 17892 4350
rect 17500 3602 17556 3612
rect 17836 3556 17892 4284
rect 17948 4116 18004 4956
rect 17948 4022 18004 4060
rect 17836 3554 18004 3556
rect 17836 3502 17838 3554
rect 17890 3502 18004 3554
rect 17836 3500 18004 3502
rect 17836 3490 17892 3500
rect 17500 3444 17556 3454
rect 17388 3442 17556 3444
rect 17388 3390 17502 3442
rect 17554 3390 17556 3442
rect 17388 3388 17556 3390
rect 17500 3378 17556 3388
rect 17724 3444 17780 3454
rect 17724 800 17780 3388
rect 17948 3444 18004 3500
rect 18060 3444 18116 5180
rect 18620 5170 18676 5182
rect 18732 6804 18788 6814
rect 18732 5124 18788 6748
rect 18844 6132 18900 6142
rect 18956 6132 19012 7756
rect 19292 6802 19348 7756
rect 19404 7698 19460 8204
rect 19404 7646 19406 7698
rect 19458 7646 19460 7698
rect 19404 7634 19460 7646
rect 19516 7364 19572 8876
rect 19628 8372 19684 11116
rect 19740 11106 19796 11116
rect 19836 11004 20100 11014
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 19836 10938 20100 10948
rect 19836 9436 20100 9446
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 19836 9370 20100 9380
rect 20076 8932 20132 8942
rect 20076 8838 20132 8876
rect 20188 8820 20244 12684
rect 20300 12674 20356 12684
rect 20412 11396 20468 12908
rect 21868 12404 21924 14812
rect 22876 14308 22932 15092
rect 24892 14868 24948 20524
rect 25228 20130 25284 20860
rect 25340 20804 25396 20814
rect 25340 20710 25396 20748
rect 25564 20580 25620 21644
rect 25676 21606 25732 21644
rect 26460 21586 26516 21598
rect 26460 21534 26462 21586
rect 26514 21534 26516 21586
rect 26012 20804 26068 20814
rect 25676 20748 26012 20804
rect 26068 20748 26292 20804
rect 25676 20690 25732 20748
rect 26012 20710 26068 20748
rect 25676 20638 25678 20690
rect 25730 20638 25732 20690
rect 25676 20626 25732 20638
rect 25564 20514 25620 20524
rect 26124 20580 26180 20590
rect 26124 20486 26180 20524
rect 25228 20078 25230 20130
rect 25282 20078 25284 20130
rect 25228 20066 25284 20078
rect 25900 20468 25956 20478
rect 25564 19906 25620 19918
rect 25564 19854 25566 19906
rect 25618 19854 25620 19906
rect 25564 19460 25620 19854
rect 25564 19394 25620 19404
rect 25452 19348 25508 19358
rect 25116 19124 25172 19134
rect 25116 19030 25172 19068
rect 25452 19122 25508 19292
rect 25452 19070 25454 19122
rect 25506 19070 25508 19122
rect 25452 19058 25508 19070
rect 25788 19124 25844 19134
rect 25340 18340 25396 18350
rect 25340 18246 25396 18284
rect 25676 18338 25732 18350
rect 25676 18286 25678 18338
rect 25730 18286 25732 18338
rect 25676 18228 25732 18286
rect 25676 18162 25732 18172
rect 24892 14802 24948 14812
rect 25116 17556 25172 17566
rect 25116 16884 25172 17500
rect 25340 16884 25396 16894
rect 25116 16882 25396 16884
rect 25116 16830 25342 16882
rect 25394 16830 25396 16882
rect 25116 16828 25396 16830
rect 22876 13970 22932 14252
rect 22876 13918 22878 13970
rect 22930 13918 22932 13970
rect 22876 13906 22932 13918
rect 24892 14532 24948 14542
rect 25116 14532 25172 16828
rect 25340 16818 25396 16828
rect 25564 16436 25620 16446
rect 25564 16210 25620 16380
rect 25564 16158 25566 16210
rect 25618 16158 25620 16210
rect 25564 16146 25620 16158
rect 25676 15876 25732 15886
rect 25676 14642 25732 15820
rect 25676 14590 25678 14642
rect 25730 14590 25732 14642
rect 25676 14578 25732 14590
rect 24892 14530 25172 14532
rect 24892 14478 24894 14530
rect 24946 14478 25172 14530
rect 24892 14476 25172 14478
rect 23548 13860 23604 13870
rect 22540 13748 22596 13758
rect 22540 12964 22596 13692
rect 21756 12348 21924 12404
rect 22428 12962 22596 12964
rect 22428 12910 22542 12962
rect 22594 12910 22596 12962
rect 22428 12908 22596 12910
rect 20748 11508 20804 11518
rect 20748 11414 20804 11452
rect 21756 11508 21812 12348
rect 21868 12180 21924 12190
rect 22428 12180 22484 12908
rect 22540 12898 22596 12908
rect 21868 12178 22484 12180
rect 21868 12126 21870 12178
rect 21922 12126 22484 12178
rect 21868 12124 22484 12126
rect 23324 12850 23380 12862
rect 23324 12798 23326 12850
rect 23378 12798 23380 12850
rect 21868 12114 21924 12124
rect 20412 11394 20580 11396
rect 20412 11342 20414 11394
rect 20466 11342 20580 11394
rect 20412 11340 20580 11342
rect 20412 11330 20468 11340
rect 20300 9828 20356 9838
rect 20300 9734 20356 9772
rect 20188 8754 20244 8764
rect 20412 8708 20468 8718
rect 19628 8260 19684 8316
rect 19964 8372 20020 8382
rect 19964 8278 20020 8316
rect 19852 8260 19908 8270
rect 19628 8258 19908 8260
rect 19628 8206 19854 8258
rect 19906 8206 19908 8258
rect 19628 8204 19908 8206
rect 19852 8194 19908 8204
rect 20076 8260 20132 8270
rect 20076 8166 20132 8204
rect 20188 8148 20244 8158
rect 19628 8036 19684 8046
rect 19628 7942 19684 7980
rect 19836 7868 20100 7878
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 19836 7802 20100 7812
rect 19740 7588 19796 7598
rect 19740 7494 19796 7532
rect 19964 7586 20020 7598
rect 19964 7534 19966 7586
rect 20018 7534 20020 7586
rect 19852 7476 19908 7486
rect 19964 7476 20020 7534
rect 20188 7588 20244 8092
rect 20300 7700 20356 7710
rect 20300 7606 20356 7644
rect 20188 7522 20244 7532
rect 20076 7476 20132 7486
rect 19964 7420 20076 7476
rect 19628 7364 19684 7374
rect 19516 7362 19684 7364
rect 19516 7310 19630 7362
rect 19682 7310 19684 7362
rect 19516 7308 19684 7310
rect 19628 7298 19684 7308
rect 19292 6750 19294 6802
rect 19346 6750 19348 6802
rect 19292 6738 19348 6750
rect 19628 6692 19684 6702
rect 19516 6468 19572 6478
rect 18844 6130 19012 6132
rect 18844 6078 18846 6130
rect 18898 6078 19012 6130
rect 18844 6076 19012 6078
rect 19068 6244 19124 6254
rect 18844 6066 18900 6076
rect 18956 5908 19012 5918
rect 18844 5124 18900 5134
rect 18732 5122 18900 5124
rect 18732 5070 18846 5122
rect 18898 5070 18900 5122
rect 18732 5068 18900 5070
rect 18844 5058 18900 5068
rect 18172 5012 18228 5050
rect 18172 4946 18228 4956
rect 18284 5012 18340 5022
rect 18508 5012 18564 5022
rect 18340 5010 18564 5012
rect 18340 4958 18510 5010
rect 18562 4958 18564 5010
rect 18340 4956 18564 4958
rect 18284 4946 18340 4956
rect 18508 4946 18564 4956
rect 18284 4788 18340 4798
rect 18284 4450 18340 4732
rect 18620 4564 18676 4574
rect 18956 4564 19012 5852
rect 19068 4788 19124 6188
rect 19516 6020 19572 6412
rect 19628 6132 19684 6636
rect 19852 6578 19908 7420
rect 20076 7410 20132 7420
rect 19852 6526 19854 6578
rect 19906 6526 19908 6578
rect 19852 6514 19908 6526
rect 20076 6690 20132 6702
rect 20076 6638 20078 6690
rect 20130 6638 20132 6690
rect 20076 6468 20132 6638
rect 20132 6412 20244 6468
rect 20076 6402 20132 6412
rect 19836 6300 20100 6310
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 19836 6234 20100 6244
rect 19852 6132 19908 6142
rect 19628 6130 19908 6132
rect 19628 6078 19854 6130
rect 19906 6078 19908 6130
rect 19628 6076 19908 6078
rect 19852 6066 19908 6076
rect 20188 6130 20244 6412
rect 20188 6078 20190 6130
rect 20242 6078 20244 6130
rect 20188 6066 20244 6078
rect 19516 5964 19684 6020
rect 19292 5796 19348 5806
rect 19068 4722 19124 4732
rect 19180 5794 19348 5796
rect 19180 5742 19294 5794
rect 19346 5742 19348 5794
rect 19180 5740 19348 5742
rect 18620 4562 19012 4564
rect 18620 4510 18622 4562
rect 18674 4510 19012 4562
rect 18620 4508 19012 4510
rect 19068 4564 19124 4574
rect 18620 4498 18676 4508
rect 18284 4398 18286 4450
rect 18338 4398 18340 4450
rect 18284 3668 18340 4398
rect 19068 4338 19124 4508
rect 19068 4286 19070 4338
rect 19122 4286 19124 4338
rect 19068 4274 19124 4286
rect 18284 3602 18340 3612
rect 18620 4116 18676 4126
rect 19180 4116 19236 5740
rect 19292 5730 19348 5740
rect 19516 5796 19572 5806
rect 19404 5684 19460 5694
rect 19292 4564 19348 4574
rect 19404 4564 19460 5628
rect 19516 5122 19572 5740
rect 19516 5070 19518 5122
rect 19570 5070 19572 5122
rect 19516 5058 19572 5070
rect 19292 4562 19460 4564
rect 19292 4510 19294 4562
rect 19346 4510 19460 4562
rect 19292 4508 19460 4510
rect 19292 4498 19348 4508
rect 19628 4450 19684 5964
rect 20412 5908 20468 8652
rect 20524 8258 20580 11340
rect 21644 10836 21700 10846
rect 21756 10836 21812 11452
rect 22540 12066 22596 12078
rect 22540 12014 22542 12066
rect 22594 12014 22596 12066
rect 22540 11506 22596 12014
rect 22540 11454 22542 11506
rect 22594 11454 22596 11506
rect 22540 11442 22596 11454
rect 23212 11508 23268 11518
rect 23324 11508 23380 12798
rect 23212 11506 23380 11508
rect 23212 11454 23214 11506
rect 23266 11454 23380 11506
rect 23212 11452 23380 11454
rect 23436 12068 23492 12078
rect 23212 11442 23268 11452
rect 22316 11396 22372 11406
rect 22988 11396 23044 11406
rect 21644 10834 21812 10836
rect 21644 10782 21646 10834
rect 21698 10782 21812 10834
rect 21644 10780 21812 10782
rect 21868 11394 22372 11396
rect 21868 11342 22318 11394
rect 22370 11342 22372 11394
rect 21868 11340 22372 11342
rect 21644 10770 21700 10780
rect 20860 9828 20916 9838
rect 20860 9734 20916 9772
rect 20524 8206 20526 8258
rect 20578 8206 20580 8258
rect 20524 8148 20580 8206
rect 21420 8932 21476 8942
rect 21308 8148 21364 8158
rect 20524 8146 21364 8148
rect 20524 8094 21310 8146
rect 21362 8094 21364 8146
rect 20524 8092 21364 8094
rect 21308 8082 21364 8092
rect 20972 7924 21028 7934
rect 21420 7924 21476 8876
rect 21868 8484 21924 11340
rect 22316 11330 22372 11340
rect 22764 11394 23044 11396
rect 22764 11342 22990 11394
rect 23042 11342 23044 11394
rect 22764 11340 23044 11342
rect 22652 11284 22708 11294
rect 22652 11190 22708 11228
rect 22764 10836 22820 11340
rect 22988 11330 23044 11340
rect 23324 11284 23380 11294
rect 23436 11284 23492 12012
rect 23324 11282 23492 11284
rect 23324 11230 23326 11282
rect 23378 11230 23492 11282
rect 23324 11228 23492 11230
rect 23324 11218 23380 11228
rect 22204 10780 22820 10836
rect 21756 8428 21924 8484
rect 22092 9044 22148 9054
rect 20860 7868 20972 7924
rect 20636 7812 20692 7822
rect 20636 7698 20692 7756
rect 20636 7646 20638 7698
rect 20690 7646 20692 7698
rect 20636 7634 20692 7646
rect 20748 7588 20804 7598
rect 20748 6802 20804 7532
rect 20748 6750 20750 6802
rect 20802 6750 20804 6802
rect 20748 6738 20804 6750
rect 20188 5852 20468 5908
rect 20636 6580 20692 6590
rect 19964 5460 20020 5470
rect 19964 5234 20020 5404
rect 19964 5182 19966 5234
rect 20018 5182 20020 5234
rect 19964 5170 20020 5182
rect 19836 4732 20100 4742
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 19836 4666 20100 4676
rect 19628 4398 19630 4450
rect 19682 4398 19684 4450
rect 19404 4228 19460 4238
rect 19292 4116 19348 4126
rect 19180 4060 19292 4116
rect 18396 3556 18452 3566
rect 18172 3444 18228 3454
rect 18060 3442 18228 3444
rect 18060 3390 18174 3442
rect 18226 3390 18228 3442
rect 18060 3388 18228 3390
rect 17948 3378 18004 3388
rect 18172 3378 18228 3388
rect 18396 800 18452 3500
rect 18620 3554 18676 4060
rect 19292 4050 19348 4060
rect 18620 3502 18622 3554
rect 18674 3502 18676 3554
rect 18620 3490 18676 3502
rect 19068 3668 19124 3678
rect 18844 3330 18900 3342
rect 18844 3278 18846 3330
rect 18898 3278 18900 3330
rect 18844 1316 18900 3278
rect 18844 1250 18900 1260
rect 19068 800 19124 3612
rect 19292 3668 19348 3678
rect 19292 3554 19348 3612
rect 19292 3502 19294 3554
rect 19346 3502 19348 3554
rect 19292 3490 19348 3502
rect 19404 980 19460 4172
rect 19628 4228 19684 4398
rect 19964 4452 20020 4462
rect 19964 4450 20132 4452
rect 19964 4398 19966 4450
rect 20018 4398 20132 4450
rect 19964 4396 20132 4398
rect 19964 4386 20020 4396
rect 19628 4162 19684 4172
rect 19628 3668 19684 3678
rect 19516 3556 19572 3566
rect 19516 3442 19572 3500
rect 19516 3390 19518 3442
rect 19570 3390 19572 3442
rect 19516 3378 19572 3390
rect 19628 3556 19684 3612
rect 19852 3556 19908 3566
rect 19628 3554 19908 3556
rect 19628 3502 19854 3554
rect 19906 3502 19908 3554
rect 19628 3500 19908 3502
rect 19628 1764 19684 3500
rect 19852 3490 19908 3500
rect 20076 3332 20132 4396
rect 20188 3442 20244 5852
rect 20412 5012 20468 5022
rect 20412 4918 20468 4956
rect 20412 4564 20468 4574
rect 20636 4564 20692 6524
rect 20860 5124 20916 7868
rect 20972 7858 21028 7868
rect 21308 7868 21476 7924
rect 21644 8034 21700 8046
rect 21644 7982 21646 8034
rect 21698 7982 21700 8034
rect 21196 7588 21252 7598
rect 21196 7474 21252 7532
rect 21196 7422 21198 7474
rect 21250 7422 21252 7474
rect 21196 7410 21252 7422
rect 21196 5908 21252 5946
rect 21196 5842 21252 5852
rect 20748 5068 20916 5124
rect 20972 5794 21028 5806
rect 20972 5742 20974 5794
rect 21026 5742 21028 5794
rect 20748 4676 20804 5068
rect 20972 5012 21028 5742
rect 21308 5794 21364 7868
rect 21644 7812 21700 7982
rect 21420 7756 21644 7812
rect 21420 7698 21476 7756
rect 21644 7746 21700 7756
rect 21420 7646 21422 7698
rect 21474 7646 21476 7698
rect 21420 7634 21476 7646
rect 21532 6466 21588 6478
rect 21532 6414 21534 6466
rect 21586 6414 21588 6466
rect 21532 6244 21588 6414
rect 21532 6178 21588 6188
rect 21532 5908 21588 5918
rect 21532 5814 21588 5852
rect 21308 5742 21310 5794
rect 21362 5742 21364 5794
rect 21308 5730 21364 5742
rect 21532 5572 21588 5582
rect 21532 5234 21588 5516
rect 21756 5346 21812 8428
rect 22092 8260 22148 8988
rect 21868 8258 22148 8260
rect 21868 8206 22094 8258
rect 22146 8206 22148 8258
rect 21868 8204 22148 8206
rect 21868 7474 21924 8204
rect 22092 8194 22148 8204
rect 22204 8036 22260 10780
rect 22652 10610 22708 10622
rect 22652 10558 22654 10610
rect 22706 10558 22708 10610
rect 22316 9268 22372 9278
rect 22316 8260 22372 9212
rect 22316 8194 22372 8204
rect 21868 7422 21870 7474
rect 21922 7422 21924 7474
rect 21868 7410 21924 7422
rect 22092 7980 22260 8036
rect 21980 6466 22036 6478
rect 21980 6414 21982 6466
rect 22034 6414 22036 6466
rect 21980 6356 22036 6414
rect 21980 6290 22036 6300
rect 22092 6130 22148 7980
rect 22540 7362 22596 7374
rect 22540 7310 22542 7362
rect 22594 7310 22596 7362
rect 22428 7140 22484 7150
rect 22428 6690 22484 7084
rect 22540 6804 22596 7310
rect 22540 6738 22596 6748
rect 22428 6638 22430 6690
rect 22482 6638 22484 6690
rect 22428 6626 22484 6638
rect 22092 6078 22094 6130
rect 22146 6078 22148 6130
rect 22092 6066 22148 6078
rect 22204 6466 22260 6478
rect 22204 6414 22206 6466
rect 22258 6414 22260 6466
rect 22204 6018 22260 6414
rect 22652 6130 22708 10558
rect 22876 10498 22932 10510
rect 22876 10446 22878 10498
rect 22930 10446 22932 10498
rect 22764 9828 22820 9838
rect 22764 9734 22820 9772
rect 22876 8370 22932 10446
rect 22988 10500 23044 10510
rect 22988 10406 23044 10444
rect 23436 9604 23492 9614
rect 23212 9044 23268 9054
rect 23100 8988 23212 9044
rect 22876 8318 22878 8370
rect 22930 8318 22932 8370
rect 22876 8306 22932 8318
rect 22988 8930 23044 8942
rect 22988 8878 22990 8930
rect 23042 8878 23044 8930
rect 22652 6078 22654 6130
rect 22706 6078 22708 6130
rect 22652 6066 22708 6078
rect 22876 7140 22932 7150
rect 22204 5966 22206 6018
rect 22258 5966 22260 6018
rect 21868 5906 21924 5918
rect 21868 5854 21870 5906
rect 21922 5854 21924 5906
rect 21868 5684 21924 5854
rect 21868 5618 21924 5628
rect 22204 5908 22260 5966
rect 22764 6020 22820 6030
rect 22764 5926 22820 5964
rect 22540 5908 22596 5918
rect 22260 5906 22596 5908
rect 22260 5854 22542 5906
rect 22594 5854 22596 5906
rect 22260 5852 22596 5854
rect 21756 5294 21758 5346
rect 21810 5294 21812 5346
rect 21756 5282 21812 5294
rect 22092 5348 22148 5358
rect 22204 5348 22260 5852
rect 22540 5842 22596 5852
rect 22092 5346 22260 5348
rect 22092 5294 22094 5346
rect 22146 5294 22260 5346
rect 22092 5292 22260 5294
rect 22428 5348 22484 5358
rect 22092 5282 22148 5292
rect 21532 5182 21534 5234
rect 21586 5182 21588 5234
rect 21532 5170 21588 5182
rect 21644 5236 21700 5246
rect 20972 4956 21476 5012
rect 20860 4900 20916 4910
rect 20860 4898 21252 4900
rect 20860 4846 20862 4898
rect 20914 4846 21252 4898
rect 20860 4844 21252 4846
rect 20860 4834 20916 4844
rect 20748 4620 21140 4676
rect 20636 4508 20804 4564
rect 20300 4452 20356 4462
rect 20300 4338 20356 4396
rect 20300 4286 20302 4338
rect 20354 4286 20356 4338
rect 20300 4274 20356 4286
rect 20300 4114 20356 4126
rect 20300 4062 20302 4114
rect 20354 4062 20356 4114
rect 20300 3780 20356 4062
rect 20300 3714 20356 3724
rect 20188 3390 20190 3442
rect 20242 3390 20244 3442
rect 20188 3378 20244 3390
rect 20076 3266 20132 3276
rect 19836 3164 20100 3174
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 19836 3098 20100 3108
rect 19628 1698 19684 1708
rect 19404 924 19796 980
rect 19740 800 19796 924
rect 20412 800 20468 4508
rect 20636 4114 20692 4126
rect 20636 4062 20638 4114
rect 20690 4062 20692 4114
rect 20636 3780 20692 4062
rect 20636 3714 20692 3724
rect 20748 3668 20804 4508
rect 20972 4340 21028 4350
rect 20860 4338 21028 4340
rect 20860 4286 20974 4338
rect 21026 4286 21028 4338
rect 20860 4284 21028 4286
rect 20860 3892 20916 4284
rect 20972 4274 21028 4284
rect 21084 4226 21140 4620
rect 21084 4174 21086 4226
rect 21138 4174 21140 4226
rect 21084 4162 21140 4174
rect 20860 3826 20916 3836
rect 20972 3780 21028 3790
rect 20972 3668 21028 3724
rect 20748 3612 21028 3668
rect 20972 3554 21028 3612
rect 20972 3502 20974 3554
rect 21026 3502 21028 3554
rect 20972 3490 21028 3502
rect 21084 3444 21140 3454
rect 21084 800 21140 3388
rect 21196 3108 21252 4844
rect 21308 4452 21364 4462
rect 21308 4358 21364 4396
rect 21196 3042 21252 3052
rect 21308 3442 21364 3454
rect 21308 3390 21310 3442
rect 21362 3390 21364 3442
rect 21308 1540 21364 3390
rect 21420 3388 21476 4956
rect 21532 4228 21588 4238
rect 21532 3556 21588 4172
rect 21644 4226 21700 5180
rect 22092 5012 22148 5022
rect 21980 4956 22092 5012
rect 21868 4900 21924 4910
rect 21868 4806 21924 4844
rect 21644 4174 21646 4226
rect 21698 4174 21700 4226
rect 21644 4162 21700 4174
rect 21756 4450 21812 4462
rect 21756 4398 21758 4450
rect 21810 4398 21812 4450
rect 21756 4004 21812 4398
rect 21980 4452 22036 4956
rect 22092 4946 22148 4956
rect 22428 4788 22484 5292
rect 22876 5122 22932 7084
rect 22876 5070 22878 5122
rect 22930 5070 22932 5122
rect 22876 5058 22932 5070
rect 22540 5012 22596 5022
rect 22540 4918 22596 4956
rect 21980 4358 22036 4396
rect 22092 4732 22484 4788
rect 22652 4788 22708 4798
rect 21756 3938 21812 3948
rect 21756 3668 21812 3678
rect 21532 3500 21700 3556
rect 21644 3388 21700 3500
rect 21756 3554 21812 3612
rect 21756 3502 21758 3554
rect 21810 3502 21812 3554
rect 21756 3490 21812 3502
rect 21980 3444 22036 3454
rect 22092 3444 22148 4732
rect 22428 4564 22484 4574
rect 22428 4338 22484 4508
rect 22652 4562 22708 4732
rect 22652 4510 22654 4562
rect 22706 4510 22708 4562
rect 22652 4498 22708 4510
rect 22876 4676 22932 4686
rect 22428 4286 22430 4338
rect 22482 4286 22484 4338
rect 22428 4274 22484 4286
rect 22316 4228 22372 4238
rect 22316 3554 22372 4172
rect 22316 3502 22318 3554
rect 22370 3502 22372 3554
rect 22316 3490 22372 3502
rect 22428 4116 22484 4126
rect 21980 3442 22148 3444
rect 21980 3390 21982 3442
rect 22034 3390 22148 3442
rect 21980 3388 22148 3390
rect 21420 3332 21588 3388
rect 21644 3332 21812 3388
rect 21980 3378 22036 3388
rect 21532 2548 21588 3332
rect 21532 2482 21588 2492
rect 21308 1474 21364 1484
rect 21756 800 21812 3332
rect 22428 800 22484 4060
rect 22652 3330 22708 3342
rect 22652 3278 22654 3330
rect 22706 3278 22708 3330
rect 22652 1428 22708 3278
rect 22652 1362 22708 1372
rect 22876 980 22932 4620
rect 22988 4564 23044 8878
rect 23100 5124 23156 8988
rect 23212 8978 23268 8988
rect 23436 7028 23492 9548
rect 23548 9268 23604 13804
rect 24892 13748 24948 14476
rect 24892 13682 24948 13692
rect 24668 13636 24724 13646
rect 24668 12068 24724 13580
rect 25452 13524 25508 13534
rect 25452 13074 25508 13468
rect 25452 13022 25454 13074
rect 25506 13022 25508 13074
rect 25452 12402 25508 13022
rect 25788 12852 25844 19068
rect 25900 13860 25956 20412
rect 26236 20130 26292 20748
rect 26348 20692 26404 20702
rect 26348 20598 26404 20636
rect 26460 20580 26516 21534
rect 26572 20580 26628 20590
rect 26460 20578 26628 20580
rect 26460 20526 26574 20578
rect 26626 20526 26628 20578
rect 26460 20524 26628 20526
rect 26236 20078 26238 20130
rect 26290 20078 26292 20130
rect 26236 19236 26292 20078
rect 26348 20132 26404 20142
rect 26348 20038 26404 20076
rect 26460 19348 26516 20524
rect 26572 20514 26628 20524
rect 26684 20580 26740 26852
rect 27132 25394 27188 25406
rect 27132 25342 27134 25394
rect 27186 25342 27188 25394
rect 27020 25282 27076 25294
rect 27020 25230 27022 25282
rect 27074 25230 27076 25282
rect 27020 24724 27076 25230
rect 27020 24658 27076 24668
rect 27132 24050 27188 25342
rect 27244 24724 27300 24734
rect 28476 24724 28532 24734
rect 27244 24722 27860 24724
rect 27244 24670 27246 24722
rect 27298 24670 27860 24722
rect 27244 24668 27860 24670
rect 27244 24658 27300 24668
rect 27132 23998 27134 24050
rect 27186 23998 27188 24050
rect 27132 23986 27188 23998
rect 27468 23940 27524 23950
rect 27468 23846 27524 23884
rect 27580 23380 27636 23390
rect 27580 23286 27636 23324
rect 26908 23156 26964 23166
rect 26908 23062 26964 23100
rect 27356 23154 27412 23166
rect 27356 23102 27358 23154
rect 27410 23102 27412 23154
rect 27132 22932 27188 22942
rect 27132 22148 27188 22876
rect 27356 22596 27412 23102
rect 27804 23156 27860 24668
rect 27916 24610 27972 24622
rect 27916 24558 27918 24610
rect 27970 24558 27972 24610
rect 27916 24052 27972 24558
rect 28028 24052 28084 24062
rect 27916 24050 28084 24052
rect 27916 23998 28030 24050
rect 28082 23998 28084 24050
rect 27916 23996 28084 23998
rect 28028 23986 28084 23996
rect 27916 23828 27972 23838
rect 27916 23734 27972 23772
rect 28140 23714 28196 23726
rect 28140 23662 28142 23714
rect 28194 23662 28196 23714
rect 28140 23380 28196 23662
rect 28140 23314 28196 23324
rect 28476 23380 28532 24668
rect 28476 23314 28532 23324
rect 29932 23268 29988 31892
rect 30380 24724 30436 24734
rect 30044 24722 30436 24724
rect 30044 24670 30382 24722
rect 30434 24670 30436 24722
rect 30044 24668 30436 24670
rect 30044 24610 30100 24668
rect 30380 24658 30436 24668
rect 30492 24724 30548 24734
rect 30044 24558 30046 24610
rect 30098 24558 30100 24610
rect 30044 24546 30100 24558
rect 30492 23828 30548 24668
rect 30492 23762 30548 23772
rect 29932 23202 29988 23212
rect 27916 23156 27972 23166
rect 27804 23154 27972 23156
rect 27804 23102 27918 23154
rect 27970 23102 27972 23154
rect 27804 23100 27972 23102
rect 27468 23044 27524 23054
rect 27468 22950 27524 22988
rect 27356 22540 27748 22596
rect 27244 22484 27300 22494
rect 27244 22482 27636 22484
rect 27244 22430 27246 22482
rect 27298 22430 27636 22482
rect 27244 22428 27636 22430
rect 27244 22418 27300 22428
rect 27580 22370 27636 22428
rect 27580 22318 27582 22370
rect 27634 22318 27636 22370
rect 27580 22306 27636 22318
rect 27692 22372 27748 22540
rect 27692 22306 27748 22316
rect 27132 22082 27188 22092
rect 27692 22148 27748 22158
rect 27692 22054 27748 22092
rect 27244 20804 27300 20814
rect 27244 20710 27300 20748
rect 26684 20514 26740 20524
rect 26908 20580 26964 20590
rect 27356 20580 27412 20590
rect 26908 20578 27076 20580
rect 26908 20526 26910 20578
rect 26962 20526 27076 20578
rect 26908 20524 27076 20526
rect 26908 20514 26964 20524
rect 26908 20132 26964 20142
rect 26908 20038 26964 20076
rect 26460 19282 26516 19292
rect 26572 20018 26628 20030
rect 26572 19966 26574 20018
rect 26626 19966 26628 20018
rect 26348 19236 26404 19246
rect 26236 19234 26404 19236
rect 26236 19182 26350 19234
rect 26402 19182 26404 19234
rect 26236 19180 26404 19182
rect 26348 19170 26404 19180
rect 26460 19012 26516 19022
rect 26460 18918 26516 18956
rect 26460 18452 26516 18462
rect 26460 18358 26516 18396
rect 26572 18116 26628 19966
rect 27020 20020 27076 20524
rect 27356 20486 27412 20524
rect 27580 20578 27636 20590
rect 27580 20526 27582 20578
rect 27634 20526 27636 20578
rect 27580 20132 27636 20526
rect 27580 20066 27636 20076
rect 27132 20020 27188 20030
rect 27020 19964 27132 20020
rect 27132 19954 27188 19964
rect 27692 20020 27748 20030
rect 27468 19908 27524 19918
rect 26684 19236 26740 19246
rect 27020 19236 27076 19246
rect 26684 19234 27076 19236
rect 26684 19182 26686 19234
rect 26738 19182 27022 19234
rect 27074 19182 27076 19234
rect 26684 19180 27076 19182
rect 26684 19170 26740 19180
rect 27020 19170 27076 19180
rect 27468 19236 27524 19852
rect 27468 19170 27524 19180
rect 27692 19234 27748 19964
rect 27692 19182 27694 19234
rect 27746 19182 27748 19234
rect 27692 19170 27748 19182
rect 27804 20018 27860 23100
rect 27916 23090 27972 23100
rect 28700 23044 28756 23054
rect 28700 22950 28756 22988
rect 30828 23042 30884 23054
rect 30828 22990 30830 23042
rect 30882 22990 30884 23042
rect 30156 22596 30212 22606
rect 28252 22148 28308 22158
rect 27916 20580 27972 20590
rect 27916 20486 27972 20524
rect 27804 19966 27806 20018
rect 27858 19966 27860 20018
rect 27804 19124 27860 19966
rect 28252 19572 28308 22092
rect 30156 20916 30212 22540
rect 30828 22370 30884 22990
rect 30828 22318 30830 22370
rect 30882 22318 30884 22370
rect 30828 22306 30884 22318
rect 30940 22372 30996 22382
rect 30940 22278 30996 22316
rect 29484 20914 30212 20916
rect 29484 20862 30158 20914
rect 30210 20862 30212 20914
rect 29484 20860 30212 20862
rect 29036 20802 29092 20814
rect 29036 20750 29038 20802
rect 29090 20750 29092 20802
rect 29036 20692 29092 20750
rect 29484 20802 29540 20860
rect 30156 20850 30212 20860
rect 29484 20750 29486 20802
rect 29538 20750 29540 20802
rect 29484 20738 29540 20750
rect 30828 20802 30884 20814
rect 30828 20750 30830 20802
rect 30882 20750 30884 20802
rect 29036 20626 29092 20636
rect 30380 20692 30436 20702
rect 30380 20690 30660 20692
rect 30380 20638 30382 20690
rect 30434 20638 30660 20690
rect 30380 20636 30660 20638
rect 30380 20626 30436 20636
rect 28476 20580 28532 20590
rect 28476 20130 28532 20524
rect 29596 20580 29652 20590
rect 29596 20486 29652 20524
rect 29708 20578 29764 20590
rect 29708 20526 29710 20578
rect 29762 20526 29764 20578
rect 28476 20078 28478 20130
rect 28530 20078 28532 20130
rect 28476 20066 28532 20078
rect 29708 20020 29764 20526
rect 29708 19954 29764 19964
rect 30604 19906 30660 20636
rect 30604 19854 30606 19906
rect 30658 19854 30660 19906
rect 30604 19842 30660 19854
rect 28252 19506 28308 19516
rect 27468 19012 27524 19022
rect 27468 18918 27524 18956
rect 27580 19010 27636 19022
rect 27580 18958 27582 19010
rect 27634 18958 27636 19010
rect 27580 18676 27636 18958
rect 27132 18620 27636 18676
rect 27804 18676 27860 19068
rect 28476 19236 28532 19246
rect 28140 19012 28196 19022
rect 28476 19012 28532 19180
rect 28700 19124 28756 19134
rect 28588 19012 28644 19022
rect 28476 19010 28644 19012
rect 28476 18958 28590 19010
rect 28642 18958 28644 19010
rect 28476 18956 28644 18958
rect 28140 18918 28196 18956
rect 27132 18562 27188 18620
rect 27804 18610 27860 18620
rect 27132 18510 27134 18562
rect 27186 18510 27188 18562
rect 27132 18498 27188 18510
rect 26572 18050 26628 18060
rect 27132 18340 27188 18350
rect 26124 16772 26180 16782
rect 26124 16770 26740 16772
rect 26124 16718 26126 16770
rect 26178 16718 26740 16770
rect 26124 16716 26740 16718
rect 26124 16706 26180 16716
rect 26572 16436 26628 16446
rect 26572 16098 26628 16380
rect 26684 16210 26740 16716
rect 26684 16158 26686 16210
rect 26738 16158 26740 16210
rect 26684 16146 26740 16158
rect 26572 16046 26574 16098
rect 26626 16046 26628 16098
rect 26572 16034 26628 16046
rect 27132 15988 27188 18284
rect 28476 17892 28532 17902
rect 28140 17780 28196 17790
rect 28140 17668 28196 17724
rect 27916 17666 28196 17668
rect 27916 17614 28142 17666
rect 28194 17614 28196 17666
rect 27916 17612 28196 17614
rect 27804 16436 27860 16446
rect 27132 15922 27188 15932
rect 27356 16044 27636 16100
rect 26012 15874 26068 15886
rect 26012 15822 26014 15874
rect 26066 15822 26068 15874
rect 26012 15540 26068 15822
rect 26012 15474 26068 15484
rect 26348 15874 26404 15886
rect 26348 15822 26350 15874
rect 26402 15822 26404 15874
rect 26348 15148 26404 15822
rect 26796 15874 26852 15886
rect 26796 15822 26798 15874
rect 26850 15822 26852 15874
rect 26796 15764 26852 15822
rect 26796 15698 26852 15708
rect 27244 15874 27300 15886
rect 27244 15822 27246 15874
rect 27298 15822 27300 15874
rect 26236 15092 26404 15148
rect 26236 13970 26292 15092
rect 26236 13918 26238 13970
rect 26290 13918 26292 13970
rect 26236 13906 26292 13918
rect 27244 13970 27300 15822
rect 27356 15876 27412 16044
rect 27356 15810 27412 15820
rect 27468 15874 27524 15886
rect 27468 15822 27470 15874
rect 27522 15822 27524 15874
rect 27468 15540 27524 15822
rect 27580 15874 27636 16044
rect 27580 15822 27582 15874
rect 27634 15822 27636 15874
rect 27580 15810 27636 15822
rect 27692 15874 27748 15886
rect 27692 15822 27694 15874
rect 27746 15822 27748 15874
rect 27692 15652 27748 15822
rect 27692 15586 27748 15596
rect 27468 15474 27524 15484
rect 27804 15316 27860 16380
rect 27804 15250 27860 15260
rect 27916 15426 27972 17612
rect 28140 17602 28196 17612
rect 28140 16884 28196 16894
rect 28140 16210 28196 16828
rect 28252 16772 28308 16782
rect 28252 16770 28420 16772
rect 28252 16718 28254 16770
rect 28306 16718 28420 16770
rect 28252 16716 28420 16718
rect 28252 16706 28308 16716
rect 28140 16158 28142 16210
rect 28194 16158 28196 16210
rect 28140 16146 28196 16158
rect 28252 16548 28308 16558
rect 28252 16098 28308 16492
rect 28252 16046 28254 16098
rect 28306 16046 28308 16098
rect 28252 16034 28308 16046
rect 28028 15874 28084 15886
rect 28028 15822 28030 15874
rect 28082 15822 28084 15874
rect 28028 15652 28084 15822
rect 28028 15586 28084 15596
rect 27916 15374 27918 15426
rect 27970 15374 27972 15426
rect 27244 13918 27246 13970
rect 27298 13918 27300 13970
rect 27244 13906 27300 13918
rect 27804 14642 27860 14654
rect 27804 14590 27806 14642
rect 27858 14590 27860 14642
rect 26460 13860 26516 13870
rect 25900 13794 25956 13804
rect 26348 13858 26516 13860
rect 26348 13806 26462 13858
rect 26514 13806 26516 13858
rect 26348 13804 26516 13806
rect 25788 12786 25844 12796
rect 26348 12516 26404 13804
rect 26460 13794 26516 13804
rect 26572 13860 26628 13870
rect 27020 13860 27076 13870
rect 26572 13858 26964 13860
rect 26572 13806 26574 13858
rect 26626 13806 26964 13858
rect 26572 13804 26964 13806
rect 26572 13794 26628 13804
rect 26908 13746 26964 13804
rect 27020 13766 27076 13804
rect 26908 13694 26910 13746
rect 26962 13694 26964 13746
rect 26908 13636 26964 13694
rect 27132 13748 27188 13758
rect 27132 13636 27188 13692
rect 27804 13746 27860 14590
rect 27804 13694 27806 13746
rect 27858 13694 27860 13746
rect 27804 13682 27860 13694
rect 26908 13580 27188 13636
rect 27692 13636 27748 13646
rect 25452 12350 25454 12402
rect 25506 12350 25508 12402
rect 25452 12338 25508 12350
rect 25564 12460 26404 12516
rect 25228 12178 25284 12190
rect 25228 12126 25230 12178
rect 25282 12126 25284 12178
rect 24668 12066 25060 12068
rect 24668 12014 24670 12066
rect 24722 12014 25060 12066
rect 24668 12012 25060 12014
rect 24668 12002 24724 12012
rect 25004 11394 25060 12012
rect 25004 11342 25006 11394
rect 25058 11342 25060 11394
rect 25004 11330 25060 11342
rect 24892 11284 24948 11294
rect 24892 11190 24948 11228
rect 24780 11170 24836 11182
rect 24780 11118 24782 11170
rect 24834 11118 24836 11170
rect 24780 11060 24836 11118
rect 25228 11060 25284 12126
rect 25340 12068 25396 12078
rect 25340 11974 25396 12012
rect 25564 11788 25620 12460
rect 25340 11732 25620 11788
rect 25676 12290 25732 12302
rect 26460 12292 26516 12302
rect 25676 12238 25678 12290
rect 25730 12238 25732 12290
rect 25340 11172 25396 11732
rect 25452 11396 25508 11406
rect 25676 11396 25732 12238
rect 26124 12290 26516 12292
rect 26124 12238 26462 12290
rect 26514 12238 26516 12290
rect 26124 12236 26516 12238
rect 25452 11394 25732 11396
rect 25452 11342 25454 11394
rect 25506 11342 25732 11394
rect 25452 11340 25732 11342
rect 25788 11396 25844 11406
rect 25788 11394 25956 11396
rect 25788 11342 25790 11394
rect 25842 11342 25956 11394
rect 25788 11340 25956 11342
rect 25452 11330 25508 11340
rect 25340 11116 25508 11172
rect 24780 11004 25284 11060
rect 25228 10948 25284 11004
rect 25228 10834 25284 10892
rect 25228 10782 25230 10834
rect 25282 10782 25284 10834
rect 25228 10770 25284 10782
rect 25452 10610 25508 11116
rect 25452 10558 25454 10610
rect 25506 10558 25508 10610
rect 25340 10500 25396 10510
rect 25340 10406 25396 10444
rect 25452 10276 25508 10558
rect 25116 10220 25508 10276
rect 25564 10724 25620 11340
rect 25788 11330 25844 11340
rect 25676 10724 25732 10734
rect 25564 10722 25844 10724
rect 25564 10670 25678 10722
rect 25730 10670 25844 10722
rect 25564 10668 25844 10670
rect 24668 9940 24724 9950
rect 23548 9202 23604 9212
rect 23660 9714 23716 9726
rect 23660 9662 23662 9714
rect 23714 9662 23716 9714
rect 23660 9044 23716 9662
rect 24668 9268 24724 9884
rect 24668 9174 24724 9212
rect 23660 8978 23716 8988
rect 23548 8930 23604 8942
rect 23548 8878 23550 8930
rect 23602 8878 23604 8930
rect 23548 7140 23604 8878
rect 24332 8932 24388 8942
rect 24332 8930 24612 8932
rect 24332 8878 24334 8930
rect 24386 8878 24612 8930
rect 24332 8876 24612 8878
rect 24332 8866 24388 8876
rect 23548 7084 24388 7140
rect 23436 6962 23492 6972
rect 24108 6916 24164 6926
rect 23884 6804 23940 6814
rect 23212 6802 23940 6804
rect 23212 6750 23886 6802
rect 23938 6750 23940 6802
rect 23212 6748 23940 6750
rect 23212 6578 23268 6748
rect 23884 6738 23940 6748
rect 23212 6526 23214 6578
rect 23266 6526 23268 6578
rect 23212 6514 23268 6526
rect 23324 6580 23380 6590
rect 23324 6486 23380 6524
rect 23436 6580 23492 6590
rect 23660 6580 23716 6590
rect 23436 6578 23660 6580
rect 23436 6526 23438 6578
rect 23490 6526 23660 6578
rect 23436 6524 23660 6526
rect 23436 6514 23492 6524
rect 23660 6514 23716 6524
rect 23772 6578 23828 6590
rect 23772 6526 23774 6578
rect 23826 6526 23828 6578
rect 23548 6356 23604 6366
rect 23772 6356 23828 6526
rect 23996 6468 24052 6478
rect 23548 6130 23604 6300
rect 23548 6078 23550 6130
rect 23602 6078 23604 6130
rect 23548 6066 23604 6078
rect 23660 6300 23828 6356
rect 23884 6466 24052 6468
rect 23884 6414 23998 6466
rect 24050 6414 24052 6466
rect 23884 6412 24052 6414
rect 23436 5684 23492 5694
rect 23660 5684 23716 6300
rect 23884 6244 23940 6412
rect 23996 6402 24052 6412
rect 23212 5124 23268 5134
rect 23100 5122 23268 5124
rect 23100 5070 23214 5122
rect 23266 5070 23268 5122
rect 23100 5068 23268 5070
rect 23212 5058 23268 5068
rect 23324 5124 23380 5134
rect 23212 4900 23268 4910
rect 22988 4498 23044 4508
rect 23100 4844 23212 4900
rect 22988 4340 23044 4350
rect 22988 4246 23044 4284
rect 23100 3666 23156 4844
rect 23212 4834 23268 4844
rect 23324 4450 23380 5068
rect 23324 4398 23326 4450
rect 23378 4398 23380 4450
rect 23324 4386 23380 4398
rect 23212 4228 23268 4238
rect 23212 4134 23268 4172
rect 23324 3780 23380 3790
rect 23436 3780 23492 5628
rect 23548 5628 23716 5684
rect 23772 6188 23940 6244
rect 23548 5012 23604 5628
rect 23548 4946 23604 4956
rect 23660 5460 23716 5470
rect 23660 4452 23716 5404
rect 23324 3778 23492 3780
rect 23324 3726 23326 3778
rect 23378 3726 23492 3778
rect 23324 3724 23492 3726
rect 23548 4450 23716 4452
rect 23548 4398 23662 4450
rect 23714 4398 23716 4450
rect 23548 4396 23716 4398
rect 23324 3714 23380 3724
rect 23100 3614 23102 3666
rect 23154 3614 23156 3666
rect 23100 3602 23156 3614
rect 22988 3556 23044 3566
rect 22988 3462 23044 3500
rect 23548 3444 23604 4396
rect 23660 4386 23716 4396
rect 23548 3378 23604 3388
rect 23660 3554 23716 3566
rect 23660 3502 23662 3554
rect 23714 3502 23716 3554
rect 23660 3332 23716 3502
rect 23772 3388 23828 6188
rect 23884 6018 23940 6030
rect 23884 5966 23886 6018
rect 23938 5966 23940 6018
rect 23884 5236 23940 5966
rect 24108 6018 24164 6860
rect 24108 5966 24110 6018
rect 24162 5966 24164 6018
rect 24108 5954 24164 5966
rect 23884 5170 23940 5180
rect 23996 5794 24052 5806
rect 23996 5742 23998 5794
rect 24050 5742 24052 5794
rect 23996 5234 24052 5742
rect 23996 5182 23998 5234
rect 24050 5182 24052 5234
rect 23996 5170 24052 5182
rect 24220 5796 24276 5806
rect 23996 4452 24052 4462
rect 23996 4450 24164 4452
rect 23996 4398 23998 4450
rect 24050 4398 24164 4450
rect 23996 4396 24164 4398
rect 23996 4386 24052 4396
rect 23996 3892 24052 3902
rect 23996 3442 24052 3836
rect 23996 3390 23998 3442
rect 24050 3390 24052 3442
rect 23772 3332 23940 3388
rect 23996 3378 24052 3390
rect 23660 3266 23716 3276
rect 23884 2324 23940 3332
rect 23884 2258 23940 2268
rect 24108 2212 24164 4396
rect 24220 3332 24276 5740
rect 24332 4450 24388 7084
rect 24556 5348 24612 8876
rect 25004 8372 25060 8382
rect 25116 8372 25172 10220
rect 25228 9268 25284 9278
rect 25228 9174 25284 9212
rect 25564 9266 25620 10668
rect 25676 10658 25732 10668
rect 25788 10498 25844 10668
rect 25788 10446 25790 10498
rect 25842 10446 25844 10498
rect 25788 10434 25844 10446
rect 25564 9214 25566 9266
rect 25618 9214 25620 9266
rect 25564 9202 25620 9214
rect 25788 10276 25844 10286
rect 25340 9044 25396 9054
rect 25340 8372 25396 8988
rect 25004 8370 25172 8372
rect 25004 8318 25006 8370
rect 25058 8318 25172 8370
rect 25004 8316 25172 8318
rect 25228 8316 25396 8372
rect 25004 8306 25060 8316
rect 24668 8148 24724 8158
rect 24668 7362 24724 8092
rect 24668 7310 24670 7362
rect 24722 7310 24724 7362
rect 24668 7298 24724 7310
rect 24780 7028 24836 7038
rect 24668 6468 24724 6478
rect 24668 6374 24724 6412
rect 24780 6130 24836 6972
rect 25116 6468 25172 6478
rect 24780 6078 24782 6130
rect 24834 6078 24836 6130
rect 24780 6066 24836 6078
rect 25004 6466 25172 6468
rect 25004 6414 25118 6466
rect 25170 6414 25172 6466
rect 25004 6412 25172 6414
rect 24556 5292 24836 5348
rect 24332 4398 24334 4450
rect 24386 4398 24388 4450
rect 24332 4116 24388 4398
rect 24332 4050 24388 4060
rect 24444 4564 24500 4574
rect 24220 2772 24276 3276
rect 24220 2706 24276 2716
rect 24108 2146 24164 2156
rect 23772 1764 23828 1774
rect 22876 924 23156 980
rect 23100 800 23156 924
rect 23772 800 23828 1708
rect 24444 800 24500 4508
rect 24668 4452 24724 4462
rect 24668 4358 24724 4396
rect 24556 3780 24612 3790
rect 24556 3556 24612 3724
rect 24556 3490 24612 3500
rect 24780 3780 24836 5292
rect 24780 3554 24836 3724
rect 24780 3502 24782 3554
rect 24834 3502 24836 3554
rect 24780 3490 24836 3502
rect 25004 3332 25060 6412
rect 25116 6402 25172 6412
rect 25228 4338 25284 8316
rect 25564 8260 25620 8270
rect 25564 8166 25620 8204
rect 25788 8258 25844 10220
rect 25900 9044 25956 11340
rect 26012 10610 26068 10622
rect 26012 10558 26014 10610
rect 26066 10558 26068 10610
rect 26012 10498 26068 10558
rect 26124 10612 26180 12236
rect 26460 12226 26516 12236
rect 26460 12066 26516 12078
rect 26460 12014 26462 12066
rect 26514 12014 26516 12066
rect 26236 11956 26292 11966
rect 26236 11954 26404 11956
rect 26236 11902 26238 11954
rect 26290 11902 26404 11954
rect 26236 11900 26404 11902
rect 26236 11890 26292 11900
rect 26236 11620 26292 11630
rect 26236 10836 26292 11564
rect 26348 11172 26404 11900
rect 26460 11506 26516 12014
rect 26460 11454 26462 11506
rect 26514 11454 26516 11506
rect 26460 11442 26516 11454
rect 27132 11172 27188 11182
rect 26348 11116 26628 11172
rect 26460 10836 26516 10846
rect 26236 10834 26516 10836
rect 26236 10782 26462 10834
rect 26514 10782 26516 10834
rect 26236 10780 26516 10782
rect 26460 10770 26516 10780
rect 26572 10834 26628 11116
rect 26572 10782 26574 10834
rect 26626 10782 26628 10834
rect 26572 10770 26628 10782
rect 26684 10948 26740 10958
rect 26124 10556 26404 10612
rect 26012 10446 26014 10498
rect 26066 10446 26068 10498
rect 26012 10434 26068 10446
rect 26236 10388 26292 10398
rect 25900 8950 25956 8988
rect 26124 10332 26236 10388
rect 25788 8206 25790 8258
rect 25842 8206 25844 8258
rect 25788 8148 25844 8206
rect 25788 8082 25844 8092
rect 25900 8484 25956 8494
rect 25676 8034 25732 8046
rect 25676 7982 25678 8034
rect 25730 7982 25732 8034
rect 25340 7812 25396 7822
rect 25340 7698 25396 7756
rect 25340 7646 25342 7698
rect 25394 7646 25396 7698
rect 25340 7634 25396 7646
rect 25564 7364 25620 7374
rect 25452 7252 25508 7262
rect 25340 6578 25396 6590
rect 25340 6526 25342 6578
rect 25394 6526 25396 6578
rect 25340 6468 25396 6526
rect 25340 5460 25396 6412
rect 25452 6356 25508 7196
rect 25564 6580 25620 7308
rect 25676 6804 25732 7982
rect 25788 7476 25844 7486
rect 25788 7362 25844 7420
rect 25788 7310 25790 7362
rect 25842 7310 25844 7362
rect 25788 7028 25844 7310
rect 25788 6962 25844 6972
rect 25676 6738 25732 6748
rect 25676 6580 25732 6590
rect 25564 6578 25732 6580
rect 25564 6526 25678 6578
rect 25730 6526 25732 6578
rect 25564 6524 25732 6526
rect 25676 6514 25732 6524
rect 25452 6300 25732 6356
rect 25676 5906 25732 6300
rect 25676 5854 25678 5906
rect 25730 5854 25732 5906
rect 25676 5842 25732 5854
rect 25788 6132 25844 6142
rect 25452 5796 25508 5806
rect 25452 5702 25508 5740
rect 25452 5460 25508 5470
rect 25340 5404 25452 5460
rect 25452 5394 25508 5404
rect 25788 4564 25844 6076
rect 25900 6130 25956 8428
rect 26012 8260 26068 8270
rect 26012 6804 26068 8204
rect 26124 7364 26180 10332
rect 26236 10322 26292 10332
rect 26348 8932 26404 10556
rect 26684 10610 26740 10892
rect 26684 10558 26686 10610
rect 26738 10558 26740 10610
rect 26684 9716 26740 10558
rect 26908 9716 26964 9726
rect 26684 9714 26964 9716
rect 26684 9662 26910 9714
rect 26962 9662 26964 9714
rect 26684 9660 26964 9662
rect 26908 9650 26964 9660
rect 26796 9044 26852 9054
rect 26348 8866 26404 8876
rect 26684 8932 26740 8942
rect 26684 8838 26740 8876
rect 26572 8820 26628 8830
rect 26460 8764 26572 8820
rect 26236 8258 26292 8270
rect 26236 8206 26238 8258
rect 26290 8206 26292 8258
rect 26236 8148 26292 8206
rect 26236 8082 26292 8092
rect 26460 7812 26516 8764
rect 26572 8754 26628 8764
rect 26796 8258 26852 8988
rect 26908 8372 26964 8382
rect 26908 8278 26964 8316
rect 26796 8206 26798 8258
rect 26850 8206 26852 8258
rect 26796 8194 26852 8206
rect 27020 8260 27076 8270
rect 26572 8148 26628 8158
rect 26628 8092 26740 8148
rect 26572 8054 26628 8092
rect 26348 7700 26404 7710
rect 26460 7700 26516 7756
rect 26572 7700 26628 7710
rect 26460 7698 26628 7700
rect 26460 7646 26574 7698
rect 26626 7646 26628 7698
rect 26460 7644 26628 7646
rect 26348 7606 26404 7644
rect 26572 7634 26628 7644
rect 26684 7588 26740 8092
rect 27020 8034 27076 8204
rect 27020 7982 27022 8034
rect 27074 7982 27076 8034
rect 26908 7588 26964 7598
rect 26684 7586 26964 7588
rect 26684 7534 26910 7586
rect 26962 7534 26964 7586
rect 26684 7532 26964 7534
rect 26124 7308 26292 7364
rect 26012 6690 26068 6748
rect 26124 6916 26180 6926
rect 26124 6802 26180 6860
rect 26124 6750 26126 6802
rect 26178 6750 26180 6802
rect 26124 6738 26180 6750
rect 26012 6638 26014 6690
rect 26066 6638 26068 6690
rect 26012 6626 26068 6638
rect 26236 6690 26292 7308
rect 26236 6638 26238 6690
rect 26290 6638 26292 6690
rect 25900 6078 25902 6130
rect 25954 6078 25956 6130
rect 25900 6066 25956 6078
rect 26012 5684 26068 5694
rect 26012 5236 26068 5628
rect 26012 5170 26068 5180
rect 26124 5236 26180 5246
rect 26236 5236 26292 6638
rect 26348 6804 26404 6814
rect 26348 6130 26404 6748
rect 26684 6692 26740 6702
rect 26908 6692 26964 7532
rect 26684 6690 26964 6692
rect 26684 6638 26686 6690
rect 26738 6638 26964 6690
rect 26684 6636 26964 6638
rect 26684 6626 26740 6636
rect 26348 6078 26350 6130
rect 26402 6078 26404 6130
rect 26348 6066 26404 6078
rect 26796 6130 26852 6636
rect 26908 6468 26964 6478
rect 27020 6468 27076 7982
rect 26908 6466 27076 6468
rect 26908 6414 26910 6466
rect 26962 6414 27076 6466
rect 26908 6412 27076 6414
rect 26908 6402 26964 6412
rect 26796 6078 26798 6130
rect 26850 6078 26852 6130
rect 26796 6066 26852 6078
rect 26572 5908 26628 5918
rect 26572 5814 26628 5852
rect 26460 5794 26516 5806
rect 26460 5742 26462 5794
rect 26514 5742 26516 5794
rect 26124 5234 26292 5236
rect 26124 5182 26126 5234
rect 26178 5182 26292 5234
rect 26124 5180 26292 5182
rect 26348 5460 26404 5470
rect 26124 5170 26180 5180
rect 25788 4508 26180 4564
rect 25228 4286 25230 4338
rect 25282 4286 25284 4338
rect 25228 4274 25284 4286
rect 26012 4228 26068 4238
rect 26012 4134 26068 4172
rect 26124 3780 26180 4508
rect 26236 3780 26292 3790
rect 26124 3724 26236 3780
rect 25788 3668 25844 3678
rect 25004 3266 25060 3276
rect 25116 3556 25172 3566
rect 25116 800 25172 3500
rect 25340 3554 25396 3566
rect 25340 3502 25342 3554
rect 25394 3502 25396 3554
rect 25340 2100 25396 3502
rect 25340 2034 25396 2044
rect 25788 800 25844 3612
rect 26124 3554 26180 3724
rect 26236 3714 26292 3724
rect 26124 3502 26126 3554
rect 26178 3502 26180 3554
rect 26124 3490 26180 3502
rect 25900 3330 25956 3342
rect 25900 3278 25902 3330
rect 25954 3278 25956 3330
rect 25900 1652 25956 3278
rect 26348 1764 26404 5404
rect 26460 5124 26516 5742
rect 26684 5460 26740 5470
rect 26684 5234 26740 5404
rect 26684 5182 26686 5234
rect 26738 5182 26740 5234
rect 26684 5170 26740 5182
rect 27132 5234 27188 11116
rect 27692 9716 27748 13580
rect 27916 10836 27972 15374
rect 28140 15540 28196 15550
rect 28140 15148 28196 15484
rect 28364 15148 28420 16716
rect 28476 16100 28532 17836
rect 28588 17780 28644 18956
rect 28588 17686 28644 17724
rect 28700 16884 28756 19068
rect 29148 19122 29204 19134
rect 29148 19070 29150 19122
rect 29202 19070 29204 19122
rect 29148 18340 29204 19070
rect 29484 19122 29540 19134
rect 29484 19070 29486 19122
rect 29538 19070 29540 19122
rect 29484 19012 29540 19070
rect 30268 19124 30324 19134
rect 30268 19030 30324 19068
rect 30828 19124 30884 20750
rect 30940 20132 30996 20142
rect 30940 20018 30996 20076
rect 30940 19966 30942 20018
rect 30994 19966 30996 20018
rect 30940 19954 30996 19966
rect 30828 19058 30884 19068
rect 29484 18788 29540 18956
rect 29484 18722 29540 18732
rect 29708 18450 29764 18462
rect 29708 18398 29710 18450
rect 29762 18398 29764 18450
rect 29260 18340 29316 18350
rect 29148 18338 29316 18340
rect 29148 18286 29262 18338
rect 29314 18286 29316 18338
rect 29148 18284 29316 18286
rect 29260 18274 29316 18284
rect 29260 17442 29316 17454
rect 29260 17390 29262 17442
rect 29314 17390 29316 17442
rect 29260 17332 29316 17390
rect 28700 16882 29204 16884
rect 28700 16830 28702 16882
rect 28754 16830 29204 16882
rect 28700 16828 29204 16830
rect 28700 16818 28756 16828
rect 28476 16034 28532 16044
rect 28700 16098 28756 16110
rect 28700 16046 28702 16098
rect 28754 16046 28756 16098
rect 28588 15988 28644 15998
rect 28028 15092 28196 15148
rect 28252 15092 28420 15148
rect 28476 15316 28532 15326
rect 28028 13858 28084 15092
rect 28252 14530 28308 15092
rect 28476 14642 28532 15260
rect 28588 14756 28644 15932
rect 28700 15148 28756 16046
rect 29148 16098 29204 16828
rect 29260 16548 29316 17276
rect 29708 17108 29764 18398
rect 30380 18338 30436 18350
rect 30380 18286 30382 18338
rect 30434 18286 30436 18338
rect 30380 17556 30436 18286
rect 30716 18116 30772 18126
rect 30716 17666 30772 18060
rect 30716 17614 30718 17666
rect 30770 17614 30772 17666
rect 30716 17602 30772 17614
rect 30380 17490 30436 17500
rect 31052 17220 31108 74732
rect 33516 27860 33572 75404
rect 34412 67228 34468 75630
rect 34636 75122 34692 75852
rect 34748 75684 34804 79200
rect 35084 76466 35140 76478
rect 35084 76414 35086 76466
rect 35138 76414 35140 76466
rect 34748 75590 34804 75628
rect 34972 75908 35028 75918
rect 34636 75070 34638 75122
rect 34690 75070 34692 75122
rect 34636 75058 34692 75070
rect 34412 67172 34804 67228
rect 34748 28082 34804 67172
rect 34972 29204 35028 75852
rect 35084 74788 35140 76414
rect 35420 76468 35476 79200
rect 36092 76804 36148 79200
rect 36764 76804 36820 79200
rect 37212 77026 37268 77038
rect 37212 76974 37214 77026
rect 37266 76974 37268 77026
rect 36092 76748 36484 76804
rect 36764 76748 36932 76804
rect 36204 76580 36260 76590
rect 36092 76578 36260 76580
rect 36092 76526 36206 76578
rect 36258 76526 36260 76578
rect 36092 76524 36260 76526
rect 35420 76412 35700 76468
rect 35196 76076 35460 76086
rect 35252 76020 35300 76076
rect 35356 76020 35404 76076
rect 35196 76010 35460 76020
rect 35196 75796 35252 75806
rect 35196 75702 35252 75740
rect 35532 75684 35588 75694
rect 35532 75122 35588 75628
rect 35644 75684 35700 76412
rect 35644 75682 36036 75684
rect 35644 75630 35646 75682
rect 35698 75630 36036 75682
rect 35644 75628 36036 75630
rect 35644 75618 35700 75628
rect 35532 75070 35534 75122
rect 35586 75070 35588 75122
rect 35532 75058 35588 75070
rect 35980 75122 36036 75628
rect 35980 75070 35982 75122
rect 36034 75070 36036 75122
rect 35980 75058 36036 75070
rect 35084 74694 35140 74732
rect 35196 74508 35460 74518
rect 35252 74452 35300 74508
rect 35356 74452 35404 74508
rect 35196 74442 35460 74452
rect 35196 72940 35460 72950
rect 35252 72884 35300 72940
rect 35356 72884 35404 72940
rect 35196 72874 35460 72884
rect 35196 71372 35460 71382
rect 35252 71316 35300 71372
rect 35356 71316 35404 71372
rect 35196 71306 35460 71316
rect 35196 69804 35460 69814
rect 35252 69748 35300 69804
rect 35356 69748 35404 69804
rect 35196 69738 35460 69748
rect 35196 68236 35460 68246
rect 35252 68180 35300 68236
rect 35356 68180 35404 68236
rect 35196 68170 35460 68180
rect 35196 66668 35460 66678
rect 35252 66612 35300 66668
rect 35356 66612 35404 66668
rect 35196 66602 35460 66612
rect 35196 65100 35460 65110
rect 35252 65044 35300 65100
rect 35356 65044 35404 65100
rect 35196 65034 35460 65044
rect 35196 63532 35460 63542
rect 35252 63476 35300 63532
rect 35356 63476 35404 63532
rect 35196 63466 35460 63476
rect 35196 61964 35460 61974
rect 35252 61908 35300 61964
rect 35356 61908 35404 61964
rect 35196 61898 35460 61908
rect 35196 60396 35460 60406
rect 35252 60340 35300 60396
rect 35356 60340 35404 60396
rect 35196 60330 35460 60340
rect 35196 58828 35460 58838
rect 35252 58772 35300 58828
rect 35356 58772 35404 58828
rect 35196 58762 35460 58772
rect 35196 57260 35460 57270
rect 35252 57204 35300 57260
rect 35356 57204 35404 57260
rect 35196 57194 35460 57204
rect 35196 55692 35460 55702
rect 35252 55636 35300 55692
rect 35356 55636 35404 55692
rect 35196 55626 35460 55636
rect 36092 55468 36148 76524
rect 36204 76514 36260 76524
rect 36428 76468 36484 76748
rect 36876 76690 36932 76748
rect 36876 76638 36878 76690
rect 36930 76638 36932 76690
rect 36428 76466 36820 76468
rect 36428 76414 36430 76466
rect 36482 76414 36820 76466
rect 36428 76412 36820 76414
rect 36428 76402 36484 76412
rect 36204 75682 36260 75694
rect 36204 75630 36206 75682
rect 36258 75630 36260 75682
rect 36204 67228 36260 75630
rect 36764 75122 36820 76412
rect 36764 75070 36766 75122
rect 36818 75070 36820 75122
rect 36764 75058 36820 75070
rect 36876 75124 36932 76638
rect 37212 75794 37268 76974
rect 37436 76580 37492 79200
rect 37212 75742 37214 75794
rect 37266 75742 37268 75794
rect 37212 75730 37268 75742
rect 37324 76524 37492 76580
rect 38108 77026 38164 79200
rect 38108 76974 38110 77026
rect 38162 76974 38164 77026
rect 37324 75684 37380 76524
rect 37436 76356 37492 76366
rect 37436 76354 37604 76356
rect 37436 76302 37438 76354
rect 37490 76302 37604 76354
rect 37436 76300 37604 76302
rect 37436 76290 37492 76300
rect 37436 75684 37492 75694
rect 37324 75682 37492 75684
rect 37324 75630 37438 75682
rect 37490 75630 37492 75682
rect 37324 75628 37492 75630
rect 36876 75058 36932 75068
rect 37436 74674 37492 75628
rect 37436 74622 37438 74674
rect 37490 74622 37492 74674
rect 37436 74610 37492 74622
rect 37548 73948 37604 76300
rect 37884 76354 37940 76366
rect 37884 76302 37886 76354
rect 37938 76302 37940 76354
rect 37660 75124 37716 75134
rect 37660 75030 37716 75068
rect 37436 73892 37604 73948
rect 37884 73948 37940 76302
rect 37996 75908 38052 75918
rect 37996 75682 38052 75852
rect 37996 75630 37998 75682
rect 38050 75630 38052 75682
rect 37996 75618 38052 75630
rect 38108 75684 38164 76974
rect 38332 76692 38388 76702
rect 38780 76692 38836 79200
rect 38332 76690 38836 76692
rect 38332 76638 38334 76690
rect 38386 76638 38836 76690
rect 38332 76636 38836 76638
rect 39228 76692 39284 76702
rect 39452 76692 39508 79200
rect 39228 76690 39508 76692
rect 39228 76638 39230 76690
rect 39282 76638 39508 76690
rect 39228 76636 39508 76638
rect 38332 76626 38388 76636
rect 38332 75684 38388 75694
rect 38108 75682 38388 75684
rect 38108 75630 38334 75682
rect 38386 75630 38388 75682
rect 38108 75628 38388 75630
rect 38332 75618 38388 75628
rect 38220 74786 38276 74798
rect 38220 74734 38222 74786
rect 38274 74734 38276 74786
rect 38220 74674 38276 74734
rect 38668 74788 38724 76636
rect 39228 76626 39284 76636
rect 38780 76354 38836 76366
rect 38780 76302 38782 76354
rect 38834 76302 38836 76354
rect 38780 75012 38836 76302
rect 39452 75794 39508 76636
rect 39452 75742 39454 75794
rect 39506 75742 39508 75794
rect 39452 75730 39508 75742
rect 40124 76690 40180 79200
rect 40124 76638 40126 76690
rect 40178 76638 40180 76690
rect 38892 75684 38948 75694
rect 40124 75684 40180 76638
rect 40796 76692 40852 79200
rect 41020 76692 41076 76702
rect 40796 76636 41020 76692
rect 41020 76598 41076 76636
rect 41468 76580 41524 79200
rect 42028 76692 42084 76702
rect 42140 76692 42196 79200
rect 42812 77138 42868 79200
rect 43484 77364 43540 79200
rect 43484 77308 43764 77364
rect 42812 77086 42814 77138
rect 42866 77086 42868 77138
rect 42812 77074 42868 77086
rect 43596 77138 43652 77150
rect 43596 77086 43598 77138
rect 43650 77086 43652 77138
rect 42364 76692 42420 76702
rect 43596 76692 43652 77086
rect 43708 77026 43764 77308
rect 43708 76974 43710 77026
rect 43762 76974 43764 77026
rect 43708 76962 43764 76974
rect 43932 77026 43988 77038
rect 43932 76974 43934 77026
rect 43986 76974 43988 77026
rect 42140 76690 42532 76692
rect 42140 76638 42366 76690
rect 42418 76638 42532 76690
rect 42140 76636 42532 76638
rect 42028 76598 42084 76636
rect 42364 76626 42420 76636
rect 41468 76524 41748 76580
rect 38892 75682 39284 75684
rect 38892 75630 38894 75682
rect 38946 75630 39284 75682
rect 38892 75628 39284 75630
rect 38892 75618 38948 75628
rect 38780 74956 38948 75012
rect 38780 74788 38836 74798
rect 38668 74786 38836 74788
rect 38668 74734 38782 74786
rect 38834 74734 38836 74786
rect 38668 74732 38836 74734
rect 38780 74722 38836 74732
rect 38220 74622 38222 74674
rect 38274 74622 38276 74674
rect 38220 74610 38276 74622
rect 37884 73892 38612 73948
rect 37436 67228 37492 73892
rect 36204 67172 36596 67228
rect 37436 67172 38388 67228
rect 35756 55412 36148 55468
rect 35196 54124 35460 54134
rect 35252 54068 35300 54124
rect 35356 54068 35404 54124
rect 35196 54058 35460 54068
rect 35196 52556 35460 52566
rect 35252 52500 35300 52556
rect 35356 52500 35404 52556
rect 35196 52490 35460 52500
rect 35196 50988 35460 50998
rect 35252 50932 35300 50988
rect 35356 50932 35404 50988
rect 35196 50922 35460 50932
rect 35196 49420 35460 49430
rect 35252 49364 35300 49420
rect 35356 49364 35404 49420
rect 35196 49354 35460 49364
rect 35196 47852 35460 47862
rect 35252 47796 35300 47852
rect 35356 47796 35404 47852
rect 35196 47786 35460 47796
rect 35196 46284 35460 46294
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35196 46218 35460 46228
rect 35196 44716 35460 44726
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35196 44650 35460 44660
rect 35196 43148 35460 43158
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35196 43082 35460 43092
rect 35196 41580 35460 41590
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35196 41514 35460 41524
rect 35196 40012 35460 40022
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35196 39946 35460 39956
rect 35196 38444 35460 38454
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35196 38378 35460 38388
rect 35196 36876 35460 36886
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35196 36810 35460 36820
rect 35196 35308 35460 35318
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35196 35242 35460 35252
rect 35196 33740 35460 33750
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35196 33674 35460 33684
rect 35196 32172 35460 32182
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35196 32106 35460 32116
rect 35196 30604 35460 30614
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35196 30538 35460 30548
rect 34972 29138 35028 29148
rect 35196 29036 35460 29046
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35196 28970 35460 28980
rect 34748 28030 34750 28082
rect 34802 28030 34804 28082
rect 33516 27794 33572 27804
rect 34524 27972 34580 27982
rect 33404 27748 33460 27758
rect 31836 24836 31892 24846
rect 31836 22820 31892 24780
rect 33180 24612 33236 24622
rect 31836 22754 31892 22764
rect 33068 24556 33180 24612
rect 32956 21924 33012 21934
rect 31388 20916 31444 20926
rect 31388 20130 31444 20860
rect 31500 20690 31556 20702
rect 31500 20638 31502 20690
rect 31554 20638 31556 20690
rect 31500 20242 31556 20638
rect 31500 20190 31502 20242
rect 31554 20190 31556 20242
rect 31500 20178 31556 20190
rect 31388 20078 31390 20130
rect 31442 20078 31444 20130
rect 31388 20066 31444 20078
rect 31612 20020 31668 20030
rect 31164 18116 31220 18126
rect 31164 17666 31220 18060
rect 31164 17614 31166 17666
rect 31218 17614 31220 17666
rect 31164 17602 31220 17614
rect 31388 17668 31444 17678
rect 31612 17668 31668 19964
rect 32172 19906 32228 19918
rect 32620 19908 32676 19918
rect 32172 19854 32174 19906
rect 32226 19854 32228 19906
rect 32172 19796 32228 19854
rect 32172 19730 32228 19740
rect 32396 19852 32620 19908
rect 31836 19348 31892 19358
rect 31388 17666 31668 17668
rect 31388 17614 31390 17666
rect 31442 17614 31668 17666
rect 31388 17612 31668 17614
rect 31724 19292 31836 19348
rect 31388 17602 31444 17612
rect 31276 17556 31332 17566
rect 31276 17462 31332 17500
rect 29708 17042 29764 17052
rect 30940 17164 31108 17220
rect 29484 16884 29540 16894
rect 29484 16790 29540 16828
rect 29260 16482 29316 16492
rect 29148 16046 29150 16098
rect 29202 16046 29204 16098
rect 29148 16034 29204 16046
rect 29932 15988 29988 15998
rect 29596 15986 29988 15988
rect 29596 15934 29934 15986
rect 29986 15934 29988 15986
rect 29596 15932 29988 15934
rect 28700 15092 29428 15148
rect 28588 14690 28644 14700
rect 28476 14590 28478 14642
rect 28530 14590 28532 14642
rect 28476 14578 28532 14590
rect 29036 14532 29092 14542
rect 28252 14478 28254 14530
rect 28306 14478 28308 14530
rect 28252 14466 28308 14478
rect 28812 14530 29092 14532
rect 28812 14478 29038 14530
rect 29090 14478 29092 14530
rect 28812 14476 29092 14478
rect 28812 13970 28868 14476
rect 29036 14466 29092 14476
rect 29372 14084 29428 15092
rect 29596 14642 29652 15932
rect 29932 15922 29988 15932
rect 29596 14590 29598 14642
rect 29650 14590 29652 14642
rect 29596 14578 29652 14590
rect 29708 15652 29764 15662
rect 29484 14532 29540 14542
rect 29484 14438 29540 14476
rect 29708 14532 29764 15596
rect 30828 14754 30884 14766
rect 30828 14702 30830 14754
rect 30882 14702 30884 14754
rect 30828 14642 30884 14702
rect 30828 14590 30830 14642
rect 30882 14590 30884 14642
rect 30828 14532 30884 14590
rect 29708 14530 30100 14532
rect 29708 14478 29710 14530
rect 29762 14478 30100 14530
rect 29708 14476 30100 14478
rect 29708 14466 29764 14476
rect 30044 14418 30100 14476
rect 30940 14532 30996 17164
rect 31724 16996 31780 19292
rect 31836 19282 31892 19292
rect 31500 16940 31780 16996
rect 32284 17332 32340 17342
rect 32284 16994 32340 17276
rect 32284 16942 32286 16994
rect 32338 16942 32340 16994
rect 31500 15428 31556 16940
rect 32284 16930 32340 16942
rect 31612 16772 31668 16782
rect 31948 16772 32004 16782
rect 31612 16770 32004 16772
rect 31612 16718 31614 16770
rect 31666 16718 31950 16770
rect 32002 16718 32004 16770
rect 31612 16716 32004 16718
rect 31612 16706 31668 16716
rect 31948 16706 32004 16716
rect 32396 16548 32452 19852
rect 32620 19814 32676 19852
rect 32508 18340 32564 18350
rect 32508 18246 32564 18284
rect 32732 17442 32788 17454
rect 32732 17390 32734 17442
rect 32786 17390 32788 17442
rect 32732 17108 32788 17390
rect 32284 16492 32452 16548
rect 32508 17052 32732 17108
rect 32060 16210 32116 16222
rect 32060 16158 32062 16210
rect 32114 16158 32116 16210
rect 31836 16100 31892 16110
rect 31612 15428 31668 15438
rect 31500 15426 31668 15428
rect 31500 15374 31614 15426
rect 31666 15374 31668 15426
rect 31500 15372 31668 15374
rect 31052 15314 31108 15326
rect 31052 15262 31054 15314
rect 31106 15262 31108 15314
rect 31052 15148 31108 15262
rect 31052 15092 31332 15148
rect 30940 14476 31108 14532
rect 30828 14466 30884 14476
rect 30044 14366 30046 14418
rect 30098 14366 30100 14418
rect 30044 14354 30100 14366
rect 30380 14306 30436 14318
rect 30380 14254 30382 14306
rect 30434 14254 30436 14306
rect 29372 14028 29652 14084
rect 28812 13918 28814 13970
rect 28866 13918 28868 13970
rect 28812 13906 28868 13918
rect 29596 13970 29652 14028
rect 29596 13918 29598 13970
rect 29650 13918 29652 13970
rect 29596 13906 29652 13918
rect 29708 13972 29764 13982
rect 28028 13806 28030 13858
rect 28082 13806 28084 13858
rect 28028 13794 28084 13806
rect 28476 13860 28532 13870
rect 28476 13766 28532 13804
rect 28588 13858 28644 13870
rect 28588 13806 28590 13858
rect 28642 13806 28644 13858
rect 28588 13524 28644 13806
rect 29036 13860 29092 13870
rect 29036 13766 29092 13804
rect 28588 13458 28644 13468
rect 29372 13746 29428 13758
rect 29372 13694 29374 13746
rect 29426 13694 29428 13746
rect 28364 12962 28420 12974
rect 28364 12910 28366 12962
rect 28418 12910 28420 12962
rect 28364 12852 28420 12910
rect 28364 12786 28420 12796
rect 28588 12738 28644 12750
rect 28588 12686 28590 12738
rect 28642 12686 28644 12738
rect 28588 12628 28644 12686
rect 28588 12562 28644 12572
rect 29372 12628 29428 13694
rect 29372 12562 29428 12572
rect 29484 12852 29540 12862
rect 29484 12404 29540 12796
rect 29708 12740 29764 13916
rect 30268 13972 30324 13982
rect 30380 13972 30436 14254
rect 30324 13916 30436 13972
rect 30940 14308 30996 14318
rect 30940 13970 30996 14252
rect 30940 13918 30942 13970
rect 30994 13918 30996 13970
rect 30268 13906 30324 13916
rect 30940 13906 30996 13918
rect 29820 13858 29876 13870
rect 29820 13806 29822 13858
rect 29874 13806 29876 13858
rect 29820 12964 29876 13806
rect 29932 13860 29988 13870
rect 29932 13766 29988 13804
rect 29820 12908 29988 12964
rect 29820 12740 29876 12750
rect 29708 12738 29876 12740
rect 29708 12686 29822 12738
rect 29874 12686 29876 12738
rect 29708 12684 29876 12686
rect 29820 12674 29876 12684
rect 29036 12348 29540 12404
rect 28588 11732 28644 11742
rect 28588 11506 28644 11676
rect 28588 11454 28590 11506
rect 28642 11454 28644 11506
rect 28588 11442 28644 11454
rect 27804 9940 27860 9950
rect 27916 9940 27972 10780
rect 28476 10612 28532 10622
rect 28476 10518 28532 10556
rect 27860 9884 27972 9940
rect 28028 10164 28084 10174
rect 27804 9846 27860 9884
rect 27692 9660 27972 9716
rect 27244 9602 27300 9614
rect 27244 9550 27246 9602
rect 27298 9550 27300 9602
rect 27244 6692 27300 9550
rect 27804 9492 27860 9502
rect 27468 8932 27524 8942
rect 27356 8372 27412 8382
rect 27356 8278 27412 8316
rect 27468 8370 27524 8876
rect 27468 8318 27470 8370
rect 27522 8318 27524 8370
rect 27468 8306 27524 8318
rect 27580 8036 27636 8046
rect 27580 7942 27636 7980
rect 27804 7812 27860 9436
rect 27244 6598 27300 6636
rect 27580 7756 27860 7812
rect 27580 6130 27636 7756
rect 27692 7588 27748 7598
rect 27692 7494 27748 7532
rect 27804 7474 27860 7486
rect 27804 7422 27806 7474
rect 27858 7422 27860 7474
rect 27692 7252 27748 7262
rect 27692 7158 27748 7196
rect 27804 6916 27860 7422
rect 27916 7364 27972 9660
rect 28028 7700 28084 10108
rect 28588 9602 28644 9614
rect 28588 9550 28590 9602
rect 28642 9550 28644 9602
rect 28588 9156 28644 9550
rect 28140 8484 28196 8494
rect 28140 8390 28196 8428
rect 28140 8148 28196 8158
rect 28140 8054 28196 8092
rect 28252 8146 28308 8158
rect 28252 8094 28254 8146
rect 28306 8094 28308 8146
rect 28140 7700 28196 7710
rect 28028 7698 28196 7700
rect 28028 7646 28142 7698
rect 28194 7646 28196 7698
rect 28028 7644 28196 7646
rect 28140 7634 28196 7644
rect 27916 7308 28196 7364
rect 27804 6850 27860 6860
rect 27916 6692 27972 6702
rect 27804 6466 27860 6478
rect 27804 6414 27806 6466
rect 27858 6414 27860 6466
rect 27804 6356 27860 6414
rect 27804 6290 27860 6300
rect 27580 6078 27582 6130
rect 27634 6078 27636 6130
rect 27580 6066 27636 6078
rect 27916 6132 27972 6636
rect 28028 6580 28084 6590
rect 28028 6486 28084 6524
rect 28028 6132 28084 6142
rect 27916 6130 28084 6132
rect 27916 6078 28030 6130
rect 28082 6078 28084 6130
rect 27916 6076 28084 6078
rect 28028 6066 28084 6076
rect 28140 6132 28196 7308
rect 28252 6916 28308 8094
rect 28588 8148 28644 9100
rect 28812 8932 28868 8942
rect 28812 8838 28868 8876
rect 28364 7588 28420 7598
rect 28364 7140 28420 7532
rect 28476 7364 28532 7374
rect 28476 7270 28532 7308
rect 28364 7084 28532 7140
rect 28252 6850 28308 6860
rect 28364 6690 28420 6702
rect 28364 6638 28366 6690
rect 28418 6638 28420 6690
rect 28364 6468 28420 6638
rect 27468 6018 27524 6030
rect 27468 5966 27470 6018
rect 27522 5966 27524 6018
rect 27132 5182 27134 5234
rect 27186 5182 27188 5234
rect 27132 5170 27188 5182
rect 27244 5684 27300 5694
rect 27244 5346 27300 5628
rect 27244 5294 27246 5346
rect 27298 5294 27300 5346
rect 27244 5236 27300 5294
rect 27244 5170 27300 5180
rect 26460 5058 26516 5068
rect 27020 4898 27076 4910
rect 27020 4846 27022 4898
rect 27074 4846 27076 4898
rect 26460 4340 26516 4350
rect 26460 3442 26516 4284
rect 26460 3390 26462 3442
rect 26514 3390 26516 3442
rect 26460 3378 26516 3390
rect 26796 3442 26852 3454
rect 26796 3390 26798 3442
rect 26850 3390 26852 3442
rect 26796 3388 26852 3390
rect 26684 3332 26852 3388
rect 26908 3444 26964 3454
rect 26684 3220 26740 3332
rect 26684 2660 26740 3164
rect 26684 2594 26740 2604
rect 26348 1708 26516 1764
rect 25900 1586 25956 1596
rect 26460 800 26516 1708
rect 26908 1316 26964 3388
rect 27020 1540 27076 4846
rect 27132 4564 27188 4574
rect 27132 3442 27188 4508
rect 27468 3892 27524 5966
rect 27916 5908 27972 5918
rect 27692 5684 27748 5694
rect 27580 5628 27692 5684
rect 27580 5010 27636 5628
rect 27692 5590 27748 5628
rect 27580 4958 27582 5010
rect 27634 4958 27636 5010
rect 27580 4946 27636 4958
rect 27804 5572 27860 5582
rect 27804 4116 27860 5516
rect 27916 5122 27972 5852
rect 27916 5070 27918 5122
rect 27970 5070 27972 5122
rect 27916 5058 27972 5070
rect 28140 4226 28196 6076
rect 28252 6244 28308 6254
rect 28252 5124 28308 6188
rect 28364 5906 28420 6412
rect 28476 6244 28532 7084
rect 28588 6690 28644 8092
rect 29036 7698 29092 12348
rect 29708 12178 29764 12190
rect 29708 12126 29710 12178
rect 29762 12126 29764 12178
rect 29708 10612 29764 12126
rect 29932 11732 29988 12908
rect 30380 12068 30436 12078
rect 29932 11666 29988 11676
rect 30156 12066 30436 12068
rect 30156 12014 30382 12066
rect 30434 12014 30436 12066
rect 30156 12012 30436 12014
rect 30156 11506 30212 12012
rect 30380 12002 30436 12012
rect 30156 11454 30158 11506
rect 30210 11454 30212 11506
rect 30156 11442 30212 11454
rect 30380 11284 30436 11294
rect 30380 11190 30436 11228
rect 30156 11172 30212 11182
rect 30156 11078 30212 11116
rect 31052 11060 31108 14476
rect 31276 14306 31332 15092
rect 31500 14754 31556 15372
rect 31612 15362 31668 15372
rect 31500 14702 31502 14754
rect 31554 14702 31556 14754
rect 31500 14690 31556 14702
rect 31836 14530 31892 16044
rect 31948 15428 32004 15438
rect 32060 15428 32116 16158
rect 31948 15426 32116 15428
rect 31948 15374 31950 15426
rect 32002 15374 32116 15426
rect 31948 15372 32116 15374
rect 31948 15362 32004 15372
rect 32284 14644 32340 16492
rect 32508 16100 32564 17052
rect 32732 17042 32788 17052
rect 32508 16006 32564 16044
rect 32956 15652 33012 21868
rect 33068 15764 33124 24556
rect 33180 24546 33236 24556
rect 33404 23044 33460 27692
rect 34076 27076 34132 27086
rect 34076 26982 34132 27020
rect 33964 26852 34020 26862
rect 33628 26850 34020 26852
rect 33628 26798 33966 26850
rect 34018 26798 34020 26850
rect 33628 26796 34020 26798
rect 33628 24500 33684 26796
rect 33964 26786 34020 26796
rect 33404 22978 33460 22988
rect 33516 24444 33684 24500
rect 33516 22258 33572 24444
rect 34300 23714 34356 23726
rect 34300 23662 34302 23714
rect 34354 23662 34356 23714
rect 34300 23604 34356 23662
rect 34300 23538 34356 23548
rect 33740 23380 33796 23390
rect 34524 23380 34580 27916
rect 34748 27074 34804 28030
rect 35756 28084 35812 55412
rect 36540 31948 36596 67172
rect 35084 27970 35140 27982
rect 35084 27918 35086 27970
rect 35138 27918 35140 27970
rect 34972 27300 35028 27310
rect 34748 27022 34750 27074
rect 34802 27022 34804 27074
rect 34748 27010 34804 27022
rect 34860 27244 34972 27300
rect 34748 23940 34804 23950
rect 34748 23846 34804 23884
rect 33740 23378 34580 23380
rect 33740 23326 33742 23378
rect 33794 23326 34526 23378
rect 34578 23326 34580 23378
rect 33740 23324 34580 23326
rect 33740 23314 33796 23324
rect 34524 23314 34580 23324
rect 34860 23380 34916 27244
rect 34972 27234 35028 27244
rect 34972 26964 35028 26974
rect 35084 26964 35140 27918
rect 35308 27860 35364 27870
rect 35308 27766 35364 27804
rect 35532 27746 35588 27758
rect 35532 27694 35534 27746
rect 35586 27694 35588 27746
rect 35196 27468 35460 27478
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35196 27402 35460 27412
rect 35028 26908 35140 26964
rect 34972 26870 35028 26908
rect 35420 26852 35476 26862
rect 35196 26516 35252 26526
rect 35196 26422 35252 26460
rect 35420 26068 35476 26796
rect 35532 26628 35588 27694
rect 35756 27074 35812 28028
rect 35756 27022 35758 27074
rect 35810 27022 35812 27074
rect 35756 27010 35812 27022
rect 35980 31892 36596 31948
rect 35644 26964 35700 26974
rect 35644 26852 35924 26908
rect 35532 26572 35700 26628
rect 35420 26012 35588 26068
rect 35196 25900 35460 25910
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35196 25834 35460 25844
rect 35532 25732 35588 26012
rect 35308 25676 35588 25732
rect 34972 24948 35028 24958
rect 35308 24948 35364 25676
rect 35532 25508 35588 25518
rect 35532 25284 35588 25452
rect 34972 24946 35364 24948
rect 34972 24894 34974 24946
rect 35026 24894 35310 24946
rect 35362 24894 35364 24946
rect 34972 24892 35364 24894
rect 34972 24882 35028 24892
rect 35308 24882 35364 24892
rect 35420 25282 35588 25284
rect 35420 25230 35534 25282
rect 35586 25230 35588 25282
rect 35420 25228 35588 25230
rect 35420 24948 35476 25228
rect 35532 25218 35588 25228
rect 35420 24882 35476 24892
rect 35084 24722 35140 24734
rect 35084 24670 35086 24722
rect 35138 24670 35140 24722
rect 35084 23940 35140 24670
rect 35420 24724 35476 24734
rect 35420 24722 35588 24724
rect 35420 24670 35422 24722
rect 35474 24670 35588 24722
rect 35420 24668 35588 24670
rect 35420 24658 35476 24668
rect 35196 24332 35460 24342
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35196 24266 35460 24276
rect 35084 23884 35252 23940
rect 35084 23716 35140 23726
rect 35084 23622 35140 23660
rect 35196 23492 35252 23884
rect 35196 23436 35364 23492
rect 35084 23380 35140 23390
rect 34860 23378 35140 23380
rect 34860 23326 35086 23378
rect 35138 23326 35140 23378
rect 34860 23324 35140 23326
rect 34188 23156 34244 23166
rect 34188 23062 34244 23100
rect 34300 23154 34356 23166
rect 34636 23156 34692 23166
rect 34300 23102 34302 23154
rect 34354 23102 34356 23154
rect 34300 22370 34356 23102
rect 34300 22318 34302 22370
rect 34354 22318 34356 22370
rect 34300 22306 34356 22318
rect 34412 23154 34692 23156
rect 34412 23102 34638 23154
rect 34690 23102 34692 23154
rect 34412 23100 34692 23102
rect 33516 22206 33518 22258
rect 33570 22206 33572 22258
rect 33516 22194 33572 22206
rect 34300 22146 34356 22158
rect 34300 22094 34302 22146
rect 34354 22094 34356 22146
rect 33292 21474 33348 21486
rect 33292 21422 33294 21474
rect 33346 21422 33348 21474
rect 33292 20916 33348 21422
rect 33292 20850 33348 20860
rect 33628 21474 33684 21486
rect 33628 21422 33630 21474
rect 33682 21422 33684 21474
rect 33628 20914 33684 21422
rect 33628 20862 33630 20914
rect 33682 20862 33684 20914
rect 33628 20850 33684 20862
rect 34188 20804 34244 20814
rect 33964 20802 34244 20804
rect 33964 20750 34190 20802
rect 34242 20750 34244 20802
rect 33964 20748 34244 20750
rect 33516 20692 33572 20702
rect 33516 20130 33572 20636
rect 33964 20242 34020 20748
rect 34188 20738 34244 20748
rect 33964 20190 33966 20242
rect 34018 20190 34020 20242
rect 33964 20178 34020 20190
rect 34300 20132 34356 22094
rect 34412 20914 34468 23100
rect 34636 23090 34692 23100
rect 34860 23156 34916 23324
rect 35084 23314 35140 23324
rect 35196 23156 35252 23166
rect 34860 23090 34916 23100
rect 34972 23154 35252 23156
rect 34972 23102 35198 23154
rect 35250 23102 35252 23154
rect 34972 23100 35252 23102
rect 34748 21588 34804 21598
rect 34524 21476 34580 21486
rect 34524 21382 34580 21420
rect 34412 20862 34414 20914
rect 34466 20862 34468 20914
rect 34412 20850 34468 20862
rect 34636 20690 34692 20702
rect 34636 20638 34638 20690
rect 34690 20638 34692 20690
rect 34636 20468 34692 20638
rect 34636 20402 34692 20412
rect 34412 20244 34468 20254
rect 34412 20150 34468 20188
rect 34748 20244 34804 21532
rect 34860 21474 34916 21486
rect 34860 21422 34862 21474
rect 34914 21422 34916 21474
rect 34860 21364 34916 21422
rect 34860 21298 34916 21308
rect 34972 21252 35028 23100
rect 35196 23090 35252 23100
rect 35308 23156 35364 23436
rect 35308 23090 35364 23100
rect 35084 22930 35140 22942
rect 35084 22878 35086 22930
rect 35138 22878 35140 22930
rect 35084 22484 35140 22878
rect 35532 22932 35588 24668
rect 35644 24612 35700 26572
rect 35868 26402 35924 26852
rect 35868 26350 35870 26402
rect 35922 26350 35924 26402
rect 35756 26178 35812 26190
rect 35756 26126 35758 26178
rect 35810 26126 35812 26178
rect 35756 24834 35812 26126
rect 35868 25618 35924 26350
rect 35980 26516 36036 31892
rect 38332 28868 38388 67172
rect 37548 28812 38388 28868
rect 37548 28754 37604 28812
rect 37548 28702 37550 28754
rect 37602 28702 37604 28754
rect 37548 28690 37604 28702
rect 37884 28644 37940 28654
rect 37884 28642 38164 28644
rect 37884 28590 37886 28642
rect 37938 28590 38164 28642
rect 37884 28588 38164 28590
rect 37660 28532 37716 28542
rect 36652 28420 36708 28430
rect 36540 28364 36652 28420
rect 36204 27858 36260 27870
rect 36204 27806 36206 27858
rect 36258 27806 36260 27858
rect 36204 27076 36260 27806
rect 36260 27020 36372 27076
rect 36204 27010 36260 27020
rect 35980 26290 36036 26460
rect 35980 26238 35982 26290
rect 36034 26238 36036 26290
rect 35980 26226 36036 26238
rect 36204 26850 36260 26862
rect 36204 26798 36206 26850
rect 36258 26798 36260 26850
rect 35868 25566 35870 25618
rect 35922 25566 35924 25618
rect 35868 25554 35924 25566
rect 35756 24782 35758 24834
rect 35810 24782 35812 24834
rect 35756 24770 35812 24782
rect 35980 24722 36036 24734
rect 35980 24670 35982 24722
rect 36034 24670 36036 24722
rect 35644 24556 35812 24612
rect 35644 23828 35700 23838
rect 35644 23734 35700 23772
rect 35756 23604 35812 24556
rect 35980 24162 36036 24670
rect 35980 24110 35982 24162
rect 36034 24110 36036 24162
rect 35980 24098 36036 24110
rect 35868 23940 35924 23950
rect 35868 23938 36148 23940
rect 35868 23886 35870 23938
rect 35922 23886 36148 23938
rect 35868 23884 36148 23886
rect 35868 23874 35924 23884
rect 35980 23714 36036 23726
rect 35980 23662 35982 23714
rect 36034 23662 36036 23714
rect 35980 23604 36036 23662
rect 35756 23548 35924 23604
rect 35868 23266 35924 23548
rect 35980 23538 36036 23548
rect 35868 23214 35870 23266
rect 35922 23214 35924 23266
rect 35868 23202 35924 23214
rect 35756 23156 35812 23166
rect 35756 23062 35812 23100
rect 36092 23044 36148 23884
rect 36204 23380 36260 26798
rect 36316 26290 36372 27020
rect 36316 26238 36318 26290
rect 36370 26238 36372 26290
rect 36316 26226 36372 26238
rect 36428 25396 36484 25406
rect 36428 25302 36484 25340
rect 36540 23604 36596 28364
rect 36652 28354 36708 28364
rect 37100 28084 37156 28094
rect 37100 27990 37156 28028
rect 37660 28082 37716 28476
rect 37660 28030 37662 28082
rect 37714 28030 37716 28082
rect 37660 28018 37716 28030
rect 36652 27860 36708 27870
rect 37884 27860 37940 28588
rect 36652 27766 36708 27804
rect 37772 27858 37940 27860
rect 37772 27806 37886 27858
rect 37938 27806 37940 27858
rect 37772 27804 37940 27806
rect 36988 27076 37044 27086
rect 37436 27076 37492 27086
rect 36988 26982 37044 27020
rect 37324 27074 37492 27076
rect 37324 27022 37438 27074
rect 37490 27022 37492 27074
rect 37324 27020 37492 27022
rect 37324 26290 37380 27020
rect 37436 27010 37492 27020
rect 37324 26238 37326 26290
rect 37378 26238 37380 26290
rect 37324 25732 37380 26238
rect 37772 26290 37828 27804
rect 37884 27794 37940 27804
rect 37996 28418 38052 28430
rect 37996 28366 37998 28418
rect 38050 28366 38052 28418
rect 37772 26238 37774 26290
rect 37826 26238 37828 26290
rect 37772 26226 37828 26238
rect 37324 25666 37380 25676
rect 37772 25620 37828 25630
rect 37772 25526 37828 25564
rect 37324 25506 37380 25518
rect 37324 25454 37326 25506
rect 37378 25454 37380 25506
rect 37324 25396 37380 25454
rect 37996 25508 38052 28366
rect 38108 27074 38164 28588
rect 38332 28642 38388 28812
rect 38332 28590 38334 28642
rect 38386 28590 38388 28642
rect 38332 28578 38388 28590
rect 38556 28532 38612 73892
rect 38892 38668 38948 74956
rect 39228 67228 39284 75628
rect 40124 75618 40180 75628
rect 40684 76354 40740 76366
rect 40684 76302 40686 76354
rect 40738 76302 40740 76354
rect 39228 67172 39956 67228
rect 38892 38612 39172 38668
rect 38892 29204 38948 29214
rect 38948 29148 39060 29204
rect 38892 29138 38948 29148
rect 38612 28476 38724 28532
rect 38556 28466 38612 28476
rect 38108 27022 38110 27074
rect 38162 27022 38164 27074
rect 38108 26290 38164 27022
rect 38556 27746 38612 27758
rect 38556 27694 38558 27746
rect 38610 27694 38612 27746
rect 38108 26238 38110 26290
rect 38162 26238 38164 26290
rect 38108 26226 38164 26238
rect 38332 26850 38388 26862
rect 38332 26798 38334 26850
rect 38386 26798 38388 26850
rect 38332 26180 38388 26798
rect 38556 26404 38612 27694
rect 38668 27074 38724 28476
rect 38668 27022 38670 27074
rect 38722 27022 38724 27074
rect 38668 27010 38724 27022
rect 38780 28530 38836 28542
rect 38780 28478 38782 28530
rect 38834 28478 38836 28530
rect 38780 27970 38836 28478
rect 38780 27918 38782 27970
rect 38834 27918 38836 27970
rect 38780 26962 38836 27918
rect 39004 27860 39060 29148
rect 39116 28084 39172 38612
rect 39900 28084 39956 67172
rect 40684 38668 40740 76302
rect 41468 75794 41524 76524
rect 41468 75742 41470 75794
rect 41522 75742 41524 75794
rect 41468 75730 41524 75742
rect 41580 76354 41636 76366
rect 41580 76302 41582 76354
rect 41634 76302 41636 76354
rect 40908 75684 40964 75694
rect 40908 75590 40964 75628
rect 41580 43708 41636 76302
rect 41692 75682 41748 76524
rect 42476 75794 42532 76636
rect 43372 76690 43652 76692
rect 43372 76638 43598 76690
rect 43650 76638 43652 76690
rect 43372 76636 43652 76638
rect 42476 75742 42478 75794
rect 42530 75742 42532 75794
rect 42476 75730 42532 75742
rect 42924 76354 42980 76366
rect 42924 76302 42926 76354
rect 42978 76302 42980 76354
rect 41692 75630 41694 75682
rect 41746 75630 41748 75682
rect 41692 75618 41748 75630
rect 42028 75458 42084 75470
rect 42028 75406 42030 75458
rect 42082 75406 42084 75458
rect 42028 43708 42084 75406
rect 42924 43708 42980 76302
rect 43372 75794 43428 76636
rect 43596 76626 43652 76636
rect 43372 75742 43374 75794
rect 43426 75742 43428 75794
rect 43372 75730 43428 75742
rect 43932 75794 43988 76974
rect 44156 76692 44212 79200
rect 44156 76626 44212 76636
rect 44492 77026 44548 77038
rect 44492 76974 44494 77026
rect 44546 76974 44548 77026
rect 44492 76690 44548 76974
rect 44828 76804 44884 79200
rect 45500 77026 45556 79200
rect 45500 76974 45502 77026
rect 45554 76974 45556 77026
rect 45500 76962 45556 76974
rect 44492 76638 44494 76690
rect 44546 76638 44548 76690
rect 44492 76626 44548 76638
rect 44604 76748 45108 76804
rect 43932 75742 43934 75794
rect 43986 75742 43988 75794
rect 43932 75730 43988 75742
rect 44044 76354 44100 76366
rect 44604 76356 44660 76748
rect 44044 76302 44046 76354
rect 44098 76302 44100 76354
rect 44044 55468 44100 76302
rect 44380 76300 44660 76356
rect 44940 76354 44996 76366
rect 44940 76302 44942 76354
rect 44994 76302 44996 76354
rect 44380 75794 44436 76300
rect 44380 75742 44382 75794
rect 44434 75742 44436 75794
rect 44380 75730 44436 75742
rect 44940 55468 44996 76302
rect 45052 75682 45108 76748
rect 45836 76692 45892 76702
rect 46172 76692 46228 79200
rect 45892 76636 46004 76692
rect 45836 76626 45892 76636
rect 45948 76580 46004 76636
rect 46172 76626 46228 76636
rect 46732 77026 46788 77038
rect 46732 76974 46734 77026
rect 46786 76974 46788 77026
rect 45948 76578 46116 76580
rect 45948 76526 45950 76578
rect 46002 76526 46116 76578
rect 45948 76524 46116 76526
rect 45948 76514 46004 76524
rect 45500 76356 45556 76366
rect 45500 76354 45892 76356
rect 45500 76302 45502 76354
rect 45554 76302 45892 76354
rect 45500 76300 45892 76302
rect 45500 76290 45556 76300
rect 45836 75906 45892 76300
rect 45836 75854 45838 75906
rect 45890 75854 45892 75906
rect 45836 75842 45892 75854
rect 46060 75794 46116 76524
rect 46732 76466 46788 76974
rect 46844 76692 46900 79200
rect 47516 77026 47572 79200
rect 47516 76974 47518 77026
rect 47570 76974 47572 77026
rect 47516 76962 47572 76974
rect 47852 76692 47908 76702
rect 46844 76636 47124 76692
rect 46732 76414 46734 76466
rect 46786 76414 46788 76466
rect 46060 75742 46062 75794
rect 46114 75742 46116 75794
rect 46060 75730 46116 75742
rect 46284 76354 46340 76366
rect 46284 76302 46286 76354
rect 46338 76302 46340 76354
rect 45052 75630 45054 75682
rect 45106 75630 45108 75682
rect 45052 75618 45108 75630
rect 45612 75572 45668 75582
rect 43932 55412 44100 55468
rect 44268 55412 44996 55468
rect 45500 75570 45668 75572
rect 45500 75518 45614 75570
rect 45666 75518 45668 75570
rect 45500 75516 45668 75518
rect 41580 43652 41860 43708
rect 42028 43652 42532 43708
rect 42924 43652 43092 43708
rect 41132 39060 41188 39070
rect 40796 38948 40852 38958
rect 40796 38836 40852 38892
rect 40908 38836 40964 38846
rect 40796 38834 40964 38836
rect 40796 38782 40910 38834
rect 40962 38782 40964 38834
rect 40796 38780 40964 38782
rect 40908 38770 40964 38780
rect 41132 38724 41188 39004
rect 41244 38948 41300 38958
rect 41244 38946 41748 38948
rect 41244 38894 41246 38946
rect 41298 38894 41748 38946
rect 41244 38892 41748 38894
rect 41244 38882 41300 38892
rect 41692 38836 41748 38892
rect 41580 38724 41636 38734
rect 41132 38668 41524 38724
rect 40684 38612 40964 38668
rect 40908 28756 40964 38612
rect 41468 38162 41524 38668
rect 41580 38630 41636 38668
rect 41468 38110 41470 38162
rect 41522 38110 41524 38162
rect 41468 38098 41524 38110
rect 40684 28754 40964 28756
rect 40684 28702 40910 28754
rect 40962 28702 40964 28754
rect 40684 28700 40964 28702
rect 39116 28018 39172 28028
rect 39676 28082 39956 28084
rect 39676 28030 39902 28082
rect 39954 28030 39956 28082
rect 39676 28028 39956 28030
rect 39452 27860 39508 27870
rect 39004 27858 39508 27860
rect 39004 27806 39006 27858
rect 39058 27806 39454 27858
rect 39506 27806 39508 27858
rect 39004 27804 39508 27806
rect 39004 27794 39060 27804
rect 39452 27794 39508 27804
rect 38780 26910 38782 26962
rect 38834 26910 38836 26962
rect 38556 26348 38724 26404
rect 38332 26114 38388 26124
rect 38556 26178 38612 26190
rect 38556 26126 38558 26178
rect 38610 26126 38612 26178
rect 38444 25956 38500 25966
rect 38332 25844 38388 25854
rect 38220 25788 38332 25844
rect 38108 25508 38164 25518
rect 37996 25506 38164 25508
rect 37996 25454 38110 25506
rect 38162 25454 38164 25506
rect 37996 25452 38164 25454
rect 38108 25442 38164 25452
rect 37324 25330 37380 25340
rect 37436 24946 37492 24958
rect 37436 24894 37438 24946
rect 37490 24894 37492 24946
rect 37436 24612 37492 24894
rect 37436 24546 37492 24556
rect 37548 24722 37604 24734
rect 37548 24670 37550 24722
rect 37602 24670 37604 24722
rect 37212 24388 37268 24398
rect 37212 23940 37268 24332
rect 37548 23940 37604 24670
rect 37884 24724 37940 24734
rect 37884 24630 37940 24668
rect 37884 24276 37940 24286
rect 37100 23826 37156 23838
rect 37100 23774 37102 23826
rect 37154 23774 37156 23826
rect 36540 23538 36596 23548
rect 36764 23604 36820 23614
rect 36204 23324 36372 23380
rect 35532 22866 35588 22876
rect 35868 22988 36148 23044
rect 35196 22764 35460 22774
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35196 22698 35460 22708
rect 35868 22596 35924 22988
rect 35420 22540 35924 22596
rect 36204 22932 36260 22942
rect 35084 22428 35252 22484
rect 35084 21588 35140 21598
rect 35084 21494 35140 21532
rect 35196 21364 35252 22428
rect 35308 22372 35364 22382
rect 35308 22278 35364 22316
rect 35420 21810 35476 22540
rect 35756 22372 35812 22382
rect 35756 22258 35812 22316
rect 35756 22206 35758 22258
rect 35810 22206 35812 22258
rect 35756 22194 35812 22206
rect 35420 21758 35422 21810
rect 35474 21758 35476 21810
rect 35420 21746 35476 21758
rect 36204 21810 36260 22876
rect 36204 21758 36206 21810
rect 36258 21758 36260 21810
rect 36204 21746 36260 21758
rect 35532 21586 35588 21598
rect 35532 21534 35534 21586
rect 35586 21534 35588 21586
rect 35308 21364 35364 21374
rect 35196 21308 35308 21364
rect 35308 21298 35364 21308
rect 34972 21196 35140 21252
rect 35084 20916 35140 21196
rect 35196 21196 35460 21206
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35196 21130 35460 21140
rect 35420 21028 35476 21038
rect 35308 20916 35364 20926
rect 35084 20914 35364 20916
rect 35084 20862 35310 20914
rect 35362 20862 35364 20914
rect 35084 20860 35364 20862
rect 35308 20850 35364 20860
rect 34860 20804 34916 20814
rect 34860 20710 34916 20748
rect 35196 20692 35252 20702
rect 35196 20598 35252 20636
rect 35420 20468 35476 20972
rect 35532 20692 35588 21534
rect 35756 21588 35812 21598
rect 35756 20804 35812 21532
rect 35980 21586 36036 21598
rect 35980 21534 35982 21586
rect 36034 21534 36036 21586
rect 35980 21028 36036 21534
rect 35980 20962 36036 20972
rect 36204 21364 36260 21374
rect 35812 20748 36148 20804
rect 35756 20710 35812 20748
rect 35532 20598 35588 20636
rect 36092 20690 36148 20748
rect 36092 20638 36094 20690
rect 36146 20638 36148 20690
rect 36092 20626 36148 20638
rect 34748 20178 34804 20188
rect 34860 20412 35476 20468
rect 35644 20468 35700 20478
rect 33516 20078 33518 20130
rect 33570 20078 33572 20130
rect 33516 20066 33572 20078
rect 34188 20076 34356 20132
rect 34860 20130 34916 20412
rect 34860 20078 34862 20130
rect 34914 20078 34916 20130
rect 33404 19906 33460 19918
rect 33404 19854 33406 19906
rect 33458 19854 33460 19906
rect 33180 18340 33236 18350
rect 33404 18340 33460 19854
rect 33852 19906 33908 19918
rect 33852 19854 33854 19906
rect 33906 19854 33908 19906
rect 33852 19796 33908 19854
rect 33852 19730 33908 19740
rect 33740 19684 33796 19694
rect 33180 18338 33460 18340
rect 33180 18286 33182 18338
rect 33234 18286 33460 18338
rect 33180 18284 33460 18286
rect 33516 18340 33572 18350
rect 33740 18340 33796 19628
rect 34076 19124 34132 19134
rect 33180 17892 33236 18284
rect 33516 18246 33572 18284
rect 33628 18338 33796 18340
rect 33628 18286 33742 18338
rect 33794 18286 33796 18338
rect 33628 18284 33796 18286
rect 33628 18116 33684 18284
rect 33740 18274 33796 18284
rect 33964 19068 34076 19124
rect 33628 18050 33684 18060
rect 33180 17826 33236 17836
rect 33740 18004 33796 18014
rect 33404 17780 33460 17790
rect 33740 17780 33796 17948
rect 33852 17892 33908 17902
rect 33964 17892 34020 19068
rect 34076 19058 34132 19068
rect 33852 17890 34020 17892
rect 33852 17838 33854 17890
rect 33906 17838 34020 17890
rect 33852 17836 34020 17838
rect 33852 17826 33908 17836
rect 34188 17780 34244 20076
rect 34860 20066 34916 20078
rect 35308 20132 35364 20142
rect 34748 20020 34804 20030
rect 35308 20020 35364 20076
rect 35532 20132 35588 20142
rect 35532 20038 35588 20076
rect 35420 20020 35476 20030
rect 35308 19964 35420 20020
rect 34300 19908 34356 19918
rect 34300 19814 34356 19852
rect 34748 19906 34804 19964
rect 35420 19926 35476 19964
rect 34748 19854 34750 19906
rect 34802 19854 34804 19906
rect 33404 17686 33460 17724
rect 33516 17778 33796 17780
rect 33516 17726 33742 17778
rect 33794 17726 33796 17778
rect 33516 17724 33796 17726
rect 33404 17108 33460 17118
rect 33516 17108 33572 17724
rect 33740 17714 33796 17724
rect 33964 17724 34244 17780
rect 34412 19234 34468 19246
rect 34412 19182 34414 19234
rect 34466 19182 34468 19234
rect 34412 18450 34468 19182
rect 34412 18398 34414 18450
rect 34466 18398 34468 18450
rect 34412 17780 34468 18398
rect 34748 18452 34804 19854
rect 35644 19684 35700 20412
rect 36204 20018 36260 21308
rect 36316 20130 36372 23324
rect 36652 23378 36708 23390
rect 36652 23326 36654 23378
rect 36706 23326 36708 23378
rect 36652 21924 36708 23326
rect 36652 21858 36708 21868
rect 36428 21586 36484 21598
rect 36428 21534 36430 21586
rect 36482 21534 36484 21586
rect 36428 21028 36484 21534
rect 36540 21588 36596 21598
rect 36540 21494 36596 21532
rect 36428 20972 36596 21028
rect 36428 20804 36484 20814
rect 36428 20710 36484 20748
rect 36540 20692 36596 20972
rect 36540 20626 36596 20636
rect 36316 20078 36318 20130
rect 36370 20078 36372 20130
rect 36316 20066 36372 20078
rect 36204 19966 36206 20018
rect 36258 19966 36260 20018
rect 36204 19954 36260 19966
rect 36428 20020 36484 20030
rect 36484 19964 36596 20020
rect 36428 19954 36484 19964
rect 35196 19628 35460 19638
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35196 19562 35460 19572
rect 35532 19628 35700 19684
rect 35756 19684 35812 19694
rect 35532 19346 35588 19628
rect 35532 19294 35534 19346
rect 35586 19294 35588 19346
rect 35532 19282 35588 19294
rect 35756 19348 35812 19628
rect 36428 19572 36484 19582
rect 35756 19282 35812 19292
rect 36316 19516 36428 19572
rect 35644 19234 35700 19246
rect 35644 19182 35646 19234
rect 35698 19182 35700 19234
rect 35420 19124 35476 19134
rect 35420 19030 35476 19068
rect 34748 18386 34804 18396
rect 35532 19012 35588 19022
rect 35196 18060 35460 18070
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35196 17994 35460 18004
rect 35532 17892 35588 18956
rect 35308 17836 35588 17892
rect 33964 17332 34020 17724
rect 34412 17714 34468 17724
rect 34748 17780 34804 17790
rect 34748 17686 34804 17724
rect 35084 17780 35140 17790
rect 35084 17666 35140 17724
rect 35308 17778 35364 17836
rect 35308 17726 35310 17778
rect 35362 17726 35364 17778
rect 35308 17714 35364 17726
rect 35084 17614 35086 17666
rect 35138 17614 35140 17666
rect 35084 17602 35140 17614
rect 35532 17668 35588 17678
rect 35644 17668 35700 19182
rect 35868 19234 35924 19246
rect 35868 19182 35870 19234
rect 35922 19182 35924 19234
rect 35532 17666 35700 17668
rect 35532 17614 35534 17666
rect 35586 17614 35700 17666
rect 35532 17612 35700 17614
rect 35532 17602 35588 17612
rect 33404 17106 33572 17108
rect 33404 17054 33406 17106
rect 33458 17054 33572 17106
rect 33404 17052 33572 17054
rect 33740 17276 34020 17332
rect 34188 17554 34244 17566
rect 34188 17502 34190 17554
rect 34242 17502 34244 17554
rect 33404 17042 33460 17052
rect 33180 15988 33236 15998
rect 33180 15986 33572 15988
rect 33180 15934 33182 15986
rect 33234 15934 33572 15986
rect 33180 15932 33572 15934
rect 33180 15922 33236 15932
rect 33068 15708 33348 15764
rect 32956 15596 33124 15652
rect 32956 15314 33012 15326
rect 32956 15262 32958 15314
rect 33010 15262 33012 15314
rect 32956 15148 33012 15262
rect 32284 14578 32340 14588
rect 32844 15092 33012 15148
rect 31836 14478 31838 14530
rect 31890 14478 31892 14530
rect 31836 14466 31892 14478
rect 32508 14420 32564 14430
rect 32508 14326 32564 14364
rect 31276 14254 31278 14306
rect 31330 14254 31332 14306
rect 31276 14084 31332 14254
rect 31276 14028 31556 14084
rect 31164 13858 31220 13870
rect 31164 13806 31166 13858
rect 31218 13806 31220 13858
rect 31164 13636 31220 13806
rect 31276 13748 31332 13758
rect 31276 13654 31332 13692
rect 31164 13570 31220 13580
rect 31500 12740 31556 14028
rect 31724 13858 31780 13870
rect 31724 13806 31726 13858
rect 31778 13806 31780 13858
rect 31612 13748 31668 13758
rect 31612 13654 31668 13692
rect 31500 12674 31556 12684
rect 31612 12962 31668 12974
rect 31612 12910 31614 12962
rect 31666 12910 31668 12962
rect 31612 12628 31668 12910
rect 31612 12562 31668 12572
rect 31724 11396 31780 13806
rect 32284 13860 32340 13870
rect 32284 13858 32452 13860
rect 32284 13806 32286 13858
rect 32338 13806 32452 13858
rect 32284 13804 32452 13806
rect 32284 13794 32340 13804
rect 31948 13748 32004 13758
rect 31948 13654 32004 13692
rect 32172 13746 32228 13758
rect 32172 13694 32174 13746
rect 32226 13694 32228 13746
rect 32172 13636 32228 13694
rect 32396 13748 32452 13804
rect 32508 13804 32788 13860
rect 32508 13748 32564 13804
rect 32396 13692 32564 13748
rect 32172 12964 32228 13580
rect 32620 13636 32676 13646
rect 32284 13524 32340 13534
rect 32508 13524 32564 13534
rect 32284 13522 32508 13524
rect 32284 13470 32286 13522
rect 32338 13470 32508 13522
rect 32284 13468 32508 13470
rect 32284 13458 32340 13468
rect 32508 13458 32564 13468
rect 31836 12962 32228 12964
rect 31836 12910 32174 12962
rect 32226 12910 32228 12962
rect 31836 12908 32228 12910
rect 31836 12850 31892 12908
rect 32172 12898 32228 12908
rect 31836 12798 31838 12850
rect 31890 12798 31892 12850
rect 31836 12786 31892 12798
rect 32284 12738 32340 12750
rect 32284 12686 32286 12738
rect 32338 12686 32340 12738
rect 31052 10994 31108 11004
rect 31612 11340 31780 11396
rect 31948 11956 32004 11966
rect 31948 11394 32004 11900
rect 32284 11788 32340 12686
rect 32508 12738 32564 12750
rect 32508 12686 32510 12738
rect 32562 12686 32564 12738
rect 32508 12404 32564 12686
rect 32508 12338 32564 12348
rect 32508 12068 32564 12078
rect 32620 12068 32676 13580
rect 32564 12012 32676 12068
rect 32508 11974 32564 12012
rect 31948 11342 31950 11394
rect 32002 11342 32004 11394
rect 29148 10498 29204 10510
rect 29148 10446 29150 10498
rect 29202 10446 29204 10498
rect 29148 10050 29204 10446
rect 29148 9998 29150 10050
rect 29202 9998 29204 10050
rect 29148 9986 29204 9998
rect 29484 9716 29540 9726
rect 29484 9622 29540 9660
rect 29260 9604 29316 9614
rect 29260 9510 29316 9548
rect 29708 9380 29764 10556
rect 31276 10500 31332 10510
rect 31276 10406 31332 10444
rect 31612 10276 31668 11340
rect 31948 11330 32004 11342
rect 32060 11732 32340 11788
rect 32508 11844 32564 11854
rect 31836 11284 31892 11294
rect 31836 11190 31892 11228
rect 31612 10210 31668 10220
rect 31724 11170 31780 11182
rect 31724 11118 31726 11170
rect 31778 11118 31780 11170
rect 31724 10164 31780 11118
rect 32060 10388 32116 11732
rect 32396 11506 32452 11518
rect 32396 11454 32398 11506
rect 32450 11454 32452 11506
rect 32396 11394 32452 11454
rect 32396 11342 32398 11394
rect 32450 11342 32452 11394
rect 32396 11330 32452 11342
rect 32508 11060 32564 11788
rect 32060 10322 32116 10332
rect 32396 11004 32564 11060
rect 32620 11506 32676 11518
rect 32620 11454 32622 11506
rect 32674 11454 32676 11506
rect 32620 11394 32676 11454
rect 32620 11342 32622 11394
rect 32674 11342 32676 11394
rect 31724 10098 31780 10108
rect 32172 10164 32228 10174
rect 29932 9604 29988 9614
rect 29932 9602 30100 9604
rect 29932 9550 29934 9602
rect 29986 9550 30100 9602
rect 29932 9548 30100 9550
rect 29932 9538 29988 9548
rect 29596 9044 29652 9054
rect 29708 9044 29764 9324
rect 29596 9042 29764 9044
rect 29596 8990 29598 9042
rect 29650 8990 29764 9042
rect 29596 8988 29764 8990
rect 29596 8978 29652 8988
rect 29932 8484 29988 8494
rect 29036 7646 29038 7698
rect 29090 7646 29092 7698
rect 29036 7634 29092 7646
rect 29596 8372 29652 8382
rect 29596 7924 29652 8316
rect 29932 8258 29988 8428
rect 30044 8372 30100 9548
rect 30380 9602 30436 9614
rect 30380 9550 30382 9602
rect 30434 9550 30436 9602
rect 30268 8932 30324 8942
rect 30044 8306 30100 8316
rect 30156 8930 30324 8932
rect 30156 8878 30270 8930
rect 30322 8878 30324 8930
rect 30156 8876 30324 8878
rect 30156 8370 30212 8876
rect 30268 8866 30324 8876
rect 30156 8318 30158 8370
rect 30210 8318 30212 8370
rect 30156 8306 30212 8318
rect 30268 8484 30324 8494
rect 30268 8370 30324 8428
rect 30268 8318 30270 8370
rect 30322 8318 30324 8370
rect 30268 8306 30324 8318
rect 29932 8206 29934 8258
rect 29986 8206 29988 8258
rect 29932 8194 29988 8206
rect 29484 7476 29540 7486
rect 28588 6638 28590 6690
rect 28642 6638 28644 6690
rect 28588 6626 28644 6638
rect 28700 7362 28756 7374
rect 28700 7310 28702 7362
rect 28754 7310 28756 7362
rect 28700 6580 28756 7310
rect 29372 7364 29428 7374
rect 29372 7270 29428 7308
rect 28700 6356 28756 6524
rect 29148 6916 29204 6926
rect 29036 6468 29092 6478
rect 28700 6290 28756 6300
rect 28812 6466 29092 6468
rect 28812 6414 29038 6466
rect 29090 6414 29092 6466
rect 28812 6412 29092 6414
rect 28588 6244 28644 6254
rect 28476 6188 28588 6244
rect 28364 5854 28366 5906
rect 28418 5854 28420 5906
rect 28364 5842 28420 5854
rect 28588 5906 28644 6188
rect 28588 5854 28590 5906
rect 28642 5854 28644 5906
rect 28588 5842 28644 5854
rect 28588 5460 28644 5470
rect 28364 5124 28420 5134
rect 28252 5122 28420 5124
rect 28252 5070 28366 5122
rect 28418 5070 28420 5122
rect 28252 5068 28420 5070
rect 28140 4174 28142 4226
rect 28194 4174 28196 4226
rect 28140 4162 28196 4174
rect 27132 3390 27134 3442
rect 27186 3390 27188 3442
rect 27132 3378 27188 3390
rect 27356 3836 27524 3892
rect 27580 4060 27860 4116
rect 27356 3388 27412 3836
rect 27580 3554 27636 4060
rect 27580 3502 27582 3554
rect 27634 3502 27636 3554
rect 27356 3332 27524 3388
rect 27468 2996 27524 3332
rect 27468 2930 27524 2940
rect 27580 1876 27636 3502
rect 27916 4004 27972 4014
rect 27804 3330 27860 3342
rect 27804 3278 27806 3330
rect 27858 3278 27860 3330
rect 27804 2884 27860 3278
rect 27804 2818 27860 2828
rect 27580 1810 27636 1820
rect 27916 1764 27972 3948
rect 28364 4004 28420 5068
rect 28588 5010 28644 5404
rect 28588 4958 28590 5010
rect 28642 4958 28644 5010
rect 28588 4946 28644 4958
rect 28700 4340 28756 4350
rect 28700 4246 28756 4284
rect 28364 3938 28420 3948
rect 27804 1708 27972 1764
rect 28476 3668 28532 3678
rect 27020 1484 27300 1540
rect 27244 1316 27300 1484
rect 26908 1260 27188 1316
rect 27132 800 27188 1260
rect 27244 1250 27300 1260
rect 27804 800 27860 1708
rect 28476 800 28532 3612
rect 28588 3444 28644 3482
rect 28588 2548 28644 3388
rect 28588 2482 28644 2492
rect 28812 2436 28868 6412
rect 29036 6402 29092 6412
rect 29148 6244 29204 6860
rect 29260 6580 29316 6590
rect 29260 6486 29316 6524
rect 29372 6578 29428 6590
rect 29372 6526 29374 6578
rect 29426 6526 29428 6578
rect 29372 6468 29428 6526
rect 29372 6402 29428 6412
rect 29484 6244 29540 7420
rect 29596 7474 29652 7868
rect 29596 7422 29598 7474
rect 29650 7422 29652 7474
rect 29596 7410 29652 7422
rect 29708 8034 29764 8046
rect 29708 7982 29710 8034
rect 29762 7982 29764 8034
rect 29708 7476 29764 7982
rect 30380 7812 30436 9550
rect 31836 9602 31892 9614
rect 32172 9604 32228 10108
rect 32396 9826 32452 11004
rect 32508 10836 32564 10846
rect 32508 10742 32564 10780
rect 32396 9774 32398 9826
rect 32450 9774 32452 9826
rect 31836 9550 31838 9602
rect 31890 9550 31892 9602
rect 30156 7756 30436 7812
rect 30492 9380 30548 9390
rect 29932 7476 29988 7486
rect 29708 7474 29988 7476
rect 29708 7422 29934 7474
rect 29986 7422 29988 7474
rect 29708 7420 29988 7422
rect 29820 7252 29876 7262
rect 29708 6916 29764 6926
rect 28924 6188 29204 6244
rect 29260 6188 29540 6244
rect 29596 6860 29708 6916
rect 28924 6018 28980 6188
rect 29260 6130 29316 6188
rect 28924 5966 28926 6018
rect 28978 5966 28980 6018
rect 28924 5954 28980 5966
rect 29036 6074 29092 6086
rect 29036 6022 29038 6074
rect 29090 6022 29092 6074
rect 29260 6078 29262 6130
rect 29314 6078 29316 6130
rect 29036 6020 29092 6022
rect 29148 6020 29204 6030
rect 29036 5964 29148 6020
rect 29148 5954 29204 5964
rect 29260 5908 29316 6078
rect 29260 5842 29316 5852
rect 29372 6020 29428 6030
rect 29260 5684 29316 5694
rect 29148 5628 29260 5684
rect 28924 3330 28980 3342
rect 28924 3278 28926 3330
rect 28978 3278 28980 3330
rect 28924 2996 28980 3278
rect 28924 2930 28980 2940
rect 28812 2370 28868 2380
rect 29148 1652 29204 5628
rect 29260 5618 29316 5628
rect 29260 5124 29316 5134
rect 29260 5030 29316 5068
rect 29372 4676 29428 5964
rect 29484 6020 29540 6030
rect 29596 6020 29652 6860
rect 29708 6850 29764 6860
rect 29820 6690 29876 7196
rect 29820 6638 29822 6690
rect 29874 6638 29876 6690
rect 29708 6356 29764 6366
rect 29708 6132 29764 6300
rect 29708 6066 29764 6076
rect 29820 6130 29876 6638
rect 29820 6078 29822 6130
rect 29874 6078 29876 6130
rect 29820 6066 29876 6078
rect 29484 6018 29652 6020
rect 29484 5966 29486 6018
rect 29538 5966 29652 6018
rect 29484 5964 29652 5966
rect 29484 5954 29540 5964
rect 29708 5572 29764 5582
rect 29596 5348 29652 5358
rect 29596 5254 29652 5292
rect 29484 5124 29540 5134
rect 29708 5124 29764 5516
rect 29484 5122 29764 5124
rect 29484 5070 29486 5122
rect 29538 5070 29764 5122
rect 29484 5068 29764 5070
rect 29484 5058 29540 5068
rect 29932 5012 29988 7420
rect 30156 6580 30212 7756
rect 30268 7588 30324 7598
rect 30268 7586 30436 7588
rect 30268 7534 30270 7586
rect 30322 7534 30436 7586
rect 30268 7532 30436 7534
rect 30268 7522 30324 7532
rect 30156 6514 30212 6524
rect 30044 6468 30100 6478
rect 30044 5908 30100 6412
rect 30044 5842 30100 5852
rect 30156 5906 30212 5918
rect 30156 5854 30158 5906
rect 30210 5854 30212 5906
rect 30156 5684 30212 5854
rect 30268 5796 30324 5806
rect 30268 5702 30324 5740
rect 30156 5618 30212 5628
rect 30268 5348 30324 5358
rect 30268 5254 30324 5292
rect 30156 5124 30212 5134
rect 30156 5030 30212 5068
rect 29708 4956 29988 5012
rect 29372 4620 29652 4676
rect 29260 4450 29316 4462
rect 29260 4398 29262 4450
rect 29314 4398 29316 4450
rect 29260 3892 29316 4398
rect 29260 3826 29316 3836
rect 29260 3442 29316 3454
rect 29260 3390 29262 3442
rect 29314 3390 29316 3442
rect 29260 3332 29316 3390
rect 29596 3442 29652 4620
rect 29596 3390 29598 3442
rect 29650 3390 29652 3442
rect 29596 3378 29652 3390
rect 29260 2324 29316 3276
rect 29260 2258 29316 2268
rect 29148 1586 29204 1596
rect 29148 1426 29204 1438
rect 29148 1374 29150 1426
rect 29202 1374 29204 1426
rect 29148 800 29204 1374
rect 29708 1426 29764 4956
rect 30044 4900 30100 4910
rect 30044 4806 30100 4844
rect 30380 4340 30436 7532
rect 30492 6692 30548 9324
rect 31164 9268 31220 9278
rect 31164 8370 31220 9212
rect 31836 9268 31892 9550
rect 31836 9202 31892 9212
rect 32060 9602 32228 9604
rect 32060 9550 32174 9602
rect 32226 9550 32228 9602
rect 32060 9548 32228 9550
rect 31164 8318 31166 8370
rect 31218 8318 31220 8370
rect 31164 8306 31220 8318
rect 31948 8148 32004 8158
rect 32060 8148 32116 9548
rect 32172 9538 32228 9548
rect 32284 9602 32340 9614
rect 32284 9550 32286 9602
rect 32338 9550 32340 9602
rect 32284 8484 32340 9550
rect 32396 8930 32452 9774
rect 32620 9828 32676 11342
rect 32620 9714 32676 9772
rect 32620 9662 32622 9714
rect 32674 9662 32676 9714
rect 32620 9650 32676 9662
rect 32396 8878 32398 8930
rect 32450 8878 32452 8930
rect 32396 8866 32452 8878
rect 32508 9604 32564 9614
rect 32284 8418 32340 8428
rect 32396 8708 32452 8718
rect 31948 8146 32116 8148
rect 31948 8094 31950 8146
rect 32002 8094 32116 8146
rect 31948 8092 32116 8094
rect 32172 8258 32228 8270
rect 32396 8260 32452 8652
rect 32172 8206 32174 8258
rect 32226 8206 32228 8258
rect 31948 8082 32004 8092
rect 30828 8034 30884 8046
rect 30828 7982 30830 8034
rect 30882 7982 30884 8034
rect 30828 7812 30884 7982
rect 30492 6690 30660 6692
rect 30492 6638 30494 6690
rect 30546 6638 30660 6690
rect 30492 6636 30660 6638
rect 30492 6626 30548 6636
rect 30492 6132 30548 6142
rect 30492 6018 30548 6076
rect 30492 5966 30494 6018
rect 30546 5966 30548 6018
rect 30492 5348 30548 5966
rect 30492 5282 30548 5292
rect 30604 5012 30660 6636
rect 30828 6356 30884 7756
rect 31724 8034 31780 8046
rect 31724 7982 31726 8034
rect 31778 7982 31780 8034
rect 31276 7588 31332 7598
rect 31052 7532 31276 7588
rect 30940 7476 30996 7486
rect 30940 7382 30996 7420
rect 30828 5906 30884 6300
rect 30828 5854 30830 5906
rect 30882 5854 30884 5906
rect 30828 5842 30884 5854
rect 30940 6468 30996 6478
rect 30940 5346 30996 6412
rect 31052 6132 31108 7532
rect 31276 7494 31332 7532
rect 31724 7476 31780 7982
rect 32060 7588 32116 7598
rect 32060 7494 32116 7532
rect 31724 7410 31780 7420
rect 31836 7362 31892 7374
rect 31836 7310 31838 7362
rect 31890 7310 31892 7362
rect 31052 6066 31108 6076
rect 31164 6578 31220 6590
rect 31164 6526 31166 6578
rect 31218 6526 31220 6578
rect 31052 5908 31108 5918
rect 31052 5814 31108 5852
rect 31164 5684 31220 6526
rect 31388 6356 31444 6366
rect 31388 6130 31444 6300
rect 31836 6244 31892 7310
rect 32172 6356 32228 8206
rect 32284 8204 32452 8260
rect 32284 7586 32340 8204
rect 32284 7534 32286 7586
rect 32338 7534 32340 7586
rect 32284 7522 32340 7534
rect 32396 7364 32452 7374
rect 32508 7364 32564 9548
rect 32732 8932 32788 13804
rect 32844 13524 32900 15092
rect 32956 13748 33012 13758
rect 32956 13654 33012 13692
rect 32844 13458 32900 13468
rect 33068 12964 33124 15596
rect 33292 13188 33348 15708
rect 33404 15652 33460 15662
rect 33404 15538 33460 15596
rect 33404 15486 33406 15538
rect 33458 15486 33460 15538
rect 33404 15474 33460 15486
rect 33516 15538 33572 15932
rect 33516 15486 33518 15538
rect 33570 15486 33572 15538
rect 33516 15474 33572 15486
rect 33628 15314 33684 15326
rect 33628 15262 33630 15314
rect 33682 15262 33684 15314
rect 33404 14420 33460 14430
rect 33460 14364 33572 14420
rect 33404 14354 33460 14364
rect 33404 14084 33460 14094
rect 33404 13970 33460 14028
rect 33404 13918 33406 13970
rect 33458 13918 33460 13970
rect 33404 13906 33460 13918
rect 33516 13970 33572 14364
rect 33516 13918 33518 13970
rect 33570 13918 33572 13970
rect 33516 13906 33572 13918
rect 33628 13972 33684 15262
rect 33628 13878 33684 13916
rect 33292 13122 33348 13132
rect 33068 12908 33460 12964
rect 32956 11396 33012 11406
rect 32956 11302 33012 11340
rect 33068 11170 33124 11182
rect 33068 11118 33070 11170
rect 33122 11118 33124 11170
rect 32956 10164 33012 10174
rect 32956 9828 33012 10108
rect 33068 10052 33124 11118
rect 33180 11170 33236 11182
rect 33180 11118 33182 11170
rect 33234 11118 33236 11170
rect 33180 10164 33236 11118
rect 33180 10098 33236 10108
rect 33292 11172 33348 11182
rect 33292 10500 33348 11116
rect 33404 10724 33460 12908
rect 33628 12962 33684 12974
rect 33628 12910 33630 12962
rect 33682 12910 33684 12962
rect 33628 11394 33684 12910
rect 33740 11508 33796 17276
rect 33852 16884 33908 16894
rect 34188 16884 34244 17502
rect 34300 17556 34356 17566
rect 34300 17462 34356 17500
rect 34636 17554 34692 17566
rect 34636 17502 34638 17554
rect 34690 17502 34692 17554
rect 33852 16882 34244 16884
rect 33852 16830 33854 16882
rect 33906 16830 34244 16882
rect 33852 16828 34244 16830
rect 34300 16884 34356 16894
rect 34636 16884 34692 17502
rect 35644 17444 35700 17612
rect 35756 17668 35812 17678
rect 35868 17668 35924 19182
rect 35756 17666 36260 17668
rect 35756 17614 35758 17666
rect 35810 17614 36260 17666
rect 35756 17612 36260 17614
rect 35756 17602 35812 17612
rect 36092 17444 36148 17454
rect 35644 17388 36092 17444
rect 35980 17220 36036 17230
rect 35420 17108 35476 17118
rect 34300 16882 34692 16884
rect 34300 16830 34302 16882
rect 34354 16830 34692 16882
rect 34300 16828 34692 16830
rect 35308 17052 35420 17108
rect 33852 14868 33908 16828
rect 33852 14802 33908 14812
rect 34076 14084 34132 14094
rect 34076 13970 34132 14028
rect 34076 13918 34078 13970
rect 34130 13918 34132 13970
rect 34076 13906 34132 13918
rect 34300 13076 34356 16828
rect 35308 16772 35364 17052
rect 35420 17014 35476 17052
rect 35980 17106 36036 17164
rect 35980 17054 35982 17106
rect 36034 17054 36036 17106
rect 35980 17042 36036 17054
rect 36092 16994 36148 17388
rect 36092 16942 36094 16994
rect 36146 16942 36148 16994
rect 36092 16930 36148 16942
rect 36204 16996 36260 17612
rect 36316 17220 36372 19516
rect 36428 19506 36484 19516
rect 36428 19348 36484 19358
rect 36540 19348 36596 19964
rect 36428 19346 36596 19348
rect 36428 19294 36430 19346
rect 36482 19294 36596 19346
rect 36428 19292 36596 19294
rect 36428 19282 36484 19292
rect 36764 19012 36820 23548
rect 37100 21812 37156 23774
rect 37212 23826 37268 23884
rect 37212 23774 37214 23826
rect 37266 23774 37268 23826
rect 37212 23762 37268 23774
rect 37324 23884 37604 23940
rect 37772 24164 37828 24174
rect 37324 23154 37380 23884
rect 37660 23826 37716 23838
rect 37660 23774 37662 23826
rect 37714 23774 37716 23826
rect 37436 23716 37492 23726
rect 37436 23714 37604 23716
rect 37436 23662 37438 23714
rect 37490 23662 37604 23714
rect 37436 23660 37604 23662
rect 37436 23650 37492 23660
rect 37324 23102 37326 23154
rect 37378 23102 37380 23154
rect 37324 22482 37380 23102
rect 37324 22430 37326 22482
rect 37378 22430 37380 22482
rect 37324 22372 37380 22430
rect 37100 21756 37268 21812
rect 36988 20692 37044 20702
rect 36988 20598 37044 20636
rect 36764 18946 36820 18956
rect 36428 18900 36484 18910
rect 36428 17666 36484 18844
rect 36428 17614 36430 17666
rect 36482 17614 36484 17666
rect 36428 17602 36484 17614
rect 37100 17780 37156 17790
rect 36988 17556 37044 17566
rect 36988 17462 37044 17500
rect 36316 17154 36372 17164
rect 36988 17220 37044 17230
rect 35644 16884 35700 16894
rect 35644 16882 35812 16884
rect 35644 16830 35646 16882
rect 35698 16830 35812 16882
rect 35644 16828 35812 16830
rect 35644 16818 35700 16828
rect 35084 16716 35364 16772
rect 35084 15314 35140 16716
rect 35196 16492 35460 16502
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35196 16426 35460 16436
rect 35308 16212 35364 16222
rect 35644 16212 35700 16222
rect 35308 16210 35700 16212
rect 35308 16158 35310 16210
rect 35362 16158 35646 16210
rect 35698 16158 35700 16210
rect 35308 16156 35700 16158
rect 35308 16146 35364 16156
rect 35644 16146 35700 16156
rect 35756 16100 35812 16828
rect 36204 16882 36260 16940
rect 36988 16996 37044 17164
rect 36988 16902 37044 16940
rect 36204 16830 36206 16882
rect 36258 16830 36260 16882
rect 36204 16818 36260 16830
rect 36540 16884 36596 16894
rect 36540 16210 36596 16828
rect 37100 16772 37156 17724
rect 37212 17442 37268 21756
rect 37324 21476 37380 22316
rect 37436 22932 37492 22942
rect 37436 21698 37492 22876
rect 37436 21646 37438 21698
rect 37490 21646 37492 21698
rect 37436 21634 37492 21646
rect 37548 21586 37604 23660
rect 37660 23604 37716 23774
rect 37772 23828 37828 24108
rect 37772 23734 37828 23772
rect 37660 23538 37716 23548
rect 37660 23380 37716 23390
rect 37660 23154 37716 23324
rect 37660 23102 37662 23154
rect 37714 23102 37716 23154
rect 37660 23090 37716 23102
rect 37772 22372 37828 22382
rect 37772 22278 37828 22316
rect 37548 21534 37550 21586
rect 37602 21534 37604 21586
rect 37548 21522 37604 21534
rect 37324 21420 37492 21476
rect 37324 20580 37380 20590
rect 37324 19010 37380 20524
rect 37436 20020 37492 21420
rect 37884 21028 37940 24220
rect 38220 23938 38276 25788
rect 38332 25778 38388 25788
rect 38220 23886 38222 23938
rect 38274 23886 38276 23938
rect 38220 23874 38276 23886
rect 38332 25506 38388 25518
rect 38332 25454 38334 25506
rect 38386 25454 38388 25506
rect 37996 23716 38052 23726
rect 38332 23716 38388 25454
rect 37996 23714 38388 23716
rect 37996 23662 37998 23714
rect 38050 23662 38388 23714
rect 37996 23660 38388 23662
rect 37996 23650 38052 23660
rect 38444 23548 38500 25900
rect 38332 23492 38500 23548
rect 38108 23380 38164 23390
rect 37884 20972 38052 21028
rect 37884 20802 37940 20814
rect 37884 20750 37886 20802
rect 37938 20750 37940 20802
rect 37884 20132 37940 20750
rect 37996 20692 38052 20972
rect 38108 20914 38164 23324
rect 38332 22260 38388 23492
rect 38556 22932 38612 26126
rect 38668 25844 38724 26348
rect 38668 25778 38724 25788
rect 38780 26402 38836 26910
rect 39676 26908 39732 28028
rect 39900 28018 39956 28028
rect 40348 28084 40404 28094
rect 40348 27990 40404 28028
rect 40012 27412 40068 27422
rect 39788 27076 39844 27086
rect 39788 27074 39956 27076
rect 39788 27022 39790 27074
rect 39842 27022 39956 27074
rect 39788 27020 39956 27022
rect 39788 27010 39844 27020
rect 38780 26350 38782 26402
rect 38834 26350 38836 26402
rect 38780 25620 38836 26350
rect 39228 26852 39732 26908
rect 39228 26290 39284 26852
rect 39228 26238 39230 26290
rect 39282 26238 39284 26290
rect 39228 26226 39284 26238
rect 39788 26850 39844 26862
rect 39788 26798 39790 26850
rect 39842 26798 39844 26850
rect 38780 25554 38836 25564
rect 38892 26180 38948 26190
rect 38892 24388 38948 26124
rect 39452 25284 39508 25294
rect 39452 24946 39508 25228
rect 39452 24894 39454 24946
rect 39506 24894 39508 24946
rect 39452 24882 39508 24894
rect 39340 24724 39396 24734
rect 39340 24722 39620 24724
rect 39340 24670 39342 24722
rect 39394 24670 39620 24722
rect 39340 24668 39620 24670
rect 39340 24658 39396 24668
rect 38892 24322 38948 24332
rect 39452 24498 39508 24510
rect 39452 24446 39454 24498
rect 39506 24446 39508 24498
rect 39452 23938 39508 24446
rect 39452 23886 39454 23938
rect 39506 23886 39508 23938
rect 39452 23874 39508 23886
rect 39340 23716 39396 23726
rect 38556 22866 38612 22876
rect 38668 23714 39396 23716
rect 38668 23662 39342 23714
rect 39394 23662 39396 23714
rect 38668 23660 39396 23662
rect 38556 22708 38612 22718
rect 38332 22194 38388 22204
rect 38444 22652 38556 22708
rect 38108 20862 38110 20914
rect 38162 20862 38164 20914
rect 38108 20850 38164 20862
rect 38220 21810 38276 21822
rect 38220 21758 38222 21810
rect 38274 21758 38276 21810
rect 37996 20636 38164 20692
rect 37884 20066 37940 20076
rect 37660 20020 37716 20030
rect 37436 20018 37716 20020
rect 37436 19966 37662 20018
rect 37714 19966 37716 20018
rect 37436 19964 37716 19966
rect 37660 19954 37716 19964
rect 37996 20018 38052 20030
rect 37996 19966 37998 20018
rect 38050 19966 38052 20018
rect 37996 19796 38052 19966
rect 37996 19730 38052 19740
rect 38108 19346 38164 20636
rect 38108 19294 38110 19346
rect 38162 19294 38164 19346
rect 38108 19282 38164 19294
rect 37660 19236 37716 19246
rect 37660 19122 37716 19180
rect 37660 19070 37662 19122
rect 37714 19070 37716 19122
rect 37660 19058 37716 19070
rect 37996 19122 38052 19134
rect 37996 19070 37998 19122
rect 38050 19070 38052 19122
rect 37324 18958 37326 19010
rect 37378 18958 37380 19010
rect 37324 18900 37380 18958
rect 37324 18834 37380 18844
rect 37772 18340 37828 18350
rect 37436 18228 37492 18238
rect 37212 17390 37214 17442
rect 37266 17390 37268 17442
rect 37212 17378 37268 17390
rect 37324 17554 37380 17566
rect 37324 17502 37326 17554
rect 37378 17502 37380 17554
rect 37324 17444 37380 17502
rect 37324 17378 37380 17388
rect 37324 16996 37380 17006
rect 37436 16996 37492 18172
rect 37548 17554 37604 17566
rect 37548 17502 37550 17554
rect 37602 17502 37604 17554
rect 37548 17220 37604 17502
rect 37548 17154 37604 17164
rect 37772 17106 37828 18284
rect 37996 17890 38052 19070
rect 38220 18452 38276 21758
rect 38332 20690 38388 20702
rect 38332 20638 38334 20690
rect 38386 20638 38388 20690
rect 38332 19236 38388 20638
rect 38332 19142 38388 19180
rect 37996 17838 37998 17890
rect 38050 17838 38052 17890
rect 37996 17826 38052 17838
rect 38108 18396 38276 18452
rect 37772 17054 37774 17106
rect 37826 17054 37828 17106
rect 37772 17042 37828 17054
rect 37884 17668 37940 17678
rect 37324 16994 37492 16996
rect 37324 16942 37326 16994
rect 37378 16942 37492 16994
rect 37324 16940 37492 16942
rect 37324 16930 37380 16940
rect 37660 16884 37716 16894
rect 37548 16882 37716 16884
rect 37548 16830 37662 16882
rect 37714 16830 37716 16882
rect 37548 16828 37716 16830
rect 37548 16772 37604 16828
rect 37660 16818 37716 16828
rect 37100 16716 37492 16772
rect 36540 16158 36542 16210
rect 36594 16158 36596 16210
rect 36540 16146 36596 16158
rect 36764 16324 36820 16334
rect 35756 16044 35924 16100
rect 35868 15652 35924 16044
rect 35084 15262 35086 15314
rect 35138 15262 35140 15314
rect 34636 14642 34692 14654
rect 34636 14590 34638 14642
rect 34690 14590 34692 14642
rect 34636 13858 34692 14590
rect 35084 14644 35140 15262
rect 35644 15596 35924 15652
rect 35980 15986 36036 15998
rect 35980 15934 35982 15986
rect 36034 15934 36036 15986
rect 35980 15652 36036 15934
rect 35196 14924 35460 14934
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35196 14858 35460 14868
rect 35196 14644 35252 14654
rect 35084 14642 35252 14644
rect 35084 14590 35198 14642
rect 35250 14590 35252 14642
rect 35084 14588 35252 14590
rect 35196 14578 35252 14588
rect 35532 14308 35588 14318
rect 35532 14214 35588 14252
rect 34636 13806 34638 13858
rect 34690 13806 34692 13858
rect 34636 13794 34692 13806
rect 34972 14084 35028 14094
rect 34972 13858 35028 14028
rect 35308 13972 35364 13982
rect 35644 13972 35700 15596
rect 35980 15586 36036 15596
rect 35756 15316 35812 15326
rect 35756 14530 35812 15260
rect 35868 15202 35924 15214
rect 35868 15150 35870 15202
rect 35922 15150 35924 15202
rect 35868 14642 35924 15150
rect 35868 14590 35870 14642
rect 35922 14590 35924 14642
rect 35868 14578 35924 14590
rect 35756 14478 35758 14530
rect 35810 14478 35812 14530
rect 35756 14466 35812 14478
rect 35980 14306 36036 14318
rect 35980 14254 35982 14306
rect 36034 14254 36036 14306
rect 35980 13972 36036 14254
rect 36764 14308 36820 16268
rect 37436 16322 37492 16716
rect 37548 16706 37604 16716
rect 37436 16270 37438 16322
rect 37490 16270 37492 16322
rect 37436 16258 37492 16270
rect 37324 16212 37380 16222
rect 37324 15148 37380 16156
rect 37884 16210 37940 17612
rect 37996 16996 38052 17006
rect 37996 16324 38052 16940
rect 37996 16230 38052 16268
rect 37884 16158 37886 16210
rect 37938 16158 37940 16210
rect 37884 16146 37940 16158
rect 37212 15092 37380 15148
rect 37996 15204 38052 15242
rect 37996 15138 38052 15148
rect 37212 14642 37268 15092
rect 37996 14756 38052 14766
rect 37212 14590 37214 14642
rect 37266 14590 37268 14642
rect 37212 14578 37268 14590
rect 37884 14700 37996 14756
rect 36764 14242 36820 14252
rect 35364 13916 35588 13972
rect 35644 13916 35812 13972
rect 35308 13878 35364 13916
rect 34972 13806 34974 13858
rect 35026 13806 35028 13858
rect 34972 13794 35028 13806
rect 35196 13356 35460 13366
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35196 13290 35460 13300
rect 35532 13188 35588 13916
rect 35644 13748 35700 13758
rect 35644 13654 35700 13692
rect 34300 13010 34356 13020
rect 35308 13132 35588 13188
rect 34300 12852 34356 12862
rect 34300 12850 35252 12852
rect 34300 12798 34302 12850
rect 34354 12798 35252 12850
rect 34300 12796 35252 12798
rect 34300 12786 34356 12796
rect 34636 12404 34692 12414
rect 34636 12178 34692 12348
rect 35084 12404 35140 12414
rect 35084 12310 35140 12348
rect 35196 12402 35252 12796
rect 35196 12350 35198 12402
rect 35250 12350 35252 12402
rect 35196 12338 35252 12350
rect 35308 12402 35364 13132
rect 35308 12350 35310 12402
rect 35362 12350 35364 12402
rect 35308 12338 35364 12350
rect 35756 12402 35812 13916
rect 35980 13906 36036 13916
rect 37660 13860 37716 13870
rect 37660 13746 37716 13804
rect 37660 13694 37662 13746
rect 37714 13694 37716 13746
rect 36988 13300 37044 13310
rect 36428 13076 36484 13086
rect 36428 12982 36484 13020
rect 35756 12350 35758 12402
rect 35810 12350 35812 12402
rect 35756 12338 35812 12350
rect 35644 12292 35700 12302
rect 35644 12198 35700 12236
rect 36204 12292 36260 12302
rect 36204 12198 36260 12236
rect 34636 12126 34638 12178
rect 34690 12126 34692 12178
rect 34636 12114 34692 12126
rect 36988 11956 37044 13244
rect 37436 12852 37492 12862
rect 37660 12852 37716 13694
rect 37772 13858 37828 13870
rect 37772 13806 37774 13858
rect 37826 13806 37828 13858
rect 37772 13300 37828 13806
rect 37772 13234 37828 13244
rect 37772 13076 37828 13086
rect 37884 13076 37940 14700
rect 37996 14690 38052 14700
rect 37996 13748 38052 13758
rect 37996 13654 38052 13692
rect 37884 13020 38052 13076
rect 37772 12982 37828 13020
rect 37436 12850 37716 12852
rect 37436 12798 37438 12850
rect 37490 12798 37716 12850
rect 37436 12796 37716 12798
rect 37884 12852 37940 12862
rect 37436 12786 37492 12796
rect 36988 11890 37044 11900
rect 37100 12738 37156 12750
rect 37100 12686 37102 12738
rect 37154 12686 37156 12738
rect 37100 12628 37156 12686
rect 35196 11788 35460 11798
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35196 11722 35460 11732
rect 33740 11442 33796 11452
rect 36428 11620 36484 11630
rect 36428 11506 36484 11564
rect 36428 11454 36430 11506
rect 36482 11454 36484 11506
rect 33628 11342 33630 11394
rect 33682 11342 33684 11394
rect 33516 10724 33572 10734
rect 33404 10668 33516 10724
rect 33516 10658 33572 10668
rect 33628 10500 33684 11342
rect 36428 11396 36484 11454
rect 36428 11330 36484 11340
rect 37100 11394 37156 12572
rect 37884 12738 37940 12796
rect 37884 12686 37886 12738
rect 37938 12686 37940 12738
rect 37884 12404 37940 12686
rect 37884 12338 37940 12348
rect 37548 12180 37604 12190
rect 37996 12180 38052 13020
rect 37100 11342 37102 11394
rect 37154 11342 37156 11394
rect 37100 11330 37156 11342
rect 37212 12066 37268 12078
rect 37212 12014 37214 12066
rect 37266 12014 37268 12066
rect 34300 11284 34356 11294
rect 34188 11282 34356 11284
rect 34188 11230 34302 11282
rect 34354 11230 34356 11282
rect 34188 11228 34356 11230
rect 34076 10500 34132 10510
rect 33628 10498 34132 10500
rect 33628 10446 34078 10498
rect 34130 10446 34132 10498
rect 33628 10444 34132 10446
rect 33068 9986 33124 9996
rect 33068 9828 33124 9838
rect 32956 9826 33124 9828
rect 32956 9774 33070 9826
rect 33122 9774 33124 9826
rect 32956 9772 33124 9774
rect 33068 9762 33124 9772
rect 33292 9826 33348 10444
rect 33964 10052 34020 10062
rect 33964 9958 34020 9996
rect 33292 9774 33294 9826
rect 33346 9774 33348 9826
rect 33292 9762 33348 9774
rect 33516 9828 33572 9838
rect 33180 9716 33236 9726
rect 33180 9622 33236 9660
rect 33516 9714 33572 9772
rect 33516 9662 33518 9714
rect 33570 9662 33572 9714
rect 33292 9380 33348 9390
rect 32732 8866 32788 8876
rect 32956 9268 33012 9278
rect 32956 9044 33012 9212
rect 33180 9044 33236 9054
rect 32956 9042 33236 9044
rect 32956 8990 33182 9042
rect 33234 8990 33236 9042
rect 32956 8988 33236 8990
rect 32956 8258 33012 8988
rect 33180 8978 33236 8988
rect 33292 8260 33348 9324
rect 33516 9266 33572 9662
rect 33516 9214 33518 9266
rect 33570 9214 33572 9266
rect 33516 9202 33572 9214
rect 34076 9044 34132 10444
rect 34188 9938 34244 11228
rect 34300 11218 34356 11228
rect 37212 10948 37268 12014
rect 37212 10882 37268 10892
rect 37324 11170 37380 11182
rect 37324 11118 37326 11170
rect 37378 11118 37380 11170
rect 36988 10836 37044 10846
rect 36988 10610 37044 10780
rect 36988 10558 36990 10610
rect 37042 10558 37044 10610
rect 36988 10546 37044 10558
rect 35196 10220 35460 10230
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35196 10154 35460 10164
rect 35756 10052 35812 10062
rect 35756 9958 35812 9996
rect 34188 9886 34190 9938
rect 34242 9886 34244 9938
rect 34188 9874 34244 9886
rect 34972 9938 35028 9950
rect 34972 9886 34974 9938
rect 35026 9886 35028 9938
rect 34636 9714 34692 9726
rect 34636 9662 34638 9714
rect 34690 9662 34692 9714
rect 34188 9602 34244 9614
rect 34188 9550 34190 9602
rect 34242 9550 34244 9602
rect 34188 9492 34244 9550
rect 34188 9426 34244 9436
rect 34188 9044 34244 9054
rect 34076 9042 34244 9044
rect 34076 8990 34190 9042
rect 34242 8990 34244 9042
rect 34076 8988 34244 8990
rect 32956 8206 32958 8258
rect 33010 8206 33012 8258
rect 32956 8194 33012 8206
rect 33180 8204 33348 8260
rect 33852 8260 33908 8270
rect 32396 7362 32564 7364
rect 32396 7310 32398 7362
rect 32450 7310 32564 7362
rect 32396 7308 32564 7310
rect 32956 7476 33012 7486
rect 32396 7298 32452 7308
rect 32172 6290 32228 6300
rect 31836 6188 32004 6244
rect 31388 6078 31390 6130
rect 31442 6078 31444 6130
rect 31388 6066 31444 6078
rect 31836 6018 31892 6030
rect 31836 5966 31838 6018
rect 31890 5966 31892 6018
rect 31836 5796 31892 5966
rect 31836 5730 31892 5740
rect 31724 5684 31780 5694
rect 31164 5682 31780 5684
rect 31164 5630 31726 5682
rect 31778 5630 31780 5682
rect 31164 5628 31780 5630
rect 31724 5618 31780 5628
rect 30940 5294 30942 5346
rect 30994 5294 30996 5346
rect 30940 5282 30996 5294
rect 31276 5348 31332 5358
rect 31052 5236 31108 5246
rect 30604 4946 30660 4956
rect 30716 5124 30772 5134
rect 30716 5010 30772 5068
rect 30828 5124 30884 5134
rect 31052 5124 31108 5180
rect 30828 5122 31108 5124
rect 30828 5070 30830 5122
rect 30882 5070 31108 5122
rect 30828 5068 31108 5070
rect 31276 5124 31332 5292
rect 31836 5348 31892 5358
rect 31836 5234 31892 5292
rect 31836 5182 31838 5234
rect 31890 5182 31892 5234
rect 31836 5170 31892 5182
rect 30828 5058 30884 5068
rect 31276 5030 31332 5068
rect 31948 5012 32004 6188
rect 32172 6132 32228 6142
rect 32060 6076 32172 6132
rect 32060 6018 32116 6076
rect 32172 6066 32228 6076
rect 32060 5966 32062 6018
rect 32114 5966 32116 6018
rect 32060 5954 32116 5966
rect 32620 5908 32676 5918
rect 32620 5814 32676 5852
rect 30716 4958 30718 5010
rect 30770 4958 30772 5010
rect 30716 4946 30772 4958
rect 31836 4956 32004 5012
rect 32172 5796 32228 5806
rect 30940 4788 30996 4798
rect 30828 4732 30940 4788
rect 30716 4340 30772 4350
rect 30380 4338 30772 4340
rect 30380 4286 30718 4338
rect 30770 4286 30772 4338
rect 30380 4284 30772 4286
rect 30716 4274 30772 4284
rect 30044 4116 30100 4126
rect 29932 3556 29988 3566
rect 29932 3442 29988 3500
rect 29932 3390 29934 3442
rect 29986 3390 29988 3442
rect 29932 3108 29988 3390
rect 29932 3042 29988 3052
rect 30044 1764 30100 4060
rect 30268 3780 30324 3790
rect 30268 3442 30324 3724
rect 30716 3556 30772 3566
rect 30828 3556 30884 4732
rect 30940 4722 30996 4732
rect 31836 4788 31892 4956
rect 31836 4722 31892 4732
rect 31276 4452 31332 4462
rect 31276 4358 31332 4396
rect 31388 4340 31444 4350
rect 30716 3554 30884 3556
rect 30716 3502 30718 3554
rect 30770 3502 30884 3554
rect 30716 3500 30884 3502
rect 30940 4116 30996 4126
rect 30716 3490 30772 3500
rect 30268 3390 30270 3442
rect 30322 3390 30324 3442
rect 30268 3378 30324 3390
rect 30940 3442 30996 4060
rect 30940 3390 30942 3442
rect 30994 3390 30996 3442
rect 30940 3378 30996 3390
rect 31164 3668 31220 3678
rect 29708 1374 29710 1426
rect 29762 1374 29764 1426
rect 29708 1362 29764 1374
rect 29820 1708 30100 1764
rect 30492 2772 30548 2782
rect 29820 800 29876 1708
rect 30492 800 30548 2716
rect 31164 800 31220 3612
rect 31388 3554 31444 4284
rect 31836 4228 31892 4238
rect 31836 4134 31892 4172
rect 31388 3502 31390 3554
rect 31442 3502 31444 3554
rect 31388 3490 31444 3502
rect 31836 4004 31892 4014
rect 31612 3332 31668 3342
rect 31612 3238 31668 3276
rect 31836 800 31892 3948
rect 32172 3442 32228 5740
rect 32620 5460 32676 5470
rect 32396 5122 32452 5134
rect 32396 5070 32398 5122
rect 32450 5070 32452 5122
rect 32396 4340 32452 5070
rect 32620 5122 32676 5404
rect 32620 5070 32622 5122
rect 32674 5070 32676 5122
rect 32620 5058 32676 5070
rect 32732 5010 32788 5022
rect 32732 4958 32734 5010
rect 32786 4958 32788 5010
rect 32396 4274 32452 4284
rect 32508 4676 32564 4686
rect 32508 3666 32564 4620
rect 32732 4564 32788 4958
rect 32732 4498 32788 4508
rect 32508 3614 32510 3666
rect 32562 3614 32564 3666
rect 32508 3602 32564 3614
rect 32172 3390 32174 3442
rect 32226 3390 32228 3442
rect 32172 1652 32228 3390
rect 32956 3388 33012 7420
rect 33068 7474 33124 7486
rect 33068 7422 33070 7474
rect 33122 7422 33124 7474
rect 33068 6356 33124 7422
rect 33180 6804 33236 8204
rect 33852 8166 33908 8204
rect 33292 8034 33348 8046
rect 33292 7982 33294 8034
rect 33346 7982 33348 8034
rect 33292 7924 33348 7982
rect 33292 7858 33348 7868
rect 33404 8036 33460 8046
rect 33404 7698 33460 7980
rect 34188 7812 34244 8988
rect 34636 8370 34692 9662
rect 34860 9604 34916 9614
rect 34860 9510 34916 9548
rect 34972 9154 35028 9886
rect 35868 9828 35924 9838
rect 36204 9828 36260 9838
rect 35868 9826 36204 9828
rect 35868 9774 35870 9826
rect 35922 9774 36204 9826
rect 35868 9772 36204 9774
rect 35868 9762 35924 9772
rect 36204 9734 36260 9772
rect 37324 9828 37380 11118
rect 37436 10612 37492 10622
rect 37436 10050 37492 10556
rect 37436 9998 37438 10050
rect 37490 9998 37492 10050
rect 37436 9986 37492 9998
rect 37324 9734 37380 9772
rect 36540 9716 36596 9726
rect 36540 9622 36596 9660
rect 34972 9102 34974 9154
rect 35026 9102 35028 9154
rect 34972 9090 35028 9102
rect 35756 9602 35812 9614
rect 36316 9604 36372 9614
rect 35756 9550 35758 9602
rect 35810 9550 35812 9602
rect 34636 8318 34638 8370
rect 34690 8318 34692 8370
rect 34636 8306 34692 8318
rect 34748 8820 34804 8830
rect 34748 8258 34804 8764
rect 35196 8652 35460 8662
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35196 8586 35460 8596
rect 34748 8206 34750 8258
rect 34802 8206 34804 8258
rect 34748 8194 34804 8206
rect 35420 8260 35476 8270
rect 35756 8260 35812 9550
rect 36204 9602 36372 9604
rect 36204 9550 36318 9602
rect 36370 9550 36372 9602
rect 36204 9548 36372 9550
rect 34300 8148 34356 8158
rect 34300 8054 34356 8092
rect 35420 8146 35476 8204
rect 35420 8094 35422 8146
rect 35474 8094 35476 8146
rect 34524 8036 34580 8046
rect 34580 7980 34692 8036
rect 34524 7942 34580 7980
rect 33404 7646 33406 7698
rect 33458 7646 33460 7698
rect 33292 6804 33348 6814
rect 33180 6802 33348 6804
rect 33180 6750 33294 6802
rect 33346 6750 33348 6802
rect 33180 6748 33348 6750
rect 33068 6290 33124 6300
rect 33180 6132 33236 6142
rect 33180 6038 33236 6076
rect 33292 6130 33348 6748
rect 33292 6078 33294 6130
rect 33346 6078 33348 6130
rect 33292 6066 33348 6078
rect 33404 6580 33460 7646
rect 33964 7756 34580 7812
rect 33740 7476 33796 7486
rect 33740 7382 33796 7420
rect 33964 6804 34020 7756
rect 33068 5908 33124 5918
rect 33404 5908 33460 6524
rect 33068 5906 33460 5908
rect 33068 5854 33070 5906
rect 33122 5854 33460 5906
rect 33068 5852 33460 5854
rect 33516 6748 34020 6804
rect 34076 7586 34132 7598
rect 34076 7534 34078 7586
rect 34130 7534 34132 7586
rect 33068 5842 33124 5852
rect 33516 5012 33572 6748
rect 33740 6580 33796 6590
rect 33740 6486 33796 6524
rect 33964 6580 34020 6590
rect 33964 6486 34020 6524
rect 33852 6468 33908 6478
rect 33852 6374 33908 6412
rect 34076 6468 34132 7534
rect 34524 7474 34580 7756
rect 34524 7422 34526 7474
rect 34578 7422 34580 7474
rect 34524 7410 34580 7422
rect 34412 7364 34468 7374
rect 34412 6916 34468 7308
rect 34412 6860 34580 6916
rect 34076 6402 34132 6412
rect 34412 6690 34468 6702
rect 34412 6638 34414 6690
rect 34466 6638 34468 6690
rect 34412 6580 34468 6638
rect 33740 6132 33796 6142
rect 33740 5906 33796 6076
rect 34412 6132 34468 6524
rect 34412 6066 34468 6076
rect 33740 5854 33742 5906
rect 33794 5854 33796 5906
rect 33740 5842 33796 5854
rect 34412 5906 34468 5918
rect 34412 5854 34414 5906
rect 34466 5854 34468 5906
rect 34188 5794 34244 5806
rect 34188 5742 34190 5794
rect 34242 5742 34244 5794
rect 33404 4340 33460 4350
rect 33516 4340 33572 4956
rect 33404 4338 33572 4340
rect 33404 4286 33406 4338
rect 33458 4286 33572 4338
rect 33404 4284 33572 4286
rect 33740 5684 33796 5694
rect 34188 5684 34244 5742
rect 34300 5684 34356 5694
rect 34188 5628 34300 5684
rect 33404 4274 33460 4284
rect 33628 4228 33684 4238
rect 33628 3442 33684 4172
rect 33628 3390 33630 3442
rect 33682 3390 33684 3442
rect 32956 3332 33236 3388
rect 33628 3378 33684 3390
rect 32172 1586 32228 1596
rect 32508 2660 32564 2670
rect 32508 800 32564 2604
rect 33180 800 33236 3332
rect 33740 1428 33796 5628
rect 34300 5618 34356 5628
rect 34412 5572 34468 5854
rect 34524 5794 34580 6860
rect 34636 6690 34692 7980
rect 34972 8034 35028 8046
rect 34972 7982 34974 8034
rect 35026 7982 35028 8034
rect 34972 7924 35028 7982
rect 34636 6638 34638 6690
rect 34690 6638 34692 6690
rect 34636 6626 34692 6638
rect 34860 7252 34916 7262
rect 34860 6690 34916 7196
rect 34860 6638 34862 6690
rect 34914 6638 34916 6690
rect 34860 6626 34916 6638
rect 34972 6580 35028 7868
rect 35308 7476 35364 7486
rect 35196 7474 35364 7476
rect 35196 7422 35310 7474
rect 35362 7422 35364 7474
rect 35196 7420 35364 7422
rect 35196 7364 35252 7420
rect 35308 7410 35364 7420
rect 35196 7298 35252 7308
rect 35420 7364 35476 8094
rect 35420 7298 35476 7308
rect 35532 8204 35812 8260
rect 35868 8932 35924 8942
rect 35532 7252 35588 8204
rect 35756 8036 35812 8046
rect 35532 7186 35588 7196
rect 35644 8034 35812 8036
rect 35644 7982 35758 8034
rect 35810 7982 35812 8034
rect 35644 7980 35812 7982
rect 35196 7084 35460 7094
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35196 7018 35460 7028
rect 35084 6580 35140 6590
rect 35028 6578 35140 6580
rect 35028 6526 35086 6578
rect 35138 6526 35140 6578
rect 35028 6524 35140 6526
rect 34972 6486 35028 6524
rect 35084 6514 35140 6524
rect 34748 6466 34804 6478
rect 34748 6414 34750 6466
rect 34802 6414 34804 6466
rect 34748 6018 34804 6414
rect 35196 6130 35252 6142
rect 35196 6078 35198 6130
rect 35250 6078 35252 6130
rect 34748 5966 34750 6018
rect 34802 5966 34804 6018
rect 34748 5954 34804 5966
rect 35084 6020 35140 6030
rect 35084 5906 35140 5964
rect 35084 5854 35086 5906
rect 35138 5854 35140 5906
rect 35084 5842 35140 5854
rect 34524 5742 34526 5794
rect 34578 5742 34580 5794
rect 34524 5730 34580 5742
rect 35196 5684 35252 6078
rect 35644 6018 35700 7980
rect 35756 7970 35812 7980
rect 35868 7588 35924 8876
rect 36092 8146 36148 8158
rect 36092 8094 36094 8146
rect 36146 8094 36148 8146
rect 36092 7700 36148 8094
rect 36092 7634 36148 7644
rect 35644 5966 35646 6018
rect 35698 5966 35700 6018
rect 35644 5954 35700 5966
rect 35756 7364 35812 7374
rect 34412 5506 34468 5516
rect 35084 5628 35252 5684
rect 34076 5236 34132 5246
rect 33740 1362 33796 1372
rect 33852 5124 33908 5134
rect 33852 800 33908 5068
rect 33964 4898 34020 4910
rect 33964 4846 33966 4898
rect 34018 4846 34020 4898
rect 33964 3554 34020 4846
rect 34076 4450 34132 5180
rect 34076 4398 34078 4450
rect 34130 4398 34132 4450
rect 34076 4386 34132 4398
rect 33964 3502 33966 3554
rect 34018 3502 34020 3554
rect 33964 3490 34020 3502
rect 35084 4228 35140 5628
rect 35196 5516 35460 5526
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35196 5450 35460 5460
rect 35084 3554 35140 4172
rect 35196 3948 35460 3958
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35196 3882 35460 3892
rect 35084 3502 35086 3554
rect 35138 3502 35140 3554
rect 35084 3490 35140 3502
rect 34972 3444 35028 3454
rect 35308 3444 35364 3482
rect 34972 3332 35252 3388
rect 35308 3378 35364 3388
rect 35756 3388 35812 7308
rect 35868 6690 35924 7532
rect 35868 6638 35870 6690
rect 35922 6638 35924 6690
rect 35868 6626 35924 6638
rect 36204 6692 36260 9548
rect 36316 9538 36372 9548
rect 37436 9602 37492 9614
rect 37436 9550 37438 9602
rect 37490 9550 37492 9602
rect 37436 9268 37492 9550
rect 37212 9212 37492 9268
rect 37100 8932 37156 8942
rect 37212 8932 37268 9212
rect 37436 9044 37492 9054
rect 37548 9044 37604 12124
rect 37772 12124 38052 12180
rect 37772 11618 37828 12124
rect 37772 11566 37774 11618
rect 37826 11566 37828 11618
rect 37772 11554 37828 11566
rect 38108 11396 38164 18396
rect 38444 18340 38500 22652
rect 38556 22642 38612 22652
rect 38556 20690 38612 20702
rect 38556 20638 38558 20690
rect 38610 20638 38612 20690
rect 38556 19236 38612 20638
rect 38556 19142 38612 19180
rect 38332 18338 38500 18340
rect 38332 18286 38446 18338
rect 38498 18286 38500 18338
rect 38332 18284 38500 18286
rect 38332 17108 38388 18284
rect 38444 18274 38500 18284
rect 38444 17554 38500 17566
rect 38444 17502 38446 17554
rect 38498 17502 38500 17554
rect 38444 17108 38500 17502
rect 38556 17444 38612 17454
rect 38556 17350 38612 17388
rect 38668 17332 38724 23660
rect 39340 23650 39396 23660
rect 39452 23604 39508 23614
rect 39340 23268 39396 23278
rect 39004 22370 39060 22382
rect 39004 22318 39006 22370
rect 39058 22318 39060 22370
rect 39004 22036 39060 22318
rect 39004 21970 39060 21980
rect 39228 21586 39284 21598
rect 39228 21534 39230 21586
rect 39282 21534 39284 21586
rect 39228 21476 39284 21534
rect 39228 21410 39284 21420
rect 39004 20804 39060 20814
rect 39004 20690 39060 20748
rect 39340 20802 39396 23212
rect 39452 23042 39508 23548
rect 39452 22990 39454 23042
rect 39506 22990 39508 23042
rect 39452 22258 39508 22990
rect 39452 22206 39454 22258
rect 39506 22206 39508 22258
rect 39452 21698 39508 22206
rect 39452 21646 39454 21698
rect 39506 21646 39508 21698
rect 39452 21634 39508 21646
rect 39340 20750 39342 20802
rect 39394 20750 39396 20802
rect 39340 20738 39396 20750
rect 39004 20638 39006 20690
rect 39058 20638 39060 20690
rect 39004 20626 39060 20638
rect 39564 20468 39620 24668
rect 39788 24052 39844 26798
rect 39900 26292 39956 27020
rect 39900 26178 39956 26236
rect 39900 26126 39902 26178
rect 39954 26126 39956 26178
rect 39900 26114 39956 26126
rect 40012 25282 40068 27356
rect 40684 27074 40740 28700
rect 40908 28690 40964 28700
rect 41468 28084 41524 28094
rect 40684 27022 40686 27074
rect 40738 27022 40740 27074
rect 40684 27010 40740 27022
rect 41020 27858 41076 27870
rect 41020 27806 41022 27858
rect 41074 27806 41076 27858
rect 41020 27074 41076 27806
rect 41468 27858 41524 28028
rect 41468 27806 41470 27858
rect 41522 27806 41524 27858
rect 41468 27794 41524 27806
rect 41020 27022 41022 27074
rect 41074 27022 41076 27074
rect 40572 26964 40628 27002
rect 40572 26898 40628 26908
rect 40348 26290 40404 26302
rect 40348 26238 40350 26290
rect 40402 26238 40404 26290
rect 40348 25732 40404 26238
rect 41020 26292 41076 27022
rect 41356 27746 41412 27758
rect 41692 27748 41748 38780
rect 41356 27694 41358 27746
rect 41410 27694 41412 27746
rect 41020 26198 41076 26236
rect 41132 26850 41188 26862
rect 41132 26798 41134 26850
rect 41186 26798 41188 26850
rect 40348 25666 40404 25676
rect 40348 25508 40404 25518
rect 40348 25414 40404 25452
rect 40012 25230 40014 25282
rect 40066 25230 40068 25282
rect 40012 25218 40068 25230
rect 40236 25396 40292 25406
rect 40236 25284 40292 25340
rect 40460 25394 40516 25406
rect 40460 25342 40462 25394
rect 40514 25342 40516 25394
rect 40236 25228 40404 25284
rect 40348 24946 40404 25228
rect 40348 24894 40350 24946
rect 40402 24894 40404 24946
rect 40348 24882 40404 24894
rect 39788 23986 39844 23996
rect 40124 24722 40180 24734
rect 40124 24670 40126 24722
rect 40178 24670 40180 24722
rect 40124 23268 40180 24670
rect 40348 23938 40404 23950
rect 40348 23886 40350 23938
rect 40402 23886 40404 23938
rect 40348 23716 40404 23886
rect 40348 23650 40404 23660
rect 40460 23826 40516 25342
rect 40908 24724 40964 24734
rect 40460 23774 40462 23826
rect 40514 23774 40516 23826
rect 40460 23604 40516 23774
rect 40460 23538 40516 23548
rect 40796 24722 40964 24724
rect 40796 24670 40910 24722
rect 40962 24670 40964 24722
rect 40796 24668 40964 24670
rect 40124 23202 40180 23212
rect 39788 23154 39844 23166
rect 39788 23102 39790 23154
rect 39842 23102 39844 23154
rect 39788 22372 39844 23102
rect 40348 23044 40404 23054
rect 40796 23044 40852 24668
rect 40908 24658 40964 24668
rect 41020 24052 41076 24062
rect 40908 23156 40964 23166
rect 40908 23062 40964 23100
rect 40348 23042 40852 23044
rect 40348 22990 40350 23042
rect 40402 22990 40852 23042
rect 40348 22988 40852 22990
rect 40348 22708 40404 22988
rect 40348 22642 40404 22652
rect 40908 22708 40964 22718
rect 39788 21924 39844 22316
rect 40572 22484 40628 22494
rect 40572 22146 40628 22428
rect 40572 22094 40574 22146
rect 40626 22094 40628 22146
rect 40572 22082 40628 22094
rect 39788 21858 39844 21868
rect 40348 21924 40404 21934
rect 40124 20804 40180 20814
rect 40012 20692 40068 20702
rect 40012 20598 40068 20636
rect 39676 20580 39732 20590
rect 39676 20486 39732 20524
rect 39564 20402 39620 20412
rect 38780 20244 38836 20254
rect 38780 20130 38836 20188
rect 39676 20242 39732 20254
rect 39676 20190 39678 20242
rect 39730 20190 39732 20242
rect 39676 20188 39732 20190
rect 39676 20132 39844 20188
rect 38780 20078 38782 20130
rect 38834 20078 38836 20130
rect 38780 20066 38836 20078
rect 39340 20020 39396 20030
rect 39676 20020 39732 20030
rect 39004 20018 39396 20020
rect 39004 19966 39342 20018
rect 39394 19966 39396 20018
rect 39004 19964 39396 19966
rect 38780 19234 38836 19246
rect 38780 19182 38782 19234
rect 38834 19182 38836 19234
rect 38780 17780 38836 19182
rect 39004 18340 39060 19964
rect 39340 19954 39396 19964
rect 39564 20018 39732 20020
rect 39564 19966 39678 20018
rect 39730 19966 39732 20018
rect 39564 19964 39732 19966
rect 39564 19460 39620 19964
rect 39676 19954 39732 19964
rect 39788 19796 39844 20132
rect 39228 19404 39620 19460
rect 39676 19740 39844 19796
rect 39900 20018 39956 20030
rect 39900 19966 39902 20018
rect 39954 19966 39956 20018
rect 39228 19348 39284 19404
rect 39228 19234 39284 19292
rect 39228 19182 39230 19234
rect 39282 19182 39284 19234
rect 39228 19170 39284 19182
rect 39340 19236 39396 19246
rect 39340 19142 39396 19180
rect 39564 19124 39620 19134
rect 39116 19012 39172 19022
rect 39116 18918 39172 18956
rect 39004 18274 39060 18284
rect 38780 17714 38836 17724
rect 39004 17668 39060 17678
rect 39564 17668 39620 19068
rect 39676 18116 39732 19740
rect 39900 19236 39956 19966
rect 39956 19180 40068 19236
rect 39900 19170 39956 19180
rect 39676 18050 39732 18060
rect 39788 19010 39844 19022
rect 39788 18958 39790 19010
rect 39842 18958 39844 19010
rect 39004 17574 39060 17612
rect 39452 17612 39620 17668
rect 39788 17668 39844 18958
rect 40012 18674 40068 19180
rect 40124 19124 40180 20748
rect 40348 20690 40404 21868
rect 40348 20638 40350 20690
rect 40402 20638 40404 20690
rect 40348 20626 40404 20638
rect 40460 20692 40516 20702
rect 40460 20188 40516 20636
rect 40908 20692 40964 22652
rect 40908 20626 40964 20636
rect 40348 20132 40516 20188
rect 40572 20580 40628 20590
rect 40124 19122 40292 19124
rect 40124 19070 40126 19122
rect 40178 19070 40292 19122
rect 40124 19068 40292 19070
rect 40124 19058 40180 19068
rect 40012 18622 40014 18674
rect 40066 18622 40068 18674
rect 40012 18610 40068 18622
rect 40236 18450 40292 19068
rect 40348 18676 40404 20132
rect 40572 19236 40628 20524
rect 40684 20578 40740 20590
rect 40684 20526 40686 20578
rect 40738 20526 40740 20578
rect 40684 20468 40740 20526
rect 40684 20402 40740 20412
rect 40572 19170 40628 19180
rect 40684 20020 40740 20030
rect 40460 19124 40516 19134
rect 40460 19030 40516 19068
rect 40572 19010 40628 19022
rect 40572 18958 40574 19010
rect 40626 18958 40628 19010
rect 40572 18900 40628 18958
rect 40572 18834 40628 18844
rect 40348 18620 40516 18676
rect 40236 18398 40238 18450
rect 40290 18398 40292 18450
rect 40236 18228 40292 18398
rect 40236 18162 40292 18172
rect 38780 17556 38836 17566
rect 39340 17556 39396 17566
rect 38780 17462 38836 17500
rect 39116 17554 39396 17556
rect 39116 17502 39342 17554
rect 39394 17502 39396 17554
rect 39116 17500 39396 17502
rect 38668 17276 38836 17332
rect 38780 17220 38836 17276
rect 38780 17164 38948 17220
rect 38668 17108 38724 17118
rect 38444 17106 38724 17108
rect 38444 17054 38670 17106
rect 38722 17054 38724 17106
rect 38444 17052 38724 17054
rect 38220 16882 38276 16894
rect 38220 16830 38222 16882
rect 38274 16830 38276 16882
rect 38220 15988 38276 16830
rect 38332 16884 38388 17052
rect 38668 17042 38724 17052
rect 38780 16996 38836 17006
rect 38780 16902 38836 16940
rect 38556 16884 38612 16894
rect 38332 16828 38500 16884
rect 38332 16660 38388 16670
rect 38332 16566 38388 16604
rect 38332 16322 38388 16334
rect 38332 16270 38334 16322
rect 38386 16270 38388 16322
rect 38332 16210 38388 16270
rect 38332 16158 38334 16210
rect 38386 16158 38388 16210
rect 38332 16146 38388 16158
rect 38220 15922 38276 15932
rect 38444 15652 38500 16828
rect 38332 15596 38500 15652
rect 38332 14642 38388 15596
rect 38556 15538 38612 16828
rect 38780 16212 38836 16222
rect 38780 16118 38836 16156
rect 38556 15486 38558 15538
rect 38610 15486 38612 15538
rect 38556 15474 38612 15486
rect 38332 14590 38334 14642
rect 38386 14590 38388 14642
rect 38332 14578 38388 14590
rect 38444 15428 38500 15438
rect 38892 15428 38948 17164
rect 38892 15372 39060 15428
rect 38444 15202 38500 15372
rect 38444 15150 38446 15202
rect 38498 15150 38500 15202
rect 38444 14644 38500 15150
rect 38892 15204 38948 15214
rect 38892 15110 38948 15148
rect 39004 15092 39060 15372
rect 39004 15026 39060 15036
rect 39116 14756 39172 17500
rect 39340 17490 39396 17500
rect 39452 17106 39508 17612
rect 39676 17556 39732 17566
rect 39564 17442 39620 17454
rect 39564 17390 39566 17442
rect 39618 17390 39620 17442
rect 39564 17220 39620 17390
rect 39564 17154 39620 17164
rect 39452 17054 39454 17106
rect 39506 17054 39508 17106
rect 39452 17042 39508 17054
rect 39676 16994 39732 17500
rect 39676 16942 39678 16994
rect 39730 16942 39732 16994
rect 39228 16884 39284 16922
rect 39228 16818 39284 16828
rect 39564 16884 39620 16894
rect 39228 16660 39284 16670
rect 39228 16098 39284 16604
rect 39228 16046 39230 16098
rect 39282 16046 39284 16098
rect 39228 16034 39284 16046
rect 39452 15988 39508 15998
rect 39340 15932 39452 15988
rect 39228 15428 39284 15438
rect 39340 15428 39396 15932
rect 39452 15922 39508 15932
rect 39564 15874 39620 16828
rect 39676 16098 39732 16942
rect 39676 16046 39678 16098
rect 39730 16046 39732 16098
rect 39676 16034 39732 16046
rect 39788 16882 39844 17612
rect 40236 17554 40292 17566
rect 40236 17502 40238 17554
rect 40290 17502 40292 17554
rect 39900 17220 39956 17230
rect 40236 17220 40292 17502
rect 39956 17164 40292 17220
rect 40348 17442 40404 17454
rect 40348 17390 40350 17442
rect 40402 17390 40404 17442
rect 40348 17220 40404 17390
rect 39900 17154 39956 17164
rect 39788 16830 39790 16882
rect 39842 16830 39844 16882
rect 39788 16098 39844 16830
rect 39788 16046 39790 16098
rect 39842 16046 39844 16098
rect 39788 16034 39844 16046
rect 40348 15988 40404 17164
rect 40460 17106 40516 18620
rect 40572 17668 40628 17678
rect 40684 17668 40740 19964
rect 40796 19684 40852 19694
rect 40796 19234 40852 19628
rect 41020 19460 41076 23996
rect 41132 20690 41188 26798
rect 41356 24052 41412 27694
rect 41580 27692 41748 27748
rect 41580 27300 41636 27692
rect 41468 27244 41636 27300
rect 41468 26908 41524 27244
rect 41692 26964 41748 27002
rect 41468 26852 41636 26908
rect 41356 23986 41412 23996
rect 41468 26178 41524 26190
rect 41468 26126 41470 26178
rect 41522 26126 41524 26178
rect 41244 23268 41300 23278
rect 41244 22820 41300 23212
rect 41244 22754 41300 22764
rect 41356 22932 41412 22942
rect 41356 22370 41412 22876
rect 41356 22318 41358 22370
rect 41410 22318 41412 22370
rect 41356 22306 41412 22318
rect 41244 22260 41300 22270
rect 41244 22166 41300 22204
rect 41244 21924 41300 21934
rect 41244 21810 41300 21868
rect 41244 21758 41246 21810
rect 41298 21758 41300 21810
rect 41244 21700 41300 21758
rect 41244 21634 41300 21644
rect 41132 20638 41134 20690
rect 41186 20638 41188 20690
rect 41132 20626 41188 20638
rect 41244 20802 41300 20814
rect 41244 20750 41246 20802
rect 41298 20750 41300 20802
rect 41132 20020 41188 20030
rect 41132 19926 41188 19964
rect 41244 19684 41300 20750
rect 41356 20132 41412 20142
rect 41356 20038 41412 20076
rect 41244 19618 41300 19628
rect 41020 19404 41300 19460
rect 40796 19182 40798 19234
rect 40850 19182 40852 19234
rect 40796 19170 40852 19182
rect 41132 19236 41188 19246
rect 40572 17666 40740 17668
rect 40572 17614 40574 17666
rect 40626 17614 40740 17666
rect 40572 17612 40740 17614
rect 40796 18676 40852 18686
rect 40572 17602 40628 17612
rect 40460 17054 40462 17106
rect 40514 17054 40516 17106
rect 40460 17042 40516 17054
rect 40684 16212 40740 16222
rect 40796 16212 40852 18620
rect 40908 18562 40964 18574
rect 40908 18510 40910 18562
rect 40962 18510 40964 18562
rect 40908 17556 40964 18510
rect 40908 17490 40964 17500
rect 41020 18564 41076 18574
rect 41020 17332 41076 18508
rect 41132 18450 41188 19180
rect 41244 19122 41300 19404
rect 41244 19070 41246 19122
rect 41298 19070 41300 19122
rect 41244 19058 41300 19070
rect 41132 18398 41134 18450
rect 41186 18398 41188 18450
rect 41132 18386 41188 18398
rect 41244 18900 41300 18910
rect 40908 17276 41076 17332
rect 40908 16996 40964 17276
rect 41132 16996 41188 17006
rect 40908 16994 41188 16996
rect 40908 16942 41134 16994
rect 41186 16942 41188 16994
rect 40908 16940 41188 16942
rect 41132 16930 41188 16940
rect 40684 16210 40852 16212
rect 40684 16158 40686 16210
rect 40738 16158 40852 16210
rect 40684 16156 40852 16158
rect 41132 16212 41188 16222
rect 41244 16212 41300 18844
rect 41468 17554 41524 26126
rect 41580 24836 41636 26852
rect 41692 26402 41748 26908
rect 41692 26350 41694 26402
rect 41746 26350 41748 26402
rect 41692 26338 41748 26350
rect 41804 26516 41860 43652
rect 42252 40404 42308 40414
rect 42252 38946 42308 40348
rect 42252 38894 42254 38946
rect 42306 38894 42308 38946
rect 42252 38882 42308 38894
rect 42476 28084 42532 43652
rect 42924 39396 42980 39406
rect 42924 39058 42980 39340
rect 42924 39006 42926 39058
rect 42978 39006 42980 39058
rect 42924 38994 42980 39006
rect 42700 38948 42756 38958
rect 42700 38854 42756 38892
rect 42588 38836 42644 38846
rect 42588 38742 42644 38780
rect 43036 38668 43092 43652
rect 43260 41860 43316 41870
rect 43260 40404 43316 41804
rect 43260 39058 43316 40348
rect 43260 39006 43262 39058
rect 43314 39006 43316 39058
rect 43260 38994 43316 39006
rect 43708 38836 43764 38846
rect 43708 38742 43764 38780
rect 43932 38668 43988 55412
rect 44268 38668 44324 55412
rect 42140 28082 42532 28084
rect 42140 28030 42478 28082
rect 42530 28030 42532 28082
rect 42140 28028 42532 28030
rect 41916 27970 41972 27982
rect 41916 27918 41918 27970
rect 41970 27918 41972 27970
rect 41916 26964 41972 27918
rect 42140 27074 42196 28028
rect 42476 28018 42532 28028
rect 42924 38612 43092 38668
rect 43708 38612 43988 38668
rect 44156 38612 44324 38668
rect 42140 27022 42142 27074
rect 42194 27022 42196 27074
rect 42140 27010 42196 27022
rect 42924 27188 42980 38612
rect 41916 26898 41972 26908
rect 42924 26908 42980 27132
rect 43036 27076 43092 27114
rect 43036 27010 43092 27020
rect 42476 26852 42532 26862
rect 42924 26852 43092 26908
rect 41804 26290 41860 26460
rect 41804 26238 41806 26290
rect 41858 26238 41860 26290
rect 41804 26226 41860 26238
rect 42364 26850 42532 26852
rect 42364 26798 42478 26850
rect 42530 26798 42532 26850
rect 42364 26796 42532 26798
rect 41916 25732 41972 25742
rect 41804 25508 41860 25518
rect 41692 25452 41804 25508
rect 41692 25396 41748 25452
rect 41804 25442 41860 25452
rect 41692 25060 41748 25340
rect 41916 25396 41972 25676
rect 42364 25508 42420 26796
rect 42476 26786 42532 26796
rect 43036 26740 43092 26852
rect 42700 26684 43092 26740
rect 42588 26516 42644 26526
rect 42588 26422 42644 26460
rect 42700 26292 42756 26684
rect 43708 26516 43764 38612
rect 43820 27188 43876 27198
rect 43820 27094 43876 27132
rect 44156 26740 44212 38612
rect 45052 36372 45108 36382
rect 45052 36278 45108 36316
rect 44716 36260 44772 36270
rect 44716 35924 44772 36204
rect 45164 36258 45220 36270
rect 45164 36206 45166 36258
rect 45218 36206 45220 36258
rect 44716 35922 45108 35924
rect 44716 35870 44718 35922
rect 44770 35870 45108 35922
rect 44716 35868 45108 35870
rect 44716 35858 44772 35868
rect 45052 35810 45108 35868
rect 45052 35758 45054 35810
rect 45106 35758 45108 35810
rect 45052 35746 45108 35758
rect 45164 35700 45220 36206
rect 45164 35634 45220 35644
rect 45164 35474 45220 35486
rect 45164 35422 45166 35474
rect 45218 35422 45220 35474
rect 45164 35140 45220 35422
rect 45164 35074 45220 35084
rect 45164 34802 45220 34814
rect 45164 34750 45166 34802
rect 45218 34750 45220 34802
rect 44380 34692 44436 34702
rect 44380 34598 44436 34636
rect 45164 34692 45220 34750
rect 45276 34804 45332 34814
rect 45276 34710 45332 34748
rect 45164 34626 45220 34636
rect 45276 34132 45332 34142
rect 45276 33570 45332 34076
rect 45276 33518 45278 33570
rect 45330 33518 45332 33570
rect 45276 33506 45332 33518
rect 45164 33236 45220 33246
rect 45164 33142 45220 33180
rect 45500 33012 45556 75516
rect 45612 75506 45668 75516
rect 46284 55468 46340 76302
rect 45724 55412 46340 55468
rect 46508 75906 46564 75918
rect 46508 75854 46510 75906
rect 46562 75854 46564 75906
rect 45724 43708 45780 55412
rect 46508 43708 46564 75854
rect 46620 75796 46676 75806
rect 46732 75796 46788 76414
rect 46620 75794 46788 75796
rect 46620 75742 46622 75794
rect 46674 75742 46788 75794
rect 46620 75740 46788 75742
rect 46620 75730 46676 75740
rect 47068 75684 47124 76636
rect 47852 76468 47908 76636
rect 48188 76692 48244 79200
rect 48188 76626 48244 76636
rect 48300 77026 48356 77038
rect 48300 76974 48302 77026
rect 48354 76974 48356 77026
rect 48300 76692 48356 76974
rect 48860 77026 48916 79200
rect 48860 76974 48862 77026
rect 48914 76974 48916 77026
rect 48860 76962 48916 76974
rect 49532 76804 49588 79200
rect 50092 77026 50148 77038
rect 50092 76974 50094 77026
rect 50146 76974 50148 77026
rect 49532 76748 49812 76804
rect 49196 76692 49252 76702
rect 48300 76690 48580 76692
rect 48300 76638 48302 76690
rect 48354 76638 48580 76690
rect 48300 76636 48580 76638
rect 48300 76626 48356 76636
rect 47852 76466 48132 76468
rect 47852 76414 47854 76466
rect 47906 76414 48132 76466
rect 47852 76412 48132 76414
rect 47852 76402 47908 76412
rect 47404 76356 47460 76366
rect 47404 76262 47460 76300
rect 48076 75794 48132 76412
rect 48076 75742 48078 75794
rect 48130 75742 48132 75794
rect 48076 75730 48132 75742
rect 48524 75794 48580 76636
rect 48524 75742 48526 75794
rect 48578 75742 48580 75794
rect 48524 75730 48580 75742
rect 48636 76356 48692 76366
rect 46844 75682 47124 75684
rect 46844 75630 47070 75682
rect 47122 75630 47124 75682
rect 46844 75628 47124 75630
rect 46844 75122 46900 75628
rect 47068 75618 47124 75628
rect 47628 75684 47684 75694
rect 47628 75590 47684 75628
rect 46844 75070 46846 75122
rect 46898 75070 46900 75122
rect 46844 75058 46900 75070
rect 45724 43652 45892 43708
rect 46508 43652 46900 43708
rect 45612 36372 45668 36382
rect 45612 36278 45668 36316
rect 45724 35700 45780 35710
rect 45724 35606 45780 35644
rect 45836 35364 45892 43652
rect 46844 38668 46900 43652
rect 46732 38612 46900 38668
rect 46620 36260 46676 36270
rect 46508 36204 46620 36260
rect 45948 35700 46004 35710
rect 45948 35606 46004 35644
rect 46172 35698 46228 35710
rect 46172 35646 46174 35698
rect 46226 35646 46228 35698
rect 45836 35308 46004 35364
rect 45724 35140 45780 35150
rect 45724 34914 45780 35084
rect 45724 34862 45726 34914
rect 45778 34862 45780 34914
rect 45724 34850 45780 34862
rect 45948 34580 46004 35308
rect 46060 35252 46116 35262
rect 46060 34690 46116 35196
rect 46172 34916 46228 35646
rect 46396 35698 46452 35710
rect 46396 35646 46398 35698
rect 46450 35646 46452 35698
rect 46284 35028 46340 35038
rect 46284 34916 46340 34972
rect 46172 34914 46340 34916
rect 46172 34862 46174 34914
rect 46226 34862 46340 34914
rect 46172 34860 46340 34862
rect 46172 34850 46228 34860
rect 46060 34638 46062 34690
rect 46114 34638 46116 34690
rect 46060 34626 46116 34638
rect 45276 32956 45556 33012
rect 45612 34524 46004 34580
rect 44940 31778 44996 31790
rect 44940 31726 44942 31778
rect 44994 31726 44996 31778
rect 44828 31668 44884 31678
rect 44940 31668 44996 31726
rect 44884 31612 44996 31668
rect 45052 31668 45108 31678
rect 44828 31602 44884 31612
rect 45052 31574 45108 31612
rect 44268 31556 44324 31566
rect 44268 31220 44324 31500
rect 44268 31218 44660 31220
rect 44268 31166 44270 31218
rect 44322 31166 44660 31218
rect 44268 31164 44660 31166
rect 44268 31154 44324 31164
rect 44604 31106 44660 31164
rect 44604 31054 44606 31106
rect 44658 31054 44660 31106
rect 44604 31042 44660 31054
rect 44716 30996 44772 31006
rect 44716 30902 44772 30940
rect 44940 30548 44996 30558
rect 44940 30210 44996 30492
rect 44940 30158 44942 30210
rect 44994 30158 44996 30210
rect 44940 30146 44996 30158
rect 45276 30212 45332 32956
rect 45612 32900 45668 34524
rect 45724 34356 45780 34366
rect 45724 33460 45780 34300
rect 46284 34242 46340 34860
rect 46284 34190 46286 34242
rect 46338 34190 46340 34242
rect 45836 34132 45892 34142
rect 45836 34038 45892 34076
rect 46060 34018 46116 34030
rect 46060 33966 46062 34018
rect 46114 33966 46116 34018
rect 45724 33404 45892 33460
rect 45724 33236 45780 33246
rect 45724 33142 45780 33180
rect 45388 32844 45668 32900
rect 45388 31220 45444 32844
rect 45500 32676 45556 32686
rect 45836 32676 45892 33404
rect 46060 33348 46116 33966
rect 46060 33282 46116 33292
rect 46284 33236 46340 34190
rect 46396 34802 46452 35646
rect 46396 34750 46398 34802
rect 46450 34750 46452 34802
rect 46396 34132 46452 34750
rect 46508 34356 46564 36204
rect 46620 36194 46676 36204
rect 46620 34914 46676 34926
rect 46620 34862 46622 34914
rect 46674 34862 46676 34914
rect 46620 34804 46676 34862
rect 46620 34738 46676 34748
rect 46508 34290 46564 34300
rect 46508 34132 46564 34142
rect 46396 34076 46508 34132
rect 46508 34038 46564 34076
rect 46396 33236 46452 33246
rect 46284 33234 46452 33236
rect 46284 33182 46398 33234
rect 46450 33182 46452 33234
rect 46284 33180 46452 33182
rect 46396 33170 46452 33180
rect 45500 32674 45892 32676
rect 45500 32622 45502 32674
rect 45554 32622 45838 32674
rect 45890 32622 45892 32674
rect 45500 32620 45892 32622
rect 45500 32610 45556 32620
rect 45500 31556 45556 31566
rect 45500 31462 45556 31500
rect 45388 31164 45668 31220
rect 45500 30994 45556 31006
rect 45500 30942 45502 30994
rect 45554 30942 45556 30994
rect 45500 30434 45556 30942
rect 45500 30382 45502 30434
rect 45554 30382 45556 30434
rect 45500 30370 45556 30382
rect 45276 30156 45556 30212
rect 44828 30100 44884 30110
rect 44828 30006 44884 30044
rect 45164 30100 45220 30110
rect 45164 29650 45220 30044
rect 45388 29988 45444 29998
rect 45388 29894 45444 29932
rect 45164 29598 45166 29650
rect 45218 29598 45220 29650
rect 45164 29586 45220 29598
rect 44828 29540 44884 29550
rect 45052 29540 45108 29550
rect 44884 29538 45108 29540
rect 44884 29486 45054 29538
rect 45106 29486 45108 29538
rect 44884 29484 45108 29486
rect 44828 29446 44884 29484
rect 45052 29474 45108 29484
rect 44604 28644 44660 28654
rect 44604 28084 44660 28588
rect 44604 28082 44996 28084
rect 44604 28030 44606 28082
rect 44658 28030 44996 28082
rect 44604 28028 44996 28030
rect 44604 28018 44660 28028
rect 44940 27970 44996 28028
rect 44940 27918 44942 27970
rect 44994 27918 44996 27970
rect 44940 27906 44996 27918
rect 44828 27636 44884 27646
rect 44828 27188 44884 27580
rect 45052 27636 45108 27646
rect 45052 27542 45108 27580
rect 45388 27188 45444 27198
rect 44828 27186 45444 27188
rect 44828 27134 44830 27186
rect 44882 27134 45390 27186
rect 45442 27134 45444 27186
rect 44828 27132 45444 27134
rect 44828 27122 44884 27132
rect 45388 27122 45444 27132
rect 44940 26964 44996 27002
rect 44940 26898 44996 26908
rect 44156 26674 44212 26684
rect 44380 26850 44436 26862
rect 44380 26798 44382 26850
rect 44434 26798 44436 26850
rect 42364 25442 42420 25452
rect 42476 26236 42756 26292
rect 43036 26402 43092 26414
rect 43708 26404 43764 26460
rect 44044 26516 44100 26526
rect 44044 26514 44324 26516
rect 44044 26462 44046 26514
rect 44098 26462 44324 26514
rect 44044 26460 44324 26462
rect 44044 26450 44100 26460
rect 43036 26350 43038 26402
rect 43090 26350 43092 26402
rect 42476 25506 42532 26236
rect 42476 25454 42478 25506
rect 42530 25454 42532 25506
rect 42476 25442 42532 25454
rect 41916 25340 42084 25396
rect 41804 25284 41860 25294
rect 41916 25284 41972 25340
rect 41804 25282 41972 25284
rect 41804 25230 41806 25282
rect 41858 25230 41972 25282
rect 41804 25228 41972 25230
rect 41804 25218 41860 25228
rect 41692 25004 41860 25060
rect 41692 24836 41748 24846
rect 41580 24834 41748 24836
rect 41580 24782 41694 24834
rect 41746 24782 41748 24834
rect 41580 24780 41748 24782
rect 41580 23380 41636 24780
rect 41692 24770 41748 24780
rect 41692 24052 41748 24062
rect 41692 23492 41748 23996
rect 41804 23938 41860 25004
rect 41804 23886 41806 23938
rect 41858 23886 41860 23938
rect 41804 23874 41860 23886
rect 42028 23940 42084 25340
rect 42140 25394 42196 25406
rect 42140 25342 42142 25394
rect 42194 25342 42196 25394
rect 42140 23940 42196 25342
rect 42588 25396 42644 25406
rect 43036 25396 43092 26350
rect 43596 26348 43764 26404
rect 43596 26290 43652 26348
rect 43596 26238 43598 26290
rect 43650 26238 43652 26290
rect 43596 26226 43652 26238
rect 44156 26290 44212 26302
rect 44156 26238 44158 26290
rect 44210 26238 44212 26290
rect 43708 25620 43764 25630
rect 43372 25508 43428 25518
rect 42588 25394 43036 25396
rect 42588 25342 42590 25394
rect 42642 25342 43036 25394
rect 42588 25340 43036 25342
rect 42364 24052 42420 24062
rect 42588 24052 42644 25340
rect 43036 25302 43092 25340
rect 43260 25452 43372 25508
rect 42364 24050 42644 24052
rect 42364 23998 42366 24050
rect 42418 23998 42644 24050
rect 42364 23996 42644 23998
rect 43260 24050 43316 25452
rect 43372 25414 43428 25452
rect 43484 25282 43540 25294
rect 43484 25230 43486 25282
rect 43538 25230 43540 25282
rect 43260 23998 43262 24050
rect 43314 23998 43316 24050
rect 42364 23986 42420 23996
rect 43260 23986 43316 23998
rect 43372 25172 43428 25182
rect 42700 23940 42756 23950
rect 42140 23884 42308 23940
rect 42028 23874 42084 23884
rect 42252 23828 42308 23884
rect 42700 23846 42756 23884
rect 42252 23772 42532 23828
rect 41692 23436 41972 23492
rect 41580 23314 41636 23324
rect 41692 23268 41748 23278
rect 41692 23174 41748 23212
rect 41580 23154 41636 23166
rect 41580 23102 41582 23154
rect 41634 23102 41636 23154
rect 41580 19572 41636 23102
rect 41804 23156 41860 23166
rect 41692 22932 41748 22942
rect 41692 22838 41748 22876
rect 41804 22260 41860 23100
rect 41804 22194 41860 22204
rect 41916 20132 41972 23436
rect 42028 23380 42084 23390
rect 42028 22482 42084 23324
rect 42364 23154 42420 23166
rect 42364 23102 42366 23154
rect 42418 23102 42420 23154
rect 42252 23044 42308 23054
rect 42252 22950 42308 22988
rect 42028 22430 42030 22482
rect 42082 22430 42084 22482
rect 42028 22418 42084 22430
rect 42364 22372 42420 23102
rect 42476 23156 42532 23772
rect 43372 23380 43428 25116
rect 43372 23286 43428 23324
rect 42476 23090 42532 23100
rect 42812 23268 42868 23278
rect 42476 22372 42532 22382
rect 42364 22370 42532 22372
rect 42364 22318 42478 22370
rect 42530 22318 42532 22370
rect 42364 22316 42532 22318
rect 42028 21362 42084 21374
rect 42028 21310 42030 21362
rect 42082 21310 42084 21362
rect 42028 20804 42084 21310
rect 42028 20738 42084 20748
rect 41916 20066 41972 20076
rect 42140 20468 42196 20478
rect 41580 19506 41636 19516
rect 41804 19460 41860 19470
rect 41692 19348 41748 19358
rect 41580 19012 41636 19022
rect 41580 18562 41636 18956
rect 41692 18674 41748 19292
rect 41692 18622 41694 18674
rect 41746 18622 41748 18674
rect 41692 18610 41748 18622
rect 41580 18510 41582 18562
rect 41634 18510 41636 18562
rect 41580 18498 41636 18510
rect 41468 17502 41470 17554
rect 41522 17502 41524 17554
rect 41468 17490 41524 17502
rect 41580 18004 41636 18014
rect 41356 17444 41412 17454
rect 41356 16994 41412 17388
rect 41356 16942 41358 16994
rect 41410 16942 41412 16994
rect 41356 16930 41412 16942
rect 41468 16996 41524 17006
rect 41468 16902 41524 16940
rect 41580 16436 41636 17948
rect 41692 17666 41748 17678
rect 41692 17614 41694 17666
rect 41746 17614 41748 17666
rect 41692 17106 41748 17614
rect 41692 17054 41694 17106
rect 41746 17054 41748 17106
rect 41692 17042 41748 17054
rect 41132 16210 41300 16212
rect 41132 16158 41134 16210
rect 41186 16158 41300 16210
rect 41132 16156 41300 16158
rect 41468 16380 41636 16436
rect 40684 16146 40740 16156
rect 41132 16146 41188 16156
rect 40348 15932 41188 15988
rect 39564 15822 39566 15874
rect 39618 15822 39620 15874
rect 39564 15810 39620 15822
rect 40236 15876 40292 15886
rect 39228 15426 39396 15428
rect 39228 15374 39230 15426
rect 39282 15374 39396 15426
rect 39228 15372 39396 15374
rect 39228 15316 39284 15372
rect 39452 15316 39508 15326
rect 39228 15250 39284 15260
rect 39340 15314 39508 15316
rect 39340 15262 39454 15314
rect 39506 15262 39508 15314
rect 39340 15260 39508 15262
rect 39116 14690 39172 14700
rect 38668 14644 38724 14654
rect 38444 14642 38724 14644
rect 38444 14590 38670 14642
rect 38722 14590 38724 14642
rect 38444 14588 38724 14590
rect 38668 14578 38724 14588
rect 39004 14530 39060 14542
rect 39004 14478 39006 14530
rect 39058 14478 39060 14530
rect 38556 14308 38612 14318
rect 38444 13972 38500 13982
rect 38220 13860 38276 13870
rect 38220 13524 38276 13804
rect 38332 13858 38388 13870
rect 38332 13806 38334 13858
rect 38386 13806 38388 13858
rect 38332 13636 38388 13806
rect 38332 13570 38388 13580
rect 38220 13458 38276 13468
rect 38444 12962 38500 13916
rect 38556 13970 38612 14252
rect 38556 13918 38558 13970
rect 38610 13918 38612 13970
rect 38556 13906 38612 13918
rect 38780 13860 38836 13870
rect 38780 13766 38836 13804
rect 38444 12910 38446 12962
rect 38498 12910 38500 12962
rect 38444 12898 38500 12910
rect 39004 12964 39060 14478
rect 39116 14196 39172 14206
rect 39116 13970 39172 14140
rect 39116 13918 39118 13970
rect 39170 13918 39172 13970
rect 39116 13906 39172 13918
rect 39340 13970 39396 15260
rect 39452 15250 39508 15260
rect 39900 15316 39956 15326
rect 39900 15222 39956 15260
rect 40124 15314 40180 15326
rect 40124 15262 40126 15314
rect 40178 15262 40180 15314
rect 40012 15202 40068 15214
rect 40012 15150 40014 15202
rect 40066 15150 40068 15202
rect 40012 15148 40068 15150
rect 39788 15092 40068 15148
rect 39788 14642 39844 15092
rect 39788 14590 39790 14642
rect 39842 14590 39844 14642
rect 39788 14578 39844 14590
rect 40124 14196 40180 15262
rect 40124 14130 40180 14140
rect 39340 13918 39342 13970
rect 39394 13918 39396 13970
rect 39340 13906 39396 13918
rect 39564 13858 39620 13870
rect 40236 13860 40292 15820
rect 41132 15538 41188 15932
rect 41132 15486 41134 15538
rect 41186 15486 41188 15538
rect 41132 15474 41188 15486
rect 41468 15540 41524 16380
rect 41804 16324 41860 19404
rect 42140 18562 42196 20412
rect 42140 18510 42142 18562
rect 42194 18510 42196 18562
rect 41916 18452 41972 18462
rect 41916 18358 41972 18396
rect 42028 17780 42084 17790
rect 42028 17106 42084 17724
rect 42028 17054 42030 17106
rect 42082 17054 42084 17106
rect 42028 17042 42084 17054
rect 41916 16884 41972 16894
rect 41916 16790 41972 16828
rect 41580 16268 41860 16324
rect 41580 16210 41636 16268
rect 41580 16158 41582 16210
rect 41634 16158 41636 16210
rect 41580 16146 41636 16158
rect 42140 16100 42196 18510
rect 42252 19234 42308 19246
rect 42252 19182 42254 19234
rect 42306 19182 42308 19234
rect 42252 17106 42308 19182
rect 42252 17054 42254 17106
rect 42306 17054 42308 17106
rect 42252 17042 42308 17054
rect 42140 16034 42196 16044
rect 42252 16884 42308 16894
rect 41916 15986 41972 15998
rect 41916 15934 41918 15986
rect 41970 15934 41972 15986
rect 41804 15874 41860 15886
rect 41804 15822 41806 15874
rect 41858 15822 41860 15874
rect 41580 15540 41636 15550
rect 41468 15538 41636 15540
rect 41468 15486 41582 15538
rect 41634 15486 41636 15538
rect 41468 15484 41636 15486
rect 41580 15474 41636 15484
rect 41804 15316 41860 15822
rect 41580 14868 41636 14878
rect 41244 14644 41300 14654
rect 41244 13970 41300 14588
rect 41244 13918 41246 13970
rect 41298 13918 41300 13970
rect 41244 13906 41300 13918
rect 41468 14196 41524 14206
rect 41468 13970 41524 14140
rect 41468 13918 41470 13970
rect 41522 13918 41524 13970
rect 41468 13906 41524 13918
rect 39564 13806 39566 13858
rect 39618 13806 39620 13858
rect 39564 13188 39620 13806
rect 40124 13804 40292 13860
rect 39676 13746 39732 13758
rect 39676 13694 39678 13746
rect 39730 13694 39732 13746
rect 39676 13524 39732 13694
rect 39676 13458 39732 13468
rect 39564 13132 39732 13188
rect 39116 12964 39172 12974
rect 39004 12908 39116 12964
rect 39116 12898 39172 12908
rect 39564 12964 39620 12974
rect 38780 12740 38836 12750
rect 38780 12738 39508 12740
rect 38780 12686 38782 12738
rect 38834 12686 39508 12738
rect 38780 12684 39508 12686
rect 38108 11330 38164 11340
rect 38220 12066 38276 12078
rect 38220 12014 38222 12066
rect 38274 12014 38276 12066
rect 37660 11282 37716 11294
rect 37660 11230 37662 11282
rect 37714 11230 37716 11282
rect 37660 10948 37716 11230
rect 38220 11284 38276 12014
rect 38668 11396 38724 11406
rect 38220 11218 38276 11228
rect 38556 11394 38724 11396
rect 38556 11342 38670 11394
rect 38722 11342 38724 11394
rect 38556 11340 38724 11342
rect 37660 10882 37716 10892
rect 38332 11172 38388 11182
rect 38556 11172 38612 11340
rect 38668 11330 38724 11340
rect 38332 11170 38612 11172
rect 38332 11118 38334 11170
rect 38386 11118 38612 11170
rect 38332 11116 38612 11118
rect 38332 10836 38388 11116
rect 38332 10770 38388 10780
rect 38780 9940 38836 12684
rect 39452 11508 39508 12684
rect 39564 12180 39620 12908
rect 39564 12114 39620 12124
rect 39452 11452 39620 11508
rect 39452 11284 39508 11294
rect 39340 10836 39396 10846
rect 39340 10742 39396 10780
rect 39452 10834 39508 11228
rect 39452 10782 39454 10834
rect 39506 10782 39508 10834
rect 39452 10770 39508 10782
rect 39564 10834 39620 11452
rect 39676 11172 39732 13132
rect 39676 11106 39732 11116
rect 39564 10782 39566 10834
rect 39618 10782 39620 10834
rect 39564 10770 39620 10782
rect 38892 10612 38948 10622
rect 38892 10518 38948 10556
rect 38108 9826 38164 9838
rect 38108 9774 38110 9826
rect 38162 9774 38164 9826
rect 37100 8930 37268 8932
rect 37100 8878 37102 8930
rect 37154 8878 37268 8930
rect 37100 8876 37268 8878
rect 37324 9042 37604 9044
rect 37324 8990 37438 9042
rect 37490 8990 37604 9042
rect 37324 8988 37604 8990
rect 37884 9602 37940 9614
rect 37884 9550 37886 9602
rect 37938 9550 37940 9602
rect 37100 8820 37156 8876
rect 37100 8754 37156 8764
rect 36428 8372 36484 8382
rect 36428 8370 36708 8372
rect 36428 8318 36430 8370
rect 36482 8318 36708 8370
rect 36428 8316 36708 8318
rect 36428 8306 36484 8316
rect 36092 6580 36148 6590
rect 35868 6468 35924 6478
rect 35868 5010 35924 6412
rect 36092 5908 36148 6524
rect 36092 5842 36148 5852
rect 35868 4958 35870 5010
rect 35922 4958 35924 5010
rect 35868 4946 35924 4958
rect 36204 4226 36260 6636
rect 36316 8034 36372 8046
rect 36316 7982 36318 8034
rect 36370 7982 36372 8034
rect 36316 5460 36372 7982
rect 36428 6468 36484 6478
rect 36428 6466 36596 6468
rect 36428 6414 36430 6466
rect 36482 6414 36596 6466
rect 36428 6412 36596 6414
rect 36428 6402 36484 6412
rect 36316 5394 36372 5404
rect 36428 5348 36484 5358
rect 36428 5122 36484 5292
rect 36428 5070 36430 5122
rect 36482 5070 36484 5122
rect 36428 5058 36484 5070
rect 36540 4452 36596 6412
rect 36540 4386 36596 4396
rect 36204 4174 36206 4226
rect 36258 4174 36260 4226
rect 36204 4162 36260 4174
rect 36092 3668 36148 3678
rect 36092 3388 36148 3612
rect 35756 3332 35924 3388
rect 34524 1876 34580 1886
rect 34524 800 34580 1820
rect 35196 800 35252 3332
rect 35868 800 35924 3332
rect 35980 3332 36148 3388
rect 36652 3442 36708 8316
rect 37100 8148 37156 8158
rect 37100 8054 37156 8092
rect 36988 7700 37044 7710
rect 36876 5460 36932 5470
rect 36652 3390 36654 3442
rect 36706 3390 36708 3442
rect 36652 3378 36708 3390
rect 36764 5404 36876 5460
rect 36764 3388 36820 5404
rect 36876 5394 36932 5404
rect 36988 5348 37044 7644
rect 37324 6690 37380 8988
rect 37436 8978 37492 8988
rect 37772 8146 37828 8158
rect 37772 8094 37774 8146
rect 37826 8094 37828 8146
rect 37436 8036 37492 8046
rect 37436 8034 37604 8036
rect 37436 7982 37438 8034
rect 37490 7982 37604 8034
rect 37436 7980 37604 7982
rect 37436 7970 37492 7980
rect 37436 7362 37492 7374
rect 37436 7310 37438 7362
rect 37490 7310 37492 7362
rect 37436 7252 37492 7310
rect 37436 7186 37492 7196
rect 37548 6804 37604 7980
rect 37772 7028 37828 8094
rect 37772 6962 37828 6972
rect 37548 6748 37828 6804
rect 37324 6638 37326 6690
rect 37378 6638 37380 6690
rect 37324 6626 37380 6638
rect 37660 6020 37716 6030
rect 37324 6018 37716 6020
rect 37324 5966 37662 6018
rect 37714 5966 37716 6018
rect 37324 5964 37716 5966
rect 37100 5908 37156 5918
rect 37100 5906 37268 5908
rect 37100 5854 37102 5906
rect 37154 5854 37268 5906
rect 37100 5852 37268 5854
rect 37100 5842 37156 5852
rect 37100 5348 37156 5358
rect 36988 5346 37156 5348
rect 36988 5294 37102 5346
rect 37154 5294 37156 5346
rect 36988 5292 37156 5294
rect 37100 5282 37156 5292
rect 37100 5124 37156 5134
rect 36876 5122 37156 5124
rect 36876 5070 37102 5122
rect 37154 5070 37156 5122
rect 36876 5068 37156 5070
rect 36876 3668 36932 5068
rect 37100 5058 37156 5068
rect 37212 4676 37268 5852
rect 36876 3554 36932 3612
rect 36876 3502 36878 3554
rect 36930 3502 36932 3554
rect 36876 3490 36932 3502
rect 36988 4620 37268 4676
rect 36764 3332 36932 3388
rect 35980 2100 36036 3332
rect 35980 2034 36036 2044
rect 36540 2324 36596 2334
rect 36540 800 36596 2268
rect 36876 2212 36932 3332
rect 36988 2884 37044 4620
rect 37100 4450 37156 4462
rect 37100 4398 37102 4450
rect 37154 4398 37156 4450
rect 37100 4116 37156 4398
rect 37100 4050 37156 4060
rect 36988 2818 37044 2828
rect 37212 3556 37268 3566
rect 36876 2146 36932 2156
rect 37212 800 37268 3500
rect 37324 2996 37380 5964
rect 37660 5954 37716 5964
rect 37548 5460 37604 5470
rect 37436 5346 37492 5358
rect 37436 5294 37438 5346
rect 37490 5294 37492 5346
rect 37436 5122 37492 5294
rect 37436 5070 37438 5122
rect 37490 5070 37492 5122
rect 37436 5058 37492 5070
rect 37548 5122 37604 5404
rect 37548 5070 37550 5122
rect 37602 5070 37604 5122
rect 37548 5058 37604 5070
rect 37660 5236 37716 5246
rect 37660 3442 37716 5180
rect 37772 4340 37828 6748
rect 37884 6692 37940 9550
rect 38108 8260 38164 9774
rect 38668 9828 38724 9838
rect 38780 9828 38836 9884
rect 38668 9826 38836 9828
rect 38668 9774 38670 9826
rect 38722 9774 38836 9826
rect 38668 9772 38836 9774
rect 39228 9828 39284 9838
rect 39452 9828 39508 9838
rect 39228 9826 39508 9828
rect 39228 9774 39230 9826
rect 39282 9774 39454 9826
rect 39506 9774 39508 9826
rect 39228 9772 39508 9774
rect 38668 9762 38724 9772
rect 39228 9762 39284 9772
rect 39452 9762 39508 9772
rect 39788 9828 39844 9838
rect 39788 9734 39844 9772
rect 38780 9602 38836 9614
rect 38780 9550 38782 9602
rect 38834 9550 38836 9602
rect 38668 9268 38724 9278
rect 38220 9156 38276 9166
rect 38220 9062 38276 9100
rect 38668 9044 38724 9212
rect 38780 9156 38836 9550
rect 38892 9602 38948 9614
rect 38892 9550 38894 9602
rect 38946 9550 38948 9602
rect 38892 9268 38948 9550
rect 39676 9604 39732 9614
rect 39676 9510 39732 9548
rect 38892 9202 38948 9212
rect 38780 9090 38836 9100
rect 38668 8978 38724 8988
rect 38780 8370 38836 8382
rect 38780 8318 38782 8370
rect 38834 8318 38836 8370
rect 38108 8204 38276 8260
rect 38108 8034 38164 8046
rect 38108 7982 38110 8034
rect 38162 7982 38164 8034
rect 37996 6692 38052 6702
rect 37884 6690 38052 6692
rect 37884 6638 37998 6690
rect 38050 6638 38052 6690
rect 37884 6636 38052 6638
rect 37996 6626 38052 6636
rect 38108 5124 38164 7982
rect 38220 7698 38276 8204
rect 38780 7812 38836 8318
rect 40124 8370 40180 13804
rect 40796 13748 40852 13758
rect 40796 13654 40852 13692
rect 40236 13636 40292 13646
rect 40236 13074 40292 13580
rect 41356 13636 41412 13646
rect 41356 13542 41412 13580
rect 40236 13022 40238 13074
rect 40290 13022 40292 13074
rect 40236 13010 40292 13022
rect 40908 13412 40964 13422
rect 40908 12290 40964 13356
rect 41244 12404 41300 12414
rect 41580 12404 41636 14812
rect 41804 13748 41860 15260
rect 41916 14642 41972 15934
rect 42140 15316 42196 15326
rect 42028 15314 42196 15316
rect 42028 15262 42142 15314
rect 42194 15262 42196 15314
rect 42028 15260 42196 15262
rect 42028 15148 42084 15260
rect 42140 15250 42196 15260
rect 42028 15092 42196 15148
rect 41916 14590 41918 14642
rect 41970 14590 41972 14642
rect 41916 14578 41972 14590
rect 41804 13682 41860 13692
rect 42140 13746 42196 15092
rect 42140 13694 42142 13746
rect 42194 13694 42196 13746
rect 41916 12964 41972 12974
rect 42140 12964 42196 13694
rect 41972 12908 42196 12964
rect 41916 12898 41972 12908
rect 41244 12310 41300 12348
rect 41356 12402 41636 12404
rect 41356 12350 41582 12402
rect 41634 12350 41636 12402
rect 41356 12348 41636 12350
rect 40908 12238 40910 12290
rect 40962 12238 40964 12290
rect 40908 12226 40964 12238
rect 41020 12290 41076 12302
rect 41020 12238 41022 12290
rect 41074 12238 41076 12290
rect 40348 12066 40404 12078
rect 40348 12014 40350 12066
rect 40402 12014 40404 12066
rect 40236 11732 40292 11742
rect 40236 10836 40292 11676
rect 40236 10500 40292 10780
rect 40348 10722 40404 12014
rect 41020 11620 41076 12238
rect 41020 11554 41076 11564
rect 41356 11508 41412 12348
rect 41580 12338 41636 12348
rect 40348 10670 40350 10722
rect 40402 10670 40404 10722
rect 40348 10658 40404 10670
rect 41132 11452 41412 11508
rect 41020 10500 41076 10510
rect 40236 10444 40404 10500
rect 40348 9938 40404 10444
rect 40348 9886 40350 9938
rect 40402 9886 40404 9938
rect 40348 9874 40404 9886
rect 40908 10498 41076 10500
rect 40908 10446 41022 10498
rect 41074 10446 41076 10498
rect 40908 10444 41076 10446
rect 40684 9716 40740 9726
rect 40460 9714 40740 9716
rect 40460 9662 40686 9714
rect 40738 9662 40740 9714
rect 40460 9660 40740 9662
rect 40348 8932 40404 8942
rect 40460 8932 40516 9660
rect 40684 9650 40740 9660
rect 40348 8930 40516 8932
rect 40348 8878 40350 8930
rect 40402 8878 40516 8930
rect 40348 8876 40516 8878
rect 40348 8866 40404 8876
rect 40124 8318 40126 8370
rect 40178 8318 40180 8370
rect 40124 8306 40180 8318
rect 38220 7646 38222 7698
rect 38274 7646 38276 7698
rect 38220 7634 38276 7646
rect 38668 7756 38836 7812
rect 38892 8258 38948 8270
rect 38892 8206 38894 8258
rect 38946 8206 38948 8258
rect 38556 7250 38612 7262
rect 38556 7198 38558 7250
rect 38610 7198 38612 7250
rect 38556 6916 38612 7198
rect 38556 6850 38612 6860
rect 38108 5058 38164 5068
rect 38220 6580 38276 6590
rect 38108 4340 38164 4350
rect 37772 4338 38164 4340
rect 37772 4286 38110 4338
rect 38162 4286 38164 4338
rect 37772 4284 38164 4286
rect 38108 4274 38164 4284
rect 37660 3390 37662 3442
rect 37714 3390 37716 3442
rect 37660 3378 37716 3390
rect 38220 3388 38276 6524
rect 38668 5348 38724 7756
rect 38780 7588 38836 7598
rect 38780 7494 38836 7532
rect 38780 6132 38836 6142
rect 38892 6132 38948 8206
rect 40684 8258 40740 8270
rect 40684 8206 40686 8258
rect 40738 8206 40740 8258
rect 39228 8146 39284 8158
rect 39228 8094 39230 8146
rect 39282 8094 39284 8146
rect 39228 6916 39284 8094
rect 39564 8148 39620 8158
rect 39228 6850 39284 6860
rect 39340 7586 39396 7598
rect 39340 7534 39342 7586
rect 39394 7534 39396 7586
rect 39340 6804 39396 7534
rect 39340 6738 39396 6748
rect 38836 6076 38948 6132
rect 38780 6066 38836 6076
rect 39340 6018 39396 6030
rect 39340 5966 39342 6018
rect 39394 5966 39396 6018
rect 39228 5908 39284 5918
rect 38668 5282 38724 5292
rect 38892 5906 39284 5908
rect 38892 5854 39230 5906
rect 39282 5854 39284 5906
rect 38892 5852 39284 5854
rect 38892 5124 38948 5852
rect 39228 5842 39284 5852
rect 38332 5122 38948 5124
rect 38332 5070 38894 5122
rect 38946 5070 38948 5122
rect 38332 5068 38948 5070
rect 38332 5010 38388 5068
rect 38892 5058 38948 5068
rect 39004 5684 39060 5694
rect 38332 4958 38334 5010
rect 38386 4958 38388 5010
rect 38332 4946 38388 4958
rect 39004 5012 39060 5628
rect 39340 5124 39396 5966
rect 39004 4918 39060 4956
rect 39228 5068 39396 5124
rect 37324 2930 37380 2940
rect 37884 3332 38276 3388
rect 38556 4788 38612 4798
rect 37884 800 37940 3332
rect 38556 800 38612 4732
rect 39228 4564 39284 5068
rect 39116 4452 39172 4462
rect 39116 4358 39172 4396
rect 38668 4338 38724 4350
rect 38668 4286 38670 4338
rect 38722 4286 38724 4338
rect 38668 3668 38724 4286
rect 39116 3780 39172 3790
rect 39116 3686 39172 3724
rect 38668 3602 38724 3612
rect 39228 3554 39284 4508
rect 39228 3502 39230 3554
rect 39282 3502 39284 3554
rect 39228 3490 39284 3502
rect 39564 3388 39620 8092
rect 39900 7700 39956 7710
rect 39900 7364 39956 7644
rect 39676 7362 39956 7364
rect 39676 7310 39902 7362
rect 39954 7310 39956 7362
rect 39676 7308 39956 7310
rect 39676 5010 39732 7308
rect 39900 7298 39956 7308
rect 40236 7474 40292 7486
rect 40236 7422 40238 7474
rect 40290 7422 40292 7474
rect 39676 4958 39678 5010
rect 39730 4958 39732 5010
rect 39676 4946 39732 4958
rect 39900 7028 39956 7038
rect 39452 3332 39620 3388
rect 39228 3276 39508 3332
rect 39228 800 39284 3276
rect 39900 800 39956 6972
rect 40124 6804 40180 6814
rect 40124 6710 40180 6748
rect 40124 6132 40180 6142
rect 40236 6132 40292 7422
rect 40460 6692 40516 6702
rect 40180 6076 40292 6132
rect 40348 6690 40516 6692
rect 40348 6638 40462 6690
rect 40514 6638 40516 6690
rect 40348 6636 40516 6638
rect 40124 6018 40180 6076
rect 40124 5966 40126 6018
rect 40178 5966 40180 6018
rect 40124 5236 40180 5966
rect 40124 5170 40180 5180
rect 40012 5010 40068 5022
rect 40012 4958 40014 5010
rect 40066 4958 40068 5010
rect 40012 4900 40068 4958
rect 40012 4834 40068 4844
rect 40348 4676 40404 6636
rect 40460 6626 40516 6636
rect 40460 5796 40516 5806
rect 40460 5702 40516 5740
rect 40236 4562 40292 4574
rect 40236 4510 40238 4562
rect 40290 4510 40292 4562
rect 40236 3556 40292 4510
rect 40348 3668 40404 4620
rect 40348 3602 40404 3612
rect 40572 5010 40628 5022
rect 40572 4958 40574 5010
rect 40626 4958 40628 5010
rect 40236 3490 40292 3500
rect 40572 3388 40628 4958
rect 40684 4900 40740 8206
rect 40796 8258 40852 8270
rect 40796 8206 40798 8258
rect 40850 8206 40852 8258
rect 40796 5908 40852 8206
rect 40908 7028 40964 10444
rect 41020 10434 41076 10444
rect 41020 9940 41076 9950
rect 41132 9940 41188 11452
rect 41020 9938 41188 9940
rect 41020 9886 41022 9938
rect 41074 9886 41188 9938
rect 41020 9884 41188 9886
rect 41020 9874 41076 9884
rect 41132 9268 41188 9884
rect 41356 11284 41412 11294
rect 41356 10610 41412 11228
rect 42140 11284 42196 12908
rect 42140 11218 42196 11228
rect 42252 11060 42308 16828
rect 42364 15148 42420 22316
rect 42476 22306 42532 22316
rect 42588 22260 42644 22270
rect 42476 21700 42532 21710
rect 42476 21606 42532 21644
rect 42476 18450 42532 18462
rect 42476 18398 42478 18450
rect 42530 18398 42532 18450
rect 42476 16884 42532 18398
rect 42476 16818 42532 16828
rect 42588 16994 42644 22204
rect 42588 16942 42590 16994
rect 42642 16942 42644 16994
rect 42588 16212 42644 16942
rect 42700 22148 42756 22158
rect 42700 16882 42756 22092
rect 42812 21924 42868 23212
rect 43372 22708 43428 22718
rect 43372 22482 43428 22652
rect 43372 22430 43374 22482
rect 43426 22430 43428 22482
rect 43372 22418 43428 22430
rect 42812 21858 42868 21868
rect 43260 21476 43316 21486
rect 43260 21382 43316 21420
rect 42924 21140 42980 21150
rect 42812 21084 42924 21140
rect 42812 20242 42868 21084
rect 42924 21074 42980 21084
rect 42812 20190 42814 20242
rect 42866 20190 42868 20242
rect 42812 20178 42868 20190
rect 42924 20804 42980 20814
rect 42924 20130 42980 20748
rect 43260 20802 43316 20814
rect 43260 20750 43262 20802
rect 43314 20750 43316 20802
rect 43036 20580 43092 20590
rect 43036 20578 43204 20580
rect 43036 20526 43038 20578
rect 43090 20526 43204 20578
rect 43036 20524 43204 20526
rect 43036 20514 43092 20524
rect 42924 20078 42926 20130
rect 42978 20078 42980 20130
rect 42700 16830 42702 16882
rect 42754 16830 42756 16882
rect 42700 16818 42756 16830
rect 42812 19348 42868 19358
rect 42588 16146 42644 16156
rect 42812 16100 42868 19292
rect 42924 19122 42980 20078
rect 42924 19070 42926 19122
rect 42978 19070 42980 19122
rect 42924 17666 42980 19070
rect 43036 20018 43092 20030
rect 43036 19966 43038 20018
rect 43090 19966 43092 20018
rect 43036 18676 43092 19966
rect 43036 18610 43092 18620
rect 43148 18228 43204 20524
rect 43260 19684 43316 20750
rect 43484 20132 43540 25230
rect 43596 25284 43652 25294
rect 43708 25284 43764 25564
rect 44044 25620 44100 25630
rect 44044 25526 44100 25564
rect 43652 25228 43764 25284
rect 44156 25508 44212 26238
rect 43596 25218 43652 25228
rect 44044 24948 44100 24958
rect 43820 24610 43876 24622
rect 43820 24558 43822 24610
rect 43874 24558 43876 24610
rect 43596 24276 43652 24286
rect 43596 23826 43652 24220
rect 43596 23774 43598 23826
rect 43650 23774 43652 23826
rect 43596 23762 43652 23774
rect 43708 24052 43764 24062
rect 43708 23826 43764 23996
rect 43708 23774 43710 23826
rect 43762 23774 43764 23826
rect 43708 23762 43764 23774
rect 43596 23380 43652 23390
rect 43596 23156 43652 23324
rect 43596 20468 43652 23100
rect 43820 22370 43876 24558
rect 44044 24276 44100 24892
rect 44156 24722 44212 25452
rect 44268 25172 44324 26460
rect 44380 26404 44436 26798
rect 44828 26740 44884 26750
rect 44604 26516 44660 26526
rect 44604 26422 44660 26460
rect 44380 26338 44436 26348
rect 44828 25844 44884 26684
rect 44940 26404 44996 26414
rect 44940 26310 44996 26348
rect 45052 26292 45108 26302
rect 45052 26198 45108 26236
rect 44828 25506 44884 25788
rect 44828 25454 44830 25506
rect 44882 25454 44884 25506
rect 44828 25442 44884 25454
rect 45388 25732 45444 25742
rect 44940 25396 44996 25406
rect 44268 25116 44660 25172
rect 44156 24670 44158 24722
rect 44210 24670 44212 24722
rect 44156 24658 44212 24670
rect 44380 24946 44436 24958
rect 44380 24894 44382 24946
rect 44434 24894 44436 24946
rect 44156 24276 44212 24286
rect 44044 24220 44156 24276
rect 44156 24050 44212 24220
rect 44156 23998 44158 24050
rect 44210 23998 44212 24050
rect 44156 23986 44212 23998
rect 43932 23716 43988 23726
rect 43932 23714 44100 23716
rect 43932 23662 43934 23714
rect 43986 23662 44100 23714
rect 43932 23660 44100 23662
rect 43932 23650 43988 23660
rect 44044 23156 44100 23660
rect 44268 23714 44324 23726
rect 44268 23662 44270 23714
rect 44322 23662 44324 23714
rect 44044 23090 44100 23100
rect 44156 23154 44212 23166
rect 44156 23102 44158 23154
rect 44210 23102 44212 23154
rect 44156 22596 44212 23102
rect 44268 22932 44324 23662
rect 44268 22866 44324 22876
rect 44156 22530 44212 22540
rect 44380 22484 44436 24894
rect 44268 22428 44436 22484
rect 44492 23266 44548 23278
rect 44492 23214 44494 23266
rect 44546 23214 44548 23266
rect 44268 22372 44324 22428
rect 43820 22318 43822 22370
rect 43874 22318 43876 22370
rect 43820 22148 43876 22318
rect 43820 22082 43876 22092
rect 44044 22316 44324 22372
rect 44044 21698 44100 22316
rect 44268 22148 44324 22158
rect 44268 22054 44324 22092
rect 44044 21646 44046 21698
rect 44098 21646 44100 21698
rect 44044 21634 44100 21646
rect 44156 21924 44212 21934
rect 43596 20402 43652 20412
rect 43708 20916 43764 20926
rect 43708 20188 43764 20860
rect 44156 20188 44212 21868
rect 44492 21476 44548 23214
rect 44492 21410 44548 21420
rect 44604 20188 44660 25116
rect 44940 24834 44996 25340
rect 44940 24782 44942 24834
rect 44994 24782 44996 24834
rect 44940 24770 44996 24782
rect 45276 24948 45332 24958
rect 45276 24722 45332 24892
rect 45276 24670 45278 24722
rect 45330 24670 45332 24722
rect 45276 24658 45332 24670
rect 45388 24052 45444 25676
rect 45500 24276 45556 30156
rect 45612 25284 45668 31164
rect 45724 31108 45780 31118
rect 45724 31014 45780 31052
rect 45836 30884 45892 32620
rect 46060 33122 46116 33134
rect 46060 33070 46062 33122
rect 46114 33070 46116 33122
rect 46060 32676 46116 33070
rect 46172 32676 46228 32686
rect 46060 32674 46228 32676
rect 46060 32622 46174 32674
rect 46226 32622 46228 32674
rect 46060 32620 46228 32622
rect 45948 31778 46004 31790
rect 45948 31726 45950 31778
rect 46002 31726 46004 31778
rect 45948 31668 46004 31726
rect 45948 31602 46004 31612
rect 45948 30996 46004 31006
rect 45948 30902 46004 30940
rect 45724 30828 45892 30884
rect 45724 25732 45780 30828
rect 46060 30772 46116 32620
rect 46172 32610 46228 32620
rect 46172 31780 46228 31790
rect 46172 31686 46228 31724
rect 46396 31666 46452 31678
rect 46396 31614 46398 31666
rect 46450 31614 46452 31666
rect 46396 31108 46452 31614
rect 46172 30996 46228 31006
rect 46172 30902 46228 30940
rect 45836 30716 46116 30772
rect 45836 30434 45892 30716
rect 45836 30382 45838 30434
rect 45890 30382 45892 30434
rect 45836 26290 45892 30382
rect 46172 30212 46228 30222
rect 46172 30118 46228 30156
rect 46396 30210 46452 31052
rect 46396 30158 46398 30210
rect 46450 30158 46452 30210
rect 46396 30146 46452 30158
rect 46620 31666 46676 31678
rect 46620 31614 46622 31666
rect 46674 31614 46676 31666
rect 46620 31106 46676 31614
rect 46620 31054 46622 31106
rect 46674 31054 46676 31106
rect 46620 30324 46676 31054
rect 46620 30210 46676 30268
rect 46620 30158 46622 30210
rect 46674 30158 46676 30210
rect 46620 30146 46676 30158
rect 46060 30100 46116 30110
rect 46060 30006 46116 30044
rect 46060 29876 46116 29886
rect 46060 26740 46116 29820
rect 46732 28196 46788 38612
rect 46956 35028 47012 35038
rect 46844 34916 46900 34926
rect 46844 34822 46900 34860
rect 46956 34914 47012 34972
rect 46956 34862 46958 34914
rect 47010 34862 47012 34914
rect 46956 34850 47012 34862
rect 47180 34914 47236 34926
rect 47180 34862 47182 34914
rect 47234 34862 47236 34914
rect 47068 34132 47124 34142
rect 47180 34132 47236 34862
rect 47124 34076 47236 34132
rect 46844 33346 46900 33358
rect 46844 33294 46846 33346
rect 46898 33294 46900 33346
rect 46844 30324 46900 33294
rect 47068 33234 47124 34076
rect 47068 33182 47070 33234
rect 47122 33182 47124 33234
rect 47068 33170 47124 33182
rect 47292 31108 47348 31118
rect 47292 31014 47348 31052
rect 46956 30994 47012 31006
rect 46956 30942 46958 30994
rect 47010 30942 47012 30994
rect 46956 30548 47012 30942
rect 47404 30994 47460 31006
rect 47404 30942 47406 30994
rect 47458 30942 47460 30994
rect 47068 30884 47124 30894
rect 47068 30790 47124 30828
rect 46956 30482 47012 30492
rect 47292 30324 47348 30334
rect 47404 30324 47460 30942
rect 46844 30268 47124 30324
rect 47068 30212 47124 30268
rect 47348 30268 47460 30324
rect 47068 30210 47236 30212
rect 47068 30158 47070 30210
rect 47122 30158 47236 30210
rect 47068 30156 47236 30158
rect 47068 30146 47124 30156
rect 46508 28140 46788 28196
rect 46172 27636 46228 27646
rect 46172 27074 46228 27580
rect 46396 27188 46452 27198
rect 46396 27094 46452 27132
rect 46172 27022 46174 27074
rect 46226 27022 46228 27074
rect 46172 27010 46228 27022
rect 46060 26674 46116 26684
rect 46508 26516 46564 28140
rect 47068 27074 47124 27086
rect 47068 27022 47070 27074
rect 47122 27022 47124 27074
rect 46620 26962 46676 26974
rect 46620 26910 46622 26962
rect 46674 26910 46676 26962
rect 46620 26908 46676 26910
rect 46844 26962 46900 26974
rect 46844 26910 46846 26962
rect 46898 26910 46900 26962
rect 46620 26852 46788 26908
rect 46508 26460 46676 26516
rect 46060 26404 46116 26414
rect 46060 26310 46116 26348
rect 45836 26238 45838 26290
rect 45890 26238 45892 26290
rect 45836 26068 45892 26238
rect 46284 26292 46340 26302
rect 46284 26198 46340 26236
rect 46508 26292 46564 26302
rect 46508 26198 46564 26236
rect 45836 26012 46452 26068
rect 45724 25666 45780 25676
rect 45724 25508 45780 25518
rect 45724 25414 45780 25452
rect 46284 25394 46340 25406
rect 46284 25342 46286 25394
rect 46338 25342 46340 25394
rect 45836 25284 45892 25294
rect 45612 25228 45780 25284
rect 45612 24722 45668 24734
rect 45612 24670 45614 24722
rect 45666 24670 45668 24722
rect 45612 24500 45668 24670
rect 45724 24724 45780 25228
rect 45836 25282 46228 25284
rect 45836 25230 45838 25282
rect 45890 25230 46228 25282
rect 45836 25228 46228 25230
rect 45836 25218 45892 25228
rect 45948 25060 46004 25070
rect 45948 24946 46004 25004
rect 45948 24894 45950 24946
rect 46002 24894 46004 24946
rect 45948 24882 46004 24894
rect 45724 24668 46004 24724
rect 45612 24434 45668 24444
rect 45500 24220 45892 24276
rect 45276 23996 45444 24052
rect 44828 23828 44884 23838
rect 44828 23734 44884 23772
rect 44940 23714 44996 23726
rect 45164 23716 45220 23726
rect 44940 23662 44942 23714
rect 44994 23662 44996 23714
rect 44940 23604 44996 23662
rect 44940 23538 44996 23548
rect 45052 23714 45220 23716
rect 45052 23662 45166 23714
rect 45218 23662 45220 23714
rect 45052 23660 45220 23662
rect 44828 23492 44884 23502
rect 44828 22708 44884 23436
rect 44828 22482 44884 22652
rect 44828 22430 44830 22482
rect 44882 22430 44884 22482
rect 44828 22418 44884 22430
rect 44940 22260 44996 22270
rect 44940 22166 44996 22204
rect 44940 21588 44996 21598
rect 45052 21588 45108 23660
rect 45164 23650 45220 23660
rect 45276 22596 45332 23996
rect 45388 23828 45444 23838
rect 45388 23734 45444 23772
rect 45500 23716 45556 23726
rect 45500 23622 45556 23660
rect 45724 23380 45780 23390
rect 45500 23378 45780 23380
rect 45500 23326 45726 23378
rect 45778 23326 45780 23378
rect 45500 23324 45780 23326
rect 45276 22530 45332 22540
rect 45388 22820 45444 22830
rect 45388 22370 45444 22764
rect 45388 22318 45390 22370
rect 45442 22318 45444 22370
rect 45388 22306 45444 22318
rect 44940 21586 45108 21588
rect 44940 21534 44942 21586
rect 44994 21534 45108 21586
rect 44940 21532 45108 21534
rect 44940 21522 44996 21532
rect 45276 21252 45332 21262
rect 44828 20804 44884 20814
rect 44828 20710 44884 20748
rect 45276 20802 45332 21196
rect 45276 20750 45278 20802
rect 45330 20750 45332 20802
rect 45276 20738 45332 20750
rect 43708 20132 44100 20188
rect 44156 20132 44436 20188
rect 43484 20066 43540 20076
rect 43932 19796 43988 19806
rect 43260 19628 43540 19684
rect 43372 19460 43428 19470
rect 43372 19234 43428 19404
rect 43372 19182 43374 19234
rect 43426 19182 43428 19234
rect 43372 19170 43428 19182
rect 43372 18564 43428 18574
rect 43484 18564 43540 19628
rect 43932 19346 43988 19740
rect 43932 19294 43934 19346
rect 43986 19294 43988 19346
rect 43932 19282 43988 19294
rect 43428 18508 43540 18564
rect 44044 18562 44100 20132
rect 44044 18510 44046 18562
rect 44098 18510 44100 18562
rect 43372 18498 43428 18508
rect 43932 18450 43988 18462
rect 43932 18398 43934 18450
rect 43986 18398 43988 18450
rect 43708 18228 43764 18238
rect 43148 18172 43316 18228
rect 42924 17614 42926 17666
rect 42978 17614 42980 17666
rect 42924 17602 42980 17614
rect 43148 18004 43204 18014
rect 43148 17666 43204 17948
rect 43148 17614 43150 17666
rect 43202 17614 43204 17666
rect 43148 17602 43204 17614
rect 43036 17444 43092 17454
rect 43036 17350 43092 17388
rect 43036 17108 43092 17118
rect 43036 16884 43092 17052
rect 43036 16818 43092 16828
rect 42700 16044 42868 16100
rect 42924 16772 42980 16782
rect 42476 15988 42532 15998
rect 42700 15988 42756 16044
rect 42476 15986 42756 15988
rect 42476 15934 42478 15986
rect 42530 15934 42756 15986
rect 42476 15932 42756 15934
rect 42476 15922 42532 15932
rect 42812 15876 42868 15886
rect 42924 15876 42980 16716
rect 42868 15820 42980 15876
rect 42812 15782 42868 15820
rect 43260 15540 43316 18172
rect 43708 18226 43876 18228
rect 43708 18174 43710 18226
rect 43762 18174 43876 18226
rect 43708 18172 43876 18174
rect 43708 18162 43764 18172
rect 43372 18116 43428 18126
rect 43372 16098 43428 18060
rect 43596 17668 43652 17678
rect 43372 16046 43374 16098
rect 43426 16046 43428 16098
rect 43372 16034 43428 16046
rect 43484 16324 43540 16334
rect 43484 15986 43540 16268
rect 43596 16100 43652 17612
rect 43708 16100 43764 16110
rect 43596 16098 43764 16100
rect 43596 16046 43710 16098
rect 43762 16046 43764 16098
rect 43596 16044 43764 16046
rect 43708 16034 43764 16044
rect 43484 15934 43486 15986
rect 43538 15934 43540 15986
rect 43484 15922 43540 15934
rect 43260 15484 43540 15540
rect 42924 15202 42980 15214
rect 42924 15150 42926 15202
rect 42978 15150 42980 15202
rect 42924 15148 42980 15150
rect 42364 15092 42644 15148
rect 42364 14420 42420 14430
rect 42364 13074 42420 14364
rect 42476 14308 42532 14318
rect 42476 14214 42532 14252
rect 42588 13412 42644 15092
rect 42812 15092 42980 15148
rect 42812 14642 42868 15092
rect 42812 14590 42814 14642
rect 42866 14590 42868 14642
rect 42812 14578 42868 14590
rect 43372 14644 43428 14654
rect 43372 14550 43428 14588
rect 42700 14532 42756 14542
rect 42700 14438 42756 14476
rect 43260 14420 43316 14430
rect 43260 14326 43316 14364
rect 42924 14306 42980 14318
rect 42924 14254 42926 14306
rect 42978 14254 42980 14306
rect 42924 14196 42980 14254
rect 42924 14130 42980 14140
rect 43260 14196 43316 14206
rect 42812 13636 42868 13646
rect 42812 13634 43204 13636
rect 42812 13582 42814 13634
rect 42866 13582 43204 13634
rect 42812 13580 43204 13582
rect 42812 13570 42868 13580
rect 43036 13412 43092 13422
rect 42588 13356 42868 13412
rect 42364 13022 42366 13074
rect 42418 13022 42420 13074
rect 42364 13010 42420 13022
rect 42588 12962 42644 12974
rect 42588 12910 42590 12962
rect 42642 12910 42644 12962
rect 42588 12404 42644 12910
rect 42588 12338 42644 12348
rect 41356 10558 41358 10610
rect 41410 10558 41412 10610
rect 41356 9826 41412 10558
rect 42028 11004 42308 11060
rect 42588 11060 42644 11070
rect 42644 11004 42756 11060
rect 42028 10276 42084 11004
rect 42588 10994 42644 11004
rect 42140 10500 42196 10510
rect 42140 10406 42196 10444
rect 42028 10220 42644 10276
rect 41356 9774 41358 9826
rect 41410 9774 41412 9826
rect 41356 9762 41412 9774
rect 42140 9716 42196 9726
rect 42140 9622 42196 9660
rect 41132 9202 41188 9212
rect 41020 9156 41076 9166
rect 41020 9042 41076 9100
rect 41356 9156 41412 9166
rect 41020 8990 41022 9042
rect 41074 8990 41076 9042
rect 41020 8978 41076 8990
rect 41132 9042 41188 9054
rect 41132 8990 41134 9042
rect 41186 8990 41188 9042
rect 41132 8484 41188 8990
rect 41132 8418 41188 8428
rect 41244 9042 41300 9054
rect 41244 8990 41246 9042
rect 41298 8990 41300 9042
rect 40908 6962 40964 6972
rect 41132 8146 41188 8158
rect 41132 8094 41134 8146
rect 41186 8094 41188 8146
rect 41132 6020 41188 8094
rect 41244 8036 41300 8990
rect 41244 7970 41300 7980
rect 41356 7812 41412 9100
rect 41244 7756 41412 7812
rect 41468 9042 41524 9054
rect 41468 8990 41470 9042
rect 41522 8990 41524 9042
rect 41244 7700 41300 7756
rect 41244 7586 41300 7644
rect 41468 7700 41524 8990
rect 41916 9044 41972 9054
rect 42140 9044 42196 9054
rect 41916 9042 42196 9044
rect 41916 8990 41918 9042
rect 41970 8990 42142 9042
rect 42194 8990 42196 9042
rect 41916 8988 42196 8990
rect 41916 8978 41972 8988
rect 42140 8978 42196 8988
rect 42588 8370 42644 10220
rect 42700 9154 42756 11004
rect 42700 9102 42702 9154
rect 42754 9102 42756 9154
rect 42700 9090 42756 9102
rect 42588 8318 42590 8370
rect 42642 8318 42644 8370
rect 42588 8306 42644 8318
rect 41804 8258 41860 8270
rect 41804 8206 41806 8258
rect 41858 8206 41860 8258
rect 41468 7634 41524 7644
rect 41580 8036 41636 8046
rect 41244 7534 41246 7586
rect 41298 7534 41300 7586
rect 41244 7522 41300 7534
rect 41580 7474 41636 7980
rect 41580 7422 41582 7474
rect 41634 7422 41636 7474
rect 41468 7364 41524 7374
rect 41468 6580 41524 7308
rect 41580 7140 41636 7422
rect 41580 7074 41636 7084
rect 41692 7588 41748 7598
rect 41580 6580 41636 6590
rect 41468 6578 41636 6580
rect 41468 6526 41582 6578
rect 41634 6526 41636 6578
rect 41468 6524 41636 6526
rect 41580 6514 41636 6524
rect 41132 5954 41188 5964
rect 40908 5908 40964 5918
rect 40796 5852 40908 5908
rect 40908 5842 40964 5852
rect 41020 5794 41076 5806
rect 41020 5742 41022 5794
rect 41074 5742 41076 5794
rect 41020 5684 41076 5742
rect 41020 5618 41076 5628
rect 41468 5794 41524 5806
rect 41468 5742 41470 5794
rect 41522 5742 41524 5794
rect 40684 4834 40740 4844
rect 41020 5012 41076 5022
rect 41468 5012 41524 5742
rect 41076 4956 41524 5012
rect 40908 4564 40964 4574
rect 40908 4470 40964 4508
rect 41020 4450 41076 4956
rect 41020 4398 41022 4450
rect 41074 4398 41076 4450
rect 41020 4386 41076 4398
rect 41132 4340 41188 4350
rect 41132 3444 41188 4284
rect 41468 4228 41524 4238
rect 41692 4228 41748 7532
rect 41468 4226 41748 4228
rect 41468 4174 41470 4226
rect 41522 4174 41748 4226
rect 41468 4172 41748 4174
rect 41356 3668 41412 3678
rect 41356 3554 41412 3612
rect 41356 3502 41358 3554
rect 41410 3502 41412 3554
rect 41356 3490 41412 3502
rect 41132 3388 41300 3444
rect 40460 3332 40628 3388
rect 40460 3266 40516 3276
rect 40572 2548 40628 2558
rect 40572 800 40628 2492
rect 41244 800 41300 3388
rect 41468 3442 41524 4172
rect 41804 3668 41860 8206
rect 42812 7700 42868 13356
rect 43036 12962 43092 13356
rect 43148 13074 43204 13580
rect 43148 13022 43150 13074
rect 43202 13022 43204 13074
rect 43148 13010 43204 13022
rect 43036 12910 43038 12962
rect 43090 12910 43092 12962
rect 43036 12898 43092 12910
rect 43260 12962 43316 14140
rect 43260 12910 43262 12962
rect 43314 12910 43316 12962
rect 43260 12898 43316 12910
rect 43484 12964 43540 15484
rect 43820 15148 43876 18172
rect 43932 17106 43988 18398
rect 43932 17054 43934 17106
rect 43986 17054 43988 17106
rect 43932 17042 43988 17054
rect 43932 16772 43988 16782
rect 44044 16772 44100 18510
rect 43988 16716 44100 16772
rect 44156 17780 44212 17790
rect 43932 16706 43988 16716
rect 43932 16548 43988 16558
rect 43932 16210 43988 16492
rect 43932 16158 43934 16210
rect 43986 16158 43988 16210
rect 43932 16146 43988 16158
rect 44044 15876 44100 15886
rect 44044 15782 44100 15820
rect 44156 15148 44212 17724
rect 43484 12898 43540 12908
rect 43708 15092 43876 15148
rect 43932 15092 44212 15148
rect 44268 16548 44324 16558
rect 44268 15204 44324 16492
rect 43372 10500 43428 10510
rect 43428 10444 43540 10500
rect 43372 10434 43428 10444
rect 43372 10164 43428 10174
rect 42924 9604 42980 9614
rect 42924 9042 42980 9548
rect 43372 9266 43428 10108
rect 43372 9214 43374 9266
rect 43426 9214 43428 9266
rect 43372 9202 43428 9214
rect 43484 9266 43540 10444
rect 43484 9214 43486 9266
rect 43538 9214 43540 9266
rect 43484 9202 43540 9214
rect 43596 9940 43652 9950
rect 43596 9268 43652 9884
rect 43596 9174 43652 9212
rect 42924 8990 42926 9042
rect 42978 8990 42980 9042
rect 42924 8978 42980 8990
rect 43596 8820 43652 8830
rect 42924 8484 42980 8494
rect 42924 8146 42980 8428
rect 43036 8260 43092 8270
rect 43036 8258 43204 8260
rect 43036 8206 43038 8258
rect 43090 8206 43204 8258
rect 43036 8204 43204 8206
rect 43036 8194 43092 8204
rect 42924 8094 42926 8146
rect 42978 8094 42980 8146
rect 42924 8036 42980 8094
rect 42924 7970 42980 7980
rect 42924 7700 42980 7710
rect 42812 7698 42980 7700
rect 42812 7646 42926 7698
rect 42978 7646 42980 7698
rect 42812 7644 42980 7646
rect 42924 7634 42980 7644
rect 43036 7700 43092 7710
rect 43036 7586 43092 7644
rect 43036 7534 43038 7586
rect 43090 7534 43092 7586
rect 41916 7474 41972 7486
rect 41916 7422 41918 7474
rect 41970 7422 41972 7474
rect 41916 7364 41972 7422
rect 41916 7298 41972 7308
rect 42252 7476 42308 7486
rect 42252 6802 42308 7420
rect 43036 7028 43092 7534
rect 43148 7140 43204 8204
rect 43596 8258 43652 8764
rect 43596 8206 43598 8258
rect 43650 8206 43652 8258
rect 43596 8194 43652 8206
rect 43708 7476 43764 15092
rect 43932 14642 43988 15092
rect 43932 14590 43934 14642
rect 43986 14590 43988 14642
rect 43932 14578 43988 14590
rect 44268 14642 44324 15148
rect 44268 14590 44270 14642
rect 44322 14590 44324 14642
rect 44268 14578 44324 14590
rect 43708 7410 43764 7420
rect 43820 13636 43876 13646
rect 43148 7074 43204 7084
rect 43036 6962 43092 6972
rect 42252 6750 42254 6802
rect 42306 6750 42308 6802
rect 42252 6738 42308 6750
rect 42588 6018 42644 6030
rect 42588 5966 42590 6018
rect 42642 5966 42644 6018
rect 42476 5908 42532 5918
rect 42252 5796 42308 5806
rect 42140 5794 42308 5796
rect 42140 5742 42254 5794
rect 42306 5742 42308 5794
rect 42140 5740 42308 5742
rect 41916 5348 41972 5358
rect 41916 5124 41972 5292
rect 42028 5124 42084 5134
rect 41916 5122 42084 5124
rect 41916 5070 42030 5122
rect 42082 5070 42084 5122
rect 41916 5068 42084 5070
rect 42028 5058 42084 5068
rect 41916 4340 41972 4350
rect 42140 4340 42196 5740
rect 42252 5730 42308 5740
rect 42476 5460 42532 5852
rect 41972 4284 42196 4340
rect 42252 5404 42476 5460
rect 42252 4338 42308 5404
rect 42476 5366 42532 5404
rect 42476 5124 42532 5134
rect 42476 5030 42532 5068
rect 42252 4286 42254 4338
rect 42306 4286 42308 4338
rect 41916 4246 41972 4284
rect 41804 3602 41860 3612
rect 41916 3892 41972 3902
rect 41468 3390 41470 3442
rect 41522 3390 41524 3442
rect 41468 3378 41524 3390
rect 41916 800 41972 3836
rect 42252 3444 42308 4286
rect 42588 3780 42644 5966
rect 42700 5796 42756 5806
rect 42756 5740 42868 5796
rect 42700 5730 42756 5740
rect 42812 4450 42868 5740
rect 43596 5010 43652 5022
rect 43596 4958 43598 5010
rect 43650 4958 43652 5010
rect 42812 4398 42814 4450
rect 42866 4398 42868 4450
rect 42812 4386 42868 4398
rect 42924 4898 42980 4910
rect 42924 4846 42926 4898
rect 42978 4846 42980 4898
rect 42588 3714 42644 3724
rect 42700 4116 42756 4126
rect 42252 3378 42308 3388
rect 42476 3556 42532 3566
rect 42476 3442 42532 3500
rect 42476 3390 42478 3442
rect 42530 3390 42532 3442
rect 42476 3378 42532 3390
rect 42700 3388 42756 4060
rect 42812 3780 42868 3790
rect 42812 3666 42868 3724
rect 42812 3614 42814 3666
rect 42866 3614 42868 3666
rect 42812 3602 42868 3614
rect 42924 3556 42980 4846
rect 43260 4340 43316 4350
rect 43036 3556 43092 3566
rect 42924 3554 43092 3556
rect 42924 3502 43038 3554
rect 43090 3502 43092 3554
rect 42924 3500 43092 3502
rect 42588 3332 42756 3388
rect 43036 3444 43092 3500
rect 43036 3378 43092 3388
rect 42588 800 42644 3332
rect 43260 800 43316 4284
rect 43596 4340 43652 4958
rect 43820 4562 43876 13580
rect 44380 11396 44436 20132
rect 44492 20132 44548 20142
rect 44604 20132 44884 20188
rect 44492 20038 44548 20076
rect 44716 20018 44772 20030
rect 44716 19966 44718 20018
rect 44770 19966 44772 20018
rect 44716 18452 44772 19966
rect 44828 19234 44884 20132
rect 44828 19182 44830 19234
rect 44882 19182 44884 19234
rect 44828 19170 44884 19182
rect 45388 19234 45444 19246
rect 45388 19182 45390 19234
rect 45442 19182 45444 19234
rect 44716 18386 44772 18396
rect 44828 18450 44884 18462
rect 44828 18398 44830 18450
rect 44882 18398 44884 18450
rect 44828 15876 44884 18398
rect 45276 18452 45332 18462
rect 45276 18358 45332 18396
rect 45052 17892 45108 17902
rect 44940 17780 44996 17790
rect 44940 17556 44996 17724
rect 44940 17490 44996 17500
rect 45052 16996 45108 17836
rect 45276 17780 45332 17790
rect 45276 17666 45332 17724
rect 45276 17614 45278 17666
rect 45330 17614 45332 17666
rect 45276 17602 45332 17614
rect 45388 17668 45444 19182
rect 45388 17602 45444 17612
rect 45052 16210 45108 16940
rect 45276 16996 45332 17006
rect 45276 16902 45332 16940
rect 45500 16436 45556 23324
rect 45724 23314 45780 23324
rect 45612 23156 45668 23166
rect 45612 23062 45668 23100
rect 45836 23044 45892 24220
rect 45836 22978 45892 22988
rect 45612 22146 45668 22158
rect 45612 22094 45614 22146
rect 45666 22094 45668 22146
rect 45612 21924 45668 22094
rect 45836 21924 45892 21934
rect 45612 21868 45836 21924
rect 45724 20802 45780 21868
rect 45836 21858 45892 21868
rect 45836 21588 45892 21598
rect 45836 21494 45892 21532
rect 45724 20750 45726 20802
rect 45778 20750 45780 20802
rect 45724 20738 45780 20750
rect 45052 16158 45054 16210
rect 45106 16158 45108 16210
rect 45052 16146 45108 16158
rect 45388 16380 45556 16436
rect 45724 20244 45780 20254
rect 44828 15810 44884 15820
rect 45388 15764 45444 16380
rect 45500 16212 45556 16222
rect 45500 16118 45556 16156
rect 45500 15764 45556 15774
rect 45388 15708 45500 15764
rect 45500 15698 45556 15708
rect 45388 15316 45444 15326
rect 45052 15314 45444 15316
rect 45052 15262 45390 15314
rect 45442 15262 45444 15314
rect 45052 15260 45444 15262
rect 44828 15204 44884 15214
rect 44828 11732 44884 15148
rect 45052 15202 45108 15260
rect 45388 15250 45444 15260
rect 45500 15316 45556 15326
rect 45052 15150 45054 15202
rect 45106 15150 45108 15202
rect 45052 15138 45108 15150
rect 45388 14980 45444 14990
rect 45388 13970 45444 14924
rect 45500 14532 45556 15260
rect 45500 14466 45556 14476
rect 45388 13918 45390 13970
rect 45442 13918 45444 13970
rect 45276 13748 45332 13758
rect 44940 13746 45332 13748
rect 44940 13694 45278 13746
rect 45330 13694 45332 13746
rect 44940 13692 45332 13694
rect 44940 13634 44996 13692
rect 45276 13682 45332 13692
rect 44940 13582 44942 13634
rect 44994 13582 44996 13634
rect 44940 13570 44996 13582
rect 45388 13524 45444 13918
rect 45388 13458 45444 13468
rect 44828 11676 45220 11732
rect 44156 11340 44436 11396
rect 44044 9716 44100 9726
rect 43932 9268 43988 9278
rect 43932 9174 43988 9212
rect 44044 9266 44100 9660
rect 44156 9492 44212 11340
rect 44828 11284 44884 11294
rect 44268 11282 44884 11284
rect 44268 11230 44830 11282
rect 44882 11230 44884 11282
rect 44268 11228 44884 11230
rect 44268 10498 44324 11228
rect 44828 11218 44884 11228
rect 44940 11172 44996 11182
rect 44940 11170 45108 11172
rect 44940 11118 44942 11170
rect 44994 11118 45108 11170
rect 44940 11116 45108 11118
rect 44940 11106 44996 11116
rect 45052 11060 45108 11116
rect 45052 10994 45108 11004
rect 44268 10446 44270 10498
rect 44322 10446 44324 10498
rect 44268 10434 44324 10446
rect 44268 9940 44324 9950
rect 44940 9940 44996 9950
rect 44268 9938 44996 9940
rect 44268 9886 44270 9938
rect 44322 9886 44942 9938
rect 44994 9886 44996 9938
rect 44268 9884 44996 9886
rect 44268 9874 44324 9884
rect 44940 9874 44996 9884
rect 44380 9604 44436 9614
rect 44156 9436 44324 9492
rect 44044 9214 44046 9266
rect 44098 9214 44100 9266
rect 44044 9202 44100 9214
rect 44156 9268 44212 9278
rect 44156 9174 44212 9212
rect 44268 8484 44324 9436
rect 44380 9266 44436 9548
rect 44380 9214 44382 9266
rect 44434 9214 44436 9266
rect 44380 9202 44436 9214
rect 44604 9324 45108 9380
rect 44268 8428 44436 8484
rect 44380 8260 44436 8428
rect 44380 8194 44436 8204
rect 44268 8146 44324 8158
rect 44268 8094 44270 8146
rect 44322 8094 44324 8146
rect 44156 8036 44212 8046
rect 43932 7476 43988 7486
rect 43932 7382 43988 7420
rect 44156 6578 44212 7980
rect 44268 7588 44324 8094
rect 44492 7588 44548 7598
rect 44324 7586 44548 7588
rect 44324 7534 44494 7586
rect 44546 7534 44548 7586
rect 44324 7532 44548 7534
rect 44268 7494 44324 7532
rect 44492 7522 44548 7532
rect 44604 7364 44660 9324
rect 44940 9156 44996 9166
rect 44940 9062 44996 9100
rect 45052 9154 45108 9324
rect 45052 9102 45054 9154
rect 45106 9102 45108 9154
rect 45052 9090 45108 9102
rect 44940 8820 44996 8830
rect 44940 8726 44996 8764
rect 44828 8034 44884 8046
rect 44828 7982 44830 8034
rect 44882 7982 44884 8034
rect 44828 7924 44884 7982
rect 44828 7858 44884 7868
rect 44268 7308 44660 7364
rect 44268 6804 44324 7308
rect 44268 6690 44324 6748
rect 44268 6638 44270 6690
rect 44322 6638 44324 6690
rect 44268 6626 44324 6638
rect 44380 6916 44436 6926
rect 44156 6526 44158 6578
rect 44210 6526 44212 6578
rect 44156 6514 44212 6526
rect 43820 4510 43822 4562
rect 43874 4510 43876 4562
rect 43820 4498 43876 4510
rect 44268 5908 44324 5918
rect 44268 5124 44324 5852
rect 43596 4274 43652 4284
rect 44268 4338 44324 5068
rect 44268 4286 44270 4338
rect 44322 4286 44324 4338
rect 43708 4228 43764 4238
rect 43708 3554 43764 4172
rect 44268 3780 44324 4286
rect 44268 3714 44324 3724
rect 43708 3502 43710 3554
rect 43762 3502 43764 3554
rect 43708 3490 43764 3502
rect 43932 3668 43988 3678
rect 43932 800 43988 3612
rect 44380 3442 44436 6860
rect 44940 6132 44996 6142
rect 45164 6132 45220 11676
rect 45612 11060 45668 11070
rect 45612 10164 45668 11004
rect 45276 9714 45332 9726
rect 45276 9662 45278 9714
rect 45330 9662 45332 9714
rect 45276 9268 45332 9662
rect 45276 9202 45332 9212
rect 45612 9266 45668 10108
rect 45724 9940 45780 20188
rect 45948 17666 46004 24668
rect 46060 23938 46116 23950
rect 46060 23886 46062 23938
rect 46114 23886 46116 23938
rect 46060 23716 46116 23886
rect 46060 23650 46116 23660
rect 46172 23492 46228 25228
rect 46284 25172 46340 25342
rect 46284 25106 46340 25116
rect 46396 24722 46452 26012
rect 46620 25620 46676 26460
rect 46732 26404 46788 26852
rect 46732 26310 46788 26348
rect 46844 26740 46900 26910
rect 47068 26964 47124 27022
rect 47068 26898 47124 26908
rect 46508 25564 46676 25620
rect 46844 26290 46900 26684
rect 46844 26238 46846 26290
rect 46898 26238 46900 26290
rect 46508 24948 46564 25564
rect 46620 25396 46676 25406
rect 46844 25396 46900 26238
rect 46956 26628 47012 26638
rect 46956 25732 47012 26572
rect 47180 26516 47236 30156
rect 47292 30098 47348 30268
rect 47292 30046 47294 30098
rect 47346 30046 47348 30098
rect 47292 30034 47348 30046
rect 47292 27076 47348 27086
rect 47292 26982 47348 27020
rect 47516 26962 47572 26974
rect 47516 26910 47518 26962
rect 47570 26910 47572 26962
rect 47516 26908 47572 26910
rect 47740 26962 47796 26974
rect 47740 26910 47742 26962
rect 47794 26910 47796 26962
rect 47516 26852 47684 26908
rect 47516 26516 47572 26526
rect 47180 26460 47348 26516
rect 47180 26292 47236 26302
rect 46956 25618 47012 25676
rect 47068 26290 47236 26292
rect 47068 26238 47182 26290
rect 47234 26238 47236 26290
rect 47068 26236 47236 26238
rect 47068 25730 47124 26236
rect 47180 26226 47236 26236
rect 47068 25678 47070 25730
rect 47122 25678 47124 25730
rect 47068 25666 47124 25678
rect 46956 25566 46958 25618
rect 47010 25566 47012 25618
rect 46956 25554 47012 25566
rect 46620 25394 46900 25396
rect 46620 25342 46622 25394
rect 46674 25342 46900 25394
rect 46620 25340 46900 25342
rect 46620 25330 46676 25340
rect 46508 24882 46564 24892
rect 46956 25172 47012 25182
rect 46396 24670 46398 24722
rect 46450 24670 46452 24722
rect 46396 24658 46452 24670
rect 46620 24834 46676 24846
rect 46620 24782 46622 24834
rect 46674 24782 46676 24834
rect 46508 23940 46564 23950
rect 46620 23940 46676 24782
rect 46956 24834 47012 25116
rect 47292 25172 47348 26460
rect 47516 26422 47572 26460
rect 47628 26404 47684 26852
rect 47628 26310 47684 26348
rect 47740 26740 47796 26910
rect 47740 26290 47796 26684
rect 47740 26238 47742 26290
rect 47794 26238 47796 26290
rect 47740 26226 47796 26238
rect 47516 25844 47572 25854
rect 47516 25618 47572 25788
rect 47516 25566 47518 25618
rect 47570 25566 47572 25618
rect 47516 25554 47572 25566
rect 47964 25732 48020 25742
rect 47964 25618 48020 25676
rect 47964 25566 47966 25618
rect 48018 25566 48020 25618
rect 47964 25554 48020 25566
rect 47292 25106 47348 25116
rect 48188 24948 48244 24958
rect 48188 24854 48244 24892
rect 48636 24948 48692 76300
rect 48860 76354 48916 76366
rect 48860 76302 48862 76354
rect 48914 76302 48916 76354
rect 48860 67228 48916 76302
rect 49084 75796 49140 75806
rect 49196 75796 49252 76636
rect 49644 76356 49700 76366
rect 49084 75794 49252 75796
rect 49084 75742 49086 75794
rect 49138 75742 49252 75794
rect 49084 75740 49252 75742
rect 49420 76354 49700 76356
rect 49420 76302 49646 76354
rect 49698 76302 49700 76354
rect 49420 76300 49700 76302
rect 49084 75730 49140 75740
rect 48860 67172 49140 67228
rect 49084 43708 49140 67172
rect 48860 43652 49140 43708
rect 48860 26740 48916 43652
rect 49420 38668 49476 76300
rect 49644 76290 49700 76300
rect 49532 75796 49588 75806
rect 49756 75796 49812 76748
rect 50092 76690 50148 76974
rect 50092 76638 50094 76690
rect 50146 76638 50148 76690
rect 49532 75794 49812 75796
rect 49532 75742 49534 75794
rect 49586 75742 49812 75794
rect 49532 75740 49812 75742
rect 49532 75730 49588 75740
rect 49756 75682 49812 75740
rect 49756 75630 49758 75682
rect 49810 75630 49812 75682
rect 49756 75618 49812 75630
rect 49980 76244 50036 76254
rect 49980 55468 50036 76188
rect 50092 75796 50148 76638
rect 50204 76692 50260 79200
rect 50876 77138 50932 79200
rect 50876 77086 50878 77138
rect 50930 77086 50932 77138
rect 50876 77074 50932 77086
rect 51548 77026 51604 79200
rect 51548 76974 51550 77026
rect 51602 76974 51604 77026
rect 51548 76962 51604 76974
rect 51772 77138 51828 77150
rect 51772 77086 51774 77138
rect 51826 77086 51828 77138
rect 50556 76860 50820 76870
rect 50612 76804 50660 76860
rect 50716 76804 50764 76860
rect 50556 76794 50820 76804
rect 50204 76626 50260 76636
rect 51212 76692 51268 76702
rect 50540 76356 50596 76366
rect 50540 76262 50596 76300
rect 50092 75730 50148 75740
rect 50764 75796 50820 75806
rect 50764 75702 50820 75740
rect 51212 75794 51268 76636
rect 51212 75742 51214 75794
rect 51266 75742 51268 75794
rect 51212 75730 51268 75742
rect 51660 76354 51716 76366
rect 51660 76302 51662 76354
rect 51714 76302 51716 76354
rect 50316 75684 50372 75694
rect 50316 75590 50372 75628
rect 50556 75292 50820 75302
rect 50612 75236 50660 75292
rect 50716 75236 50764 75292
rect 50556 75226 50820 75236
rect 50556 73724 50820 73734
rect 50612 73668 50660 73724
rect 50716 73668 50764 73724
rect 50556 73658 50820 73668
rect 50556 72156 50820 72166
rect 50612 72100 50660 72156
rect 50716 72100 50764 72156
rect 50556 72090 50820 72100
rect 50556 70588 50820 70598
rect 50612 70532 50660 70588
rect 50716 70532 50764 70588
rect 50556 70522 50820 70532
rect 50556 69020 50820 69030
rect 50612 68964 50660 69020
rect 50716 68964 50764 69020
rect 50556 68954 50820 68964
rect 50556 67452 50820 67462
rect 50612 67396 50660 67452
rect 50716 67396 50764 67452
rect 50556 67386 50820 67396
rect 50556 65884 50820 65894
rect 50612 65828 50660 65884
rect 50716 65828 50764 65884
rect 50556 65818 50820 65828
rect 50556 64316 50820 64326
rect 50612 64260 50660 64316
rect 50716 64260 50764 64316
rect 50556 64250 50820 64260
rect 50556 62748 50820 62758
rect 50612 62692 50660 62748
rect 50716 62692 50764 62748
rect 50556 62682 50820 62692
rect 50556 61180 50820 61190
rect 50612 61124 50660 61180
rect 50716 61124 50764 61180
rect 50556 61114 50820 61124
rect 50556 59612 50820 59622
rect 50612 59556 50660 59612
rect 50716 59556 50764 59612
rect 50556 59546 50820 59556
rect 50556 58044 50820 58054
rect 50612 57988 50660 58044
rect 50716 57988 50764 58044
rect 50556 57978 50820 57988
rect 50556 56476 50820 56486
rect 50612 56420 50660 56476
rect 50716 56420 50764 56476
rect 50556 56410 50820 56420
rect 48972 38612 49476 38668
rect 49532 55412 50036 55468
rect 48972 26852 49028 38612
rect 49532 29876 49588 55412
rect 50556 54908 50820 54918
rect 50612 54852 50660 54908
rect 50716 54852 50764 54908
rect 50556 54842 50820 54852
rect 50556 53340 50820 53350
rect 50612 53284 50660 53340
rect 50716 53284 50764 53340
rect 50556 53274 50820 53284
rect 50556 51772 50820 51782
rect 50612 51716 50660 51772
rect 50716 51716 50764 51772
rect 50556 51706 50820 51716
rect 50556 50204 50820 50214
rect 50612 50148 50660 50204
rect 50716 50148 50764 50204
rect 50556 50138 50820 50148
rect 50556 48636 50820 48646
rect 50612 48580 50660 48636
rect 50716 48580 50764 48636
rect 50556 48570 50820 48580
rect 50556 47068 50820 47078
rect 50612 47012 50660 47068
rect 50716 47012 50764 47068
rect 50556 47002 50820 47012
rect 50556 45500 50820 45510
rect 50612 45444 50660 45500
rect 50716 45444 50764 45500
rect 50556 45434 50820 45444
rect 50556 43932 50820 43942
rect 50612 43876 50660 43932
rect 50716 43876 50764 43932
rect 50556 43866 50820 43876
rect 50556 42364 50820 42374
rect 50612 42308 50660 42364
rect 50716 42308 50764 42364
rect 50556 42298 50820 42308
rect 50556 40796 50820 40806
rect 50612 40740 50660 40796
rect 50716 40740 50764 40796
rect 50556 40730 50820 40740
rect 50556 39228 50820 39238
rect 50612 39172 50660 39228
rect 50716 39172 50764 39228
rect 50556 39162 50820 39172
rect 50316 38724 50372 38734
rect 50204 38612 50372 38668
rect 51660 38724 51716 76302
rect 51772 75794 51828 77086
rect 52108 77138 52164 77150
rect 52108 77086 52110 77138
rect 52162 77086 52164 77138
rect 52108 76690 52164 77086
rect 52108 76638 52110 76690
rect 52162 76638 52164 76690
rect 52108 76626 52164 76638
rect 51772 75742 51774 75794
rect 51826 75742 51828 75794
rect 51772 75730 51828 75742
rect 52220 76580 52276 79200
rect 52892 76692 52948 79200
rect 52892 76626 52948 76636
rect 53004 77026 53060 77038
rect 53004 76974 53006 77026
rect 53058 76974 53060 77026
rect 53004 76690 53060 76974
rect 53004 76638 53006 76690
rect 53058 76638 53060 76690
rect 52220 76524 52724 76580
rect 52220 75794 52276 76524
rect 52220 75742 52222 75794
rect 52274 75742 52276 75794
rect 52220 75730 52276 75742
rect 52556 76354 52612 76366
rect 52556 76302 52558 76354
rect 52610 76302 52612 76354
rect 52556 55468 52612 76302
rect 52668 75682 52724 76524
rect 53004 76468 53060 76638
rect 52668 75630 52670 75682
rect 52722 75630 52724 75682
rect 52668 75618 52724 75630
rect 52780 76412 53060 76468
rect 52780 75122 52836 76412
rect 53452 76354 53508 76366
rect 53452 76302 53454 76354
rect 53506 76302 53508 76354
rect 52780 75070 52782 75122
rect 52834 75070 52836 75122
rect 52780 75058 52836 75070
rect 53228 75682 53284 75694
rect 53228 75630 53230 75682
rect 53282 75630 53284 75682
rect 52444 55412 52612 55468
rect 51996 40292 52052 40302
rect 51660 38658 51716 38668
rect 51884 40068 51940 40078
rect 51884 39060 51940 40012
rect 49532 29810 49588 29820
rect 49868 30324 49924 30334
rect 49308 28644 49364 28654
rect 49084 27076 49140 27086
rect 49084 26982 49140 27020
rect 49196 26852 49252 26862
rect 49308 26852 49364 28588
rect 49644 27188 49700 27198
rect 49644 27074 49700 27132
rect 49644 27022 49646 27074
rect 49698 27022 49700 27074
rect 49644 27010 49700 27022
rect 49756 26964 49812 27002
rect 49756 26898 49812 26908
rect 48972 26796 49140 26852
rect 48860 26674 48916 26684
rect 48860 26404 48916 26414
rect 48860 26310 48916 26348
rect 48748 26292 48804 26302
rect 48748 26198 48804 26236
rect 48860 26068 48916 26078
rect 48860 26066 49028 26068
rect 48860 26014 48862 26066
rect 48914 26014 49028 26066
rect 48860 26012 49028 26014
rect 48860 26002 48916 26012
rect 48636 24882 48692 24892
rect 46956 24782 46958 24834
rect 47010 24782 47012 24834
rect 46956 24770 47012 24782
rect 47292 24834 47348 24846
rect 47292 24782 47294 24834
rect 47346 24782 47348 24834
rect 47292 24052 47348 24782
rect 46508 23938 46676 23940
rect 46508 23886 46510 23938
rect 46562 23886 46676 23938
rect 46508 23884 46676 23886
rect 46508 23874 46564 23884
rect 46396 23716 46452 23726
rect 46396 23622 46452 23660
rect 46172 23436 46564 23492
rect 46508 23266 46564 23436
rect 46508 23214 46510 23266
rect 46562 23214 46564 23266
rect 46508 23202 46564 23214
rect 46060 23156 46116 23166
rect 46396 23156 46452 23166
rect 46116 23100 46228 23156
rect 46060 23090 46116 23100
rect 46060 22932 46116 22942
rect 46060 22370 46116 22876
rect 46060 22318 46062 22370
rect 46114 22318 46116 22370
rect 46060 22306 46116 22318
rect 46172 22148 46228 23100
rect 46060 22092 46228 22148
rect 46284 23044 46340 23054
rect 46060 18452 46116 22092
rect 46172 21698 46228 21710
rect 46172 21646 46174 21698
rect 46226 21646 46228 21698
rect 46172 21588 46228 21646
rect 46172 21522 46228 21532
rect 46060 18386 46116 18396
rect 46172 20914 46228 20926
rect 46172 20862 46174 20914
rect 46226 20862 46228 20914
rect 45948 17614 45950 17666
rect 46002 17614 46004 17666
rect 45836 16324 45892 16334
rect 45836 16210 45892 16268
rect 45836 16158 45838 16210
rect 45890 16158 45892 16210
rect 45836 16146 45892 16158
rect 45724 9874 45780 9884
rect 45836 15764 45892 15774
rect 45836 9604 45892 15708
rect 45948 14756 46004 17614
rect 46060 17778 46116 17790
rect 46060 17726 46062 17778
rect 46114 17726 46116 17778
rect 46060 14980 46116 17726
rect 46172 17556 46228 20862
rect 46284 20188 46340 22988
rect 46396 22146 46452 23100
rect 46508 22372 46564 22382
rect 46620 22372 46676 23884
rect 46508 22370 46620 22372
rect 46508 22318 46510 22370
rect 46562 22318 46620 22370
rect 46508 22316 46620 22318
rect 46508 22306 46564 22316
rect 46620 22278 46676 22316
rect 46732 23996 47348 24052
rect 47740 24724 47796 24734
rect 46732 23938 46788 23996
rect 46732 23886 46734 23938
rect 46786 23886 46788 23938
rect 46732 22370 46788 23886
rect 47180 23884 47572 23940
rect 47068 23826 47124 23838
rect 47068 23774 47070 23826
rect 47122 23774 47124 23826
rect 47068 23716 47124 23774
rect 47180 23826 47236 23884
rect 47180 23774 47182 23826
rect 47234 23774 47236 23826
rect 47180 23762 47236 23774
rect 47404 23716 47460 23726
rect 47068 23650 47124 23660
rect 47292 23714 47460 23716
rect 47292 23662 47406 23714
rect 47458 23662 47460 23714
rect 47292 23660 47460 23662
rect 47180 23380 47236 23390
rect 47180 23286 47236 23324
rect 47068 22708 47124 22718
rect 47068 22484 47124 22652
rect 46732 22318 46734 22370
rect 46786 22318 46788 22370
rect 46396 22094 46398 22146
rect 46450 22094 46452 22146
rect 46396 22082 46452 22094
rect 46732 22036 46788 22318
rect 46956 22428 47124 22484
rect 46956 22036 47012 22428
rect 47292 22372 47348 23660
rect 47404 23650 47460 23660
rect 47516 23716 47572 23884
rect 47516 23650 47572 23660
rect 47628 23826 47684 23838
rect 47628 23774 47630 23826
rect 47682 23774 47684 23826
rect 47516 23266 47572 23278
rect 47516 23214 47518 23266
rect 47570 23214 47572 23266
rect 47516 22708 47572 23214
rect 47516 22642 47572 22652
rect 47628 22596 47684 23774
rect 47740 23826 47796 24668
rect 48860 24724 48916 24734
rect 48860 24630 48916 24668
rect 47852 24610 47908 24622
rect 47852 24558 47854 24610
rect 47906 24558 47908 24610
rect 47852 23940 47908 24558
rect 48300 24276 48356 24286
rect 48300 24050 48356 24220
rect 48300 23998 48302 24050
rect 48354 23998 48356 24050
rect 48300 23986 48356 23998
rect 47852 23874 47908 23884
rect 47740 23774 47742 23826
rect 47794 23774 47796 23826
rect 47740 23762 47796 23774
rect 48748 23828 48804 23838
rect 48748 23734 48804 23772
rect 47964 23716 48020 23726
rect 47852 23714 48020 23716
rect 47852 23662 47966 23714
rect 48018 23662 48020 23714
rect 47852 23660 48020 23662
rect 47852 23380 47908 23660
rect 47964 23650 48020 23660
rect 47740 23324 47908 23380
rect 47740 22708 47796 23324
rect 47964 23268 48020 23278
rect 47964 23266 48132 23268
rect 47964 23214 47966 23266
rect 48018 23214 48132 23266
rect 47964 23212 48132 23214
rect 47964 23202 48020 23212
rect 47852 23156 47908 23166
rect 47852 23062 47908 23100
rect 48076 23044 48132 23212
rect 48188 23156 48244 23166
rect 48860 23156 48916 23166
rect 48188 23154 48468 23156
rect 48188 23102 48190 23154
rect 48242 23102 48468 23154
rect 48188 23100 48468 23102
rect 48188 23090 48244 23100
rect 48076 22978 48132 22988
rect 48076 22708 48132 22718
rect 47740 22652 47908 22708
rect 47628 22540 47796 22596
rect 47180 22316 47348 22372
rect 47404 22372 47460 22382
rect 47068 22260 47124 22270
rect 47068 22166 47124 22204
rect 46956 21980 47124 22036
rect 46732 21970 46788 21980
rect 46956 21588 47012 21598
rect 46620 21476 46676 21486
rect 46620 21382 46676 21420
rect 46508 21364 46564 21374
rect 46508 20242 46564 21308
rect 46508 20190 46510 20242
rect 46562 20190 46564 20242
rect 46284 20132 46452 20188
rect 46508 20178 46564 20190
rect 46620 20804 46676 20814
rect 46620 20188 46676 20748
rect 46620 20132 46788 20188
rect 46172 17462 46228 17500
rect 46284 18452 46340 18462
rect 46396 18452 46452 20132
rect 46620 20020 46676 20030
rect 46620 18900 46676 19964
rect 46620 18834 46676 18844
rect 46620 18452 46676 18462
rect 46396 18396 46620 18452
rect 46172 16100 46228 16110
rect 46172 16006 46228 16044
rect 46172 15540 46228 15550
rect 46284 15540 46340 18396
rect 46172 15538 46340 15540
rect 46172 15486 46174 15538
rect 46226 15486 46340 15538
rect 46172 15484 46340 15486
rect 46396 16996 46452 17006
rect 46396 16882 46452 16940
rect 46396 16830 46398 16882
rect 46450 16830 46452 16882
rect 46172 15474 46228 15484
rect 46396 15148 46452 16830
rect 46508 15874 46564 15886
rect 46508 15822 46510 15874
rect 46562 15822 46564 15874
rect 46508 15540 46564 15822
rect 46508 15474 46564 15484
rect 46620 15538 46676 18396
rect 46732 18452 46788 20132
rect 46956 20130 47012 21532
rect 47068 21252 47124 21980
rect 47068 21186 47124 21196
rect 47180 21028 47236 22316
rect 47404 22278 47460 22316
rect 47516 22370 47572 22382
rect 47516 22318 47518 22370
rect 47570 22318 47572 22370
rect 47292 22148 47348 22158
rect 47292 22054 47348 22092
rect 47404 22036 47460 22046
rect 47516 22036 47572 22318
rect 47460 21980 47572 22036
rect 47628 22036 47684 22046
rect 47404 21586 47460 21980
rect 47404 21534 47406 21586
rect 47458 21534 47460 21586
rect 47404 21522 47460 21534
rect 47628 21586 47684 21980
rect 47740 21810 47796 22540
rect 47740 21758 47742 21810
rect 47794 21758 47796 21810
rect 47740 21746 47796 21758
rect 47628 21534 47630 21586
rect 47682 21534 47684 21586
rect 47628 21522 47684 21534
rect 47852 21364 47908 22652
rect 47964 22258 48020 22270
rect 47964 22206 47966 22258
rect 48018 22206 48020 22258
rect 47964 22148 48020 22206
rect 48076 22258 48132 22652
rect 48076 22206 48078 22258
rect 48130 22206 48132 22258
rect 48076 22194 48132 22206
rect 48300 22148 48356 22158
rect 47964 22082 48020 22092
rect 48188 22146 48356 22148
rect 48188 22094 48302 22146
rect 48354 22094 48356 22146
rect 48188 22092 48356 22094
rect 47516 21308 47908 21364
rect 47964 21586 48020 21598
rect 47964 21534 47966 21586
rect 48018 21534 48020 21586
rect 47516 21140 47572 21308
rect 47180 20962 47236 20972
rect 47404 21084 47572 21140
rect 47068 20914 47124 20926
rect 47068 20862 47070 20914
rect 47122 20862 47124 20914
rect 47068 20188 47124 20862
rect 47180 20804 47236 20814
rect 47180 20710 47236 20748
rect 47404 20188 47460 21084
rect 47740 21028 47796 21038
rect 47796 20972 47908 21028
rect 47740 20962 47796 20972
rect 47068 20132 47236 20188
rect 46956 20078 46958 20130
rect 47010 20078 47012 20130
rect 46956 19122 47012 20078
rect 47068 19908 47124 19918
rect 47068 19234 47124 19852
rect 47068 19182 47070 19234
rect 47122 19182 47124 19234
rect 47068 19170 47124 19182
rect 46956 19070 46958 19122
rect 47010 19070 47012 19122
rect 46956 19058 47012 19070
rect 46844 19010 46900 19022
rect 46844 18958 46846 19010
rect 46898 18958 46900 19010
rect 46844 18676 46900 18958
rect 46844 18610 46900 18620
rect 46956 18674 47012 18686
rect 46956 18622 46958 18674
rect 47010 18622 47012 18674
rect 46844 18452 46900 18462
rect 46732 18450 46900 18452
rect 46732 18398 46846 18450
rect 46898 18398 46900 18450
rect 46732 18396 46900 18398
rect 46732 17780 46788 18396
rect 46844 18386 46900 18396
rect 46732 16882 46788 17724
rect 46956 17554 47012 18622
rect 46956 17502 46958 17554
rect 47010 17502 47012 17554
rect 46956 17490 47012 17502
rect 46732 16830 46734 16882
rect 46786 16830 46788 16882
rect 46732 16818 46788 16830
rect 47180 15986 47236 20132
rect 47292 20132 47460 20188
rect 47740 20690 47796 20702
rect 47740 20638 47742 20690
rect 47794 20638 47796 20690
rect 47292 17666 47348 20132
rect 47516 18564 47572 18574
rect 47740 18564 47796 20638
rect 47516 18562 47796 18564
rect 47516 18510 47518 18562
rect 47570 18510 47796 18562
rect 47516 18508 47796 18510
rect 47404 18452 47460 18462
rect 47404 18358 47460 18396
rect 47292 17614 47294 17666
rect 47346 17614 47348 17666
rect 47292 17602 47348 17614
rect 47404 18004 47460 18014
rect 47180 15934 47182 15986
rect 47234 15934 47236 15986
rect 47180 15922 47236 15934
rect 47292 16884 47348 16894
rect 46620 15486 46622 15538
rect 46674 15486 46676 15538
rect 46620 15474 46676 15486
rect 47180 15764 47236 15774
rect 47180 15540 47236 15708
rect 47180 15446 47236 15484
rect 47292 15148 47348 16828
rect 47404 15428 47460 17948
rect 47516 17556 47572 18508
rect 47516 16994 47572 17500
rect 47516 16942 47518 16994
rect 47570 16942 47572 16994
rect 47516 16930 47572 16942
rect 47404 15362 47460 15372
rect 47740 16770 47796 16782
rect 47740 16718 47742 16770
rect 47794 16718 47796 16770
rect 47740 15428 47796 16718
rect 47852 16098 47908 20972
rect 47964 20244 48020 21534
rect 48076 21588 48132 21598
rect 48076 20468 48132 21532
rect 48188 20580 48244 22092
rect 48300 22082 48356 22092
rect 48300 21812 48356 21822
rect 48300 20802 48356 21756
rect 48300 20750 48302 20802
rect 48354 20750 48356 20802
rect 48300 20738 48356 20750
rect 48188 20524 48356 20580
rect 48076 20412 48244 20468
rect 48076 20244 48132 20254
rect 47964 20242 48132 20244
rect 47964 20190 48078 20242
rect 48130 20190 48132 20242
rect 47964 20188 48132 20190
rect 48076 20178 48132 20188
rect 48188 19908 48244 20412
rect 48188 19814 48244 19852
rect 47852 16046 47854 16098
rect 47906 16046 47908 16098
rect 47852 16034 47908 16046
rect 47964 15876 48020 15886
rect 47740 15362 47796 15372
rect 47852 15874 48020 15876
rect 47852 15822 47966 15874
rect 48018 15822 48020 15874
rect 47852 15820 48020 15822
rect 47740 15204 47796 15214
rect 46396 15092 46676 15148
rect 47292 15092 47684 15148
rect 46060 14924 46564 14980
rect 45948 14700 46340 14756
rect 46284 14642 46340 14700
rect 46284 14590 46286 14642
rect 46338 14590 46340 14642
rect 46284 14578 46340 14590
rect 46508 14530 46564 14924
rect 46508 14478 46510 14530
rect 46562 14478 46564 14530
rect 46508 14466 46564 14478
rect 46620 13636 46676 15092
rect 47628 14308 47684 15092
rect 47740 14530 47796 15148
rect 47740 14478 47742 14530
rect 47794 14478 47796 14530
rect 47740 14466 47796 14478
rect 47852 14532 47908 15820
rect 47964 15810 48020 15820
rect 47964 15540 48020 15550
rect 47964 15446 48020 15484
rect 48300 15204 48356 20524
rect 48412 20356 48468 23100
rect 48860 23062 48916 23100
rect 48748 22930 48804 22942
rect 48748 22878 48750 22930
rect 48802 22878 48804 22930
rect 48636 22482 48692 22494
rect 48636 22430 48638 22482
rect 48690 22430 48692 22482
rect 48636 21700 48692 22430
rect 48748 21812 48804 22878
rect 48748 21746 48804 21756
rect 48860 21810 48916 21822
rect 48860 21758 48862 21810
rect 48914 21758 48916 21810
rect 48412 20290 48468 20300
rect 48524 20804 48580 20814
rect 48524 19346 48580 20748
rect 48636 20690 48692 21644
rect 48748 21586 48804 21598
rect 48748 21534 48750 21586
rect 48802 21534 48804 21586
rect 48748 20804 48804 21534
rect 48748 20738 48804 20748
rect 48636 20638 48638 20690
rect 48690 20638 48692 20690
rect 48636 20626 48692 20638
rect 48860 20188 48916 21758
rect 48524 19294 48526 19346
rect 48578 19294 48580 19346
rect 48524 19282 48580 19294
rect 48748 20132 48916 20188
rect 48748 18564 48804 20132
rect 48860 20020 48916 20030
rect 48860 19926 48916 19964
rect 48860 18564 48916 18574
rect 48748 18562 48916 18564
rect 48748 18510 48862 18562
rect 48914 18510 48916 18562
rect 48748 18508 48916 18510
rect 48860 18498 48916 18508
rect 48972 18450 49028 26012
rect 49084 22372 49140 26796
rect 49196 26850 49364 26852
rect 49196 26798 49198 26850
rect 49250 26798 49364 26850
rect 49196 26796 49364 26798
rect 49420 26852 49476 26862
rect 49420 26850 49700 26852
rect 49420 26798 49422 26850
rect 49474 26798 49700 26850
rect 49420 26796 49700 26798
rect 49196 26786 49252 26796
rect 49420 26786 49476 26796
rect 49196 26628 49252 26638
rect 49196 23042 49252 26572
rect 49308 26516 49364 26526
rect 49532 26516 49588 26526
rect 49308 26402 49364 26460
rect 49308 26350 49310 26402
rect 49362 26350 49364 26402
rect 49308 26338 49364 26350
rect 49420 26460 49532 26516
rect 49420 26402 49476 26460
rect 49532 26450 49588 26460
rect 49420 26350 49422 26402
rect 49474 26350 49476 26402
rect 49420 26338 49476 26350
rect 49420 26068 49476 26078
rect 49420 26066 49588 26068
rect 49420 26014 49422 26066
rect 49474 26014 49588 26066
rect 49420 26012 49588 26014
rect 49420 26002 49476 26012
rect 49308 23716 49364 23726
rect 49308 23714 49476 23716
rect 49308 23662 49310 23714
rect 49362 23662 49476 23714
rect 49308 23660 49476 23662
rect 49308 23650 49364 23660
rect 49420 23604 49476 23660
rect 49196 22990 49198 23042
rect 49250 22990 49252 23042
rect 49196 22978 49252 22990
rect 49308 23042 49364 23054
rect 49308 22990 49310 23042
rect 49362 22990 49364 23042
rect 49308 22820 49364 22990
rect 49420 22932 49476 23548
rect 49420 22866 49476 22876
rect 49308 22754 49364 22764
rect 49420 22372 49476 22382
rect 49084 22306 49140 22316
rect 49196 22370 49476 22372
rect 49196 22318 49422 22370
rect 49474 22318 49476 22370
rect 49196 22316 49476 22318
rect 49084 22146 49140 22158
rect 49084 22094 49086 22146
rect 49138 22094 49140 22146
rect 49084 21924 49140 22094
rect 49084 21588 49140 21868
rect 49084 21522 49140 21532
rect 49196 20804 49252 22316
rect 49420 22306 49476 22316
rect 49420 22148 49476 22158
rect 49420 21586 49476 22092
rect 49420 21534 49422 21586
rect 49474 21534 49476 21586
rect 49420 21522 49476 21534
rect 49532 21028 49588 26012
rect 49644 23940 49700 26796
rect 49644 23884 49812 23940
rect 49644 23716 49700 23726
rect 49644 23622 49700 23660
rect 49756 21364 49812 23884
rect 49868 23716 49924 30268
rect 50092 29204 50148 29214
rect 49868 23650 49924 23660
rect 49980 26850 50036 26862
rect 49980 26798 49982 26850
rect 50034 26798 50036 26850
rect 49980 23548 50036 26798
rect 50092 26514 50148 29148
rect 50092 26462 50094 26514
rect 50146 26462 50148 26514
rect 50092 26404 50148 26462
rect 50092 26338 50148 26348
rect 50204 26908 50260 38612
rect 50556 37660 50820 37670
rect 50612 37604 50660 37660
rect 50716 37604 50764 37660
rect 50556 37594 50820 37604
rect 50556 36092 50820 36102
rect 50612 36036 50660 36092
rect 50716 36036 50764 36092
rect 50556 36026 50820 36036
rect 50556 34524 50820 34534
rect 50612 34468 50660 34524
rect 50716 34468 50764 34524
rect 50556 34458 50820 34468
rect 50556 32956 50820 32966
rect 50612 32900 50660 32956
rect 50716 32900 50764 32956
rect 50556 32890 50820 32900
rect 51324 32004 51380 32014
rect 51100 31780 51156 31790
rect 51100 31686 51156 31724
rect 50556 31388 50820 31398
rect 50612 31332 50660 31388
rect 50716 31332 50764 31388
rect 50556 31322 50820 31332
rect 50316 31108 50372 31118
rect 50316 31014 50372 31052
rect 50540 30994 50596 31006
rect 50540 30942 50542 30994
rect 50594 30942 50596 30994
rect 50540 30884 50596 30942
rect 51100 30996 51156 31006
rect 51100 30902 51156 30940
rect 50540 30818 50596 30828
rect 50764 30884 50820 30894
rect 50764 30882 50932 30884
rect 50764 30830 50766 30882
rect 50818 30830 50932 30882
rect 50764 30828 50932 30830
rect 50764 30818 50820 30828
rect 50652 30212 50708 30222
rect 50652 30118 50708 30156
rect 50764 30100 50820 30110
rect 50764 30006 50820 30044
rect 50556 29820 50820 29830
rect 50612 29764 50660 29820
rect 50716 29764 50764 29820
rect 50556 29754 50820 29764
rect 50316 29428 50372 29438
rect 50316 28644 50372 29372
rect 50316 27186 50372 28588
rect 50316 27134 50318 27186
rect 50370 27134 50372 27186
rect 50316 27122 50372 27134
rect 50428 29316 50484 29326
rect 50204 26796 50372 26908
rect 50204 26068 50260 26796
rect 50428 26516 50484 29260
rect 50556 28252 50820 28262
rect 50612 28196 50660 28252
rect 50716 28196 50764 28252
rect 50556 28186 50820 28196
rect 50876 27524 50932 30828
rect 51212 30772 51268 30782
rect 51212 30678 51268 30716
rect 51324 30324 51380 31948
rect 51436 31892 51492 31902
rect 51436 31666 51492 31836
rect 51436 31614 51438 31666
rect 51490 31614 51492 31666
rect 51436 31602 51492 31614
rect 51660 31554 51716 31566
rect 51660 31502 51662 31554
rect 51714 31502 51716 31554
rect 51436 31220 51492 31230
rect 51436 31106 51492 31164
rect 51436 31054 51438 31106
rect 51490 31054 51492 31106
rect 51436 31042 51492 31054
rect 50876 27458 50932 27468
rect 51212 30268 51380 30324
rect 50764 27188 50820 27198
rect 50764 27094 50820 27132
rect 51212 27188 51268 30268
rect 51324 30100 51380 30110
rect 51324 30098 51604 30100
rect 51324 30046 51326 30098
rect 51378 30046 51604 30098
rect 51324 30044 51604 30046
rect 51324 30034 51380 30044
rect 51212 27122 51268 27132
rect 51324 27524 51380 27534
rect 51212 26740 51268 26750
rect 50556 26684 50820 26694
rect 50612 26628 50660 26684
rect 50716 26628 50764 26684
rect 50556 26618 50820 26628
rect 50988 26684 51212 26740
rect 50540 26516 50596 26526
rect 50484 26514 50596 26516
rect 50484 26462 50542 26514
rect 50594 26462 50596 26514
rect 50484 26460 50596 26462
rect 50428 26422 50484 26460
rect 50540 26450 50596 26460
rect 50204 26012 50372 26068
rect 49980 23492 50148 23548
rect 50092 23426 50148 23436
rect 49868 23044 49924 23054
rect 49868 22950 49924 22988
rect 50204 23042 50260 23054
rect 50204 22990 50206 23042
rect 50258 22990 50260 23042
rect 50204 22930 50260 22990
rect 50204 22878 50206 22930
rect 50258 22878 50260 22930
rect 50204 22866 50260 22878
rect 49868 22596 49924 22606
rect 49924 22540 50036 22596
rect 49868 22530 49924 22540
rect 49980 22370 50036 22540
rect 49980 22318 49982 22370
rect 50034 22318 50036 22370
rect 49980 22306 50036 22318
rect 49868 21700 49924 21710
rect 49868 21606 49924 21644
rect 50204 21588 50260 21598
rect 50092 21586 50260 21588
rect 50092 21534 50206 21586
rect 50258 21534 50260 21586
rect 50092 21532 50260 21534
rect 49756 21308 50036 21364
rect 49196 20738 49252 20748
rect 49308 20972 49588 21028
rect 49196 20578 49252 20590
rect 49196 20526 49198 20578
rect 49250 20526 49252 20578
rect 49196 20188 49252 20526
rect 48972 18398 48974 18450
rect 49026 18398 49028 18450
rect 48972 18386 49028 18398
rect 49084 20132 49252 20188
rect 48748 17666 48804 17678
rect 48748 17614 48750 17666
rect 48802 17614 48804 17666
rect 48300 15138 48356 15148
rect 48412 17442 48468 17454
rect 48412 17390 48414 17442
rect 48466 17390 48468 17442
rect 47852 14476 48356 14532
rect 47628 14252 48132 14308
rect 48076 13970 48132 14252
rect 48076 13918 48078 13970
rect 48130 13918 48132 13970
rect 48076 13906 48132 13918
rect 48188 14306 48244 14318
rect 48188 14254 48190 14306
rect 48242 14254 48244 14306
rect 46620 13542 46676 13580
rect 45836 9538 45892 9548
rect 46956 9828 47012 9838
rect 45612 9214 45614 9266
rect 45666 9214 45668 9266
rect 45612 9202 45668 9214
rect 46060 9268 46116 9278
rect 46060 9174 46116 9212
rect 45276 8370 45332 8382
rect 45276 8318 45278 8370
rect 45330 8318 45332 8370
rect 45276 8260 45332 8318
rect 45276 8194 45332 8204
rect 45948 8034 46004 8046
rect 45948 7982 45950 8034
rect 46002 7982 46004 8034
rect 45948 7924 46004 7982
rect 45948 7858 46004 7868
rect 46284 8034 46340 8046
rect 46284 7982 46286 8034
rect 46338 7982 46340 8034
rect 46060 7586 46116 7598
rect 46060 7534 46062 7586
rect 46114 7534 46116 7586
rect 45724 7028 45780 7038
rect 44940 6130 45220 6132
rect 44940 6078 44942 6130
rect 44994 6078 45220 6130
rect 44940 6076 45220 6078
rect 45276 6356 45332 6366
rect 44940 6066 44996 6076
rect 44492 5908 44548 5918
rect 44492 5814 44548 5852
rect 44828 5460 44884 5470
rect 44828 5122 44884 5404
rect 44828 5070 44830 5122
rect 44882 5070 44884 5122
rect 44828 5058 44884 5070
rect 44380 3390 44382 3442
rect 44434 3390 44436 3442
rect 44380 3378 44436 3390
rect 44604 3780 44660 3790
rect 45276 3780 45332 6300
rect 45612 6020 45668 6030
rect 45500 5964 45612 6020
rect 45388 5010 45444 5022
rect 45388 4958 45390 5010
rect 45442 4958 45444 5010
rect 45388 4900 45444 4958
rect 45388 4834 45444 4844
rect 45500 4564 45556 5964
rect 45612 5926 45668 5964
rect 45388 4452 45444 4462
rect 45500 4452 45556 4508
rect 45388 4450 45556 4452
rect 45388 4398 45390 4450
rect 45442 4398 45556 4450
rect 45388 4396 45556 4398
rect 45388 4386 45444 4396
rect 45276 3724 45444 3780
rect 44604 800 44660 3724
rect 45276 3556 45332 3594
rect 45276 3490 45332 3500
rect 45164 3444 45220 3482
rect 45388 3388 45444 3724
rect 45724 3666 45780 6972
rect 46060 6578 46116 7534
rect 46060 6526 46062 6578
rect 46114 6526 46116 6578
rect 46060 6514 46116 6526
rect 46284 7474 46340 7982
rect 46284 7422 46286 7474
rect 46338 7422 46340 7474
rect 46284 6356 46340 7422
rect 46844 7476 46900 7486
rect 46844 7382 46900 7420
rect 46956 7140 47012 9772
rect 47516 7362 47572 7374
rect 47516 7310 47518 7362
rect 47570 7310 47572 7362
rect 46844 7084 47012 7140
rect 47404 7140 47460 7150
rect 46284 6290 46340 6300
rect 46508 6690 46564 6702
rect 46508 6638 46510 6690
rect 46562 6638 46564 6690
rect 45724 3614 45726 3666
rect 45778 3614 45780 3666
rect 45724 3602 45780 3614
rect 45948 5572 46004 5582
rect 45164 3378 45220 3388
rect 45276 3332 45444 3388
rect 45276 800 45332 3332
rect 45948 800 46004 5516
rect 46508 5012 46564 6638
rect 46508 4946 46564 4956
rect 46620 6466 46676 6478
rect 46620 6414 46622 6466
rect 46674 6414 46676 6466
rect 46396 4564 46452 4574
rect 46396 4450 46452 4508
rect 46396 4398 46398 4450
rect 46450 4398 46452 4450
rect 46396 4386 46452 4398
rect 46620 4452 46676 6414
rect 46732 6020 46788 6030
rect 46732 5794 46788 5964
rect 46732 5742 46734 5794
rect 46786 5742 46788 5794
rect 46732 5730 46788 5742
rect 46844 5684 46900 7084
rect 47068 6690 47124 6702
rect 47068 6638 47070 6690
rect 47122 6638 47124 6690
rect 46956 5908 47012 5918
rect 46956 5814 47012 5852
rect 46844 5628 47012 5684
rect 46620 4358 46676 4396
rect 46732 5460 46788 5470
rect 46732 3388 46788 5404
rect 46956 5234 47012 5628
rect 46956 5182 46958 5234
rect 47010 5182 47012 5234
rect 46956 5170 47012 5182
rect 46844 5124 46900 5134
rect 46844 5030 46900 5068
rect 47068 3444 47124 6638
rect 47404 6132 47460 7084
rect 47516 6244 47572 7310
rect 48076 7362 48132 7374
rect 48076 7310 48078 7362
rect 48130 7310 48132 7362
rect 47516 6188 47908 6244
rect 47404 6076 47684 6132
rect 47628 5796 47684 6076
rect 47740 6020 47796 6030
rect 47740 5926 47796 5964
rect 47852 5908 47908 6188
rect 47964 5908 48020 5918
rect 47852 5906 48020 5908
rect 47852 5854 47966 5906
rect 48018 5854 48020 5906
rect 47852 5852 48020 5854
rect 47628 5740 47796 5796
rect 47292 5682 47348 5694
rect 47292 5630 47294 5682
rect 47346 5630 47348 5682
rect 47292 4340 47348 5630
rect 47516 5236 47572 5246
rect 47404 5010 47460 5022
rect 47404 4958 47406 5010
rect 47458 4958 47460 5010
rect 47404 4564 47460 4958
rect 47404 4498 47460 4508
rect 47292 4338 47460 4340
rect 47292 4286 47294 4338
rect 47346 4286 47460 4338
rect 47292 4284 47460 4286
rect 47292 4274 47348 4284
rect 47404 3666 47460 4284
rect 47404 3614 47406 3666
rect 47458 3614 47460 3666
rect 47404 3602 47460 3614
rect 47180 3444 47236 3454
rect 47068 3388 47180 3444
rect 46620 3332 46788 3388
rect 47180 3378 47236 3388
rect 47516 3332 47572 5180
rect 47628 4452 47684 4462
rect 47628 3778 47684 4396
rect 47628 3726 47630 3778
rect 47682 3726 47684 3778
rect 47628 3714 47684 3726
rect 47740 3668 47796 5740
rect 47964 5572 48020 5852
rect 47964 5506 48020 5516
rect 48076 5348 48132 7310
rect 48188 6020 48244 14254
rect 48300 7252 48356 14476
rect 48412 9716 48468 17390
rect 48412 9650 48468 9660
rect 48524 17444 48580 17454
rect 48524 8260 48580 17388
rect 48748 15988 48804 17614
rect 48748 15922 48804 15932
rect 48860 17554 48916 17566
rect 48860 17502 48862 17554
rect 48914 17502 48916 17554
rect 48748 15428 48804 15438
rect 48860 15428 48916 17502
rect 49084 16994 49140 20132
rect 49308 20020 49364 20972
rect 49420 20804 49476 20814
rect 49420 20710 49476 20748
rect 49756 20804 49812 20814
rect 49756 20710 49812 20748
rect 49868 20580 49924 20590
rect 49644 20578 49924 20580
rect 49644 20526 49870 20578
rect 49922 20526 49924 20578
rect 49644 20524 49924 20526
rect 49420 20132 49476 20142
rect 49420 20038 49476 20076
rect 49084 16942 49086 16994
rect 49138 16942 49140 16994
rect 49084 16930 49140 16942
rect 49196 19964 49364 20020
rect 49196 16884 49252 19964
rect 49644 19796 49700 20524
rect 49868 20514 49924 20524
rect 49308 19740 49700 19796
rect 49756 20356 49812 20366
rect 49308 19122 49364 19740
rect 49308 19070 49310 19122
rect 49362 19070 49364 19122
rect 49308 19058 49364 19070
rect 49308 16884 49364 16894
rect 49196 16882 49364 16884
rect 49196 16830 49310 16882
rect 49362 16830 49364 16882
rect 49196 16828 49364 16830
rect 49308 16818 49364 16828
rect 48972 16098 49028 16110
rect 48972 16046 48974 16098
rect 49026 16046 49028 16098
rect 48972 15652 49028 16046
rect 48972 15586 49028 15596
rect 49420 15986 49476 15998
rect 49420 15934 49422 15986
rect 49474 15934 49476 15986
rect 48972 15428 49028 15438
rect 48860 15372 48972 15428
rect 48748 15334 48804 15372
rect 48748 14530 48804 14542
rect 48748 14478 48750 14530
rect 48802 14478 48804 14530
rect 48748 12852 48804 14478
rect 48972 14418 49028 15372
rect 49420 15428 49476 15934
rect 49420 15362 49476 15372
rect 49756 15314 49812 20300
rect 49868 19236 49924 19246
rect 49980 19236 50036 21308
rect 50092 20804 50148 21532
rect 50204 21522 50260 21532
rect 50092 20738 50148 20748
rect 50092 20020 50148 20030
rect 50092 19926 50148 19964
rect 49868 19234 50036 19236
rect 49868 19182 49870 19234
rect 49922 19182 50036 19234
rect 49868 19180 50036 19182
rect 50204 19908 50260 19918
rect 49868 19170 49924 19180
rect 49756 15262 49758 15314
rect 49810 15262 49812 15314
rect 49756 15250 49812 15262
rect 49868 18674 49924 18686
rect 49868 18622 49870 18674
rect 49922 18622 49924 18674
rect 48972 14366 48974 14418
rect 49026 14366 49028 14418
rect 48972 14354 49028 14366
rect 49084 15092 49140 15102
rect 48860 14084 48916 14094
rect 48860 13970 48916 14028
rect 48860 13918 48862 13970
rect 48914 13918 48916 13970
rect 48860 13906 48916 13918
rect 48748 12786 48804 12796
rect 48524 8194 48580 8204
rect 48412 7252 48468 7262
rect 48300 7196 48412 7252
rect 48412 7186 48468 7196
rect 49084 6692 49140 15036
rect 49868 7700 49924 18622
rect 49980 17780 50036 17790
rect 49980 17332 50036 17724
rect 50204 17778 50260 19852
rect 50204 17726 50206 17778
rect 50258 17726 50260 17778
rect 50204 17714 50260 17726
rect 50316 17668 50372 26012
rect 50556 25116 50820 25126
rect 50612 25060 50660 25116
rect 50716 25060 50764 25116
rect 50556 25050 50820 25060
rect 50556 23548 50820 23558
rect 50612 23492 50660 23548
rect 50716 23492 50764 23548
rect 50556 23482 50820 23492
rect 50428 22708 50484 22718
rect 50428 22482 50484 22652
rect 50428 22430 50430 22482
rect 50482 22430 50484 22482
rect 50428 22418 50484 22430
rect 50540 22594 50596 22606
rect 50540 22542 50542 22594
rect 50594 22542 50596 22594
rect 50540 22260 50596 22542
rect 50428 22204 50596 22260
rect 50428 20802 50484 22204
rect 50876 22148 50932 22158
rect 50876 22054 50932 22092
rect 50556 21980 50820 21990
rect 50612 21924 50660 21980
rect 50716 21924 50764 21980
rect 50556 21914 50820 21924
rect 50428 20750 50430 20802
rect 50482 20750 50484 20802
rect 50428 20738 50484 20750
rect 50652 21756 50932 21812
rect 50652 21700 50708 21756
rect 50652 20690 50708 21644
rect 50876 21698 50932 21756
rect 50876 21646 50878 21698
rect 50930 21646 50932 21698
rect 50876 21634 50932 21646
rect 50652 20638 50654 20690
rect 50706 20638 50708 20690
rect 50652 20626 50708 20638
rect 50876 21474 50932 21486
rect 50876 21422 50878 21474
rect 50930 21422 50932 21474
rect 50556 20412 50820 20422
rect 50612 20356 50660 20412
rect 50716 20356 50764 20412
rect 50556 20346 50820 20356
rect 50876 20132 50932 21422
rect 50988 20580 51044 26684
rect 51212 26674 51268 26684
rect 51100 24948 51156 24958
rect 51100 23378 51156 24892
rect 51324 23548 51380 27468
rect 51100 23326 51102 23378
rect 51154 23326 51156 23378
rect 51100 22594 51156 23326
rect 51100 22542 51102 22594
rect 51154 22542 51156 22594
rect 51100 22530 51156 22542
rect 51212 23492 51380 23548
rect 51212 20804 51268 23492
rect 51324 22594 51380 22606
rect 51324 22542 51326 22594
rect 51378 22542 51380 22594
rect 51324 21586 51380 22542
rect 51324 21534 51326 21586
rect 51378 21534 51380 21586
rect 51324 21522 51380 21534
rect 51436 22146 51492 22158
rect 51436 22094 51438 22146
rect 51490 22094 51492 22146
rect 51212 20738 51268 20748
rect 51324 20916 51380 20926
rect 50988 20524 51268 20580
rect 50876 20066 50932 20076
rect 51100 20018 51156 20030
rect 51100 19966 51102 20018
rect 51154 19966 51156 20018
rect 50876 19908 50932 19918
rect 50556 18844 50820 18854
rect 50612 18788 50660 18844
rect 50716 18788 50764 18844
rect 50556 18778 50820 18788
rect 50764 17778 50820 17790
rect 50764 17726 50766 17778
rect 50818 17726 50820 17778
rect 50316 17612 50596 17668
rect 50540 17556 50596 17612
rect 50540 17490 50596 17500
rect 50764 17444 50820 17726
rect 50876 17554 50932 19852
rect 50988 19234 51044 19246
rect 50988 19182 50990 19234
rect 51042 19182 51044 19234
rect 50988 18004 51044 19182
rect 50988 17938 51044 17948
rect 51100 19122 51156 19966
rect 51100 19070 51102 19122
rect 51154 19070 51156 19122
rect 51100 18562 51156 19070
rect 51100 18510 51102 18562
rect 51154 18510 51156 18562
rect 50876 17502 50878 17554
rect 50930 17502 50932 17554
rect 50876 17490 50932 17502
rect 50988 17666 51044 17678
rect 50988 17614 50990 17666
rect 51042 17614 51044 17666
rect 50988 17556 51044 17614
rect 50764 17378 50820 17388
rect 49980 17266 50036 17276
rect 50556 17276 50820 17286
rect 50612 17220 50660 17276
rect 50716 17220 50764 17276
rect 50556 17210 50820 17220
rect 50428 17108 50484 17118
rect 50316 17106 50484 17108
rect 50316 17054 50430 17106
rect 50482 17054 50484 17106
rect 50316 17052 50484 17054
rect 50316 14420 50372 17052
rect 50428 17042 50484 17052
rect 50988 16996 51044 17500
rect 50988 16930 51044 16940
rect 51100 16994 51156 18510
rect 51212 18564 51268 20524
rect 51324 19908 51380 20860
rect 51324 19842 51380 19852
rect 51436 20018 51492 22094
rect 51436 19966 51438 20018
rect 51490 19966 51492 20018
rect 51436 19684 51492 19966
rect 51436 19618 51492 19628
rect 51548 19460 51604 30044
rect 51660 21924 51716 31502
rect 51772 30212 51828 30222
rect 51772 30118 51828 30156
rect 51772 23492 51828 23502
rect 51772 22594 51828 23436
rect 51772 22542 51774 22594
rect 51826 22542 51828 22594
rect 51772 22482 51828 22542
rect 51772 22430 51774 22482
rect 51826 22430 51828 22482
rect 51772 22418 51828 22430
rect 51660 21858 51716 21868
rect 51772 21698 51828 21710
rect 51772 21646 51774 21698
rect 51826 21646 51828 21698
rect 51660 21588 51716 21598
rect 51660 20802 51716 21532
rect 51772 20916 51828 21646
rect 51772 20850 51828 20860
rect 51660 20750 51662 20802
rect 51714 20750 51716 20802
rect 51660 20738 51716 20750
rect 51212 18498 51268 18508
rect 51436 19404 51604 19460
rect 51660 20580 51716 20590
rect 51324 18450 51380 18462
rect 51324 18398 51326 18450
rect 51378 18398 51380 18450
rect 51324 17780 51380 18398
rect 51436 18116 51492 19404
rect 51660 19348 51716 20524
rect 51436 18050 51492 18060
rect 51548 19292 51716 19348
rect 51772 19908 51828 19918
rect 51772 19346 51828 19852
rect 51772 19294 51774 19346
rect 51826 19294 51828 19346
rect 51324 17714 51380 17724
rect 51548 17556 51604 19292
rect 51772 19282 51828 19294
rect 51660 19124 51716 19134
rect 51660 17666 51716 19068
rect 51660 17614 51662 17666
rect 51714 17614 51716 17666
rect 51660 17602 51716 17614
rect 51100 16942 51102 16994
rect 51154 16942 51156 16994
rect 51100 16210 51156 16942
rect 51100 16158 51102 16210
rect 51154 16158 51156 16210
rect 51100 16146 51156 16158
rect 51212 17500 51604 17556
rect 50428 15876 50484 15886
rect 50428 15782 50484 15820
rect 50556 15708 50820 15718
rect 50612 15652 50660 15708
rect 50716 15652 50764 15708
rect 50556 15642 50820 15652
rect 50652 15428 50708 15438
rect 50652 15334 50708 15372
rect 51212 15428 51268 17500
rect 51436 16882 51492 16894
rect 51436 16830 51438 16882
rect 51490 16830 51492 16882
rect 51436 16436 51492 16830
rect 50876 15314 50932 15326
rect 50876 15262 50878 15314
rect 50930 15262 50932 15314
rect 50428 14420 50484 14430
rect 50316 14364 50428 14420
rect 50428 14354 50484 14364
rect 50876 14308 50932 15262
rect 51100 14644 51156 14654
rect 51212 14644 51268 15372
rect 51100 14642 51268 14644
rect 51100 14590 51102 14642
rect 51154 14590 51268 14642
rect 51100 14588 51268 14590
rect 51324 15876 51380 15886
rect 51436 15876 51492 16380
rect 51660 15876 51716 15886
rect 51436 15874 51716 15876
rect 51436 15822 51662 15874
rect 51714 15822 51716 15874
rect 51436 15820 51716 15822
rect 51100 14578 51156 14588
rect 51324 14532 51380 15820
rect 51660 15810 51716 15820
rect 51660 15204 51716 15242
rect 51660 15138 51716 15148
rect 51324 14438 51380 14476
rect 50876 14242 50932 14252
rect 50556 14140 50820 14150
rect 50612 14084 50660 14140
rect 50716 14084 50764 14140
rect 50556 14074 50820 14084
rect 50556 12572 50820 12582
rect 50612 12516 50660 12572
rect 50716 12516 50764 12572
rect 50556 12506 50820 12516
rect 50556 11004 50820 11014
rect 50612 10948 50660 11004
rect 50716 10948 50764 11004
rect 50556 10938 50820 10948
rect 50556 9436 50820 9446
rect 50612 9380 50660 9436
rect 50716 9380 50764 9436
rect 50556 9370 50820 9380
rect 49868 7634 49924 7644
rect 50204 9044 50260 9054
rect 49084 6626 49140 6636
rect 49532 7476 49588 7486
rect 48636 6580 48692 6590
rect 48636 6486 48692 6524
rect 49084 6466 49140 6478
rect 49084 6414 49086 6466
rect 49138 6414 49140 6466
rect 48188 5954 48244 5964
rect 48748 6132 48804 6142
rect 48748 5906 48804 6076
rect 48748 5854 48750 5906
rect 48802 5854 48804 5906
rect 48748 5842 48804 5854
rect 48972 5908 49028 5918
rect 48748 5684 48804 5694
rect 47964 5292 48132 5348
rect 48300 5348 48356 5358
rect 47964 3892 48020 5292
rect 47964 3826 48020 3836
rect 48076 5124 48132 5134
rect 47964 3668 48020 3678
rect 47740 3666 48020 3668
rect 47740 3614 47966 3666
rect 48018 3614 48020 3666
rect 47740 3612 48020 3614
rect 47964 3602 48020 3612
rect 46620 800 46676 3332
rect 47292 3276 47572 3332
rect 47292 800 47348 3276
rect 48076 3108 48132 5068
rect 48300 3442 48356 5292
rect 48748 4562 48804 5628
rect 48972 5010 49028 5852
rect 48972 4958 48974 5010
rect 49026 4958 49028 5010
rect 48972 4946 49028 4958
rect 48748 4510 48750 4562
rect 48802 4510 48804 4562
rect 48748 4498 48804 4510
rect 48972 4340 49028 4350
rect 48524 3892 48580 3902
rect 48524 3554 48580 3836
rect 48524 3502 48526 3554
rect 48578 3502 48580 3554
rect 48524 3490 48580 3502
rect 48300 3390 48302 3442
rect 48354 3390 48356 3442
rect 48300 3378 48356 3390
rect 48972 3442 49028 4284
rect 49084 4338 49140 6414
rect 49196 5906 49252 5918
rect 49196 5854 49198 5906
rect 49250 5854 49252 5906
rect 49196 5796 49252 5854
rect 49196 5124 49252 5740
rect 49196 5058 49252 5068
rect 49308 5460 49364 5470
rect 49308 5122 49364 5404
rect 49308 5070 49310 5122
rect 49362 5070 49364 5122
rect 49308 5058 49364 5070
rect 49532 5124 49588 7420
rect 50204 6692 50260 8988
rect 50556 7868 50820 7878
rect 50612 7812 50660 7868
rect 50716 7812 50764 7868
rect 50556 7802 50820 7812
rect 51100 6692 51156 6702
rect 50204 6690 50372 6692
rect 50204 6638 50206 6690
rect 50258 6638 50372 6690
rect 50204 6636 50372 6638
rect 50204 6626 50260 6636
rect 49084 4286 49086 4338
rect 49138 4286 49140 4338
rect 49084 4116 49140 4286
rect 49532 4338 49588 5068
rect 49644 6580 49700 6590
rect 49644 5010 49700 6524
rect 49756 5796 49812 5806
rect 49756 5702 49812 5740
rect 50204 5794 50260 5806
rect 50204 5742 50206 5794
rect 50258 5742 50260 5794
rect 49868 5236 49924 5246
rect 49868 5122 49924 5180
rect 49868 5070 49870 5122
rect 49922 5070 49924 5122
rect 49868 5058 49924 5070
rect 49644 4958 49646 5010
rect 49698 4958 49700 5010
rect 49644 4946 49700 4958
rect 49532 4286 49534 4338
rect 49586 4286 49588 4338
rect 49532 4274 49588 4286
rect 49084 4050 49140 4060
rect 49308 4116 49364 4126
rect 48972 3390 48974 3442
rect 49026 3390 49028 3442
rect 48972 3378 49028 3390
rect 49196 3554 49252 3566
rect 49196 3502 49198 3554
rect 49250 3502 49252 3554
rect 47964 3052 48132 3108
rect 49196 3332 49252 3502
rect 47964 800 48020 3052
rect 49196 2548 49252 3276
rect 49196 2482 49252 2492
rect 49308 800 49364 4060
rect 49868 3892 49924 3902
rect 49868 3668 49924 3836
rect 49868 3554 49924 3612
rect 49868 3502 49870 3554
rect 49922 3502 49924 3554
rect 49868 3490 49924 3502
rect 50092 3556 50148 3566
rect 49644 3444 49700 3482
rect 49644 3378 49700 3388
rect 50092 2996 50148 3500
rect 50204 3332 50260 5742
rect 50316 5346 50372 6636
rect 51100 6690 51268 6692
rect 51100 6638 51102 6690
rect 51154 6638 51268 6690
rect 51100 6636 51268 6638
rect 51100 6626 51156 6636
rect 50764 6578 50820 6590
rect 50764 6526 50766 6578
rect 50818 6526 50820 6578
rect 50764 6468 50820 6526
rect 51212 6580 51268 6636
rect 51212 6514 51268 6524
rect 51548 6690 51604 6702
rect 51548 6638 51550 6690
rect 51602 6638 51604 6690
rect 50764 6402 50820 6412
rect 51212 6356 51268 6366
rect 50556 6300 50820 6310
rect 50612 6244 50660 6300
rect 50716 6244 50764 6300
rect 50556 6234 50820 6244
rect 50988 5794 51044 5806
rect 50988 5742 50990 5794
rect 51042 5742 51044 5794
rect 50316 5294 50318 5346
rect 50370 5294 50372 5346
rect 50316 5282 50372 5294
rect 50876 5572 50932 5582
rect 50876 5234 50932 5516
rect 50988 5346 51044 5742
rect 50988 5294 50990 5346
rect 51042 5294 51044 5346
rect 50988 5282 51044 5294
rect 50876 5182 50878 5234
rect 50930 5182 50932 5234
rect 50876 5170 50932 5182
rect 50428 5124 50484 5134
rect 50428 5030 50484 5068
rect 50316 5012 50372 5022
rect 50316 3442 50372 4956
rect 50556 4732 50820 4742
rect 50612 4676 50660 4732
rect 50716 4676 50764 4732
rect 50556 4666 50820 4676
rect 50540 4116 50596 4126
rect 50540 4022 50596 4060
rect 50540 3780 50596 3790
rect 50540 3554 50596 3724
rect 50540 3502 50542 3554
rect 50594 3502 50596 3554
rect 50540 3490 50596 3502
rect 50316 3390 50318 3442
rect 50370 3390 50372 3442
rect 50316 3378 50372 3390
rect 50876 3444 50932 3454
rect 50204 3266 50260 3276
rect 50556 3164 50820 3174
rect 50612 3108 50660 3164
rect 50716 3108 50764 3164
rect 50556 3098 50820 3108
rect 50876 2996 50932 3388
rect 51212 3442 51268 6300
rect 51548 6132 51604 6638
rect 51884 6468 51940 39004
rect 51996 38836 52052 40236
rect 51996 13972 52052 38780
rect 52444 38668 52500 55412
rect 52444 38612 52612 38668
rect 52332 33460 52388 33470
rect 52220 33404 52332 33460
rect 52220 22596 52276 33404
rect 52332 33394 52388 33404
rect 52332 32340 52388 32350
rect 52332 31218 52388 32284
rect 52332 31166 52334 31218
rect 52386 31166 52388 31218
rect 52332 31108 52388 31166
rect 52332 31042 52388 31052
rect 52220 22540 52500 22596
rect 52220 22372 52276 22382
rect 52220 21586 52276 22316
rect 52220 21534 52222 21586
rect 52274 21534 52276 21586
rect 52220 21522 52276 21534
rect 52332 21474 52388 21486
rect 52332 21422 52334 21474
rect 52386 21422 52388 21474
rect 52108 21364 52164 21374
rect 52108 20130 52164 21308
rect 52108 20078 52110 20130
rect 52162 20078 52164 20130
rect 52108 20066 52164 20078
rect 52108 17780 52164 17790
rect 52108 17686 52164 17724
rect 52108 16996 52164 17006
rect 52108 16210 52164 16940
rect 52332 16994 52388 21422
rect 52444 18788 52500 22540
rect 52556 20020 52612 38612
rect 52780 36708 52836 36718
rect 52780 31892 52836 36652
rect 52780 31798 52836 31836
rect 52892 34356 52948 34366
rect 52780 31220 52836 31230
rect 52892 31220 52948 34300
rect 53116 33460 53172 33498
rect 53116 33394 53172 33404
rect 53004 33348 53060 33358
rect 53004 33254 53060 33292
rect 52836 31164 52948 31220
rect 52780 31126 52836 31164
rect 52780 22596 52836 22606
rect 52780 22372 52836 22540
rect 52556 19954 52612 19964
rect 52668 22370 52836 22372
rect 52668 22318 52782 22370
rect 52834 22318 52836 22370
rect 52668 22316 52836 22318
rect 52668 19234 52724 22316
rect 52780 22306 52836 22316
rect 53228 22484 53284 75630
rect 53452 67228 53508 76302
rect 53564 75684 53620 79200
rect 53900 76692 53956 76702
rect 53900 76598 53956 76636
rect 54236 76132 54292 79200
rect 54908 76580 54964 79200
rect 55580 77812 55636 79200
rect 55580 77756 55860 77812
rect 55132 76692 55188 76702
rect 55132 76598 55188 76636
rect 54908 76514 54964 76524
rect 55580 76580 55636 76590
rect 55636 76524 55748 76580
rect 55580 76514 55636 76524
rect 54460 76356 54516 76366
rect 54460 76354 54852 76356
rect 54460 76302 54462 76354
rect 54514 76302 54852 76354
rect 54460 76300 54852 76302
rect 54460 76290 54516 76300
rect 54236 76076 54740 76132
rect 53788 75684 53844 75694
rect 53564 75682 53844 75684
rect 53564 75630 53790 75682
rect 53842 75630 53844 75682
rect 53564 75628 53844 75630
rect 53564 75122 53620 75628
rect 53788 75618 53844 75628
rect 54348 75682 54404 75694
rect 54348 75630 54350 75682
rect 54402 75630 54404 75682
rect 53564 75070 53566 75122
rect 53618 75070 53620 75122
rect 53564 75058 53620 75070
rect 54348 71764 54404 75630
rect 54460 75122 54516 76076
rect 54684 75682 54740 76076
rect 54684 75630 54686 75682
rect 54738 75630 54740 75682
rect 54684 75618 54740 75630
rect 54460 75070 54462 75122
rect 54514 75070 54516 75122
rect 54460 75058 54516 75070
rect 54348 71708 54628 71764
rect 54460 71540 54516 71550
rect 53452 67172 53732 67228
rect 53340 33460 53396 33470
rect 53340 33234 53396 33404
rect 53340 33182 53342 33234
rect 53394 33182 53396 33234
rect 53340 33170 53396 33182
rect 52668 19182 52670 19234
rect 52722 19182 52724 19234
rect 52668 19170 52724 19182
rect 52780 21586 52836 21598
rect 52780 21534 52782 21586
rect 52834 21534 52836 21586
rect 52780 20802 52836 21534
rect 53116 21588 53172 21598
rect 53116 21494 53172 21532
rect 52780 20750 52782 20802
rect 52834 20750 52836 20802
rect 52780 20018 52836 20750
rect 53228 20802 53284 22428
rect 53676 22484 53732 67172
rect 54460 55468 54516 71484
rect 54348 55412 54516 55468
rect 54236 40180 54292 40190
rect 54124 36148 54180 36158
rect 54012 35700 54068 35710
rect 54012 35606 54068 35644
rect 53788 35028 53844 35038
rect 53788 34802 53844 34972
rect 53900 34916 53956 34926
rect 53900 34822 53956 34860
rect 53788 34750 53790 34802
rect 53842 34750 53844 34802
rect 53788 34738 53844 34750
rect 54012 34690 54068 34702
rect 54012 34638 54014 34690
rect 54066 34638 54068 34690
rect 54012 26908 54068 34638
rect 54124 33460 54180 36092
rect 54236 35812 54292 40124
rect 54236 35718 54292 35756
rect 54124 33366 54180 33404
rect 53900 26852 54068 26908
rect 53788 22484 53844 22494
rect 53676 22482 53844 22484
rect 53676 22430 53790 22482
rect 53842 22430 53844 22482
rect 53676 22428 53844 22430
rect 53340 22370 53396 22382
rect 53340 22318 53342 22370
rect 53394 22318 53396 22370
rect 53340 20916 53396 22318
rect 53676 22372 53732 22428
rect 53788 22418 53844 22428
rect 53676 22306 53732 22316
rect 53788 21924 53844 21934
rect 53676 21476 53732 21486
rect 53676 21382 53732 21420
rect 53340 20850 53396 20860
rect 53228 20750 53230 20802
rect 53282 20750 53284 20802
rect 53228 20738 53284 20750
rect 53452 20804 53508 20814
rect 53452 20690 53508 20748
rect 53452 20638 53454 20690
rect 53506 20638 53508 20690
rect 52892 20580 52948 20590
rect 52892 20578 53172 20580
rect 52892 20526 52894 20578
rect 52946 20526 53172 20578
rect 52892 20524 53172 20526
rect 52892 20514 52948 20524
rect 52780 19966 52782 20018
rect 52834 19966 52836 20018
rect 52780 19124 52836 19966
rect 52780 19058 52836 19068
rect 52892 20242 52948 20254
rect 52892 20190 52894 20242
rect 52946 20190 52948 20242
rect 52780 18788 52836 18798
rect 52444 18732 52780 18788
rect 52780 18722 52836 18732
rect 52556 18564 52612 18574
rect 52444 18338 52500 18350
rect 52444 18286 52446 18338
rect 52498 18286 52500 18338
rect 52444 18004 52500 18286
rect 52444 17938 52500 17948
rect 52332 16942 52334 16994
rect 52386 16942 52388 16994
rect 52332 16930 52388 16942
rect 52556 16882 52612 18508
rect 52892 17556 52948 20190
rect 52780 17500 52948 17556
rect 53004 18340 53060 18350
rect 52556 16830 52558 16882
rect 52610 16830 52612 16882
rect 52556 16818 52612 16830
rect 52668 17444 52724 17454
rect 52108 16158 52110 16210
rect 52162 16158 52164 16210
rect 52108 16146 52164 16158
rect 52668 16098 52724 17388
rect 52668 16046 52670 16098
rect 52722 16046 52724 16098
rect 52668 16034 52724 16046
rect 52556 15428 52612 15438
rect 52556 15314 52612 15372
rect 52780 15426 52836 17500
rect 52780 15374 52782 15426
rect 52834 15374 52836 15426
rect 52780 15362 52836 15374
rect 52556 15262 52558 15314
rect 52610 15262 52612 15314
rect 52556 15250 52612 15262
rect 52108 14756 52164 14766
rect 52108 14662 52164 14700
rect 52892 14756 52948 14766
rect 52668 14532 52724 14542
rect 52668 14438 52724 14476
rect 52668 13972 52724 13982
rect 51996 13916 52164 13972
rect 52108 13524 52164 13916
rect 52444 13970 52724 13972
rect 52444 13918 52670 13970
rect 52722 13918 52724 13970
rect 52444 13916 52724 13918
rect 52220 13748 52276 13758
rect 52220 13654 52276 13692
rect 51996 13468 52164 13524
rect 51996 6580 52052 13468
rect 51996 6514 52052 6524
rect 51884 6402 51940 6412
rect 52108 6466 52164 6478
rect 52108 6414 52110 6466
rect 52162 6414 52164 6466
rect 51548 6066 51604 6076
rect 52108 6132 52164 6414
rect 52108 6066 52164 6076
rect 51436 5794 51492 5806
rect 51436 5742 51438 5794
rect 51490 5742 51492 5794
rect 51324 5236 51380 5246
rect 51324 5142 51380 5180
rect 51436 3780 51492 5742
rect 52444 5796 52500 13916
rect 52668 13906 52724 13916
rect 52892 13746 52948 14700
rect 52892 13694 52894 13746
rect 52946 13694 52948 13746
rect 52892 13682 52948 13694
rect 52444 5730 52500 5740
rect 52556 11620 52612 11630
rect 52556 5796 52612 11564
rect 53004 11172 53060 18284
rect 53116 17444 53172 20524
rect 53452 20130 53508 20638
rect 53452 20078 53454 20130
rect 53506 20078 53508 20130
rect 53452 20066 53508 20078
rect 53564 20244 53620 20254
rect 53340 20020 53396 20030
rect 53340 19926 53396 19964
rect 53228 19234 53284 19246
rect 53228 19182 53230 19234
rect 53282 19182 53284 19234
rect 53228 19124 53284 19182
rect 53228 19058 53284 19068
rect 53228 18788 53284 18798
rect 53228 17666 53284 18732
rect 53452 18564 53508 18574
rect 53228 17614 53230 17666
rect 53282 17614 53284 17666
rect 53228 17602 53284 17614
rect 53340 18562 53508 18564
rect 53340 18510 53454 18562
rect 53506 18510 53508 18562
rect 53340 18508 53508 18510
rect 53116 17388 53284 17444
rect 53116 17220 53172 17230
rect 53116 14642 53172 17164
rect 53116 14590 53118 14642
rect 53170 14590 53172 14642
rect 53116 14578 53172 14590
rect 53228 13860 53284 17388
rect 53340 17332 53396 18508
rect 53452 18498 53508 18508
rect 53452 17556 53508 17566
rect 53564 17556 53620 20188
rect 53788 19012 53844 21868
rect 53900 19234 53956 26852
rect 54236 22484 54292 22494
rect 54236 22390 54292 22428
rect 54348 21700 54404 55412
rect 54572 21812 54628 71708
rect 54684 35586 54740 35598
rect 54684 35534 54686 35586
rect 54738 35534 54740 35586
rect 54684 31556 54740 35534
rect 54796 31668 54852 76300
rect 55244 75682 55300 75694
rect 55692 75684 55748 76524
rect 55804 76356 55860 77756
rect 56252 77364 56308 79200
rect 56252 77308 56756 77364
rect 55916 76356 55972 76366
rect 55804 76354 55972 76356
rect 55804 76302 55918 76354
rect 55970 76302 55972 76354
rect 55804 76300 55972 76302
rect 55916 76290 55972 76300
rect 56700 75906 56756 77308
rect 56924 76692 56980 79200
rect 57596 77028 57652 79200
rect 57596 76972 57764 77028
rect 56924 76626 56980 76636
rect 56700 75854 56702 75906
rect 56754 75854 56756 75906
rect 56700 75842 56756 75854
rect 57596 76468 57652 76478
rect 55244 75630 55246 75682
rect 55298 75630 55300 75682
rect 55244 71540 55300 75630
rect 55356 75682 55748 75684
rect 55356 75630 55694 75682
rect 55746 75630 55748 75682
rect 55356 75628 55748 75630
rect 55356 75122 55412 75628
rect 55692 75618 55748 75628
rect 55916 75684 55972 75694
rect 55356 75070 55358 75122
rect 55410 75070 55412 75122
rect 55356 75058 55412 75070
rect 55244 71474 55300 71484
rect 55804 45332 55860 45342
rect 55804 42866 55860 45276
rect 55804 42814 55806 42866
rect 55858 42814 55860 42866
rect 55804 42802 55860 42814
rect 55244 42532 55300 42542
rect 55020 42530 55300 42532
rect 55020 42478 55246 42530
rect 55298 42478 55300 42530
rect 55020 42476 55300 42478
rect 55020 42194 55076 42476
rect 55244 42466 55300 42476
rect 55020 42142 55022 42194
rect 55074 42142 55076 42194
rect 55020 42130 55076 42142
rect 55580 41860 55636 41870
rect 55580 41766 55636 41804
rect 55356 41748 55412 41758
rect 55468 41748 55524 41758
rect 55356 41746 55468 41748
rect 55356 41694 55358 41746
rect 55410 41694 55468 41746
rect 55356 41692 55468 41694
rect 55356 41682 55412 41692
rect 55468 41410 55524 41692
rect 55468 41358 55470 41410
rect 55522 41358 55524 41410
rect 55468 41346 55524 41358
rect 55804 41746 55860 41758
rect 55804 41694 55806 41746
rect 55858 41694 55860 41746
rect 55804 41410 55860 41694
rect 55804 41358 55806 41410
rect 55858 41358 55860 41410
rect 55804 41346 55860 41358
rect 55244 41186 55300 41198
rect 55244 41134 55246 41186
rect 55298 41134 55300 41186
rect 54908 40964 54964 40974
rect 55244 40964 55300 41134
rect 54908 40962 55300 40964
rect 54908 40910 54910 40962
rect 54962 40910 55300 40962
rect 54908 40908 55300 40910
rect 54908 40068 54964 40908
rect 55244 40628 55300 40908
rect 55244 40562 55300 40572
rect 54908 40002 54964 40012
rect 55356 35924 55412 35934
rect 54908 35812 54964 35822
rect 54908 35028 54964 35756
rect 55356 35810 55412 35868
rect 55356 35758 55358 35810
rect 55410 35758 55412 35810
rect 55356 35746 55412 35758
rect 55020 35698 55076 35710
rect 55020 35646 55022 35698
rect 55074 35646 55076 35698
rect 55020 35252 55076 35646
rect 55692 35588 55748 35598
rect 55692 35494 55748 35532
rect 55020 35186 55076 35196
rect 55020 35028 55076 35038
rect 54908 35026 55076 35028
rect 54908 34974 55022 35026
rect 55074 34974 55076 35026
rect 54908 34972 55076 34974
rect 55020 34962 55076 34972
rect 55356 35028 55412 35038
rect 55356 34934 55412 34972
rect 54796 31612 55076 31668
rect 54684 31490 54740 31500
rect 55020 23548 55076 31612
rect 54348 21586 54404 21644
rect 54348 21534 54350 21586
rect 54402 21534 54404 21586
rect 54348 21522 54404 21534
rect 54460 21698 54516 21710
rect 54460 21646 54462 21698
rect 54514 21646 54516 21698
rect 54460 21476 54516 21646
rect 54124 20916 54180 20926
rect 54124 20804 54180 20860
rect 54124 20802 54404 20804
rect 54124 20750 54126 20802
rect 54178 20750 54404 20802
rect 54124 20748 54404 20750
rect 54124 20738 54180 20748
rect 54236 20580 54292 20590
rect 53900 19182 53902 19234
rect 53954 19182 53956 19234
rect 53900 19170 53956 19182
rect 54124 20578 54292 20580
rect 54124 20526 54238 20578
rect 54290 20526 54292 20578
rect 54124 20524 54292 20526
rect 54124 19122 54180 20524
rect 54236 20514 54292 20524
rect 54348 20468 54404 20748
rect 54460 20692 54516 21420
rect 54572 20804 54628 21756
rect 54796 23492 55076 23548
rect 55132 31556 55188 31566
rect 54684 20804 54740 20814
rect 54572 20802 54740 20804
rect 54572 20750 54686 20802
rect 54738 20750 54740 20802
rect 54572 20748 54740 20750
rect 54684 20738 54740 20748
rect 54460 20626 54516 20636
rect 54348 20412 54516 20468
rect 54348 20244 54404 20254
rect 54348 20150 54404 20188
rect 54460 20018 54516 20412
rect 54460 19966 54462 20018
rect 54514 19966 54516 20018
rect 54460 19954 54516 19966
rect 54796 20132 54852 23492
rect 55020 21810 55076 21822
rect 55020 21758 55022 21810
rect 55074 21758 55076 21810
rect 54908 21586 54964 21598
rect 54908 21534 54910 21586
rect 54962 21534 54964 21586
rect 54908 20916 54964 21534
rect 54908 20850 54964 20860
rect 54796 20018 54852 20076
rect 54796 19966 54798 20018
rect 54850 19966 54852 20018
rect 54796 19954 54852 19966
rect 55020 19572 55076 21758
rect 55020 19506 55076 19516
rect 54124 19070 54126 19122
rect 54178 19070 54180 19122
rect 54124 19058 54180 19070
rect 54796 19124 54852 19134
rect 53788 18956 53956 19012
rect 53676 18450 53732 18462
rect 53676 18398 53678 18450
rect 53730 18398 53732 18450
rect 53676 18340 53732 18398
rect 53676 18274 53732 18284
rect 53452 17554 53620 17556
rect 53452 17502 53454 17554
rect 53506 17502 53620 17554
rect 53452 17500 53620 17502
rect 53676 18116 53732 18126
rect 53452 17490 53508 17500
rect 53340 17266 53396 17276
rect 53452 17108 53508 17118
rect 53228 13794 53284 13804
rect 53340 17106 53508 17108
rect 53340 17054 53454 17106
rect 53506 17054 53508 17106
rect 53340 17052 53508 17054
rect 52892 11116 53060 11172
rect 52892 9268 52948 11116
rect 52892 9202 52948 9212
rect 53004 10948 53060 10958
rect 53004 6356 53060 10892
rect 53340 10164 53396 17052
rect 53452 17042 53508 17052
rect 53676 16098 53732 18060
rect 53676 16046 53678 16098
rect 53730 16046 53732 16098
rect 53676 16034 53732 16046
rect 53788 15874 53844 15886
rect 53788 15822 53790 15874
rect 53842 15822 53844 15874
rect 53340 10098 53396 10108
rect 53452 15538 53508 15550
rect 53452 15486 53454 15538
rect 53506 15486 53508 15538
rect 53452 8428 53508 15486
rect 53452 8372 53732 8428
rect 53004 6290 53060 6300
rect 53452 8036 53508 8046
rect 53004 6132 53060 6142
rect 52556 5794 52724 5796
rect 52556 5742 52558 5794
rect 52610 5742 52724 5794
rect 52556 5740 52724 5742
rect 52556 5730 52612 5740
rect 51996 5348 52052 5358
rect 51996 5346 52164 5348
rect 51996 5294 51998 5346
rect 52050 5294 52164 5346
rect 51996 5292 52164 5294
rect 51996 5282 52052 5292
rect 51772 5122 51828 5134
rect 51772 5070 51774 5122
rect 51826 5070 51828 5122
rect 51436 3714 51492 3724
rect 51660 4900 51716 4910
rect 51212 3390 51214 3442
rect 51266 3390 51268 3442
rect 51212 3332 51268 3390
rect 51212 3266 51268 3276
rect 51324 3668 51380 3678
rect 49980 2940 50148 2996
rect 50652 2940 50932 2996
rect 49980 800 50036 2940
rect 50652 800 50708 2940
rect 51324 800 51380 3612
rect 51660 3556 51716 4844
rect 51772 3892 51828 5070
rect 51772 3826 51828 3836
rect 51660 3462 51716 3500
rect 51996 3556 52052 3566
rect 51996 800 52052 3500
rect 52108 3442 52164 5292
rect 52668 4340 52724 5740
rect 52780 5122 52836 5134
rect 52780 5070 52782 5122
rect 52834 5070 52836 5122
rect 52780 4900 52836 5070
rect 52780 4834 52836 4844
rect 52892 4340 52948 4350
rect 52668 4338 52948 4340
rect 52668 4286 52894 4338
rect 52946 4286 52948 4338
rect 52668 4284 52948 4286
rect 52892 4274 52948 4284
rect 52556 4226 52612 4238
rect 52556 4174 52558 4226
rect 52610 4174 52612 4226
rect 52108 3390 52110 3442
rect 52162 3390 52164 3442
rect 52108 3378 52164 3390
rect 52332 3556 52388 3566
rect 52556 3556 52612 4174
rect 52332 3554 52612 3556
rect 52332 3502 52334 3554
rect 52386 3502 52612 3554
rect 52332 3500 52612 3502
rect 52668 4116 52724 4126
rect 53004 4116 53060 6076
rect 53340 4900 53396 4910
rect 52332 3444 52388 3500
rect 52332 3378 52388 3388
rect 52668 800 52724 4060
rect 52780 4060 53060 4116
rect 53228 4898 53396 4900
rect 53228 4846 53342 4898
rect 53394 4846 53396 4898
rect 53228 4844 53396 4846
rect 52780 3442 52836 4060
rect 53004 3668 53060 3678
rect 53004 3554 53060 3612
rect 53004 3502 53006 3554
rect 53058 3502 53060 3554
rect 53004 3490 53060 3502
rect 53228 3556 53284 4844
rect 53340 4834 53396 4844
rect 53228 3490 53284 3500
rect 53340 3668 53396 3678
rect 52780 3390 52782 3442
rect 52834 3390 52836 3442
rect 52780 3378 52836 3390
rect 53340 800 53396 3612
rect 53452 3442 53508 7980
rect 53676 4676 53732 8372
rect 53676 4610 53732 4620
rect 53788 4228 53844 15822
rect 53900 13972 53956 18956
rect 53900 13746 53956 13916
rect 53900 13694 53902 13746
rect 53954 13694 53956 13746
rect 53900 13682 53956 13694
rect 54012 18674 54068 18686
rect 54012 18622 54014 18674
rect 54066 18622 54068 18674
rect 54012 8428 54068 18622
rect 54796 17666 54852 19068
rect 55132 18452 55188 31500
rect 55916 23492 55972 75628
rect 56140 75682 56196 75694
rect 56140 75630 56142 75682
rect 56194 75630 56196 75682
rect 56140 67228 56196 75630
rect 57036 75684 57092 75694
rect 56140 67172 56308 67228
rect 56140 42532 56196 42542
rect 56028 42530 56196 42532
rect 56028 42478 56142 42530
rect 56194 42478 56196 42530
rect 56028 42476 56196 42478
rect 56028 41746 56084 42476
rect 56140 42466 56196 42476
rect 56140 41860 56196 41870
rect 56140 41766 56196 41804
rect 56028 41694 56030 41746
rect 56082 41694 56084 41746
rect 56028 41682 56084 41694
rect 56252 41636 56308 67172
rect 57036 47012 57092 75628
rect 57036 46946 57092 46956
rect 57596 75122 57652 76412
rect 57596 75070 57598 75122
rect 57650 75070 57652 75122
rect 56700 43652 56756 43662
rect 56700 42866 56756 43596
rect 56700 42814 56702 42866
rect 56754 42814 56756 42866
rect 56700 42802 56756 42814
rect 57596 42866 57652 75070
rect 57708 74788 57764 76972
rect 58044 76804 58100 76814
rect 58044 75236 58100 76748
rect 58268 76692 58324 79200
rect 58156 76636 58324 76692
rect 58156 75460 58212 76636
rect 58268 76468 58324 76478
rect 58828 76468 58884 76478
rect 58268 76466 58548 76468
rect 58268 76414 58270 76466
rect 58322 76414 58548 76466
rect 58268 76412 58548 76414
rect 58268 76402 58324 76412
rect 58156 75394 58212 75404
rect 58044 75180 58212 75236
rect 58044 74788 58100 74798
rect 57708 74786 58100 74788
rect 57708 74734 58046 74786
rect 58098 74734 58100 74786
rect 57708 74732 58100 74734
rect 58044 74722 58100 74732
rect 57596 42814 57598 42866
rect 57650 42814 57652 42866
rect 57596 42802 57652 42814
rect 57148 42754 57204 42766
rect 57148 42702 57150 42754
rect 57202 42702 57204 42754
rect 57148 42194 57204 42702
rect 57148 42142 57150 42194
rect 57202 42142 57204 42194
rect 57148 42130 57204 42142
rect 58044 42754 58100 42766
rect 58044 42702 58046 42754
rect 58098 42702 58100 42754
rect 58044 42194 58100 42702
rect 58044 42142 58046 42194
rect 58098 42142 58100 42194
rect 58044 42130 58100 42142
rect 55916 23426 55972 23436
rect 56140 41580 56308 41636
rect 56588 41858 56644 41870
rect 56588 41806 56590 41858
rect 56642 41806 56644 41858
rect 56028 21812 56084 21822
rect 56028 21718 56084 21756
rect 55580 21700 55636 21710
rect 55580 21606 55636 21644
rect 55580 20916 55636 20926
rect 55580 20802 55636 20860
rect 55580 20750 55582 20802
rect 55634 20750 55636 20802
rect 55580 20738 55636 20750
rect 56140 20916 56196 41580
rect 56252 40962 56308 40974
rect 56252 40910 56254 40962
rect 56306 40910 56308 40962
rect 56252 40852 56308 40910
rect 56252 40292 56308 40796
rect 56588 40852 56644 41806
rect 57484 41858 57540 41870
rect 57484 41806 57486 41858
rect 57538 41806 57540 41858
rect 56812 41748 56868 41758
rect 56812 41654 56868 41692
rect 57484 41524 57540 41806
rect 57708 41748 57764 41758
rect 57708 41654 57764 41692
rect 57148 41468 57484 41524
rect 57148 41298 57204 41468
rect 57148 41246 57150 41298
rect 57202 41246 57204 41298
rect 57148 41234 57204 41246
rect 56588 40786 56644 40796
rect 56252 40226 56308 40236
rect 56812 39284 56868 39294
rect 56812 35924 56868 39228
rect 56812 35830 56868 35868
rect 56700 35588 56756 35598
rect 56700 26908 56756 35532
rect 56700 26852 56868 26908
rect 56140 20802 56196 20860
rect 56140 20750 56142 20802
rect 56194 20750 56196 20802
rect 56140 20738 56196 20750
rect 55244 20692 55300 20702
rect 55244 20130 55300 20636
rect 56252 20692 56308 20702
rect 56252 20598 56308 20636
rect 55244 20078 55246 20130
rect 55298 20078 55300 20130
rect 55244 20066 55300 20078
rect 55692 20578 55748 20590
rect 55692 20526 55694 20578
rect 55746 20526 55748 20578
rect 55468 19234 55524 19246
rect 55468 19182 55470 19234
rect 55522 19182 55524 19234
rect 55468 19124 55524 19182
rect 55468 19058 55524 19068
rect 55132 18358 55188 18396
rect 55356 19010 55412 19022
rect 55356 18958 55358 19010
rect 55410 18958 55412 19010
rect 54796 17614 54798 17666
rect 54850 17614 54852 17666
rect 54796 17332 54852 17614
rect 54796 17266 54852 17276
rect 55020 17442 55076 17454
rect 55020 17390 55022 17442
rect 55074 17390 55076 17442
rect 54572 16994 54628 17006
rect 54572 16942 54574 16994
rect 54626 16942 54628 16994
rect 54572 16098 54628 16942
rect 54572 16046 54574 16098
rect 54626 16046 54628 16098
rect 54572 15426 54628 16046
rect 54572 15374 54574 15426
rect 54626 15374 54628 15426
rect 54460 15314 54516 15326
rect 54460 15262 54462 15314
rect 54514 15262 54516 15314
rect 54460 14980 54516 15262
rect 54460 14914 54516 14924
rect 54572 14756 54628 15374
rect 54684 16882 54740 16894
rect 54684 16830 54686 16882
rect 54738 16830 54740 16882
rect 54684 15316 54740 16830
rect 54684 15250 54740 15260
rect 54796 16098 54852 16110
rect 54796 16046 54798 16098
rect 54850 16046 54852 16098
rect 54572 14690 54628 14700
rect 54796 14644 54852 16046
rect 54796 14578 54852 14588
rect 54236 13860 54292 13870
rect 54236 13766 54292 13804
rect 53900 8372 54068 8428
rect 54236 13188 54292 13198
rect 53900 7476 53956 8372
rect 53900 7410 53956 7420
rect 53900 5236 53956 5246
rect 53900 4340 53956 5180
rect 54012 5236 54068 5246
rect 54236 5236 54292 13132
rect 55020 9380 55076 17390
rect 55132 13972 55188 13982
rect 55132 13878 55188 13916
rect 55356 13748 55412 18958
rect 55692 18562 55748 20526
rect 56700 20132 56756 20142
rect 56700 20038 56756 20076
rect 55804 20020 55860 20030
rect 55804 19926 55860 19964
rect 56588 19572 56644 19582
rect 55692 18510 55694 18562
rect 55746 18510 55748 18562
rect 55692 18498 55748 18510
rect 56140 19234 56196 19246
rect 56140 19182 56142 19234
rect 56194 19182 56196 19234
rect 56140 19124 56196 19182
rect 55692 17666 55748 17678
rect 55692 17614 55694 17666
rect 55746 17614 55748 17666
rect 55692 16884 55748 17614
rect 56028 16884 56084 16894
rect 55692 16882 56084 16884
rect 55692 16830 56030 16882
rect 56082 16830 56084 16882
rect 55692 16828 56084 16830
rect 55020 9314 55076 9324
rect 55244 13692 55412 13748
rect 55244 7588 55300 13692
rect 56028 11732 56084 16828
rect 56028 11666 56084 11676
rect 55244 7522 55300 7532
rect 55356 11396 55412 11406
rect 54012 5234 54292 5236
rect 54012 5182 54014 5234
rect 54066 5182 54292 5234
rect 54012 5180 54292 5182
rect 54012 5170 54068 5180
rect 54236 5122 54292 5180
rect 55244 5236 55300 5246
rect 55244 5142 55300 5180
rect 54236 5070 54238 5122
rect 54290 5070 54292 5122
rect 54236 5058 54292 5070
rect 55356 5012 55412 11340
rect 56028 11284 56084 11294
rect 56028 6130 56084 11228
rect 56140 11172 56196 19068
rect 56588 17666 56644 19516
rect 56700 18340 56756 18350
rect 56700 18246 56756 18284
rect 56588 17614 56590 17666
rect 56642 17614 56644 17666
rect 56588 17602 56644 17614
rect 56812 17666 56868 26852
rect 57484 23156 57540 41468
rect 58156 38948 58212 75180
rect 58492 74226 58548 76412
rect 58828 76374 58884 76412
rect 58940 75348 58996 79200
rect 59612 76468 59668 79200
rect 59836 76692 59892 76702
rect 59836 76598 59892 76636
rect 59612 76402 59668 76412
rect 59052 75684 59108 75694
rect 59052 75682 59556 75684
rect 59052 75630 59054 75682
rect 59106 75630 59556 75682
rect 59052 75628 59556 75630
rect 59052 75618 59108 75628
rect 59388 75460 59444 75470
rect 58940 75282 58996 75292
rect 59164 75404 59388 75460
rect 58492 74174 58494 74226
rect 58546 74174 58548 74226
rect 58492 45332 58548 74174
rect 59164 74226 59220 75404
rect 59388 75366 59444 75404
rect 59164 74174 59166 74226
rect 59218 74174 59220 74226
rect 59164 74162 59220 74174
rect 59500 74226 59556 75628
rect 60284 75572 60340 79200
rect 60956 75572 61012 79200
rect 61628 77028 61684 79200
rect 61628 76962 61684 76972
rect 62300 77026 62356 79200
rect 62300 76974 62302 77026
rect 62354 76974 62356 77026
rect 62300 76962 62356 76974
rect 62860 77028 62916 77038
rect 61964 76916 62020 76926
rect 61740 76580 61796 76590
rect 61404 76578 61796 76580
rect 61404 76526 61742 76578
rect 61794 76526 61796 76578
rect 61404 76524 61796 76526
rect 61180 75572 61236 75582
rect 60956 75516 61124 75572
rect 60284 75506 60340 75516
rect 59500 74174 59502 74226
rect 59554 74174 59556 74226
rect 58492 45266 58548 45276
rect 58604 53844 58660 53854
rect 58492 42868 58548 42878
rect 58492 42774 58548 42812
rect 58380 41748 58436 41758
rect 58380 41074 58436 41692
rect 58380 41022 58382 41074
rect 58434 41022 58436 41074
rect 58380 41010 58436 41022
rect 58156 38882 58212 38892
rect 57484 23090 57540 23100
rect 57932 37156 57988 37166
rect 57148 20916 57204 20926
rect 57148 20822 57204 20860
rect 57372 19124 57428 19134
rect 57372 19030 57428 19068
rect 57148 18452 57204 18462
rect 57148 18358 57204 18396
rect 56812 17614 56814 17666
rect 56866 17614 56868 17666
rect 56812 17106 56868 17614
rect 56812 17054 56814 17106
rect 56866 17054 56868 17106
rect 56812 17042 56868 17054
rect 57148 17668 57204 17678
rect 57148 17106 57204 17612
rect 57148 17054 57150 17106
rect 57202 17054 57204 17106
rect 57148 14868 57204 17054
rect 57932 16996 57988 37100
rect 58604 31780 58660 53788
rect 59500 43764 59556 74174
rect 59500 43698 59556 43708
rect 59724 75458 59780 75470
rect 59724 75406 59726 75458
rect 59778 75406 59780 75458
rect 59724 41300 59780 75406
rect 60508 75458 60564 75470
rect 60508 75406 60510 75458
rect 60562 75406 60564 75458
rect 60508 75348 60564 75406
rect 60844 75460 60900 75470
rect 61068 75460 61124 75516
rect 61180 75478 61236 75516
rect 60844 75458 61012 75460
rect 60844 75406 60846 75458
rect 60898 75406 61012 75458
rect 60844 75404 61012 75406
rect 60844 75394 60900 75404
rect 60508 75282 60564 75292
rect 60396 74900 60452 74910
rect 60844 74900 60900 74910
rect 60396 74898 60900 74900
rect 60396 74846 60398 74898
rect 60450 74846 60846 74898
rect 60898 74846 60900 74898
rect 60396 74844 60900 74846
rect 60396 73948 60452 74844
rect 60844 74834 60900 74844
rect 59948 73892 60452 73948
rect 59948 42868 60004 73892
rect 60956 67284 61012 75404
rect 61068 75394 61124 75404
rect 61292 75348 61348 75358
rect 61292 75122 61348 75292
rect 61292 75070 61294 75122
rect 61346 75070 61348 75122
rect 61292 75058 61348 75070
rect 61404 67508 61460 76524
rect 61740 76514 61796 76524
rect 61740 75684 61796 75694
rect 61740 75590 61796 75628
rect 61516 75572 61572 75582
rect 61572 75516 61684 75572
rect 61516 75506 61572 75516
rect 61628 75124 61684 75516
rect 61740 75124 61796 75134
rect 61628 75122 61796 75124
rect 61628 75070 61742 75122
rect 61794 75070 61796 75122
rect 61628 75068 61796 75070
rect 61740 75058 61796 75068
rect 60956 67218 61012 67228
rect 61180 67452 61460 67508
rect 59948 42802 60004 42812
rect 59724 41234 59780 41244
rect 60508 41186 60564 41198
rect 60508 41134 60510 41186
rect 60562 41134 60564 41186
rect 58716 41074 58772 41086
rect 58716 41022 58718 41074
rect 58770 41022 58772 41074
rect 58716 40404 58772 41022
rect 59836 40516 59892 40526
rect 59836 40422 59892 40460
rect 58716 40338 58772 40348
rect 60060 40404 60116 40414
rect 60060 40310 60116 40348
rect 60508 40404 60564 41134
rect 61068 41076 61124 41086
rect 61068 40982 61124 41020
rect 60956 40516 61012 40526
rect 60508 40338 60564 40348
rect 60732 40402 60788 40414
rect 60732 40350 60734 40402
rect 60786 40350 60788 40402
rect 60172 40290 60228 40302
rect 60172 40238 60174 40290
rect 60226 40238 60228 40290
rect 58604 31714 58660 31724
rect 58828 33236 58884 33246
rect 58828 30212 58884 33180
rect 58828 30146 58884 30156
rect 58940 31668 58996 31678
rect 58940 29428 58996 31612
rect 58940 29362 58996 29372
rect 59612 30996 59668 31006
rect 58716 17668 58772 17678
rect 58716 17574 58772 17612
rect 58828 17554 58884 17566
rect 58828 17502 58830 17554
rect 58882 17502 58884 17554
rect 58380 17444 58436 17454
rect 58380 17350 58436 17388
rect 58828 17332 58884 17502
rect 58828 17266 58884 17276
rect 57932 16930 57988 16940
rect 57148 14802 57204 14812
rect 57932 15204 57988 15214
rect 56140 11106 56196 11116
rect 57148 10164 57204 10174
rect 56028 6078 56030 6130
rect 56082 6078 56084 6130
rect 56028 5908 56084 6078
rect 56028 5842 56084 5852
rect 56588 9940 56644 9950
rect 56140 5236 56196 5246
rect 55356 4956 55972 5012
rect 53900 4284 54068 4340
rect 53788 4162 53844 4172
rect 53900 4116 53956 4126
rect 53900 4022 53956 4060
rect 53676 3556 53732 3566
rect 53676 3462 53732 3500
rect 53452 3390 53454 3442
rect 53506 3390 53508 3442
rect 53452 3378 53508 3390
rect 54012 800 54068 4284
rect 54684 4116 54740 4126
rect 54236 3780 54292 3790
rect 54236 3666 54292 3724
rect 54236 3614 54238 3666
rect 54290 3614 54292 3666
rect 54236 3602 54292 3614
rect 54684 800 54740 4060
rect 55356 3556 55412 3566
rect 55356 800 55412 3500
rect 55468 3554 55524 4956
rect 55916 4562 55972 4956
rect 55916 4510 55918 4562
rect 55970 4510 55972 4562
rect 55916 4498 55972 4510
rect 56028 3668 56084 3678
rect 56028 3574 56084 3612
rect 55468 3502 55470 3554
rect 55522 3502 55524 3554
rect 55468 3490 55524 3502
rect 56140 2324 56196 5180
rect 56588 4338 56644 9884
rect 56812 6692 56868 6702
rect 56812 6466 56868 6636
rect 56812 6414 56814 6466
rect 56866 6414 56868 6466
rect 56588 4286 56590 4338
rect 56642 4286 56644 4338
rect 56588 3668 56644 4286
rect 56588 3602 56644 3612
rect 56700 5684 56756 5694
rect 56028 2268 56196 2324
rect 56028 800 56084 2268
rect 56700 800 56756 5628
rect 56812 5124 56868 6414
rect 56924 5908 56980 5918
rect 56924 5814 56980 5852
rect 57148 5908 57204 10108
rect 57932 7812 57988 15148
rect 59612 9828 59668 30940
rect 59612 9762 59668 9772
rect 59948 27412 60004 27422
rect 59948 8428 60004 27356
rect 60172 25732 60228 40238
rect 60732 40292 60788 40350
rect 60732 39618 60788 40236
rect 60732 39566 60734 39618
rect 60786 39566 60788 39618
rect 60732 39554 60788 39566
rect 60620 39394 60676 39406
rect 60620 39342 60622 39394
rect 60674 39342 60676 39394
rect 60508 37716 60564 37726
rect 60508 35028 60564 37660
rect 60508 34962 60564 34972
rect 60172 25666 60228 25676
rect 60620 23716 60676 39342
rect 60956 39058 61012 40460
rect 61068 40404 61124 40414
rect 61068 39618 61124 40348
rect 61068 39566 61070 39618
rect 61122 39566 61124 39618
rect 61068 39554 61124 39566
rect 61180 39732 61236 67452
rect 61292 67284 61348 67294
rect 61292 40516 61348 67228
rect 61964 67228 62020 76860
rect 62636 76580 62692 76590
rect 62300 76578 62692 76580
rect 62300 76526 62638 76578
rect 62690 76526 62692 76578
rect 62300 76524 62692 76526
rect 62076 76468 62132 76478
rect 62076 76374 62132 76412
rect 62076 75570 62132 75582
rect 62076 75518 62078 75570
rect 62130 75518 62132 75570
rect 62076 75460 62132 75518
rect 62076 75124 62132 75404
rect 62188 75124 62244 75134
rect 62076 75122 62244 75124
rect 62076 75070 62190 75122
rect 62242 75070 62244 75122
rect 62076 75068 62244 75070
rect 62188 75058 62244 75068
rect 61964 67172 62132 67228
rect 61852 58212 61908 58222
rect 61852 50428 61908 58156
rect 61740 50372 61908 50428
rect 61628 41970 61684 41982
rect 61628 41918 61630 41970
rect 61682 41918 61684 41970
rect 61292 40450 61348 40460
rect 61516 41300 61572 41310
rect 61516 40514 61572 41244
rect 61628 41076 61684 41918
rect 61628 41010 61684 41020
rect 61516 40462 61518 40514
rect 61570 40462 61572 40514
rect 61516 40450 61572 40462
rect 61180 39506 61236 39676
rect 61180 39454 61182 39506
rect 61234 39454 61236 39506
rect 61180 39442 61236 39454
rect 61404 40290 61460 40302
rect 61404 40238 61406 40290
rect 61458 40238 61460 40290
rect 60956 39006 60958 39058
rect 61010 39006 61012 39058
rect 60956 38994 61012 39006
rect 61404 28308 61460 40238
rect 61740 29652 61796 50372
rect 62076 42756 62132 67172
rect 62076 42690 62132 42700
rect 62188 47012 62244 47022
rect 62188 42532 62244 46956
rect 62132 42476 62244 42532
rect 62300 42532 62356 76524
rect 62636 76514 62692 76524
rect 62748 76468 62804 76478
rect 62748 75572 62804 76412
rect 62860 76466 62916 76972
rect 62972 76692 63028 79200
rect 62972 76626 63028 76636
rect 63308 77026 63364 77038
rect 63308 76974 63310 77026
rect 63362 76974 63364 77026
rect 63308 76690 63364 76974
rect 63644 77026 63700 79200
rect 64316 77138 64372 79200
rect 64316 77086 64318 77138
rect 64370 77086 64372 77138
rect 64316 77074 64372 77086
rect 63644 76974 63646 77026
rect 63698 76974 63700 77026
rect 63644 76962 63700 76974
rect 64652 77026 64708 77038
rect 64652 76974 64654 77026
rect 64706 76974 64708 77026
rect 63308 76638 63310 76690
rect 63362 76638 63364 76690
rect 62860 76414 62862 76466
rect 62914 76414 62916 76466
rect 62860 75684 62916 76414
rect 63308 75906 63364 76638
rect 63980 76692 64036 76702
rect 64036 76636 64260 76692
rect 63980 76598 64036 76636
rect 63308 75854 63310 75906
rect 63362 75854 63364 75906
rect 63308 75842 63364 75854
rect 63644 76578 63700 76590
rect 63644 76526 63646 76578
rect 63698 76526 63700 76578
rect 63308 75684 63364 75694
rect 62860 75682 63364 75684
rect 62860 75630 63310 75682
rect 63362 75630 63364 75682
rect 62860 75628 63364 75630
rect 63308 75618 63364 75628
rect 62748 75516 62916 75572
rect 62412 75460 62468 75470
rect 62412 75458 62804 75460
rect 62412 75406 62414 75458
rect 62466 75406 62804 75458
rect 62412 75404 62804 75406
rect 62412 75394 62468 75404
rect 62748 67228 62804 75404
rect 62860 75458 62916 75516
rect 62860 75406 62862 75458
rect 62914 75406 62916 75458
rect 62860 75394 62916 75406
rect 62748 67172 62916 67228
rect 62860 50428 62916 67172
rect 63644 50428 63700 76526
rect 63756 75906 63812 75918
rect 63756 75854 63758 75906
rect 63810 75854 63812 75906
rect 63756 75794 63812 75854
rect 63756 75742 63758 75794
rect 63810 75742 63812 75794
rect 63756 75730 63812 75742
rect 64204 75794 64260 76636
rect 64652 76690 64708 76974
rect 64988 76804 65044 79200
rect 65324 77138 65380 77150
rect 65324 77086 65326 77138
rect 65378 77086 65380 77138
rect 64988 76748 65156 76804
rect 64652 76638 64654 76690
rect 64706 76638 64708 76690
rect 64316 76580 64372 76590
rect 64316 76578 64596 76580
rect 64316 76526 64318 76578
rect 64370 76526 64596 76578
rect 64316 76524 64596 76526
rect 64316 76514 64372 76524
rect 64204 75742 64206 75794
rect 64258 75742 64260 75794
rect 64204 75730 64260 75742
rect 62412 50372 62916 50428
rect 63420 50372 63700 50428
rect 63756 75572 63812 75582
rect 62412 42868 62468 50372
rect 62412 42866 62916 42868
rect 62412 42814 62414 42866
rect 62466 42814 62916 42866
rect 62412 42812 62916 42814
rect 62412 42802 62468 42812
rect 62300 42476 62692 42532
rect 62132 42196 62188 42476
rect 62132 42140 62580 42196
rect 62188 41860 62244 41870
rect 61852 41858 62244 41860
rect 61852 41806 62190 41858
rect 62242 41806 62244 41858
rect 61852 41804 62244 41806
rect 61852 41186 61908 41804
rect 62188 41636 62244 41804
rect 62188 41570 62244 41580
rect 61852 41134 61854 41186
rect 61906 41134 61908 41186
rect 61852 41122 61908 41134
rect 62188 41412 62244 41422
rect 62188 41186 62244 41356
rect 62188 41134 62190 41186
rect 62242 41134 62244 41186
rect 62188 41122 62244 41134
rect 62412 41188 62468 41198
rect 62412 41094 62468 41132
rect 61740 29586 61796 29596
rect 62076 40962 62132 40974
rect 62076 40910 62078 40962
rect 62130 40910 62132 40962
rect 62076 28532 62132 40910
rect 62524 40516 62580 42140
rect 62636 41860 62692 42476
rect 62860 42082 62916 42812
rect 62860 42030 62862 42082
rect 62914 42030 62916 42082
rect 62860 42018 62916 42030
rect 62636 41412 62692 41804
rect 62636 41346 62692 41356
rect 62748 41970 62804 41982
rect 62748 41918 62750 41970
rect 62802 41918 62804 41970
rect 62748 41188 62804 41918
rect 63308 41970 63364 41982
rect 63308 41918 63310 41970
rect 63362 41918 63364 41970
rect 63084 41860 63140 41870
rect 62748 41122 62804 41132
rect 62860 41858 63140 41860
rect 62860 41806 63086 41858
rect 63138 41806 63140 41858
rect 62860 41804 63140 41806
rect 62300 40514 62580 40516
rect 62300 40462 62526 40514
rect 62578 40462 62580 40514
rect 62300 40460 62580 40462
rect 62188 40402 62244 40414
rect 62188 40350 62190 40402
rect 62242 40350 62244 40402
rect 62188 40292 62244 40350
rect 62188 40226 62244 40236
rect 62300 39730 62356 40460
rect 62524 40450 62580 40460
rect 62300 39678 62302 39730
rect 62354 39678 62356 39730
rect 62300 39666 62356 39678
rect 62636 39732 62692 39742
rect 62636 39638 62692 39676
rect 62860 38836 62916 41804
rect 63084 41794 63140 41804
rect 63308 41636 63364 41918
rect 62972 41188 63028 41226
rect 63308 41188 63364 41580
rect 62972 41122 63028 41132
rect 63084 41186 63364 41188
rect 63084 41134 63310 41186
rect 63362 41134 63364 41186
rect 63084 41132 63364 41134
rect 62972 40962 63028 40974
rect 62972 40910 62974 40962
rect 63026 40910 63028 40962
rect 62972 38948 63028 40910
rect 63084 40402 63140 41132
rect 63308 41122 63364 41132
rect 63420 41972 63476 50372
rect 63756 43316 63812 75516
rect 64540 71652 64596 76524
rect 64652 75122 64708 76638
rect 64988 76580 65044 76590
rect 64652 75070 64654 75122
rect 64706 75070 64708 75122
rect 64652 75058 64708 75070
rect 64876 76578 65044 76580
rect 64876 76526 64990 76578
rect 65042 76526 65044 76578
rect 64876 76524 65044 76526
rect 64876 72100 64932 76524
rect 64988 76514 65044 76524
rect 64988 75796 65044 75806
rect 65100 75796 65156 76748
rect 65324 76690 65380 77086
rect 65660 77026 65716 79200
rect 66332 77138 66388 79200
rect 66332 77086 66334 77138
rect 66386 77086 66388 77138
rect 66332 77074 66388 77086
rect 65660 76974 65662 77026
rect 65714 76974 65716 77026
rect 65660 76962 65716 76974
rect 66444 77026 66500 77038
rect 66444 76974 66446 77026
rect 66498 76974 66500 77026
rect 65324 76638 65326 76690
rect 65378 76638 65380 76690
rect 65324 75796 65380 76638
rect 66444 76690 66500 76974
rect 67004 77028 67060 79200
rect 67004 76962 67060 76972
rect 67116 77138 67172 77150
rect 67116 77086 67118 77138
rect 67170 77086 67172 77138
rect 67116 76692 67172 77086
rect 67676 77026 67732 79200
rect 67676 76974 67678 77026
rect 67730 76974 67732 77026
rect 67676 76962 67732 76974
rect 67788 77028 67844 77038
rect 67788 76692 67844 76972
rect 66444 76638 66446 76690
rect 66498 76638 66500 76690
rect 64988 75794 65268 75796
rect 64988 75742 64990 75794
rect 65042 75742 65268 75794
rect 64988 75740 65268 75742
rect 64988 75730 65044 75740
rect 65212 75682 65268 75740
rect 65324 75730 65380 75740
rect 65660 76578 65716 76590
rect 65660 76526 65662 76578
rect 65714 76526 65716 76578
rect 65212 75630 65214 75682
rect 65266 75630 65268 75682
rect 65212 75618 65268 75630
rect 65548 75460 65604 75470
rect 65548 75366 65604 75404
rect 65324 73444 65380 73454
rect 64876 72044 65268 72100
rect 64540 71596 65156 71652
rect 63756 43250 63812 43260
rect 64876 67284 64932 67294
rect 63420 41074 63476 41916
rect 64540 41972 64596 41982
rect 64540 41878 64596 41916
rect 64876 41972 64932 67228
rect 64876 41906 64932 41916
rect 63644 41860 63700 41870
rect 63644 41766 63700 41804
rect 63420 41022 63422 41074
rect 63474 41022 63476 41074
rect 63420 41010 63476 41022
rect 64204 41188 64260 41198
rect 63532 40628 63588 40638
rect 63532 40626 63812 40628
rect 63532 40574 63534 40626
rect 63586 40574 63812 40626
rect 63532 40572 63812 40574
rect 63532 40562 63588 40572
rect 63420 40404 63476 40414
rect 63084 40350 63086 40402
rect 63138 40350 63140 40402
rect 63084 40338 63140 40350
rect 63196 40402 63476 40404
rect 63196 40350 63422 40402
rect 63474 40350 63476 40402
rect 63196 40348 63476 40350
rect 63196 40292 63252 40348
rect 63420 40338 63476 40348
rect 63196 39730 63252 40236
rect 63196 39678 63198 39730
rect 63250 39678 63252 39730
rect 63196 39666 63252 39678
rect 63644 39396 63700 39406
rect 63308 39340 63644 39396
rect 63308 39058 63364 39340
rect 63644 39302 63700 39340
rect 63308 39006 63310 39058
rect 63362 39006 63364 39058
rect 63308 38994 63364 39006
rect 62972 38892 63140 38948
rect 62636 38780 62916 38836
rect 62636 35308 62692 38780
rect 62972 38724 63028 38734
rect 62972 38612 63028 38668
rect 62860 38556 63028 38612
rect 63084 38612 63140 38892
rect 63532 38834 63588 38846
rect 63532 38782 63534 38834
rect 63586 38782 63588 38834
rect 63532 38724 63588 38782
rect 63532 38658 63588 38668
rect 63084 38556 63364 38612
rect 62860 36596 62916 38556
rect 62860 36530 62916 36540
rect 63308 35308 63364 38556
rect 62636 35252 62804 35308
rect 62076 28466 62132 28476
rect 61404 28242 61460 28252
rect 61292 27300 61348 27310
rect 61292 24500 61348 27244
rect 62748 24722 62804 35252
rect 63084 35252 63364 35308
rect 62860 28532 62916 28542
rect 62860 25506 62916 28476
rect 63084 26292 63140 35252
rect 63084 26226 63140 26236
rect 63196 34132 63252 34142
rect 62860 25454 62862 25506
rect 62914 25454 62916 25506
rect 62860 25442 62916 25454
rect 63196 25506 63252 34076
rect 63308 25620 63364 25630
rect 63308 25526 63364 25564
rect 63196 25454 63198 25506
rect 63250 25454 63252 25506
rect 63196 25442 63252 25454
rect 63420 25284 63476 25294
rect 63420 25282 63588 25284
rect 63420 25230 63422 25282
rect 63474 25230 63588 25282
rect 63420 25228 63588 25230
rect 63420 25218 63476 25228
rect 63196 25172 63252 25182
rect 63196 24946 63252 25116
rect 63196 24894 63198 24946
rect 63250 24894 63252 24946
rect 63196 24882 63252 24894
rect 62748 24670 62750 24722
rect 62802 24670 62804 24722
rect 62748 24658 62804 24670
rect 63420 24722 63476 24734
rect 63420 24670 63422 24722
rect 63474 24670 63476 24722
rect 61292 24434 61348 24444
rect 63308 24610 63364 24622
rect 63308 24558 63310 24610
rect 63362 24558 63364 24610
rect 63308 24164 63364 24558
rect 63308 24098 63364 24108
rect 60620 23650 60676 23660
rect 63420 23604 63476 24670
rect 63420 23538 63476 23548
rect 63532 23268 63588 25228
rect 63756 24948 63812 40572
rect 64204 40404 64260 41132
rect 64428 41186 64484 41198
rect 64428 41134 64430 41186
rect 64482 41134 64484 41186
rect 64428 40964 64484 41134
rect 64876 41188 64932 41198
rect 64876 41094 64932 41132
rect 64428 40898 64484 40908
rect 65100 40516 65156 71596
rect 65212 67284 65268 72044
rect 65212 67218 65268 67228
rect 65324 67228 65380 73388
rect 65660 67228 65716 76526
rect 65916 76076 66180 76086
rect 65972 76020 66020 76076
rect 66076 76020 66124 76076
rect 65916 76010 66180 76020
rect 65996 75796 66052 75806
rect 65996 75702 66052 75740
rect 66444 75794 66500 76638
rect 67004 76690 67172 76692
rect 67004 76638 67118 76690
rect 67170 76638 67172 76690
rect 67004 76636 67172 76638
rect 66444 75742 66446 75794
rect 66498 75742 66500 75794
rect 66444 75730 66500 75742
rect 66780 76578 66836 76590
rect 66780 76526 66782 76578
rect 66834 76526 66836 76578
rect 65916 74508 66180 74518
rect 65972 74452 66020 74508
rect 66076 74452 66124 74508
rect 65916 74442 66180 74452
rect 65916 72940 66180 72950
rect 65972 72884 66020 72940
rect 66076 72884 66124 72940
rect 65916 72874 66180 72884
rect 65916 71372 66180 71382
rect 65972 71316 66020 71372
rect 66076 71316 66124 71372
rect 65916 71306 66180 71316
rect 65916 69804 66180 69814
rect 65972 69748 66020 69804
rect 66076 69748 66124 69804
rect 65916 69738 66180 69748
rect 65916 68236 66180 68246
rect 65972 68180 66020 68236
rect 66076 68180 66124 68236
rect 65916 68170 66180 68180
rect 65324 67172 65492 67228
rect 65660 67172 66388 67228
rect 65212 56196 65268 56206
rect 65212 40740 65268 56140
rect 65324 41972 65380 41982
rect 65324 41298 65380 41916
rect 65324 41246 65326 41298
rect 65378 41246 65380 41298
rect 65324 41076 65380 41246
rect 65324 41010 65380 41020
rect 65212 40684 65380 40740
rect 65100 40422 65156 40460
rect 64428 40404 64484 40414
rect 64204 40402 64484 40404
rect 64204 40350 64430 40402
rect 64482 40350 64484 40402
rect 64204 40348 64484 40350
rect 63980 39508 64036 39518
rect 64204 39508 64260 40348
rect 64428 40338 64484 40348
rect 63980 39506 64260 39508
rect 63980 39454 63982 39506
rect 64034 39454 64260 39506
rect 63980 39452 64260 39454
rect 64876 40290 64932 40302
rect 64876 40238 64878 40290
rect 64930 40238 64932 40290
rect 63980 39442 64036 39452
rect 64316 39396 64372 39406
rect 64316 38836 64372 39340
rect 64316 38770 64372 38780
rect 63868 27972 63924 27982
rect 63868 26180 63924 27916
rect 64876 27860 64932 40238
rect 65212 38836 65268 38846
rect 65212 38742 65268 38780
rect 64876 27794 64932 27804
rect 65324 27300 65380 40684
rect 65436 35812 65492 67172
rect 65916 66668 66180 66678
rect 65972 66612 66020 66668
rect 66076 66612 66124 66668
rect 65916 66602 66180 66612
rect 65916 65100 66180 65110
rect 65972 65044 66020 65100
rect 66076 65044 66124 65100
rect 65916 65034 66180 65044
rect 65916 63532 66180 63542
rect 65972 63476 66020 63532
rect 66076 63476 66124 63532
rect 65916 63466 66180 63476
rect 66332 62188 66388 67172
rect 66780 62188 66836 76526
rect 67004 75794 67060 76636
rect 67116 76626 67172 76636
rect 67564 76690 67844 76692
rect 67564 76638 67790 76690
rect 67842 76638 67844 76690
rect 67564 76636 67844 76638
rect 67004 75742 67006 75794
rect 67058 75742 67060 75794
rect 67004 75730 67060 75742
rect 67452 76578 67508 76590
rect 67452 76526 67454 76578
rect 67506 76526 67508 76578
rect 66892 75460 66948 75470
rect 66892 67228 66948 75404
rect 67452 67228 67508 76526
rect 67564 75794 67620 76636
rect 67788 76626 67844 76636
rect 68348 76692 68404 79200
rect 69020 77250 69076 79200
rect 69020 77198 69022 77250
rect 69074 77198 69076 77250
rect 69020 77186 69076 77198
rect 68348 76626 68404 76636
rect 68460 77026 68516 77038
rect 68460 76974 68462 77026
rect 68514 76974 68516 77026
rect 68460 76690 68516 76974
rect 68460 76638 68462 76690
rect 68514 76638 68516 76690
rect 67564 75742 67566 75794
rect 67618 75742 67620 75794
rect 67564 75730 67620 75742
rect 68124 76578 68180 76590
rect 68124 76526 68126 76578
rect 68178 76526 68180 76578
rect 66892 67172 67172 67228
rect 67452 67172 67732 67228
rect 66332 62132 66500 62188
rect 66780 62132 67060 62188
rect 65916 61964 66180 61974
rect 65972 61908 66020 61964
rect 66076 61908 66124 61964
rect 65916 61898 66180 61908
rect 65916 60396 66180 60406
rect 65972 60340 66020 60396
rect 66076 60340 66124 60396
rect 65916 60330 66180 60340
rect 65916 58828 66180 58838
rect 65972 58772 66020 58828
rect 66076 58772 66124 58828
rect 65916 58762 66180 58772
rect 65916 57260 66180 57270
rect 65972 57204 66020 57260
rect 66076 57204 66124 57260
rect 65916 57194 66180 57204
rect 65916 55692 66180 55702
rect 65972 55636 66020 55692
rect 66076 55636 66124 55692
rect 65916 55626 66180 55636
rect 65916 54124 66180 54134
rect 65972 54068 66020 54124
rect 66076 54068 66124 54124
rect 65916 54058 66180 54068
rect 65916 52556 66180 52566
rect 65972 52500 66020 52556
rect 66076 52500 66124 52556
rect 65916 52490 66180 52500
rect 65916 50988 66180 50998
rect 65972 50932 66020 50988
rect 66076 50932 66124 50988
rect 65916 50922 66180 50932
rect 65916 49420 66180 49430
rect 65972 49364 66020 49420
rect 66076 49364 66124 49420
rect 65916 49354 66180 49364
rect 65916 47852 66180 47862
rect 65972 47796 66020 47852
rect 66076 47796 66124 47852
rect 65916 47786 66180 47796
rect 65916 46284 66180 46294
rect 65972 46228 66020 46284
rect 66076 46228 66124 46284
rect 65916 46218 66180 46228
rect 65916 44716 66180 44726
rect 65972 44660 66020 44716
rect 66076 44660 66124 44716
rect 65916 44650 66180 44660
rect 65916 43148 66180 43158
rect 65972 43092 66020 43148
rect 66076 43092 66124 43148
rect 65916 43082 66180 43092
rect 65916 41580 66180 41590
rect 65972 41524 66020 41580
rect 66076 41524 66124 41580
rect 65916 41514 66180 41524
rect 65660 41188 65716 41198
rect 65548 40404 65604 40414
rect 65660 40404 65716 41132
rect 65772 41076 65828 41086
rect 65772 40982 65828 41020
rect 66444 40964 66500 62132
rect 66780 41186 66836 41198
rect 66780 41134 66782 41186
rect 66834 41134 66836 41186
rect 66444 40908 66612 40964
rect 66332 40628 66388 40638
rect 66332 40514 66388 40572
rect 66332 40462 66334 40514
rect 66386 40462 66388 40514
rect 66332 40450 66388 40462
rect 65884 40404 65940 40414
rect 65548 40402 65940 40404
rect 65548 40350 65550 40402
rect 65602 40350 65886 40402
rect 65938 40350 65940 40402
rect 65548 40348 65940 40350
rect 65548 40338 65604 40348
rect 65660 39620 65716 39630
rect 65772 39620 65828 40348
rect 65884 40338 65940 40348
rect 66444 40290 66500 40302
rect 66444 40238 66446 40290
rect 66498 40238 66500 40290
rect 65916 40012 66180 40022
rect 65972 39956 66020 40012
rect 66076 39956 66124 40012
rect 65916 39946 66180 39956
rect 66220 39732 66276 39742
rect 66220 39730 66388 39732
rect 66220 39678 66222 39730
rect 66274 39678 66388 39730
rect 66220 39676 66388 39678
rect 66220 39666 66276 39676
rect 66108 39620 66164 39630
rect 65772 39618 66164 39620
rect 65772 39566 66110 39618
rect 66162 39566 66164 39618
rect 65772 39564 66164 39566
rect 65660 38836 65716 39564
rect 66108 39554 66164 39564
rect 66332 39060 66388 39676
rect 66220 39004 66388 39060
rect 65772 38836 65828 38846
rect 66108 38836 66164 38846
rect 65660 38834 66164 38836
rect 65660 38782 65774 38834
rect 65826 38782 66110 38834
rect 66162 38782 66164 38834
rect 65660 38780 66164 38782
rect 65772 38770 65828 38780
rect 66108 38770 66164 38780
rect 66220 38668 66276 39004
rect 65436 35746 65492 35756
rect 65660 38612 66276 38668
rect 66332 38836 66388 38846
rect 65324 27234 65380 27244
rect 63868 26114 63924 26124
rect 63756 24882 63812 24892
rect 63980 25172 64036 25182
rect 63980 24946 64036 25116
rect 63980 24894 63982 24946
rect 64034 24894 64036 24946
rect 63980 24882 64036 24894
rect 63532 23202 63588 23212
rect 61628 22148 61684 22158
rect 61292 21476 61348 21486
rect 57932 7746 57988 7756
rect 59388 8372 60004 8428
rect 60172 19796 60228 19806
rect 59388 5908 59444 8372
rect 59500 8260 59556 8270
rect 59500 6692 59556 8204
rect 60172 7362 60228 19740
rect 60172 7310 60174 7362
rect 60226 7310 60228 7362
rect 60172 7028 60228 7310
rect 59948 6972 60228 7028
rect 60284 12964 60340 12974
rect 59500 6690 59892 6692
rect 59500 6638 59502 6690
rect 59554 6638 59892 6690
rect 59500 6636 59892 6638
rect 59500 6626 59556 6636
rect 59388 5852 59556 5908
rect 57148 5842 57204 5852
rect 57932 5684 57988 5694
rect 57932 5590 57988 5628
rect 59388 5684 59444 5694
rect 58156 5236 58212 5246
rect 58156 5142 58212 5180
rect 57148 5124 57204 5134
rect 56812 5122 57204 5124
rect 56812 5070 57150 5122
rect 57202 5070 57204 5122
rect 56812 5068 57204 5070
rect 57148 5058 57204 5068
rect 58716 4900 58772 4910
rect 57596 4116 57652 4126
rect 57596 4022 57652 4060
rect 58156 3780 58212 3790
rect 58044 3668 58100 3678
rect 58044 3574 58100 3612
rect 57372 3444 57428 3454
rect 57372 800 57428 3388
rect 58156 1652 58212 3724
rect 58044 1596 58212 1652
rect 58044 800 58100 1596
rect 58716 800 58772 4844
rect 59052 3668 59108 3678
rect 59052 3574 59108 3612
rect 59388 800 59444 5628
rect 59500 3556 59556 5852
rect 59836 5906 59892 6636
rect 59836 5854 59838 5906
rect 59890 5854 59892 5906
rect 59836 5842 59892 5854
rect 59948 5124 60004 6972
rect 60060 6692 60116 6702
rect 60284 6692 60340 12908
rect 60508 6692 60564 6702
rect 60060 6690 60564 6692
rect 60060 6638 60062 6690
rect 60114 6638 60510 6690
rect 60562 6638 60564 6690
rect 60060 6636 60564 6638
rect 60060 6626 60116 6636
rect 60508 6626 60564 6636
rect 61292 6692 61348 21420
rect 61292 6626 61348 6636
rect 59948 5058 60004 5068
rect 60060 6468 60116 6478
rect 59500 3490 59556 3500
rect 59724 4114 59780 4126
rect 59724 4062 59726 4114
rect 59778 4062 59780 4114
rect 59724 3444 59780 4062
rect 59724 3378 59780 3388
rect 60060 800 60116 6412
rect 61516 6468 61572 6478
rect 61516 6374 61572 6412
rect 60844 5684 60900 5694
rect 60844 5590 60900 5628
rect 60732 5236 60788 5246
rect 60508 5124 60564 5134
rect 60508 5030 60564 5068
rect 60732 800 60788 5180
rect 61516 4900 61572 4910
rect 61516 4806 61572 4844
rect 61628 4564 61684 22092
rect 65660 21812 65716 38612
rect 65916 38444 66180 38454
rect 65972 38388 66020 38444
rect 66076 38388 66124 38444
rect 65916 38378 66180 38388
rect 66332 38276 66388 38780
rect 66108 38220 66388 38276
rect 66108 38050 66164 38220
rect 66108 37998 66110 38050
rect 66162 37998 66164 38050
rect 66108 37986 66164 37998
rect 65916 36876 66180 36886
rect 65972 36820 66020 36876
rect 66076 36820 66124 36876
rect 65916 36810 66180 36820
rect 65916 35308 66180 35318
rect 65972 35252 66020 35308
rect 66076 35252 66124 35308
rect 65916 35242 66180 35252
rect 65916 33740 66180 33750
rect 65972 33684 66020 33740
rect 66076 33684 66124 33740
rect 65916 33674 66180 33684
rect 65916 32172 66180 32182
rect 65972 32116 66020 32172
rect 66076 32116 66124 32172
rect 65916 32106 66180 32116
rect 65916 30604 66180 30614
rect 65972 30548 66020 30604
rect 66076 30548 66124 30604
rect 65916 30538 66180 30548
rect 65916 29036 66180 29046
rect 65972 28980 66020 29036
rect 66076 28980 66124 29036
rect 65916 28970 66180 28980
rect 65916 27468 66180 27478
rect 65972 27412 66020 27468
rect 66076 27412 66124 27468
rect 65916 27402 66180 27412
rect 65916 25900 66180 25910
rect 65972 25844 66020 25900
rect 66076 25844 66124 25900
rect 65916 25834 66180 25844
rect 65916 24332 66180 24342
rect 65972 24276 66020 24332
rect 66076 24276 66124 24332
rect 65916 24266 66180 24276
rect 65916 22764 66180 22774
rect 65972 22708 66020 22764
rect 66076 22708 66124 22764
rect 65916 22698 66180 22708
rect 65660 21746 65716 21756
rect 66444 21588 66500 40238
rect 66556 39732 66612 40908
rect 66556 39506 66612 39676
rect 66556 39454 66558 39506
rect 66610 39454 66612 39506
rect 66556 39442 66612 39454
rect 66668 40962 66724 40974
rect 66668 40910 66670 40962
rect 66722 40910 66724 40962
rect 66668 39396 66724 40910
rect 66780 40402 66836 41134
rect 66780 40350 66782 40402
rect 66834 40350 66836 40402
rect 66780 39620 66836 40350
rect 66780 39554 66836 39564
rect 67004 39396 67060 62132
rect 67116 41972 67172 67172
rect 67116 41916 67508 41972
rect 67452 40628 67508 41916
rect 67452 40534 67508 40572
rect 67676 40628 67732 67172
rect 68124 58884 68180 76526
rect 68460 75794 68516 76638
rect 69020 77026 69076 77038
rect 69020 76974 69022 77026
rect 69074 76974 69076 77026
rect 69020 76354 69076 76974
rect 69692 77028 69748 79200
rect 69692 76962 69748 76972
rect 70028 77250 70084 77262
rect 70028 77198 70030 77250
rect 70082 77198 70084 77250
rect 69356 76692 69412 76702
rect 69020 76302 69022 76354
rect 69074 76302 69076 76354
rect 69020 76290 69076 76302
rect 69132 76636 69356 76692
rect 68460 75742 68462 75794
rect 68514 75742 68516 75794
rect 68460 75730 68516 75742
rect 69132 75794 69188 76636
rect 69356 76598 69412 76636
rect 69132 75742 69134 75794
rect 69186 75742 69188 75794
rect 69132 75730 69188 75742
rect 69692 76578 69748 76590
rect 69692 76526 69694 76578
rect 69746 76526 69748 76578
rect 68684 75684 68740 75694
rect 68124 58818 68180 58828
rect 68572 71876 68628 71886
rect 68572 50428 68628 71820
rect 67116 39732 67172 39742
rect 67116 39638 67172 39676
rect 66668 39340 66948 39396
rect 66556 38722 66612 38734
rect 66556 38670 66558 38722
rect 66610 38670 66612 38722
rect 66556 38668 66612 38670
rect 66556 38612 66724 38668
rect 66556 38052 66612 38062
rect 66556 37958 66612 37996
rect 66444 21522 66500 21532
rect 63420 21252 63476 21262
rect 63420 8428 63476 21196
rect 65916 21196 66180 21206
rect 63644 21140 63700 21150
rect 65972 21140 66020 21196
rect 66076 21140 66124 21196
rect 65916 21130 66180 21140
rect 63420 8372 63588 8428
rect 63420 6692 63476 6702
rect 63196 6636 63420 6692
rect 62748 6468 62804 6478
rect 61628 4338 61684 4508
rect 62524 4564 62580 4574
rect 62524 4470 62580 4508
rect 61628 4286 61630 4338
rect 61682 4286 61684 4338
rect 61628 4274 61684 4286
rect 62076 3892 62132 3902
rect 61404 3780 61460 3790
rect 60956 3556 61012 3566
rect 60956 3462 61012 3500
rect 61404 800 61460 3724
rect 61852 3556 61908 3566
rect 61852 3462 61908 3500
rect 62076 800 62132 3836
rect 62748 800 62804 6412
rect 63196 6130 63252 6636
rect 63420 6598 63476 6636
rect 63196 6078 63198 6130
rect 63250 6078 63252 6130
rect 63196 6066 63252 6078
rect 63532 5124 63588 8372
rect 63196 5122 63588 5124
rect 63196 5070 63534 5122
rect 63586 5070 63588 5122
rect 63196 5068 63588 5070
rect 63196 4562 63252 5068
rect 63532 5058 63588 5068
rect 63532 4564 63588 4574
rect 63644 4564 63700 21084
rect 66668 20804 66724 38612
rect 66892 22708 66948 39340
rect 67004 38946 67060 39340
rect 67564 39396 67620 39406
rect 67564 39302 67620 39340
rect 67004 38894 67006 38946
rect 67058 38894 67060 38946
rect 67004 38882 67060 38894
rect 67676 38946 67732 40572
rect 68012 50372 68628 50428
rect 67900 40516 67956 40526
rect 67900 40422 67956 40460
rect 67676 38894 67678 38946
rect 67730 38894 67732 38946
rect 67676 38882 67732 38894
rect 67228 38834 67284 38846
rect 67228 38782 67230 38834
rect 67282 38782 67284 38834
rect 67228 38724 67284 38782
rect 67340 38724 67396 38734
rect 67228 38668 67340 38724
rect 67340 38162 67396 38668
rect 67340 38110 67342 38162
rect 67394 38110 67396 38162
rect 67340 38098 67396 38110
rect 67676 38722 67732 38734
rect 67676 38670 67678 38722
rect 67730 38670 67732 38722
rect 66892 22642 66948 22652
rect 67676 22484 67732 38670
rect 67788 37826 67844 37838
rect 67788 37774 67790 37826
rect 67842 37774 67844 37826
rect 67788 37492 67844 37774
rect 67788 37426 67844 37436
rect 68012 35028 68068 50372
rect 68684 42868 68740 75628
rect 69692 67228 69748 76526
rect 70028 75794 70084 77198
rect 70252 77250 70308 77262
rect 70252 77198 70254 77250
rect 70306 77198 70308 77250
rect 70028 75742 70030 75794
rect 70082 75742 70084 75794
rect 70028 75730 70084 75742
rect 70140 77026 70196 77038
rect 70140 76974 70142 77026
rect 70194 76974 70196 77026
rect 68684 42802 68740 42812
rect 69468 67172 69748 67228
rect 68348 41076 68404 41086
rect 68348 40626 68404 41020
rect 68348 40574 68350 40626
rect 68402 40574 68404 40626
rect 68348 40562 68404 40574
rect 69020 40964 69076 40974
rect 69244 40964 69300 40974
rect 69020 40962 69300 40964
rect 69020 40910 69022 40962
rect 69074 40910 69246 40962
rect 69298 40910 69300 40962
rect 69020 40908 69300 40910
rect 68572 40404 68628 40414
rect 69020 40404 69076 40908
rect 69244 40898 69300 40908
rect 69132 40404 69188 40414
rect 68572 40402 69188 40404
rect 68572 40350 68574 40402
rect 68626 40350 69134 40402
rect 69186 40350 69188 40402
rect 68572 40348 69188 40350
rect 68572 40292 68628 40348
rect 69132 40338 69188 40348
rect 68236 40236 68628 40292
rect 68124 38834 68180 38846
rect 68124 38782 68126 38834
rect 68178 38782 68180 38834
rect 68124 38724 68180 38782
rect 68124 38658 68180 38668
rect 68124 37156 68180 37166
rect 68236 37156 68292 40236
rect 69020 39732 69076 39742
rect 68908 39730 69076 39732
rect 68908 39678 69022 39730
rect 69074 39678 69076 39730
rect 68908 39676 69076 39678
rect 68572 39618 68628 39630
rect 68572 39566 68574 39618
rect 68626 39566 68628 39618
rect 68572 38836 68628 39566
rect 68572 38668 68628 38780
rect 68348 38612 68628 38668
rect 68348 38052 68404 38612
rect 68348 37958 68404 37996
rect 68572 37826 68628 37838
rect 68572 37774 68574 37826
rect 68626 37774 68628 37826
rect 68460 37492 68516 37502
rect 68460 37398 68516 37436
rect 68180 37100 68292 37156
rect 68124 37062 68180 37100
rect 68012 34962 68068 34972
rect 68572 26908 68628 37774
rect 68684 37266 68740 37278
rect 68684 37214 68686 37266
rect 68738 37214 68740 37266
rect 68684 37156 68740 37214
rect 68684 37090 68740 37100
rect 68796 36596 68852 36606
rect 68796 36502 68852 36540
rect 68908 32228 68964 39676
rect 69020 39666 69076 39676
rect 69468 39732 69524 67172
rect 69916 58884 69972 58894
rect 69580 41412 69636 41422
rect 69580 41074 69636 41356
rect 69580 41022 69582 41074
rect 69634 41022 69636 41074
rect 69580 41010 69636 41022
rect 69580 40628 69636 40638
rect 69580 40534 69636 40572
rect 69804 40628 69860 40638
rect 69244 39508 69300 39518
rect 69468 39508 69524 39676
rect 69580 39620 69636 39630
rect 69580 39526 69636 39564
rect 69244 39506 69524 39508
rect 69244 39454 69246 39506
rect 69298 39454 69524 39506
rect 69244 39452 69524 39454
rect 69244 39442 69300 39452
rect 69356 38892 69636 38948
rect 69020 38836 69076 38846
rect 69020 38742 69076 38780
rect 69356 38724 69412 38892
rect 69580 38834 69636 38892
rect 69580 38782 69582 38834
rect 69634 38782 69636 38834
rect 69580 38770 69636 38782
rect 68908 32162 68964 32172
rect 69020 38612 69076 38622
rect 69020 30772 69076 38556
rect 69244 38500 69300 38510
rect 69244 37938 69300 38444
rect 69356 38050 69412 38668
rect 69468 38722 69524 38734
rect 69468 38670 69470 38722
rect 69522 38670 69524 38722
rect 69468 38668 69524 38670
rect 69804 38668 69860 40572
rect 69468 38612 69636 38668
rect 69356 37998 69358 38050
rect 69410 37998 69412 38050
rect 69356 37986 69412 37998
rect 69468 38388 69524 38398
rect 69244 37886 69246 37938
rect 69298 37886 69300 37938
rect 69132 37266 69188 37278
rect 69132 37214 69134 37266
rect 69186 37214 69188 37266
rect 69132 36596 69188 37214
rect 69132 36530 69188 36540
rect 69244 36484 69300 37886
rect 69468 37490 69524 38332
rect 69468 37438 69470 37490
rect 69522 37438 69524 37490
rect 69468 37426 69524 37438
rect 69244 36418 69300 36428
rect 69132 30772 69188 30782
rect 69020 30716 69132 30772
rect 69132 30706 69188 30716
rect 69580 29428 69636 38612
rect 69692 38612 69860 38668
rect 69916 38946 69972 58828
rect 70028 40962 70084 40974
rect 70028 40910 70030 40962
rect 70082 40910 70084 40962
rect 70028 40628 70084 40910
rect 70028 40562 70084 40572
rect 69916 38894 69918 38946
rect 69970 38894 69972 38946
rect 69692 36932 69748 38612
rect 69916 38162 69972 38894
rect 70140 38500 70196 76974
rect 70252 76690 70308 77198
rect 70252 76638 70254 76690
rect 70306 76638 70308 76690
rect 70252 76626 70308 76638
rect 70364 76580 70420 79200
rect 71036 77138 71092 79200
rect 71036 77086 71038 77138
rect 71090 77086 71092 77138
rect 71036 77074 71092 77086
rect 71708 77140 71764 79200
rect 71708 77074 71764 77084
rect 72268 77138 72324 77150
rect 72268 77086 72270 77138
rect 72322 77086 72324 77138
rect 70924 77028 70980 77038
rect 70364 76514 70420 76524
rect 70588 76578 70644 76590
rect 70924 76580 70980 76972
rect 72268 76692 72324 77086
rect 72044 76690 72324 76692
rect 72044 76638 72270 76690
rect 72322 76638 72324 76690
rect 72044 76636 72324 76638
rect 70588 76526 70590 76578
rect 70642 76526 70644 76578
rect 70476 74116 70532 74126
rect 70476 43540 70532 74060
rect 70588 67284 70644 76526
rect 70700 76578 70980 76580
rect 70700 76526 70926 76578
rect 70978 76526 70980 76578
rect 70700 76524 70980 76526
rect 70700 75794 70756 76524
rect 70924 76514 70980 76524
rect 71260 76578 71316 76590
rect 71596 76580 71652 76590
rect 71932 76580 71988 76590
rect 71260 76526 71262 76578
rect 71314 76526 71316 76578
rect 70700 75742 70702 75794
rect 70754 75742 70756 75794
rect 70700 75730 70756 75742
rect 71260 67508 71316 76526
rect 71372 76524 71596 76580
rect 71372 75794 71428 76524
rect 71596 76486 71652 76524
rect 71820 76578 71988 76580
rect 71820 76526 71934 76578
rect 71986 76526 71988 76578
rect 71820 76524 71988 76526
rect 71372 75742 71374 75794
rect 71426 75742 71428 75794
rect 71372 75730 71428 75742
rect 70588 67218 70644 67228
rect 70812 67452 71316 67508
rect 70812 50428 70868 67452
rect 71148 67284 71204 67294
rect 71148 62188 71204 67228
rect 71148 62132 71316 62188
rect 70476 43474 70532 43484
rect 70700 50372 70868 50428
rect 70588 41858 70644 41870
rect 70588 41806 70590 41858
rect 70642 41806 70644 41858
rect 70588 41748 70644 41806
rect 70588 41682 70644 41692
rect 70364 41188 70420 41198
rect 70364 40962 70420 41132
rect 70364 40910 70366 40962
rect 70418 40910 70420 40962
rect 70252 40628 70308 40638
rect 70364 40628 70420 40910
rect 70308 40572 70420 40628
rect 70252 40534 70308 40572
rect 70700 40516 70756 50372
rect 71148 45332 71204 45342
rect 70812 41860 70868 41870
rect 71036 41860 71092 41870
rect 70812 41298 70868 41804
rect 70812 41246 70814 41298
rect 70866 41246 70868 41298
rect 70812 41234 70868 41246
rect 70924 41858 71092 41860
rect 70924 41806 71038 41858
rect 71090 41806 71092 41858
rect 70924 41804 71092 41806
rect 70924 41300 70980 41804
rect 71036 41794 71092 41804
rect 70812 40852 70868 40862
rect 70924 40852 70980 41244
rect 70868 40796 70980 40852
rect 70812 40786 70868 40796
rect 70588 40460 70756 40516
rect 70140 38434 70196 38444
rect 70252 39620 70308 39630
rect 70252 38836 70308 39564
rect 70476 39394 70532 39406
rect 70476 39342 70478 39394
rect 70530 39342 70532 39394
rect 70364 38836 70420 38846
rect 70252 38834 70420 38836
rect 70252 38782 70366 38834
rect 70418 38782 70420 38834
rect 70252 38780 70420 38782
rect 69916 38110 69918 38162
rect 69970 38110 69972 38162
rect 69916 38098 69972 38110
rect 70252 38052 70308 38780
rect 70364 38770 70420 38780
rect 70476 38836 70532 39342
rect 70588 39396 70644 40460
rect 70812 40404 70868 40414
rect 70700 40348 70812 40404
rect 70700 40290 70756 40348
rect 70812 40338 70868 40348
rect 70700 40238 70702 40290
rect 70754 40238 70756 40290
rect 70700 40226 70756 40238
rect 71148 39732 71204 45276
rect 70812 39676 71204 39732
rect 70700 39620 70756 39630
rect 70700 39526 70756 39564
rect 70588 39340 70756 39396
rect 70476 38770 70532 38780
rect 70700 38836 70756 39340
rect 70700 38770 70756 38780
rect 70588 38722 70644 38734
rect 70588 38670 70590 38722
rect 70642 38670 70644 38722
rect 70588 38668 70644 38670
rect 70812 38668 70868 39676
rect 70924 39508 70980 39518
rect 70924 39414 70980 39452
rect 70028 38050 70308 38052
rect 70028 37998 70254 38050
rect 70306 37998 70308 38050
rect 70028 37996 70308 37998
rect 70028 37940 70084 37996
rect 70252 37986 70308 37996
rect 70476 38612 70644 38668
rect 70700 38612 70868 38668
rect 70924 38834 70980 38846
rect 70924 38782 70926 38834
rect 70978 38782 70980 38834
rect 70924 38724 70980 38782
rect 69804 37884 70084 37940
rect 69804 37490 69860 37884
rect 70364 37826 70420 37838
rect 70364 37774 70366 37826
rect 70418 37774 70420 37826
rect 70140 37604 70196 37614
rect 69804 37438 69806 37490
rect 69858 37438 69860 37490
rect 69804 37426 69860 37438
rect 70028 37492 70084 37502
rect 70028 37266 70084 37436
rect 70028 37214 70030 37266
rect 70082 37214 70084 37266
rect 70028 37202 70084 37214
rect 69692 36876 69860 36932
rect 69692 36484 69748 36494
rect 69692 36390 69748 36428
rect 69804 35308 69860 36876
rect 69580 29362 69636 29372
rect 69692 35252 69860 35308
rect 68796 28308 68852 28318
rect 68572 26852 68740 26908
rect 68684 23156 68740 26852
rect 68796 26068 68852 28252
rect 69692 26852 69748 35252
rect 70140 27860 70196 37548
rect 70364 29764 70420 37774
rect 70476 37604 70532 38612
rect 70588 38500 70644 38510
rect 70588 38050 70644 38444
rect 70588 37998 70590 38050
rect 70642 37998 70644 38050
rect 70588 37986 70644 37998
rect 70476 37538 70532 37548
rect 70588 37492 70644 37502
rect 70588 37266 70644 37436
rect 70588 37214 70590 37266
rect 70642 37214 70644 37266
rect 70588 37202 70644 37214
rect 70700 32788 70756 38612
rect 70812 38052 70868 38062
rect 70924 38052 70980 38668
rect 71260 38500 71316 62132
rect 71820 50428 71876 76524
rect 71932 76514 71988 76524
rect 71932 75796 71988 75806
rect 72044 75796 72100 76636
rect 72268 76626 72324 76636
rect 71932 75794 72100 75796
rect 71932 75742 71934 75794
rect 71986 75742 72100 75794
rect 71932 75740 72100 75742
rect 72380 75794 72436 79200
rect 73052 77028 73108 79200
rect 73052 76962 73108 76972
rect 73164 77140 73220 77150
rect 72604 76580 72660 76590
rect 72940 76580 72996 76590
rect 72604 76578 72772 76580
rect 72604 76526 72606 76578
rect 72658 76526 72772 76578
rect 72604 76524 72772 76526
rect 72604 76514 72660 76524
rect 72380 75742 72382 75794
rect 72434 75742 72436 75794
rect 71932 75730 71988 75740
rect 72380 75684 72436 75742
rect 72604 75684 72660 75694
rect 72380 75682 72660 75684
rect 72380 75630 72606 75682
rect 72658 75630 72660 75682
rect 72380 75628 72660 75630
rect 72604 75618 72660 75628
rect 72156 68740 72212 68750
rect 71596 50372 71876 50428
rect 72044 51492 72100 51502
rect 71372 41748 71428 41758
rect 71372 41410 71428 41692
rect 71372 41358 71374 41410
rect 71426 41358 71428 41410
rect 71372 41346 71428 41358
rect 71484 41298 71540 41310
rect 71484 41246 71486 41298
rect 71538 41246 71540 41298
rect 71484 41188 71540 41246
rect 71484 41122 71540 41132
rect 71372 39732 71428 39742
rect 71372 39638 71428 39676
rect 71596 39732 71652 50372
rect 71932 46228 71988 46238
rect 71820 46172 71932 46228
rect 71708 41186 71764 41198
rect 71708 41134 71710 41186
rect 71762 41134 71764 41186
rect 71708 40404 71764 41134
rect 71820 41076 71876 46172
rect 71932 46162 71988 46172
rect 72044 41524 72100 51436
rect 72156 42980 72212 68684
rect 72716 62132 72772 76524
rect 72828 76578 72996 76580
rect 72828 76526 72942 76578
rect 72994 76526 72996 76578
rect 72828 76524 72996 76526
rect 72828 67396 72884 76524
rect 72940 76514 72996 76524
rect 73164 76468 73220 77084
rect 73724 77140 73780 79200
rect 73724 77074 73780 77084
rect 74284 77028 74340 77038
rect 74060 76580 74116 76590
rect 74060 76486 74116 76524
rect 74284 76468 74340 76972
rect 74396 77026 74452 79200
rect 75068 77364 75124 79200
rect 75068 77308 75236 77364
rect 74396 76974 74398 77026
rect 74450 76974 74452 77026
rect 74396 76962 74452 76974
rect 74508 77140 74564 77150
rect 73164 76466 73444 76468
rect 73164 76414 73166 76466
rect 73218 76414 73444 76466
rect 73164 76412 73444 76414
rect 73164 76402 73220 76412
rect 73388 75794 73444 76412
rect 74172 76466 74340 76468
rect 74172 76414 74286 76466
rect 74338 76414 74340 76466
rect 74172 76412 74340 76414
rect 74172 76356 74228 76412
rect 74284 76402 74340 76412
rect 73388 75742 73390 75794
rect 73442 75742 73444 75794
rect 73388 75730 73444 75742
rect 73948 76300 74228 76356
rect 73948 75794 74004 76300
rect 73948 75742 73950 75794
rect 74002 75742 74004 75794
rect 73948 75730 74004 75742
rect 74508 75794 74564 77084
rect 75068 77140 75124 77150
rect 74956 77026 75012 77038
rect 74956 76974 74958 77026
rect 75010 76974 75012 77026
rect 74508 75742 74510 75794
rect 74562 75742 74564 75794
rect 74508 75730 74564 75742
rect 74620 76692 74676 76702
rect 72940 75460 72996 75470
rect 74060 75460 74116 75470
rect 72940 75458 73332 75460
rect 72940 75406 72942 75458
rect 72994 75406 73332 75458
rect 72940 75404 73332 75406
rect 72940 75394 72996 75404
rect 72828 67340 72996 67396
rect 72716 62066 72772 62076
rect 72940 50428 72996 67340
rect 73276 67228 73332 75404
rect 74060 75122 74116 75404
rect 74060 75070 74062 75122
rect 74114 75070 74116 75122
rect 74060 75058 74116 75070
rect 74508 75124 74564 75134
rect 74620 75124 74676 76636
rect 74508 75122 74676 75124
rect 74508 75070 74510 75122
rect 74562 75070 74676 75122
rect 74508 75068 74676 75070
rect 74732 76578 74788 76590
rect 74732 76526 74734 76578
rect 74786 76526 74788 76578
rect 74508 75058 74564 75068
rect 74732 73948 74788 76526
rect 74956 75796 75012 76974
rect 75068 76578 75124 77084
rect 75180 77138 75236 77308
rect 75740 77252 75796 79200
rect 76412 77476 76468 79200
rect 76412 77420 76916 77476
rect 75740 77196 76244 77252
rect 75180 77086 75182 77138
rect 75234 77086 75236 77138
rect 75180 77074 75236 77086
rect 75628 77138 75684 77150
rect 75628 77086 75630 77138
rect 75682 77086 75684 77138
rect 75404 76580 75460 76590
rect 75068 76526 75070 76578
rect 75122 76526 75124 76578
rect 75068 76514 75124 76526
rect 75180 76578 75460 76580
rect 75180 76526 75406 76578
rect 75458 76526 75460 76578
rect 75180 76524 75460 76526
rect 75068 75796 75124 75806
rect 74956 75794 75124 75796
rect 74956 75742 75070 75794
rect 75122 75742 75124 75794
rect 74956 75740 75124 75742
rect 75068 75730 75124 75740
rect 74956 75124 75012 75134
rect 74956 75030 75012 75068
rect 74620 73892 74788 73948
rect 73948 68852 74004 68862
rect 73276 67172 73668 67228
rect 72604 50372 72996 50428
rect 73052 62132 73108 62142
rect 72156 42914 72212 42924
rect 72268 44660 72324 44670
rect 72044 41458 72100 41468
rect 71932 41300 71988 41310
rect 71932 41206 71988 41244
rect 72044 41300 72100 41310
rect 72044 41298 72212 41300
rect 72044 41246 72046 41298
rect 72098 41246 72212 41298
rect 72044 41244 72212 41246
rect 72044 41234 72100 41244
rect 72156 41188 72212 41244
rect 72156 41122 72212 41132
rect 71820 41020 71988 41076
rect 71708 40338 71764 40348
rect 71820 39732 71876 39742
rect 71596 39730 71876 39732
rect 71596 39678 71822 39730
rect 71874 39678 71876 39730
rect 71596 39676 71876 39678
rect 71596 39620 71652 39676
rect 71820 39666 71876 39676
rect 71596 39554 71652 39564
rect 71372 39508 71428 39518
rect 71372 38946 71428 39452
rect 71932 39396 71988 41020
rect 71372 38894 71374 38946
rect 71426 38894 71428 38946
rect 71372 38724 71428 38894
rect 71372 38658 71428 38668
rect 71484 39340 71988 39396
rect 72044 40964 72100 40974
rect 71260 38434 71316 38444
rect 71148 38052 71204 38062
rect 70812 38050 71204 38052
rect 70812 37998 70814 38050
rect 70866 37998 71150 38050
rect 71202 37998 71204 38050
rect 70812 37996 71204 37998
rect 70812 37986 70868 37996
rect 71148 37986 71204 37996
rect 71372 38052 71428 38062
rect 71372 37958 71428 37996
rect 71484 37716 71540 39340
rect 71596 39060 71652 39070
rect 71596 38834 71652 39004
rect 71596 38782 71598 38834
rect 71650 38782 71652 38834
rect 71596 38770 71652 38782
rect 72044 38668 72100 40908
rect 71932 38612 72100 38668
rect 72156 38836 72212 38846
rect 71708 37938 71764 37950
rect 71708 37886 71710 37938
rect 71762 37886 71764 37938
rect 71372 37660 71540 37716
rect 71596 37826 71652 37838
rect 71596 37774 71598 37826
rect 71650 37774 71652 37826
rect 70812 37604 70868 37614
rect 70812 37490 70868 37548
rect 70812 37438 70814 37490
rect 70866 37438 70868 37490
rect 70812 37426 70868 37438
rect 71148 37492 71204 37502
rect 71148 37398 71204 37436
rect 71260 36596 71316 36606
rect 71260 36502 71316 36540
rect 71372 36148 71428 37660
rect 71484 37492 71540 37502
rect 71484 37398 71540 37436
rect 71372 36092 71540 36148
rect 71372 35924 71428 35934
rect 71372 35830 71428 35868
rect 71372 34916 71428 34926
rect 71148 34244 71204 34254
rect 71148 34150 71204 34188
rect 71260 34132 71316 34142
rect 70924 34020 70980 34030
rect 70924 33926 70980 33964
rect 71260 34018 71316 34076
rect 71260 33966 71262 34018
rect 71314 33966 71316 34018
rect 71260 33954 71316 33966
rect 71372 33796 71428 34860
rect 71148 33740 71428 33796
rect 71484 34242 71540 36092
rect 71596 34356 71652 37774
rect 71708 37604 71764 37886
rect 71708 37538 71764 37548
rect 71708 37268 71764 37278
rect 71708 36594 71764 37212
rect 71708 36542 71710 36594
rect 71762 36542 71764 36594
rect 71708 36530 71764 36542
rect 71708 35588 71764 35598
rect 71708 35494 71764 35532
rect 71820 34692 71876 34702
rect 71820 34598 71876 34636
rect 71596 34300 71876 34356
rect 71484 34190 71486 34242
rect 71538 34190 71540 34242
rect 71148 33458 71204 33740
rect 71484 33570 71540 34190
rect 71484 33518 71486 33570
rect 71538 33518 71540 33570
rect 71484 33506 71540 33518
rect 71708 34132 71764 34142
rect 71148 33406 71150 33458
rect 71202 33406 71204 33458
rect 71148 33394 71204 33406
rect 71596 33124 71652 33134
rect 71596 33030 71652 33068
rect 71708 33012 71764 34076
rect 70924 32788 70980 32798
rect 70700 32786 71428 32788
rect 70700 32734 70926 32786
rect 70978 32734 71428 32786
rect 70700 32732 71428 32734
rect 70924 32722 70980 32732
rect 71036 32564 71092 32574
rect 70924 32562 71092 32564
rect 70924 32510 71038 32562
rect 71090 32510 71092 32562
rect 70924 32508 71092 32510
rect 70924 31892 70980 32508
rect 71036 32498 71092 32508
rect 71372 32562 71428 32732
rect 71708 32674 71764 32956
rect 71820 32900 71876 34300
rect 71820 32834 71876 32844
rect 71708 32622 71710 32674
rect 71762 32622 71764 32674
rect 71708 32610 71764 32622
rect 71372 32510 71374 32562
rect 71426 32510 71428 32562
rect 71372 32498 71428 32510
rect 71148 32452 71204 32462
rect 71148 32340 71204 32396
rect 70924 31778 70980 31836
rect 70924 31726 70926 31778
rect 70978 31726 70980 31778
rect 70924 31714 70980 31726
rect 71036 32284 71204 32340
rect 71260 32450 71316 32462
rect 71260 32398 71262 32450
rect 71314 32398 71316 32450
rect 70924 31108 70980 31118
rect 70924 31014 70980 31052
rect 70364 29708 70644 29764
rect 70252 27860 70308 27870
rect 70140 27858 70308 27860
rect 70140 27806 70254 27858
rect 70306 27806 70308 27858
rect 70140 27804 70308 27806
rect 70252 27794 70308 27804
rect 70588 27074 70644 29708
rect 71036 29428 71092 32284
rect 71260 31892 71316 32398
rect 71708 31892 71764 31902
rect 71260 31836 71428 31892
rect 71260 31666 71316 31678
rect 71260 31614 71262 31666
rect 71314 31614 71316 31666
rect 71148 31554 71204 31566
rect 71148 31502 71150 31554
rect 71202 31502 71204 31554
rect 71148 29652 71204 31502
rect 71260 30770 71316 31614
rect 71372 31108 71428 31836
rect 71708 31780 71764 31836
rect 71596 31778 71764 31780
rect 71596 31726 71710 31778
rect 71762 31726 71764 31778
rect 71596 31724 71764 31726
rect 71484 31666 71540 31678
rect 71484 31614 71486 31666
rect 71538 31614 71540 31666
rect 71484 31556 71540 31614
rect 71484 31490 71540 31500
rect 71372 31052 71540 31108
rect 71372 30884 71428 30894
rect 71372 30790 71428 30828
rect 71260 30718 71262 30770
rect 71314 30718 71316 30770
rect 71260 30706 71316 30718
rect 71484 29764 71540 31052
rect 71596 30098 71652 31724
rect 71708 31714 71764 31724
rect 71820 31220 71876 31230
rect 71932 31220 71988 38612
rect 72156 38162 72212 38780
rect 72156 38110 72158 38162
rect 72210 38110 72212 38162
rect 72156 38098 72212 38110
rect 72268 37828 72324 44604
rect 72156 37772 72324 37828
rect 72380 39394 72436 39406
rect 72380 39342 72382 39394
rect 72434 39342 72436 39394
rect 72380 38948 72436 39342
rect 72492 38948 72548 38958
rect 72380 38946 72548 38948
rect 72380 38894 72494 38946
rect 72546 38894 72548 38946
rect 72380 38892 72548 38894
rect 72380 37828 72436 38892
rect 72492 38882 72548 38892
rect 72604 38668 72660 50372
rect 72940 40180 72996 40190
rect 72940 40086 72996 40124
rect 72940 39732 72996 39742
rect 72156 37156 72212 37772
rect 72380 37762 72436 37772
rect 72492 38612 72660 38668
rect 72828 39618 72884 39630
rect 72828 39566 72830 39618
rect 72882 39566 72884 39618
rect 72828 39058 72884 39566
rect 72940 39618 72996 39676
rect 72940 39566 72942 39618
rect 72994 39566 72996 39618
rect 72940 39554 72996 39566
rect 72828 39006 72830 39058
rect 72882 39006 72884 39058
rect 72828 38668 72884 39006
rect 72828 38612 72996 38668
rect 72268 37604 72324 37614
rect 72268 37378 72324 37548
rect 72268 37326 72270 37378
rect 72322 37326 72324 37378
rect 72268 37314 72324 37326
rect 72492 37268 72548 38612
rect 72604 38500 72660 38510
rect 72604 38162 72660 38444
rect 72604 38110 72606 38162
rect 72658 38110 72660 38162
rect 72604 38098 72660 38110
rect 72716 38274 72772 38286
rect 72716 38222 72718 38274
rect 72770 38222 72772 38274
rect 72492 37266 72660 37268
rect 72492 37214 72494 37266
rect 72546 37214 72660 37266
rect 72492 37212 72660 37214
rect 72492 37202 72548 37212
rect 72156 37100 72324 37156
rect 72156 36484 72212 36494
rect 72156 36390 72212 36428
rect 72268 35924 72324 37100
rect 72156 35868 72324 35924
rect 72380 37154 72436 37166
rect 72380 37102 72382 37154
rect 72434 37102 72436 37154
rect 72156 35700 72212 35868
rect 72156 35634 72212 35644
rect 72268 35698 72324 35710
rect 72268 35646 72270 35698
rect 72322 35646 72324 35698
rect 72268 35588 72324 35646
rect 72268 35476 72324 35532
rect 72156 35420 72324 35476
rect 72156 34692 72212 35420
rect 72044 34690 72212 34692
rect 72044 34638 72158 34690
rect 72210 34638 72212 34690
rect 72044 34636 72212 34638
rect 72044 33908 72100 34636
rect 72156 34626 72212 34636
rect 72156 34244 72212 34254
rect 72380 34244 72436 37102
rect 72492 36932 72548 36942
rect 72492 35028 72548 36876
rect 72604 36594 72660 37212
rect 72604 36542 72606 36594
rect 72658 36542 72660 36594
rect 72604 36530 72660 36542
rect 72716 36036 72772 38222
rect 72940 37828 72996 38612
rect 73052 38052 73108 62076
rect 73612 50428 73668 67172
rect 73276 50372 73668 50428
rect 73164 41076 73220 41086
rect 73164 40982 73220 41020
rect 73164 40402 73220 40414
rect 73164 40350 73166 40402
rect 73218 40350 73220 40402
rect 73164 39730 73220 40350
rect 73276 40068 73332 50372
rect 73948 41972 74004 68796
rect 74620 68068 74676 73892
rect 74284 68012 74676 68068
rect 74844 72324 74900 72334
rect 74284 67228 74340 68012
rect 74284 67172 74452 67228
rect 73500 41970 74004 41972
rect 73500 41918 73950 41970
rect 74002 41918 74004 41970
rect 73500 41916 74004 41918
rect 73500 41186 73556 41916
rect 73948 41906 74004 41916
rect 74060 45220 74116 45230
rect 74060 41412 74116 45164
rect 73500 41134 73502 41186
rect 73554 41134 73556 41186
rect 73500 41122 73556 41134
rect 73948 41356 74116 41412
rect 73724 41074 73780 41086
rect 73724 41022 73726 41074
rect 73778 41022 73780 41074
rect 73388 40962 73444 40974
rect 73388 40910 73390 40962
rect 73442 40910 73444 40962
rect 73388 40628 73444 40910
rect 73724 40628 73780 41022
rect 73388 40572 73668 40628
rect 73612 40402 73668 40572
rect 73724 40562 73780 40572
rect 73612 40350 73614 40402
rect 73666 40350 73668 40402
rect 73612 40338 73668 40350
rect 73388 40292 73444 40302
rect 73388 40198 73444 40236
rect 73276 40012 73444 40068
rect 73164 39678 73166 39730
rect 73218 39678 73220 39730
rect 73164 39666 73220 39678
rect 73276 39508 73332 39518
rect 73052 37958 73108 37996
rect 73164 38946 73220 38958
rect 73164 38894 73166 38946
rect 73218 38894 73220 38946
rect 73164 37828 73220 38894
rect 73276 38274 73332 39452
rect 73276 38222 73278 38274
rect 73330 38222 73332 38274
rect 73276 38210 73332 38222
rect 72940 37772 73108 37828
rect 73164 37772 73332 37828
rect 73052 37716 73108 37772
rect 73052 37660 73220 37716
rect 72828 37604 72884 37614
rect 72884 37548 73108 37604
rect 72828 37538 72884 37548
rect 72828 37380 72884 37390
rect 72828 37286 72884 37324
rect 72828 36484 72884 36494
rect 72940 36484 72996 37548
rect 73052 37266 73108 37548
rect 73052 37214 73054 37266
rect 73106 37214 73108 37266
rect 73052 37202 73108 37214
rect 73164 36932 73220 37660
rect 73276 37380 73332 37772
rect 73276 37314 73332 37324
rect 73388 37268 73444 40012
rect 73500 39620 73556 39630
rect 73500 39060 73556 39564
rect 73836 39508 73892 39518
rect 73836 39414 73892 39452
rect 73500 38946 73556 39004
rect 73500 38894 73502 38946
rect 73554 38894 73556 38946
rect 73500 38724 73556 38894
rect 73500 38658 73556 38668
rect 73836 37938 73892 37950
rect 73836 37886 73838 37938
rect 73890 37886 73892 37938
rect 73500 37828 73556 37838
rect 73836 37828 73892 37886
rect 73556 37772 73892 37828
rect 73500 37734 73556 37772
rect 73948 37604 74004 41356
rect 74172 41300 74228 41310
rect 74060 41244 74172 41300
rect 74060 41186 74116 41244
rect 74060 41134 74062 41186
rect 74114 41134 74116 41186
rect 74060 41122 74116 41134
rect 74172 39506 74228 41244
rect 74284 41188 74340 41198
rect 74284 41094 74340 41132
rect 74284 40402 74340 40414
rect 74284 40350 74286 40402
rect 74338 40350 74340 40402
rect 74284 39620 74340 40350
rect 74284 39554 74340 39564
rect 74172 39454 74174 39506
rect 74226 39454 74228 39506
rect 74060 39396 74116 39406
rect 74060 37828 74116 39340
rect 74172 39060 74228 39454
rect 74396 39396 74452 67172
rect 74844 55468 74900 72268
rect 75180 68740 75236 76524
rect 75404 76514 75460 76524
rect 75628 76356 75684 77086
rect 75740 77026 75796 77038
rect 75740 76974 75742 77026
rect 75794 76974 75796 77026
rect 75740 76578 75796 76974
rect 76076 76804 76132 76814
rect 76076 76690 76132 76748
rect 76076 76638 76078 76690
rect 76130 76638 76132 76690
rect 76076 76626 76132 76638
rect 75740 76526 75742 76578
rect 75794 76526 75796 76578
rect 75740 76514 75796 76526
rect 75628 76300 75796 76356
rect 75404 75682 75460 75694
rect 75404 75630 75406 75682
rect 75458 75630 75460 75682
rect 75404 75572 75460 75630
rect 75404 75506 75460 75516
rect 75628 75684 75684 75694
rect 75628 75570 75684 75628
rect 75628 75518 75630 75570
rect 75682 75518 75684 75570
rect 75628 75506 75684 75518
rect 75404 75012 75460 75022
rect 75404 74918 75460 74956
rect 75628 75010 75684 75022
rect 75628 74958 75630 75010
rect 75682 74958 75684 75010
rect 75292 74116 75348 74126
rect 75292 74022 75348 74060
rect 75628 68852 75684 74958
rect 75740 74226 75796 76300
rect 76188 75682 76244 77196
rect 76412 77138 76468 77150
rect 76412 77086 76414 77138
rect 76466 77086 76468 77138
rect 76412 76578 76468 77086
rect 76412 76526 76414 76578
rect 76466 76526 76468 76578
rect 76412 76514 76468 76526
rect 76188 75630 76190 75682
rect 76242 75630 76244 75682
rect 76076 75572 76132 75582
rect 75964 75012 76020 75022
rect 75964 74918 76020 74956
rect 76076 74338 76132 75516
rect 76188 75124 76244 75630
rect 76188 75058 76244 75068
rect 76300 76468 76356 76478
rect 76076 74286 76078 74338
rect 76130 74286 76132 74338
rect 76076 74274 76132 74286
rect 75740 74174 75742 74226
rect 75794 74174 75796 74226
rect 75740 74162 75796 74174
rect 76188 73556 76244 73566
rect 76300 73556 76356 76412
rect 76748 76356 76804 76366
rect 76748 76262 76804 76300
rect 76524 75684 76580 75694
rect 76860 75684 76916 77420
rect 76524 75570 76580 75628
rect 76524 75518 76526 75570
rect 76578 75518 76580 75570
rect 76524 75506 76580 75518
rect 76636 75682 76916 75684
rect 76636 75630 76862 75682
rect 76914 75630 76916 75682
rect 76636 75628 76916 75630
rect 76412 74788 76468 74798
rect 76412 74786 76580 74788
rect 76412 74734 76414 74786
rect 76466 74734 76580 74786
rect 76412 74732 76580 74734
rect 76412 74722 76468 74732
rect 76412 74338 76468 74350
rect 76412 74286 76414 74338
rect 76466 74286 76468 74338
rect 76412 74226 76468 74286
rect 76412 74174 76414 74226
rect 76466 74174 76468 74226
rect 76412 74162 76468 74174
rect 76188 73554 76356 73556
rect 76188 73502 76190 73554
rect 76242 73502 76356 73554
rect 76188 73500 76356 73502
rect 76188 73490 76244 73500
rect 76524 72660 76580 74732
rect 76636 73554 76692 75628
rect 76860 75618 76916 75628
rect 76972 76804 77028 76814
rect 76860 75124 76916 75134
rect 76972 75124 77028 76748
rect 77084 76468 77140 79200
rect 77308 79156 77364 79166
rect 77084 76402 77140 76412
rect 77196 76916 77252 76926
rect 77196 75570 77252 76860
rect 77308 76692 77364 79100
rect 77308 76598 77364 76636
rect 77756 76020 77812 79200
rect 78428 77476 78484 79200
rect 78764 78036 78820 78046
rect 78428 77420 78708 77476
rect 78204 76578 78260 76590
rect 78204 76526 78206 76578
rect 78258 76526 78260 76578
rect 77868 76468 77924 76478
rect 77868 76374 77924 76412
rect 78204 76132 78260 76526
rect 78204 76066 78260 76076
rect 77196 75518 77198 75570
rect 77250 75518 77252 75570
rect 77196 75506 77252 75518
rect 77308 75964 77812 76020
rect 76860 75122 77252 75124
rect 76860 75070 76862 75122
rect 76914 75070 77252 75122
rect 76860 75068 77252 75070
rect 76860 75058 76916 75068
rect 76636 73502 76638 73554
rect 76690 73502 76692 73554
rect 76636 73490 76692 73502
rect 76972 74114 77028 74126
rect 76972 74062 76974 74114
rect 77026 74062 77028 74114
rect 76524 72604 76916 72660
rect 75628 68786 75684 68796
rect 76748 72436 76804 72446
rect 75180 68674 75236 68684
rect 74508 55412 74900 55468
rect 74508 39732 74564 55412
rect 76748 43708 76804 72380
rect 76860 67228 76916 72604
rect 76972 72324 77028 74062
rect 77196 73554 77252 75068
rect 77196 73502 77198 73554
rect 77250 73502 77252 73554
rect 77196 73490 77252 73502
rect 77308 74898 77364 75964
rect 77756 75796 77812 75806
rect 77756 75794 78036 75796
rect 77756 75742 77758 75794
rect 77810 75742 78036 75794
rect 77756 75740 78036 75742
rect 77756 75730 77812 75740
rect 77308 74846 77310 74898
rect 77362 74846 77364 74898
rect 77308 73332 77364 74846
rect 77532 75124 77588 75134
rect 77532 74114 77588 75068
rect 77532 74062 77534 74114
rect 77586 74062 77588 74114
rect 77532 74050 77588 74062
rect 77756 74786 77812 74798
rect 77756 74734 77758 74786
rect 77810 74734 77812 74786
rect 77644 73556 77700 73566
rect 77644 73462 77700 73500
rect 77196 73276 77364 73332
rect 77196 72658 77252 73276
rect 77196 72606 77198 72658
rect 77250 72606 77252 72658
rect 77196 72594 77252 72606
rect 77644 72436 77700 72446
rect 77644 72342 77700 72380
rect 76972 72258 77028 72268
rect 77644 71650 77700 71662
rect 77644 71598 77646 71650
rect 77698 71598 77700 71650
rect 77644 71316 77700 71598
rect 77644 71250 77700 71260
rect 77644 70980 77700 70990
rect 77644 70886 77700 70924
rect 77420 70756 77476 70766
rect 77420 70662 77476 70700
rect 77644 69186 77700 69198
rect 77644 69134 77646 69186
rect 77698 69134 77700 69186
rect 77644 69076 77700 69134
rect 77644 69010 77700 69020
rect 77420 68628 77476 68638
rect 77420 68534 77476 68572
rect 77644 68516 77700 68526
rect 77644 68422 77700 68460
rect 76860 67172 77028 67228
rect 75404 43652 75460 43662
rect 76748 43652 76916 43708
rect 75292 42980 75348 42990
rect 75292 42868 75348 42924
rect 75068 42866 75348 42868
rect 75068 42814 75294 42866
rect 75346 42814 75348 42866
rect 75068 42812 75348 42814
rect 74956 41972 75012 41982
rect 74844 41970 75012 41972
rect 74844 41918 74958 41970
rect 75010 41918 75012 41970
rect 74844 41916 75012 41918
rect 74732 41860 74788 41870
rect 74732 41766 74788 41804
rect 74844 41524 74900 41916
rect 74956 41906 75012 41916
rect 74620 41468 74900 41524
rect 74620 41410 74676 41468
rect 75068 41412 75124 42812
rect 75292 42802 75348 42812
rect 75404 42644 75460 43596
rect 75180 42588 75460 42644
rect 76300 43540 76356 43550
rect 75180 41860 75236 42588
rect 75292 42082 75348 42094
rect 75292 42030 75294 42082
rect 75346 42030 75348 42082
rect 75292 41972 75348 42030
rect 75740 42084 75796 42094
rect 75628 41972 75684 41982
rect 75292 41970 75684 41972
rect 75292 41918 75630 41970
rect 75682 41918 75684 41970
rect 75292 41916 75684 41918
rect 75628 41906 75684 41916
rect 75180 41804 75348 41860
rect 74620 41358 74622 41410
rect 74674 41358 74676 41410
rect 74620 41346 74676 41358
rect 74844 41356 75124 41412
rect 74620 40628 74676 40638
rect 74620 40534 74676 40572
rect 74620 39732 74676 39742
rect 74564 39730 74676 39732
rect 74564 39678 74622 39730
rect 74674 39678 74676 39730
rect 74564 39676 74676 39678
rect 74508 39638 74564 39676
rect 74620 39666 74676 39676
rect 74396 39330 74452 39340
rect 74172 38994 74228 39004
rect 74508 38946 74564 38958
rect 74508 38894 74510 38946
rect 74562 38894 74564 38946
rect 74172 38834 74228 38846
rect 74172 38782 74174 38834
rect 74226 38782 74228 38834
rect 74172 38724 74228 38782
rect 74172 38658 74228 38668
rect 74508 38612 74564 38894
rect 74732 38836 74788 38846
rect 74508 38546 74564 38556
rect 74620 38834 74788 38836
rect 74620 38782 74734 38834
rect 74786 38782 74788 38834
rect 74620 38780 74788 38782
rect 74284 38052 74340 38062
rect 74172 37940 74228 37950
rect 74172 37846 74228 37884
rect 74060 37762 74116 37772
rect 73948 37548 74228 37604
rect 73724 37380 73780 37390
rect 73948 37380 74004 37390
rect 74060 37380 74116 37390
rect 73724 37378 73948 37380
rect 73724 37326 73726 37378
rect 73778 37326 73948 37378
rect 73724 37324 73948 37326
rect 74004 37378 74116 37380
rect 74004 37326 74062 37378
rect 74114 37326 74116 37378
rect 74004 37324 74116 37326
rect 73724 37314 73780 37324
rect 73388 37266 73668 37268
rect 73388 37214 73390 37266
rect 73442 37214 73668 37266
rect 73388 37212 73668 37214
rect 73388 37202 73444 37212
rect 73164 36866 73220 36876
rect 73276 37154 73332 37166
rect 73276 37102 73278 37154
rect 73330 37102 73332 37154
rect 72828 36482 72996 36484
rect 72828 36430 72830 36482
rect 72882 36430 72996 36482
rect 72828 36428 72996 36430
rect 73164 36484 73220 36494
rect 72828 36418 72884 36428
rect 73164 36390 73220 36428
rect 73052 36260 73108 36270
rect 73052 36166 73108 36204
rect 72716 35980 73220 36036
rect 72604 35924 72660 35934
rect 72716 35924 72772 35980
rect 72604 35922 72772 35924
rect 72604 35870 72606 35922
rect 72658 35870 72772 35922
rect 72604 35868 72772 35870
rect 72604 35858 72660 35868
rect 72940 35812 72996 35822
rect 72828 35810 72996 35812
rect 72828 35758 72942 35810
rect 72994 35758 72996 35810
rect 72828 35756 72996 35758
rect 72604 35028 72660 35038
rect 72492 35026 72660 35028
rect 72492 34974 72606 35026
rect 72658 34974 72660 35026
rect 72492 34972 72660 34974
rect 72380 34188 72548 34244
rect 72156 34130 72212 34188
rect 72156 34078 72158 34130
rect 72210 34078 72212 34130
rect 72156 34066 72212 34078
rect 72380 34020 72436 34030
rect 72268 34018 72436 34020
rect 72268 33966 72382 34018
rect 72434 33966 72436 34018
rect 72268 33964 72436 33966
rect 72044 33852 72212 33908
rect 72044 33570 72100 33582
rect 72044 33518 72046 33570
rect 72098 33518 72100 33570
rect 72044 33458 72100 33518
rect 72044 33406 72046 33458
rect 72098 33406 72100 33458
rect 72044 33394 72100 33406
rect 72156 32452 72212 33852
rect 72156 32386 72212 32396
rect 72268 32116 72324 33964
rect 72380 33954 72436 33964
rect 72268 32050 72324 32060
rect 72380 32674 72436 32686
rect 72380 32622 72382 32674
rect 72434 32622 72436 32674
rect 72268 31780 72324 31790
rect 72380 31780 72436 32622
rect 72268 31778 72436 31780
rect 72268 31726 72270 31778
rect 72322 31726 72436 31778
rect 72268 31724 72436 31726
rect 72156 31666 72212 31678
rect 72156 31614 72158 31666
rect 72210 31614 72212 31666
rect 71820 31218 71988 31220
rect 71820 31166 71822 31218
rect 71874 31166 71988 31218
rect 71820 31164 71988 31166
rect 72044 31554 72100 31566
rect 72044 31502 72046 31554
rect 72098 31502 72100 31554
rect 71820 30770 71876 31164
rect 71820 30718 71822 30770
rect 71874 30718 71876 30770
rect 71820 30706 71876 30718
rect 71596 30046 71598 30098
rect 71650 30046 71652 30098
rect 71596 30034 71652 30046
rect 71820 30210 71876 30222
rect 71820 30158 71822 30210
rect 71874 30158 71876 30210
rect 71484 29708 71652 29764
rect 71148 29596 71540 29652
rect 71372 29428 71428 29438
rect 71036 29426 71428 29428
rect 71036 29374 71038 29426
rect 71090 29374 71374 29426
rect 71426 29374 71428 29426
rect 71036 29372 71428 29374
rect 71036 29362 71092 29372
rect 71260 29092 71316 29102
rect 71260 28754 71316 29036
rect 71260 28702 71262 28754
rect 71314 28702 71316 28754
rect 71260 28690 71316 28702
rect 70700 28084 70756 28094
rect 70700 27990 70756 28028
rect 70588 27022 70590 27074
rect 70642 27022 70644 27074
rect 70588 27010 70644 27022
rect 70700 27860 70756 27870
rect 69580 26796 69748 26852
rect 69580 26740 69636 26796
rect 68796 26002 68852 26012
rect 69356 26684 69636 26740
rect 68684 23090 68740 23100
rect 67676 22418 67732 22428
rect 66668 20738 66724 20748
rect 67228 21700 67284 21710
rect 63756 20692 63812 20702
rect 63756 17108 63812 20636
rect 65916 19628 66180 19638
rect 65972 19572 66020 19628
rect 66076 19572 66124 19628
rect 65916 19562 66180 19572
rect 63756 17042 63812 17052
rect 64540 18676 64596 18686
rect 63868 9716 63924 9726
rect 63868 6132 63924 9660
rect 64428 6468 64484 6478
rect 64428 6374 64484 6412
rect 63868 6130 64484 6132
rect 63868 6078 63870 6130
rect 63922 6078 64484 6130
rect 63868 6076 64484 6078
rect 63868 6066 63924 6076
rect 64428 5906 64484 6076
rect 64428 5854 64430 5906
rect 64482 5854 64484 5906
rect 64428 5842 64484 5854
rect 64428 5236 64484 5246
rect 64428 5142 64484 5180
rect 63196 4510 63198 4562
rect 63250 4510 63252 4562
rect 63196 4498 63252 4510
rect 63308 4562 63700 4564
rect 63308 4510 63534 4562
rect 63586 4510 63700 4562
rect 63308 4508 63700 4510
rect 63756 5124 63812 5134
rect 63308 4340 63364 4508
rect 63532 4498 63588 4508
rect 63084 4284 63364 4340
rect 63084 3554 63140 4284
rect 63084 3502 63086 3554
rect 63138 3502 63140 3554
rect 63084 3490 63140 3502
rect 63756 980 63812 5068
rect 64540 4338 64596 18620
rect 67228 18452 67284 21644
rect 67788 20916 67844 20926
rect 67788 19012 67844 20860
rect 68908 20244 68964 20254
rect 67788 18946 67844 18956
rect 67900 19908 67956 19918
rect 67228 18386 67284 18396
rect 65916 18060 66180 18070
rect 65972 18004 66020 18060
rect 66076 18004 66124 18060
rect 65916 17994 66180 18004
rect 65916 16492 66180 16502
rect 65972 16436 66020 16492
rect 66076 16436 66124 16492
rect 65916 16426 66180 16436
rect 65916 14924 66180 14934
rect 65972 14868 66020 14924
rect 66076 14868 66124 14924
rect 65916 14858 66180 14868
rect 65916 13356 66180 13366
rect 65972 13300 66020 13356
rect 66076 13300 66124 13356
rect 65916 13290 66180 13300
rect 65916 11788 66180 11798
rect 65972 11732 66020 11788
rect 66076 11732 66124 11788
rect 65916 11722 66180 11732
rect 65916 10220 66180 10230
rect 65972 10164 66020 10220
rect 66076 10164 66124 10220
rect 65916 10154 66180 10164
rect 66556 9268 66612 9278
rect 65916 8652 66180 8662
rect 65972 8596 66020 8652
rect 66076 8596 66124 8652
rect 65916 8586 66180 8596
rect 65916 7084 66180 7094
rect 65972 7028 66020 7084
rect 66076 7028 66124 7084
rect 65916 7018 66180 7028
rect 65548 5794 65604 5806
rect 65548 5742 65550 5794
rect 65602 5742 65604 5794
rect 65548 5124 65604 5742
rect 65916 5516 66180 5526
rect 65972 5460 66020 5516
rect 66076 5460 66124 5516
rect 65916 5450 66180 5460
rect 65548 5058 65604 5068
rect 66332 5236 66388 5246
rect 64540 4286 64542 4338
rect 64594 4286 64596 4338
rect 64092 4116 64148 4126
rect 63868 3668 63924 3678
rect 63868 3574 63924 3612
rect 63420 924 63812 980
rect 63420 800 63476 924
rect 64092 800 64148 4060
rect 64540 3668 64596 4286
rect 65548 4226 65604 4238
rect 65548 4174 65550 4226
rect 65602 4174 65604 4226
rect 65548 3780 65604 4174
rect 65916 3948 66180 3958
rect 65972 3892 66020 3948
rect 66076 3892 66124 3948
rect 65916 3882 66180 3892
rect 65548 3714 65604 3724
rect 64540 3602 64596 3612
rect 65660 3668 65716 3678
rect 65660 3574 65716 3612
rect 65436 3556 65492 3566
rect 64764 3444 64820 3454
rect 64764 800 64820 3388
rect 65436 800 65492 3500
rect 66332 2660 66388 5180
rect 66444 5236 66500 5246
rect 66556 5236 66612 9212
rect 66668 7700 66724 7710
rect 66724 7644 67060 7700
rect 66668 7606 66724 7644
rect 67004 7474 67060 7644
rect 67004 7422 67006 7474
rect 67058 7422 67060 7474
rect 67004 7410 67060 7422
rect 66444 5234 66612 5236
rect 66444 5182 66446 5234
rect 66498 5182 66612 5234
rect 66444 5180 66612 5182
rect 67116 7252 67172 7262
rect 67116 6020 67172 7196
rect 67900 6692 67956 19852
rect 68796 17444 68852 17454
rect 68796 15092 68852 17388
rect 68908 16324 68964 20188
rect 68908 16258 68964 16268
rect 68796 15026 68852 15036
rect 68460 14420 68516 14430
rect 68348 6692 68404 6702
rect 67900 6690 68404 6692
rect 67900 6638 67902 6690
rect 67954 6638 68350 6690
rect 68402 6638 68404 6690
rect 67900 6636 68404 6638
rect 67900 6626 67956 6636
rect 68348 6626 68404 6636
rect 67340 6468 67396 6478
rect 67340 6466 67508 6468
rect 67340 6414 67342 6466
rect 67394 6414 67508 6466
rect 67340 6412 67508 6414
rect 67340 6402 67396 6412
rect 67116 5964 67396 6020
rect 67116 5234 67172 5964
rect 67340 5906 67396 5964
rect 67340 5854 67342 5906
rect 67394 5854 67396 5906
rect 67340 5842 67396 5854
rect 67340 5572 67396 5582
rect 67116 5182 67118 5234
rect 67170 5182 67172 5234
rect 66444 3554 66500 5180
rect 67116 5170 67172 5182
rect 67228 5516 67340 5572
rect 66444 3502 66446 3554
rect 66498 3502 66500 3554
rect 66444 3490 66500 3502
rect 66780 5124 66836 5134
rect 66108 2604 66388 2660
rect 66108 800 66164 2604
rect 66780 800 66836 5068
rect 67228 3220 67284 5516
rect 67340 5506 67396 5516
rect 67340 5346 67396 5358
rect 67340 5294 67342 5346
rect 67394 5294 67396 5346
rect 67340 4900 67396 5294
rect 67452 5124 67508 6412
rect 67564 6132 67620 6142
rect 67564 5346 67620 6076
rect 67564 5294 67566 5346
rect 67618 5294 67620 5346
rect 67564 5282 67620 5294
rect 68348 5124 68404 5134
rect 68460 5124 68516 14364
rect 69356 10948 69412 26684
rect 69580 26404 69636 26414
rect 69580 23548 69636 26348
rect 70588 26066 70644 26078
rect 70588 26014 70590 26066
rect 70642 26014 70644 26066
rect 70588 25956 70644 26014
rect 70364 25900 70644 25956
rect 70364 25508 70420 25900
rect 70700 25844 70756 27804
rect 70924 27860 70980 27870
rect 71372 27860 71428 29372
rect 71484 27972 71540 29596
rect 71596 28532 71652 29708
rect 71708 29540 71764 29550
rect 71820 29540 71876 30158
rect 71708 29538 71876 29540
rect 71708 29486 71710 29538
rect 71762 29486 71876 29538
rect 71708 29484 71876 29486
rect 71708 29474 71764 29484
rect 71708 28756 71764 28766
rect 71708 28662 71764 28700
rect 71820 28644 71876 29484
rect 71932 28644 71988 28654
rect 71820 28588 71932 28644
rect 71932 28578 71988 28588
rect 71596 28476 71876 28532
rect 71820 28420 71876 28476
rect 71820 28364 71988 28420
rect 71820 28196 71876 28206
rect 71820 28082 71876 28140
rect 71820 28030 71822 28082
rect 71874 28030 71876 28082
rect 71820 28018 71876 28030
rect 71932 27972 71988 28364
rect 71484 27916 71764 27972
rect 71372 27804 71652 27860
rect 70924 27766 70980 27804
rect 70812 27746 70868 27758
rect 70812 27694 70814 27746
rect 70866 27694 70868 27746
rect 70812 26178 70868 27694
rect 71372 27636 71428 27646
rect 71036 27076 71092 27086
rect 71372 27076 71428 27580
rect 71036 27074 71428 27076
rect 71036 27022 71038 27074
rect 71090 27022 71428 27074
rect 71036 27020 71428 27022
rect 71036 27010 71092 27020
rect 71148 26852 71204 26862
rect 71036 26850 71204 26852
rect 71036 26798 71150 26850
rect 71202 26798 71204 26850
rect 71036 26796 71204 26798
rect 70924 26516 70980 26526
rect 70924 26422 70980 26460
rect 71036 26292 71092 26796
rect 71148 26786 71204 26796
rect 71260 26850 71316 26862
rect 71260 26798 71262 26850
rect 71314 26798 71316 26850
rect 71260 26404 71316 26798
rect 71260 26338 71316 26348
rect 70812 26126 70814 26178
rect 70866 26126 70868 26178
rect 70812 26114 70868 26126
rect 70924 26236 71092 26292
rect 71148 26290 71204 26302
rect 71148 26238 71150 26290
rect 71202 26238 71204 26290
rect 70476 25788 70756 25844
rect 70476 25620 70532 25788
rect 70476 25564 70756 25620
rect 70700 25508 70756 25564
rect 70812 25508 70868 25518
rect 70364 25452 70644 25508
rect 69468 23492 69636 23548
rect 69468 23380 69524 23492
rect 69468 23314 69524 23324
rect 70588 22596 70644 25452
rect 70700 25506 70868 25508
rect 70700 25454 70814 25506
rect 70866 25454 70868 25506
rect 70700 25452 70868 25454
rect 70700 25394 70756 25452
rect 70812 25442 70868 25452
rect 70700 25342 70702 25394
rect 70754 25342 70756 25394
rect 70700 25330 70756 25342
rect 70812 24724 70868 24734
rect 70924 24724 70980 26236
rect 71148 25956 71204 26238
rect 71372 26290 71428 26302
rect 71372 26238 71374 26290
rect 71426 26238 71428 26290
rect 71148 25890 71204 25900
rect 71260 26178 71316 26190
rect 71260 26126 71262 26178
rect 71314 26126 71316 26178
rect 71036 25618 71092 25630
rect 71036 25566 71038 25618
rect 71090 25566 71092 25618
rect 71036 25284 71092 25566
rect 71036 25218 71092 25228
rect 70868 24668 70980 24724
rect 70812 24658 70868 24668
rect 71260 24500 71316 26126
rect 71372 25396 71428 26238
rect 71372 25330 71428 25340
rect 71372 24612 71428 24622
rect 71372 24518 71428 24556
rect 70700 24444 71316 24500
rect 70700 23044 70756 24444
rect 70700 22978 70756 22988
rect 71372 24388 71428 24398
rect 70588 22530 70644 22540
rect 70924 22708 70980 22718
rect 70364 22260 70420 22270
rect 70028 21812 70084 21822
rect 70084 21756 70308 21812
rect 70028 21718 70084 21756
rect 70252 21586 70308 21756
rect 70252 21534 70254 21586
rect 70306 21534 70308 21586
rect 70252 21522 70308 21534
rect 70364 19348 70420 22204
rect 70364 19282 70420 19292
rect 70588 21474 70644 21486
rect 70588 21422 70590 21474
rect 70642 21422 70644 21474
rect 70588 17780 70644 21422
rect 70924 20916 70980 22652
rect 71372 21586 71428 24332
rect 71596 23548 71652 27804
rect 71708 26908 71764 27916
rect 71932 27906 71988 27916
rect 71932 27412 71988 27422
rect 71932 27186 71988 27356
rect 71932 27134 71934 27186
rect 71986 27134 71988 27186
rect 71932 27122 71988 27134
rect 71708 26852 71876 26908
rect 71820 25506 71876 26852
rect 71820 25454 71822 25506
rect 71874 25454 71876 25506
rect 71820 25442 71876 25454
rect 71708 24948 71764 24958
rect 71708 24854 71764 24892
rect 71372 21534 71374 21586
rect 71426 21534 71428 21586
rect 71372 21522 71428 21534
rect 71484 23492 71652 23548
rect 70924 20914 71092 20916
rect 70924 20862 70926 20914
rect 70978 20862 71092 20914
rect 70924 20860 71092 20862
rect 70924 20850 70980 20860
rect 71036 20802 71092 20860
rect 71036 20750 71038 20802
rect 71090 20750 71092 20802
rect 71036 20738 71092 20750
rect 71260 20914 71316 20926
rect 71260 20862 71262 20914
rect 71314 20862 71316 20914
rect 71260 20692 71316 20862
rect 71260 20626 71316 20636
rect 71484 20356 71540 23492
rect 71708 23380 71764 23390
rect 71708 23286 71764 23324
rect 71708 23156 71764 23166
rect 71708 22482 71764 23100
rect 71708 22430 71710 22482
rect 71762 22430 71764 22482
rect 71708 22372 71764 22430
rect 71708 22306 71764 22316
rect 71596 21586 71652 21598
rect 71596 21534 71598 21586
rect 71650 21534 71652 21586
rect 71596 21476 71652 21534
rect 71596 21410 71652 21420
rect 72044 20802 72100 31502
rect 72156 31444 72212 31614
rect 72268 31556 72324 31724
rect 72268 31490 72324 31500
rect 72156 31378 72212 31388
rect 72492 30324 72548 34188
rect 72604 34242 72660 34972
rect 72828 34914 72884 35756
rect 72940 35746 72996 35756
rect 73164 35698 73220 35980
rect 73276 35924 73332 37102
rect 73612 37156 73668 37212
rect 73612 37100 73892 37156
rect 73388 37044 73444 37054
rect 73388 36482 73444 36988
rect 73388 36430 73390 36482
rect 73442 36430 73444 36482
rect 73388 36418 73444 36430
rect 73500 36932 73556 36942
rect 73276 35868 73444 35924
rect 73164 35646 73166 35698
rect 73218 35646 73220 35698
rect 73164 35634 73220 35646
rect 73276 35700 73332 35710
rect 72828 34862 72830 34914
rect 72882 34862 72884 34914
rect 72828 34468 72884 34862
rect 72828 34402 72884 34412
rect 72940 35252 72996 35262
rect 72940 34244 72996 35196
rect 73276 34914 73332 35644
rect 73276 34862 73278 34914
rect 73330 34862 73332 34914
rect 73276 34850 73332 34862
rect 73052 34692 73108 34702
rect 73052 34598 73108 34636
rect 72604 34190 72606 34242
rect 72658 34190 72660 34242
rect 72604 34178 72660 34190
rect 72828 34188 72996 34244
rect 73164 34468 73220 34478
rect 73164 34244 73220 34412
rect 72716 34132 72772 34142
rect 72716 34038 72772 34076
rect 72716 33348 72772 33358
rect 72828 33348 72884 34188
rect 73164 34150 73220 34188
rect 73276 34020 73332 34030
rect 72716 33346 72884 33348
rect 72716 33294 72718 33346
rect 72770 33294 72884 33346
rect 72716 33292 72884 33294
rect 73164 34018 73332 34020
rect 73164 33966 73278 34018
rect 73330 33966 73332 34018
rect 73164 33964 73332 33966
rect 72716 32674 72772 33292
rect 72940 33122 72996 33134
rect 72940 33070 72942 33122
rect 72994 33070 72996 33122
rect 72940 33012 72996 33070
rect 72940 32946 72996 32956
rect 72716 32622 72718 32674
rect 72770 32622 72772 32674
rect 72716 32610 72772 32622
rect 72604 31892 72660 31902
rect 72604 31778 72660 31836
rect 72604 31726 72606 31778
rect 72658 31726 72660 31778
rect 72604 31714 72660 31726
rect 73052 31780 73108 31790
rect 73052 31686 73108 31724
rect 72828 31554 72884 31566
rect 72828 31502 72830 31554
rect 72882 31502 72884 31554
rect 72716 31444 72772 31454
rect 72716 31218 72772 31388
rect 72716 31166 72718 31218
rect 72770 31166 72772 31218
rect 72716 31154 72772 31166
rect 72380 30268 72548 30324
rect 72156 29764 72212 29774
rect 72156 28754 72212 29708
rect 72380 29650 72436 30268
rect 72828 30212 72884 31502
rect 72828 30146 72884 30156
rect 72492 30098 72548 30110
rect 72492 30046 72494 30098
rect 72546 30046 72548 30098
rect 72492 29988 72548 30046
rect 72716 30100 72772 30110
rect 72716 30006 72772 30044
rect 73052 30098 73108 30110
rect 73052 30046 73054 30098
rect 73106 30046 73108 30098
rect 72604 29988 72660 29998
rect 72492 29932 72604 29988
rect 72604 29922 72660 29932
rect 72828 29988 72884 29998
rect 73052 29988 73108 30046
rect 72828 29986 72996 29988
rect 72828 29934 72830 29986
rect 72882 29934 72996 29986
rect 72828 29932 72996 29934
rect 72828 29922 72884 29932
rect 72716 29876 72772 29886
rect 72380 29598 72382 29650
rect 72434 29598 72436 29650
rect 72380 29586 72436 29598
rect 72604 29652 72660 29662
rect 72716 29652 72772 29820
rect 72604 29650 72772 29652
rect 72604 29598 72606 29650
rect 72658 29598 72772 29650
rect 72604 29596 72772 29598
rect 72604 29586 72660 29596
rect 72828 29426 72884 29438
rect 72828 29374 72830 29426
rect 72882 29374 72884 29426
rect 72716 29316 72772 29326
rect 72716 29222 72772 29260
rect 72604 28980 72660 28990
rect 72156 28702 72158 28754
rect 72210 28702 72212 28754
rect 72156 28690 72212 28702
rect 72492 28924 72604 28980
rect 72380 28644 72436 28654
rect 72380 28550 72436 28588
rect 72268 27972 72324 27982
rect 72156 25506 72212 25518
rect 72156 25454 72158 25506
rect 72210 25454 72212 25506
rect 72156 25172 72212 25454
rect 72268 25508 72324 27916
rect 72380 27076 72436 27114
rect 72380 27010 72436 27020
rect 72380 26852 72436 26862
rect 72380 26516 72436 26796
rect 72492 26740 72548 28924
rect 72604 28914 72660 28924
rect 72716 28532 72772 28542
rect 72716 28438 72772 28476
rect 72828 28196 72884 29374
rect 72940 28980 72996 29932
rect 73052 29922 73108 29932
rect 72940 28914 72996 28924
rect 72828 28130 72884 28140
rect 72940 28532 72996 28542
rect 72716 27972 72772 27982
rect 72716 27878 72772 27916
rect 72940 27970 72996 28476
rect 72940 27918 72942 27970
rect 72994 27918 72996 27970
rect 72940 27906 72996 27918
rect 73052 27748 73108 27758
rect 72716 27746 73108 27748
rect 72716 27694 73054 27746
rect 73106 27694 73108 27746
rect 72716 27692 73108 27694
rect 72604 27300 72660 27310
rect 72604 26908 72660 27244
rect 72716 27076 72772 27692
rect 73052 27682 73108 27692
rect 73164 27188 73220 33964
rect 73276 33954 73332 33964
rect 73276 31666 73332 31678
rect 73276 31614 73278 31666
rect 73330 31614 73332 31666
rect 73276 31556 73332 31614
rect 73276 30210 73332 31500
rect 73276 30158 73278 30210
rect 73330 30158 73332 30210
rect 73276 30146 73332 30158
rect 73276 29652 73332 29662
rect 73388 29652 73444 35868
rect 73500 35252 73556 36876
rect 73836 36594 73892 37100
rect 73948 37044 74004 37324
rect 74060 37314 74116 37324
rect 73948 36978 74004 36988
rect 74060 37156 74116 37166
rect 73836 36542 73838 36594
rect 73890 36542 73892 36594
rect 73836 36530 73892 36542
rect 74060 36372 74116 37100
rect 73724 36316 74116 36372
rect 73612 36260 73668 36270
rect 73612 35364 73668 36204
rect 73612 35298 73668 35308
rect 73500 35186 73556 35196
rect 73612 35140 73668 35150
rect 73500 34804 73556 34814
rect 73500 34710 73556 34748
rect 73500 34244 73556 34254
rect 73612 34244 73668 35084
rect 73724 34468 73780 36316
rect 74172 35810 74228 37548
rect 74284 37492 74340 37996
rect 74508 38052 74564 38062
rect 74620 38052 74676 38780
rect 74732 38770 74788 38780
rect 74564 37996 74676 38052
rect 74844 38050 74900 41356
rect 75180 41300 75236 41310
rect 75180 41206 75236 41244
rect 74956 41186 75012 41198
rect 74956 41134 74958 41186
rect 75010 41134 75012 41186
rect 74956 40404 75012 41134
rect 75292 41076 75348 41804
rect 75740 41748 75796 42028
rect 75516 41692 75796 41748
rect 75516 41410 75572 41692
rect 75516 41358 75518 41410
rect 75570 41358 75572 41410
rect 75516 41346 75572 41358
rect 76188 41076 76244 41086
rect 75180 41020 75348 41076
rect 75740 41074 76244 41076
rect 75740 41022 76190 41074
rect 76242 41022 76244 41074
rect 75740 41020 76244 41022
rect 74956 40338 75012 40348
rect 75068 40402 75124 40414
rect 75068 40350 75070 40402
rect 75122 40350 75124 40402
rect 75068 39844 75124 40350
rect 75068 39778 75124 39788
rect 74956 39618 75012 39630
rect 74956 39566 74958 39618
rect 75010 39566 75012 39618
rect 74956 39508 75012 39566
rect 74956 39442 75012 39452
rect 75180 39172 75236 41020
rect 75292 40514 75348 40526
rect 75292 40462 75294 40514
rect 75346 40462 75348 40514
rect 75292 39956 75348 40462
rect 75292 39890 75348 39900
rect 75404 40180 75460 40190
rect 75292 39620 75348 39630
rect 75292 39394 75348 39564
rect 75404 39618 75460 40124
rect 75404 39566 75406 39618
rect 75458 39566 75460 39618
rect 75404 39554 75460 39566
rect 75628 39732 75684 39742
rect 75628 39618 75684 39676
rect 75628 39566 75630 39618
rect 75682 39566 75684 39618
rect 75628 39554 75684 39566
rect 75292 39342 75294 39394
rect 75346 39342 75348 39394
rect 75292 39330 75348 39342
rect 75180 39116 75348 39172
rect 75068 38948 75124 38958
rect 75068 38834 75124 38892
rect 75068 38782 75070 38834
rect 75122 38782 75124 38834
rect 75068 38770 75124 38782
rect 74956 38722 75012 38734
rect 74956 38670 74958 38722
rect 75010 38670 75012 38722
rect 74956 38276 75012 38670
rect 74956 38210 75012 38220
rect 75068 38612 75124 38622
rect 74844 37998 74846 38050
rect 74898 37998 74900 38050
rect 74508 37958 74564 37996
rect 74844 37986 74900 37998
rect 75068 38050 75124 38556
rect 75068 37998 75070 38050
rect 75122 37998 75124 38050
rect 75068 37986 75124 37998
rect 74620 37828 74676 37838
rect 74620 37826 74788 37828
rect 74620 37774 74622 37826
rect 74674 37774 74788 37826
rect 74620 37772 74788 37774
rect 74620 37762 74676 37772
rect 74284 37426 74340 37436
rect 74284 37268 74340 37278
rect 74284 37174 74340 37212
rect 74620 37268 74676 37278
rect 74620 37174 74676 37212
rect 74508 37156 74564 37166
rect 74508 37062 74564 37100
rect 74284 37044 74340 37054
rect 74340 36988 74452 37044
rect 74284 36978 74340 36988
rect 74396 36594 74452 36988
rect 74732 36820 74788 37772
rect 75068 37268 75124 37278
rect 75068 37174 75124 37212
rect 75180 37154 75236 37166
rect 75180 37102 75182 37154
rect 75234 37102 75236 37154
rect 75180 37044 75236 37102
rect 75292 37044 75348 39116
rect 75740 39060 75796 41020
rect 76188 41010 76244 41020
rect 75404 39004 75796 39060
rect 75852 40180 75908 40190
rect 75404 38946 75460 39004
rect 75404 38894 75406 38946
rect 75458 38894 75460 38946
rect 75404 38612 75460 38894
rect 75404 38546 75460 38556
rect 75628 37378 75684 39004
rect 75740 38164 75796 38174
rect 75852 38164 75908 40124
rect 75964 39844 76020 39854
rect 75964 39058 76020 39788
rect 75964 39006 75966 39058
rect 76018 39006 76020 39058
rect 75964 38994 76020 39006
rect 76076 39732 76132 39742
rect 75740 38162 75908 38164
rect 75740 38110 75742 38162
rect 75794 38110 75908 38162
rect 75740 38108 75908 38110
rect 76076 38836 76132 39676
rect 76188 39508 76244 39518
rect 76188 39414 76244 39452
rect 76300 39396 76356 43484
rect 76524 42868 76580 42878
rect 76524 42774 76580 42812
rect 76412 42756 76468 42766
rect 76412 41300 76468 42700
rect 76412 41186 76468 41244
rect 76412 41134 76414 41186
rect 76466 41134 76468 41186
rect 76412 41122 76468 41134
rect 76748 42754 76804 42766
rect 76748 42702 76750 42754
rect 76802 42702 76804 42754
rect 76748 41412 76804 42702
rect 76748 41186 76804 41356
rect 76748 41134 76750 41186
rect 76802 41134 76804 41186
rect 76524 41076 76580 41086
rect 76524 40514 76580 41020
rect 76524 40462 76526 40514
rect 76578 40462 76580 40514
rect 76524 40450 76580 40462
rect 76636 40962 76692 40974
rect 76636 40910 76638 40962
rect 76690 40910 76692 40962
rect 76524 39620 76580 39630
rect 76524 39526 76580 39564
rect 76300 39340 76580 39396
rect 76412 38948 76468 38958
rect 76300 38836 76356 38846
rect 76076 38834 76356 38836
rect 76076 38782 76302 38834
rect 76354 38782 76356 38834
rect 76076 38780 76356 38782
rect 75740 38098 75796 38108
rect 75628 37326 75630 37378
rect 75682 37326 75684 37378
rect 75628 37314 75684 37326
rect 76076 37940 76132 38780
rect 76300 38770 76356 38780
rect 76412 38162 76468 38892
rect 76524 38946 76580 39340
rect 76524 38894 76526 38946
rect 76578 38894 76580 38946
rect 76524 38882 76580 38894
rect 76412 38110 76414 38162
rect 76466 38110 76468 38162
rect 76412 38098 76468 38110
rect 75404 37268 75460 37278
rect 75404 37174 75460 37212
rect 76076 37266 76132 37884
rect 76188 37940 76244 37950
rect 76188 37938 76356 37940
rect 76188 37886 76190 37938
rect 76242 37886 76356 37938
rect 76188 37884 76356 37886
rect 76188 37874 76244 37884
rect 76188 37380 76244 37390
rect 76188 37286 76244 37324
rect 76076 37214 76078 37266
rect 76130 37214 76132 37266
rect 75516 37156 75572 37166
rect 75292 36988 75460 37044
rect 75180 36978 75236 36988
rect 74396 36542 74398 36594
rect 74450 36542 74452 36594
rect 74396 36530 74452 36542
rect 74508 36764 74788 36820
rect 74172 35758 74174 35810
rect 74226 35758 74228 35810
rect 74172 35746 74228 35758
rect 74284 35922 74340 35934
rect 74508 35924 74564 36764
rect 74732 36596 74788 36606
rect 74732 36482 74788 36540
rect 75292 36484 75348 36494
rect 74732 36430 74734 36482
rect 74786 36430 74788 36482
rect 74732 36418 74788 36430
rect 74956 36482 75348 36484
rect 74956 36430 75294 36482
rect 75346 36430 75348 36482
rect 74956 36428 75348 36430
rect 74956 36370 75012 36428
rect 75292 36418 75348 36428
rect 74956 36318 74958 36370
rect 75010 36318 75012 36370
rect 74956 36306 75012 36318
rect 75404 36260 75460 36988
rect 75516 36594 75572 37100
rect 75516 36542 75518 36594
rect 75570 36542 75572 36594
rect 75516 36530 75572 36542
rect 75628 36372 75684 36382
rect 75628 36278 75684 36316
rect 75292 36204 75460 36260
rect 74284 35870 74286 35922
rect 74338 35870 74340 35922
rect 74060 35698 74116 35710
rect 74060 35646 74062 35698
rect 74114 35646 74116 35698
rect 74060 35588 74116 35646
rect 74284 35588 74340 35870
rect 74396 35868 74564 35924
rect 75068 36036 75124 36046
rect 74396 35700 74452 35868
rect 74620 35700 74676 35710
rect 74732 35700 74788 35710
rect 74396 35644 74564 35700
rect 74060 35532 74228 35588
rect 74060 35364 74116 35374
rect 73836 35252 73892 35262
rect 73836 34916 73892 35196
rect 73948 34916 74004 34926
rect 73836 34914 74004 34916
rect 73836 34862 73950 34914
rect 74002 34862 74004 34914
rect 73836 34860 74004 34862
rect 73948 34850 74004 34860
rect 73948 34468 74004 34478
rect 73724 34412 73892 34468
rect 73500 34242 73668 34244
rect 73500 34190 73502 34242
rect 73554 34190 73668 34242
rect 73500 34188 73668 34190
rect 73500 34178 73556 34188
rect 73724 34132 73780 34142
rect 73724 34038 73780 34076
rect 73836 33908 73892 34412
rect 73612 33852 73892 33908
rect 73612 32564 73668 33852
rect 73948 33572 74004 34412
rect 73948 33478 74004 33516
rect 73836 33460 73892 33470
rect 73836 33366 73892 33404
rect 73724 33122 73780 33134
rect 73724 33070 73726 33122
rect 73778 33070 73780 33122
rect 73724 32788 73780 33070
rect 73724 32722 73780 32732
rect 73948 32900 74004 32910
rect 73724 32564 73780 32574
rect 73612 32562 73780 32564
rect 73612 32510 73726 32562
rect 73778 32510 73780 32562
rect 73612 32508 73780 32510
rect 73724 32498 73780 32508
rect 73500 32452 73556 32462
rect 73500 32358 73556 32396
rect 73724 31780 73780 31790
rect 73724 31686 73780 31724
rect 73500 31332 73556 31342
rect 73500 31218 73556 31276
rect 73500 31166 73502 31218
rect 73554 31166 73556 31218
rect 73500 31154 73556 31166
rect 73836 30996 73892 31006
rect 73836 30902 73892 30940
rect 73948 30210 74004 32844
rect 74060 31778 74116 35308
rect 74172 34692 74228 35532
rect 74284 35522 74340 35532
rect 74172 34598 74228 34636
rect 74284 34130 74340 34142
rect 74284 34078 74286 34130
rect 74338 34078 74340 34130
rect 74284 33348 74340 34078
rect 74284 33282 74340 33292
rect 74396 33458 74452 33470
rect 74396 33406 74398 33458
rect 74450 33406 74452 33458
rect 74396 33236 74452 33406
rect 74508 33346 74564 35644
rect 74620 35698 74788 35700
rect 74620 35646 74622 35698
rect 74674 35646 74734 35698
rect 74786 35646 74788 35698
rect 74620 35644 74788 35646
rect 74620 35476 74676 35644
rect 74732 35634 74788 35644
rect 74956 35588 75012 35598
rect 74620 35410 74676 35420
rect 74844 35586 75012 35588
rect 74844 35534 74958 35586
rect 75010 35534 75012 35586
rect 74844 35532 75012 35534
rect 74844 35308 74900 35532
rect 74956 35522 75012 35532
rect 75068 35364 75124 35980
rect 75180 35812 75236 35822
rect 75292 35812 75348 36204
rect 76076 36036 76132 37214
rect 76300 37268 76356 37884
rect 76412 37828 76468 37838
rect 76412 37734 76468 37772
rect 76636 37716 76692 40910
rect 76748 40964 76804 41134
rect 76748 40898 76804 40908
rect 76748 39730 76804 39742
rect 76748 39678 76750 39730
rect 76802 39678 76804 39730
rect 76748 38948 76804 39678
rect 76748 38882 76804 38892
rect 76748 38722 76804 38734
rect 76748 38670 76750 38722
rect 76802 38670 76804 38722
rect 76748 38276 76804 38670
rect 76860 38388 76916 43652
rect 76972 40180 77028 67172
rect 77644 66946 77700 66958
rect 77644 66894 77646 66946
rect 77698 66894 77700 66946
rect 77644 66836 77700 66894
rect 77644 66770 77700 66780
rect 77644 66050 77700 66062
rect 77644 65998 77646 66050
rect 77698 65998 77700 66050
rect 77644 65716 77700 65998
rect 77644 65650 77700 65660
rect 77644 64708 77700 64718
rect 77644 64614 77700 64652
rect 77420 64596 77476 64606
rect 77420 64502 77476 64540
rect 77644 64036 77700 64046
rect 77420 63924 77476 63934
rect 77420 63830 77476 63868
rect 77644 63922 77700 63980
rect 77644 63870 77646 63922
rect 77698 63870 77700 63922
rect 77644 63858 77700 63870
rect 77644 62916 77700 62926
rect 77644 62822 77700 62860
rect 77644 61572 77700 61582
rect 77644 61478 77700 61516
rect 77420 61346 77476 61358
rect 77420 61294 77422 61346
rect 77474 61294 77476 61346
rect 77420 61236 77476 61294
rect 77756 61348 77812 74734
rect 77868 74004 77924 74042
rect 77868 73938 77924 73948
rect 77868 73444 77924 73454
rect 77868 73350 77924 73388
rect 77980 73220 78036 75740
rect 78204 75572 78260 75582
rect 78092 75570 78260 75572
rect 78092 75518 78206 75570
rect 78258 75518 78260 75570
rect 78092 75516 78260 75518
rect 78092 75460 78148 75516
rect 78204 75506 78260 75516
rect 78652 75572 78708 77420
rect 78652 75506 78708 75516
rect 78092 75394 78148 75404
rect 78204 75124 78260 75134
rect 78204 75030 78260 75068
rect 78764 75124 78820 77980
rect 78764 75058 78820 75068
rect 79100 75012 79156 79200
rect 79100 74946 79156 74956
rect 78316 74676 78372 74686
rect 78092 74116 78148 74126
rect 78092 74022 78148 74060
rect 78204 73556 78260 73566
rect 78316 73556 78372 74620
rect 78260 73500 78372 73556
rect 78204 73462 78260 73500
rect 77980 73164 78484 73220
rect 78204 72436 78260 72446
rect 78204 72342 78260 72380
rect 77868 72324 77924 72334
rect 77868 72230 77924 72268
rect 77868 71876 77924 71886
rect 77868 71782 77924 71820
rect 78204 71762 78260 71774
rect 78204 71710 78206 71762
rect 78258 71710 78260 71762
rect 78204 71316 78260 71710
rect 78204 71250 78260 71260
rect 78204 70756 78260 70766
rect 78204 70196 78260 70700
rect 78204 70130 78260 70140
rect 77868 69188 77924 69198
rect 77868 69094 77924 69132
rect 78204 69186 78260 69198
rect 78204 69134 78206 69186
rect 78258 69134 78260 69186
rect 78204 69076 78260 69134
rect 78204 69010 78260 69020
rect 78204 68628 78260 68638
rect 78204 67956 78260 68572
rect 78204 67890 78260 67900
rect 78428 67228 78484 73164
rect 78764 70980 78820 70990
rect 78764 67228 78820 70924
rect 77868 67172 77924 67182
rect 78428 67172 78708 67228
rect 78764 67172 78932 67228
rect 77868 67170 78148 67172
rect 77868 67118 77870 67170
rect 77922 67118 78148 67170
rect 77868 67116 78148 67118
rect 77868 67106 77924 67116
rect 77868 66052 77924 66062
rect 77868 65958 77924 65996
rect 77868 62914 77924 62926
rect 77868 62862 77870 62914
rect 77922 62862 77924 62914
rect 77868 62244 77924 62862
rect 77868 62178 77924 62188
rect 78092 61572 78148 67116
rect 78204 67058 78260 67070
rect 78204 67006 78206 67058
rect 78258 67006 78260 67058
rect 78204 66836 78260 67006
rect 78204 66770 78260 66780
rect 78204 66050 78260 66062
rect 78204 65998 78206 66050
rect 78258 65998 78260 66050
rect 78204 65716 78260 65998
rect 78204 65650 78260 65660
rect 78204 64596 78260 64606
rect 78204 64502 78260 64540
rect 78204 63924 78260 63934
rect 78204 63476 78260 63868
rect 78204 63410 78260 63420
rect 78204 63026 78260 63038
rect 78204 62974 78206 63026
rect 78258 62974 78260 63026
rect 78204 62916 78260 62974
rect 78204 62356 78260 62860
rect 78204 62290 78260 62300
rect 78092 61516 78484 61572
rect 77756 61292 78036 61348
rect 77420 61170 77476 61180
rect 77868 60900 77924 60910
rect 77868 60806 77924 60844
rect 77644 60788 77700 60798
rect 77644 60694 77700 60732
rect 77420 59106 77476 59118
rect 77420 59054 77422 59106
rect 77474 59054 77476 59106
rect 77420 58996 77476 59054
rect 77644 59108 77700 59118
rect 77644 59014 77700 59052
rect 77420 58930 77476 58940
rect 77644 58210 77700 58222
rect 77644 58158 77646 58210
rect 77698 58158 77700 58210
rect 77644 57876 77700 58158
rect 77868 58212 77924 58222
rect 77868 58118 77924 58156
rect 77644 57810 77700 57820
rect 77644 56756 77700 56766
rect 77644 56662 77700 56700
rect 77868 56644 77924 56654
rect 77756 56642 77924 56644
rect 77756 56590 77870 56642
rect 77922 56590 77924 56642
rect 77756 56588 77924 56590
rect 77756 56196 77812 56588
rect 77868 56578 77924 56588
rect 77420 56140 77812 56196
rect 77868 56196 77924 56206
rect 77308 50372 77364 50382
rect 77308 45332 77364 50316
rect 77420 46900 77476 56140
rect 77868 56102 77924 56140
rect 77644 55970 77700 55982
rect 77644 55918 77646 55970
rect 77698 55918 77700 55970
rect 77644 55636 77700 55918
rect 77644 55570 77700 55580
rect 77644 55076 77700 55086
rect 77644 54982 77700 55020
rect 77868 55074 77924 55086
rect 77868 55022 77870 55074
rect 77922 55022 77924 55074
rect 77868 54068 77924 55022
rect 77868 54002 77924 54012
rect 77868 53844 77924 53854
rect 77868 53618 77924 53788
rect 77868 53566 77870 53618
rect 77922 53566 77924 53618
rect 77868 53554 77924 53566
rect 77644 53506 77700 53518
rect 77644 53454 77646 53506
rect 77698 53454 77700 53506
rect 77644 53396 77700 53454
rect 77644 53330 77700 53340
rect 77980 53284 78036 61292
rect 78204 61346 78260 61358
rect 78204 61294 78206 61346
rect 78258 61294 78260 61346
rect 78204 61236 78260 61294
rect 78204 61170 78260 61180
rect 78204 60788 78260 60798
rect 78204 60116 78260 60732
rect 78204 60050 78260 60060
rect 78204 59218 78260 59230
rect 78204 59166 78206 59218
rect 78258 59166 78260 59218
rect 78204 58996 78260 59166
rect 78204 58930 78260 58940
rect 78204 58210 78260 58222
rect 78204 58158 78206 58210
rect 78258 58158 78260 58210
rect 78204 57876 78260 58158
rect 78204 57810 78260 57820
rect 78204 56756 78260 56766
rect 78204 56662 78260 56700
rect 78204 56082 78260 56094
rect 78204 56030 78206 56082
rect 78258 56030 78260 56082
rect 78204 55636 78260 56030
rect 78204 55570 78260 55580
rect 78204 55186 78260 55198
rect 78204 55134 78206 55186
rect 78258 55134 78260 55186
rect 78204 55076 78260 55134
rect 78204 54516 78260 55020
rect 78204 54450 78260 54460
rect 78204 53618 78260 53630
rect 78204 53566 78206 53618
rect 78258 53566 78260 53618
rect 78204 53396 78260 53566
rect 78204 53330 78260 53340
rect 77756 53228 78036 53284
rect 77644 52836 77700 52846
rect 77644 52742 77700 52780
rect 77644 51266 77700 51278
rect 77644 51214 77646 51266
rect 77698 51214 77700 51266
rect 77644 51156 77700 51214
rect 77644 51090 77700 51100
rect 77644 50484 77700 50494
rect 77644 50390 77700 50428
rect 77756 49028 77812 53228
rect 77868 53060 77924 53070
rect 77868 53058 78148 53060
rect 77868 53006 77870 53058
rect 77922 53006 78148 53058
rect 77868 53004 78148 53006
rect 77868 52994 77924 53004
rect 77868 51492 77924 51502
rect 77868 51398 77924 51436
rect 77868 50372 77924 50382
rect 77868 50278 77924 50316
rect 77756 48972 78036 49028
rect 77644 48916 77700 48926
rect 77644 48822 77700 48860
rect 77868 48802 77924 48814
rect 77868 48750 77870 48802
rect 77922 48750 77924 48802
rect 77868 48580 77924 48750
rect 77420 46834 77476 46844
rect 77532 48524 77924 48580
rect 77532 46228 77588 48524
rect 77868 48356 77924 48366
rect 77868 48262 77924 48300
rect 77644 48130 77700 48142
rect 77644 48078 77646 48130
rect 77698 48078 77700 48130
rect 77644 47796 77700 48078
rect 77644 47730 77700 47740
rect 77644 47348 77700 47358
rect 77644 47254 77700 47292
rect 77868 47236 77924 47246
rect 77868 47142 77924 47180
rect 77532 46162 77588 46172
rect 77644 45666 77700 45678
rect 77868 45668 77924 45678
rect 77644 45614 77646 45666
rect 77698 45614 77700 45666
rect 77644 45556 77700 45614
rect 77644 45490 77700 45500
rect 77756 45666 77924 45668
rect 77756 45614 77870 45666
rect 77922 45614 77924 45666
rect 77756 45612 77924 45614
rect 77308 45266 77364 45276
rect 77644 44996 77700 45006
rect 77644 44902 77700 44940
rect 77756 44660 77812 45612
rect 77868 45602 77924 45612
rect 77868 45220 77924 45230
rect 77868 45126 77924 45164
rect 77756 44594 77812 44604
rect 77980 44098 78036 48972
rect 78092 47012 78148 53004
rect 78204 52946 78260 52958
rect 78204 52894 78206 52946
rect 78258 52894 78260 52946
rect 78204 52836 78260 52894
rect 78204 52276 78260 52780
rect 78204 52210 78260 52220
rect 78204 51378 78260 51390
rect 78204 51326 78206 51378
rect 78258 51326 78260 51378
rect 78204 51156 78260 51326
rect 78204 51090 78260 51100
rect 78204 50484 78260 50494
rect 78204 50036 78260 50428
rect 78204 49970 78260 49980
rect 78204 48916 78260 48926
rect 78204 48822 78260 48860
rect 78204 48242 78260 48254
rect 78204 48190 78206 48242
rect 78258 48190 78260 48242
rect 78204 47796 78260 48190
rect 78204 47730 78260 47740
rect 78092 46946 78148 46956
rect 78204 47348 78260 47358
rect 78204 46676 78260 47292
rect 78204 46610 78260 46620
rect 78204 45778 78260 45790
rect 78204 45726 78206 45778
rect 78258 45726 78260 45778
rect 78204 45556 78260 45726
rect 78204 45490 78260 45500
rect 78204 45106 78260 45118
rect 78204 45054 78206 45106
rect 78258 45054 78260 45106
rect 78204 44996 78260 45054
rect 78204 44436 78260 44940
rect 78204 44370 78260 44380
rect 77980 44046 77982 44098
rect 78034 44046 78036 44098
rect 77868 43652 77924 43662
rect 77868 43558 77924 43596
rect 77084 43540 77140 43550
rect 77084 43446 77140 43484
rect 77644 43426 77700 43438
rect 77644 43374 77646 43426
rect 77698 43374 77700 43426
rect 77644 43316 77700 43374
rect 77644 43250 77700 43260
rect 77308 43092 77364 43102
rect 77980 43092 78036 44046
rect 78204 43538 78260 43550
rect 78204 43486 78206 43538
rect 78258 43486 78260 43538
rect 78204 43316 78260 43486
rect 78204 43250 78260 43260
rect 77084 42868 77140 42878
rect 77084 42754 77140 42812
rect 77084 42702 77086 42754
rect 77138 42702 77140 42754
rect 77084 42690 77140 42702
rect 77084 42530 77140 42542
rect 77084 42478 77086 42530
rect 77138 42478 77140 42530
rect 77084 41300 77140 42478
rect 77308 41412 77364 43036
rect 77532 43036 78036 43092
rect 77420 42644 77476 42654
rect 77420 42550 77476 42588
rect 77308 41356 77476 41412
rect 77084 41244 77364 41300
rect 76972 40114 77028 40124
rect 77084 41074 77140 41086
rect 77084 41022 77086 41074
rect 77138 41022 77140 41074
rect 77084 40964 77140 41022
rect 76972 38836 77028 38846
rect 76972 38742 77028 38780
rect 77084 38834 77140 40908
rect 77196 40962 77252 40974
rect 77196 40910 77198 40962
rect 77250 40910 77252 40962
rect 77196 39172 77252 40910
rect 77308 39618 77364 41244
rect 77308 39566 77310 39618
rect 77362 39566 77364 39618
rect 77308 39554 77364 39566
rect 77420 41186 77476 41356
rect 77420 41134 77422 41186
rect 77474 41134 77476 41186
rect 77196 39106 77252 39116
rect 77420 39060 77476 41134
rect 77420 38994 77476 39004
rect 77532 38946 77588 43036
rect 77756 42642 77812 42654
rect 77756 42590 77758 42642
rect 77810 42590 77812 42642
rect 77756 42084 77812 42590
rect 78092 42532 78148 42542
rect 78092 42530 78260 42532
rect 78092 42478 78094 42530
rect 78146 42478 78260 42530
rect 78092 42476 78260 42478
rect 78092 42466 78148 42476
rect 77756 42018 77812 42028
rect 77980 42196 78036 42206
rect 77980 41858 78036 42140
rect 77980 41806 77982 41858
rect 78034 41806 78036 41858
rect 77980 41794 78036 41806
rect 78092 41300 78148 41310
rect 78092 41206 78148 41244
rect 77532 38894 77534 38946
rect 77586 38894 77588 38946
rect 77532 38882 77588 38894
rect 77644 41074 77700 41086
rect 77644 41022 77646 41074
rect 77698 41022 77700 41074
rect 77644 40964 77700 41022
rect 77644 40628 77700 40908
rect 77084 38782 77086 38834
rect 77138 38782 77140 38834
rect 77084 38770 77140 38782
rect 77644 38834 77700 40572
rect 78204 40402 78260 42476
rect 78204 40350 78206 40402
rect 78258 40350 78260 40402
rect 78204 40338 78260 40350
rect 77980 40292 78036 40302
rect 77980 39730 78036 40236
rect 78428 40180 78484 61516
rect 78540 48356 78596 48366
rect 78540 40852 78596 48300
rect 78540 40786 78596 40796
rect 78652 40292 78708 67172
rect 78764 47236 78820 47246
rect 78764 40404 78820 47180
rect 78876 43708 78932 67172
rect 78876 43652 79044 43708
rect 78764 40348 78932 40404
rect 78652 40236 78820 40292
rect 78428 40124 78708 40180
rect 77980 39678 77982 39730
rect 78034 39678 78036 39730
rect 77980 39666 78036 39678
rect 78092 39956 78148 39966
rect 77868 39508 77924 39518
rect 77644 38782 77646 38834
rect 77698 38782 77700 38834
rect 77644 38770 77700 38782
rect 77756 39506 77924 39508
rect 77756 39454 77870 39506
rect 77922 39454 77924 39506
rect 77756 39452 77924 39454
rect 77308 38722 77364 38734
rect 77308 38670 77310 38722
rect 77362 38670 77364 38722
rect 77308 38668 77364 38670
rect 77196 38612 77364 38668
rect 76860 38332 77140 38388
rect 76748 38220 76916 38276
rect 76636 37660 76804 37716
rect 76412 37492 76468 37502
rect 76412 37398 76468 37436
rect 76300 37212 76468 37268
rect 76076 35970 76132 35980
rect 76188 37044 76244 37054
rect 75180 35810 75348 35812
rect 75180 35758 75182 35810
rect 75234 35758 75348 35810
rect 75180 35756 75348 35758
rect 75628 35812 75684 35822
rect 75180 35746 75236 35756
rect 75404 35700 75460 35710
rect 74732 35252 74900 35308
rect 74956 35308 75124 35364
rect 75292 35698 75460 35700
rect 75292 35646 75406 35698
rect 75458 35646 75460 35698
rect 75292 35644 75460 35646
rect 74620 34690 74676 34702
rect 74620 34638 74622 34690
rect 74674 34638 74676 34690
rect 74620 34468 74676 34638
rect 74620 34402 74676 34412
rect 74620 34242 74676 34254
rect 74620 34190 74622 34242
rect 74674 34190 74676 34242
rect 74620 34132 74676 34190
rect 74620 34066 74676 34076
rect 74508 33294 74510 33346
rect 74562 33294 74564 33346
rect 74508 33282 74564 33294
rect 74396 33170 74452 33180
rect 74172 33124 74228 33134
rect 74172 32786 74228 33068
rect 74172 32734 74174 32786
rect 74226 32734 74228 32786
rect 74172 32722 74228 32734
rect 74396 32562 74452 32574
rect 74396 32510 74398 32562
rect 74450 32510 74452 32562
rect 74284 32450 74340 32462
rect 74284 32398 74286 32450
rect 74338 32398 74340 32450
rect 74284 32004 74340 32398
rect 74396 32116 74452 32510
rect 74396 32050 74452 32060
rect 74284 31938 74340 31948
rect 74732 31892 74788 35252
rect 74844 34914 74900 34926
rect 74844 34862 74846 34914
rect 74898 34862 74900 34914
rect 74844 33796 74900 34862
rect 74844 33730 74900 33740
rect 74844 33460 74900 33470
rect 74844 33366 74900 33404
rect 74956 32562 75012 35308
rect 75292 34692 75348 35644
rect 75404 35634 75460 35644
rect 75292 34468 75348 34636
rect 75180 34412 75348 34468
rect 75404 34914 75460 34926
rect 75404 34862 75406 34914
rect 75458 34862 75460 34914
rect 75068 34244 75124 34254
rect 75068 34130 75124 34188
rect 75068 34078 75070 34130
rect 75122 34078 75124 34130
rect 75068 34066 75124 34078
rect 75180 33684 75236 34412
rect 75292 34242 75348 34254
rect 75292 34190 75294 34242
rect 75346 34190 75348 34242
rect 75292 33908 75348 34190
rect 75292 33842 75348 33852
rect 75180 33618 75236 33628
rect 75068 33572 75124 33582
rect 75068 32676 75124 33516
rect 75292 33348 75348 33358
rect 75292 33254 75348 33292
rect 75068 32610 75124 32620
rect 75180 33236 75236 33246
rect 74956 32510 74958 32562
rect 75010 32510 75012 32562
rect 74956 32498 75012 32510
rect 74844 32340 74900 32350
rect 74844 32246 74900 32284
rect 75068 32340 75124 32350
rect 74060 31726 74062 31778
rect 74114 31726 74116 31778
rect 74060 31714 74116 31726
rect 74396 31836 74788 31892
rect 74956 32228 75012 32238
rect 74172 30996 74228 31006
rect 74172 30902 74228 30940
rect 74060 30324 74116 30334
rect 74060 30230 74116 30268
rect 73948 30158 73950 30210
rect 74002 30158 74004 30210
rect 73948 30146 74004 30158
rect 73276 29650 73444 29652
rect 73276 29598 73278 29650
rect 73330 29598 73444 29650
rect 73276 29596 73444 29598
rect 73500 29988 73556 29998
rect 73500 29650 73556 29932
rect 74396 29764 74452 31836
rect 74620 31668 74676 31678
rect 74620 31574 74676 31612
rect 74508 31556 74564 31566
rect 74508 31462 74564 31500
rect 74732 31554 74788 31566
rect 74732 31502 74734 31554
rect 74786 31502 74788 31554
rect 74508 31108 74564 31118
rect 74508 31014 74564 31052
rect 74732 30324 74788 31502
rect 74844 30996 74900 31006
rect 74844 30902 74900 30940
rect 74956 30772 75012 32172
rect 74732 30258 74788 30268
rect 74844 30716 75012 30772
rect 74060 29708 74452 29764
rect 74508 30100 74564 30110
rect 73500 29598 73502 29650
rect 73554 29598 73556 29650
rect 73276 29586 73332 29596
rect 73500 29586 73556 29598
rect 73724 29652 73780 29662
rect 73780 29596 73892 29652
rect 73724 29586 73780 29596
rect 73724 29428 73780 29438
rect 73724 29334 73780 29372
rect 73612 29314 73668 29326
rect 73612 29262 73614 29314
rect 73666 29262 73668 29314
rect 73612 29204 73668 29262
rect 73612 29138 73668 29148
rect 73388 28980 73444 28990
rect 73388 28754 73444 28924
rect 73724 28756 73780 28766
rect 73836 28756 73892 29596
rect 73388 28702 73390 28754
rect 73442 28702 73444 28754
rect 73388 28690 73444 28702
rect 73500 28754 73892 28756
rect 73500 28702 73726 28754
rect 73778 28702 73892 28754
rect 73500 28700 73892 28702
rect 73500 28532 73556 28700
rect 73724 28690 73780 28700
rect 73276 28476 73556 28532
rect 73724 28532 73780 28542
rect 73276 27970 73332 28476
rect 73276 27918 73278 27970
rect 73330 27918 73332 27970
rect 73276 27906 73332 27918
rect 73500 27860 73556 27870
rect 73164 27122 73220 27132
rect 73388 27300 73444 27310
rect 72716 27020 72996 27076
rect 72604 26852 72884 26908
rect 72828 26850 72884 26852
rect 72828 26798 72830 26850
rect 72882 26798 72884 26850
rect 72828 26786 72884 26798
rect 72492 26684 72660 26740
rect 72380 26450 72436 26460
rect 72380 26292 72436 26302
rect 72380 25508 72436 26236
rect 72492 25508 72548 25518
rect 72380 25506 72548 25508
rect 72380 25454 72494 25506
rect 72546 25454 72548 25506
rect 72380 25452 72548 25454
rect 72268 25442 72324 25452
rect 72492 25442 72548 25452
rect 72156 25106 72212 25116
rect 72156 24948 72212 24958
rect 72156 24722 72212 24892
rect 72156 24670 72158 24722
rect 72210 24670 72212 24722
rect 72156 24658 72212 24670
rect 72380 24500 72436 24510
rect 72380 24406 72436 24444
rect 72268 23938 72324 23950
rect 72268 23886 72270 23938
rect 72322 23886 72324 23938
rect 72156 23716 72212 23726
rect 72268 23716 72324 23886
rect 72212 23660 72324 23716
rect 72156 23622 72212 23660
rect 72156 23380 72212 23390
rect 72156 23154 72212 23324
rect 72156 23102 72158 23154
rect 72210 23102 72212 23154
rect 72156 23090 72212 23102
rect 72380 22930 72436 22942
rect 72380 22878 72382 22930
rect 72434 22878 72436 22930
rect 72156 22484 72212 22494
rect 72156 22372 72212 22428
rect 72268 22372 72324 22382
rect 72156 22370 72324 22372
rect 72156 22318 72270 22370
rect 72322 22318 72324 22370
rect 72156 22316 72324 22318
rect 72268 22306 72324 22316
rect 72268 21698 72324 21710
rect 72268 21646 72270 21698
rect 72322 21646 72324 21698
rect 72044 20750 72046 20802
rect 72098 20750 72100 20802
rect 72044 20738 72100 20750
rect 72156 20914 72212 20926
rect 72156 20862 72158 20914
rect 72210 20862 72212 20914
rect 70588 17714 70644 17724
rect 70812 20300 71540 20356
rect 70812 17554 70868 20300
rect 72156 19236 72212 20862
rect 72156 19170 72212 19180
rect 70812 17502 70814 17554
rect 70866 17502 70868 17554
rect 70812 17490 70868 17502
rect 71372 18452 71428 18462
rect 70252 17444 70308 17454
rect 70476 17444 70532 17454
rect 70252 17442 70532 17444
rect 70252 17390 70254 17442
rect 70306 17390 70478 17442
rect 70530 17390 70532 17442
rect 70252 17388 70532 17390
rect 70252 16660 70308 17388
rect 70476 17378 70532 17388
rect 70252 16594 70308 16604
rect 69356 10882 69412 10892
rect 69020 9380 69076 9390
rect 67452 5122 68516 5124
rect 67452 5070 68350 5122
rect 68402 5070 68516 5122
rect 67452 5068 68516 5070
rect 68572 7362 68628 7374
rect 68572 7310 68574 7362
rect 68626 7310 68628 7362
rect 68572 5124 68628 7310
rect 68348 5058 68404 5068
rect 68572 5058 68628 5068
rect 68908 5794 68964 5806
rect 68908 5742 68910 5794
rect 68962 5742 68964 5794
rect 67452 4900 67508 4910
rect 67340 4898 67508 4900
rect 67340 4846 67454 4898
rect 67506 4846 67508 4898
rect 67340 4844 67508 4846
rect 67340 4338 67396 4844
rect 67452 4834 67508 4844
rect 68124 4900 68180 4910
rect 67340 4286 67342 4338
rect 67394 4286 67396 4338
rect 67340 4274 67396 4286
rect 67452 3780 67508 3790
rect 67452 3686 67508 3724
rect 67228 3164 67508 3220
rect 67452 800 67508 3164
rect 68124 800 68180 4844
rect 68348 4116 68404 4126
rect 68348 4022 68404 4060
rect 68796 4116 68852 4126
rect 68796 800 68852 4060
rect 68908 3556 68964 5742
rect 69020 5684 69076 9324
rect 69804 7700 69860 7710
rect 69020 5618 69076 5628
rect 69356 6466 69412 6478
rect 69356 6414 69358 6466
rect 69410 6414 69412 6466
rect 69356 5572 69412 6414
rect 69356 5506 69412 5516
rect 69356 5236 69412 5246
rect 69356 5142 69412 5180
rect 68908 3490 68964 3500
rect 69468 3780 69524 3790
rect 69468 800 69524 3724
rect 69804 3668 69860 7644
rect 71260 6690 71316 6702
rect 71260 6638 71262 6690
rect 71314 6638 71316 6690
rect 70476 6468 70532 6478
rect 70364 6412 70476 6468
rect 69804 3666 70308 3668
rect 69804 3614 69806 3666
rect 69858 3614 70308 3666
rect 69804 3612 70308 3614
rect 69804 3602 69860 3612
rect 70252 3554 70308 3612
rect 70252 3502 70254 3554
rect 70306 3502 70308 3554
rect 70252 3490 70308 3502
rect 70364 980 70420 6412
rect 70476 6402 70532 6412
rect 71036 5908 71092 5918
rect 71260 5908 71316 6638
rect 71092 5852 71316 5908
rect 71036 5814 71092 5852
rect 70476 5794 70532 5806
rect 70476 5742 70478 5794
rect 70530 5742 70532 5794
rect 70476 5572 70532 5742
rect 70476 5506 70532 5516
rect 70812 5684 70868 5694
rect 70476 4340 70532 4350
rect 70476 4226 70532 4284
rect 70476 4174 70478 4226
rect 70530 4174 70532 4226
rect 70476 4004 70532 4174
rect 70476 3938 70532 3948
rect 70140 924 70420 980
rect 70140 800 70196 924
rect 70812 800 70868 5628
rect 71372 5124 71428 18396
rect 72268 17892 72324 21646
rect 72380 20244 72436 22878
rect 72492 22482 72548 22494
rect 72492 22430 72494 22482
rect 72546 22430 72548 22482
rect 72492 22260 72548 22430
rect 72492 22194 72548 22204
rect 72604 21586 72660 26684
rect 72716 26516 72772 26526
rect 72716 25730 72772 26460
rect 72940 26404 72996 27020
rect 73388 27074 73444 27244
rect 73388 27022 73390 27074
rect 73442 27022 73444 27074
rect 73388 27010 73444 27022
rect 73500 27074 73556 27804
rect 73724 27858 73780 28476
rect 73724 27806 73726 27858
rect 73778 27806 73780 27858
rect 73724 27794 73780 27806
rect 73836 28420 73892 28430
rect 73500 27022 73502 27074
rect 73554 27022 73556 27074
rect 73500 27010 73556 27022
rect 73052 26964 73108 26974
rect 73836 26908 73892 28364
rect 73052 26870 73108 26908
rect 73164 26850 73220 26862
rect 73164 26798 73166 26850
rect 73218 26798 73220 26850
rect 72716 25678 72718 25730
rect 72770 25678 72772 25730
rect 72716 25666 72772 25678
rect 72828 26348 72996 26404
rect 73052 26628 73108 26638
rect 72828 23156 72884 26348
rect 72940 26180 72996 26190
rect 72940 26086 72996 26124
rect 73052 24722 73108 26572
rect 73052 24670 73054 24722
rect 73106 24670 73108 24722
rect 73052 24658 73108 24670
rect 72940 23156 72996 23166
rect 72828 23154 72996 23156
rect 72828 23102 72942 23154
rect 72994 23102 72996 23154
rect 72828 23100 72996 23102
rect 72940 23090 72996 23100
rect 72604 21534 72606 21586
rect 72658 21534 72660 21586
rect 72604 21522 72660 21534
rect 73052 21474 73108 21486
rect 73052 21422 73054 21474
rect 73106 21422 73108 21474
rect 72940 20916 72996 20926
rect 72940 20822 72996 20860
rect 72716 20804 72772 20814
rect 72380 20178 72436 20188
rect 72604 20748 72716 20804
rect 72604 20242 72660 20748
rect 72716 20710 72772 20748
rect 72604 20190 72606 20242
rect 72658 20190 72660 20242
rect 72604 20178 72660 20190
rect 73052 19460 73108 21422
rect 73164 20804 73220 26798
rect 73612 26852 73668 26862
rect 73500 26290 73556 26302
rect 73500 26238 73502 26290
rect 73554 26238 73556 26290
rect 73276 26178 73332 26190
rect 73276 26126 73278 26178
rect 73330 26126 73332 26178
rect 73276 26068 73332 26126
rect 73276 26002 73332 26012
rect 73500 26068 73556 26238
rect 73500 26002 73556 26012
rect 73276 25508 73332 25518
rect 73276 25414 73332 25452
rect 73500 24724 73556 24734
rect 73500 24630 73556 24668
rect 73612 24500 73668 26796
rect 73500 24444 73668 24500
rect 73724 26852 73892 26908
rect 73948 27746 74004 27758
rect 73948 27694 73950 27746
rect 74002 27694 74004 27746
rect 73948 26964 74004 27694
rect 73948 26898 74004 26908
rect 73276 23940 73332 23950
rect 73276 23846 73332 23884
rect 73500 23604 73556 24444
rect 73612 23940 73668 23950
rect 73612 23846 73668 23884
rect 73724 23826 73780 26852
rect 74060 26628 74116 29708
rect 74396 29540 74452 29550
rect 74508 29540 74564 30044
rect 74396 29538 74564 29540
rect 74396 29486 74398 29538
rect 74450 29486 74564 29538
rect 74396 29484 74564 29486
rect 74396 29474 74452 29484
rect 74620 29428 74676 29438
rect 74508 29426 74676 29428
rect 74508 29374 74622 29426
rect 74674 29374 74676 29426
rect 74508 29372 74676 29374
rect 74508 28868 74564 29372
rect 74620 29362 74676 29372
rect 74844 29204 74900 30716
rect 74956 30212 75012 30222
rect 74956 30118 75012 30156
rect 74956 29540 75012 29550
rect 74956 29446 75012 29484
rect 74284 28812 74564 28868
rect 74620 29148 74900 29204
rect 74284 28644 74340 28812
rect 74284 28550 74340 28588
rect 74396 28532 74452 28542
rect 74172 27972 74228 27982
rect 74172 27878 74228 27916
rect 74284 27860 74340 27870
rect 74284 26962 74340 27804
rect 74396 27636 74452 28476
rect 74508 28420 74564 28430
rect 74508 28326 74564 28364
rect 74620 28196 74676 29148
rect 75068 29092 75124 32284
rect 75180 31892 75236 33180
rect 75404 32676 75460 34862
rect 75628 34802 75684 35756
rect 76076 35700 76132 35710
rect 75852 35698 76132 35700
rect 75852 35646 76078 35698
rect 76130 35646 76132 35698
rect 75852 35644 76132 35646
rect 75628 34750 75630 34802
rect 75682 34750 75684 34802
rect 75628 34738 75684 34750
rect 75740 35476 75796 35486
rect 75740 34132 75796 35420
rect 75628 34130 75796 34132
rect 75628 34078 75742 34130
rect 75794 34078 75796 34130
rect 75628 34076 75796 34078
rect 75292 32620 75460 32676
rect 75516 34020 75572 34030
rect 75292 32452 75348 32620
rect 75516 32562 75572 33964
rect 75516 32510 75518 32562
rect 75570 32510 75572 32562
rect 75516 32498 75572 32510
rect 75292 32386 75348 32396
rect 75404 32450 75460 32462
rect 75404 32398 75406 32450
rect 75458 32398 75460 32450
rect 75292 31892 75348 31902
rect 75180 31890 75348 31892
rect 75180 31838 75294 31890
rect 75346 31838 75348 31890
rect 75180 31836 75348 31838
rect 75292 31826 75348 31836
rect 75180 31106 75236 31118
rect 75180 31054 75182 31106
rect 75234 31054 75236 31106
rect 75180 30996 75236 31054
rect 75180 30930 75236 30940
rect 75404 30436 75460 32398
rect 75628 31332 75684 34076
rect 75740 34066 75796 34076
rect 75852 33684 75908 35644
rect 76076 35634 76132 35644
rect 76188 34914 76244 36988
rect 76300 36708 76356 36718
rect 76300 36614 76356 36652
rect 76300 36372 76356 36382
rect 76412 36372 76468 37212
rect 76524 37266 76580 37278
rect 76748 37268 76804 37660
rect 76524 37214 76526 37266
rect 76578 37214 76580 37266
rect 76524 37044 76580 37214
rect 76524 36978 76580 36988
rect 76636 37212 76804 37268
rect 76524 36484 76580 36494
rect 76636 36484 76692 37212
rect 76524 36482 76692 36484
rect 76524 36430 76526 36482
rect 76578 36430 76692 36482
rect 76524 36428 76692 36430
rect 76748 37044 76804 37054
rect 76524 36418 76580 36428
rect 76356 36316 76468 36372
rect 76300 36306 76356 36316
rect 76300 35924 76356 35934
rect 76300 35810 76356 35868
rect 76300 35758 76302 35810
rect 76354 35758 76356 35810
rect 76300 35746 76356 35758
rect 76748 35812 76804 36988
rect 76860 36482 76916 38220
rect 77084 36820 77140 38332
rect 77196 38050 77252 38612
rect 77196 37998 77198 38050
rect 77250 37998 77252 38050
rect 77196 37986 77252 37998
rect 77308 38274 77364 38286
rect 77308 38222 77310 38274
rect 77362 38222 77364 38274
rect 77308 37716 77364 38222
rect 77308 37650 77364 37660
rect 77532 38050 77588 38062
rect 77532 37998 77534 38050
rect 77586 37998 77588 38050
rect 77532 37492 77588 37998
rect 77532 37426 77588 37436
rect 77644 37828 77700 37838
rect 77308 37266 77364 37278
rect 77308 37214 77310 37266
rect 77362 37214 77364 37266
rect 77084 36764 77252 36820
rect 76860 36430 76862 36482
rect 76914 36430 76916 36482
rect 76860 36418 76916 36430
rect 77084 36594 77140 36606
rect 77084 36542 77086 36594
rect 77138 36542 77140 36594
rect 76748 35698 76804 35756
rect 76972 36036 77028 36046
rect 76972 35810 77028 35980
rect 76972 35758 76974 35810
rect 77026 35758 77028 35810
rect 76972 35746 77028 35758
rect 76748 35646 76750 35698
rect 76802 35646 76804 35698
rect 76748 35634 76804 35646
rect 76524 35586 76580 35598
rect 76524 35534 76526 35586
rect 76578 35534 76580 35586
rect 76524 35252 76580 35534
rect 76524 35196 76916 35252
rect 76188 34862 76190 34914
rect 76242 34862 76244 34914
rect 76188 34850 76244 34862
rect 76300 35026 76356 35038
rect 76300 34974 76302 35026
rect 76354 34974 76356 35026
rect 76300 34356 76356 34974
rect 76300 34290 76356 34300
rect 76524 35028 76580 35038
rect 75740 31892 75796 31902
rect 75740 31798 75796 31836
rect 75628 31266 75684 31276
rect 75852 31218 75908 33628
rect 75964 34242 76020 34254
rect 75964 34190 75966 34242
rect 76018 34190 76020 34242
rect 75964 32788 76020 34190
rect 76300 34130 76356 34142
rect 76300 34078 76302 34130
rect 76354 34078 76356 34130
rect 76300 33236 76356 34078
rect 76524 34130 76580 34972
rect 76860 34914 76916 35196
rect 76860 34862 76862 34914
rect 76914 34862 76916 34914
rect 76860 34850 76916 34862
rect 77084 34356 77140 36542
rect 77196 35924 77252 36764
rect 77196 35858 77252 35868
rect 77308 35922 77364 37214
rect 77420 37156 77476 37166
rect 77420 37062 77476 37100
rect 77532 37042 77588 37054
rect 77532 36990 77534 37042
rect 77586 36990 77588 37042
rect 77308 35870 77310 35922
rect 77362 35870 77364 35922
rect 77308 35858 77364 35870
rect 77420 36708 77476 36718
rect 77420 36372 77476 36652
rect 77308 35700 77364 35710
rect 77308 35606 77364 35644
rect 77420 35364 77476 36316
rect 77532 36148 77588 36990
rect 77644 36372 77700 37772
rect 77756 36708 77812 39452
rect 77868 39442 77924 39452
rect 78092 39506 78148 39900
rect 78092 39454 78094 39506
rect 78146 39454 78148 39506
rect 78092 39442 78148 39454
rect 77868 39172 77924 39182
rect 77868 37266 77924 39116
rect 77980 39060 78036 39070
rect 78204 39060 78260 39070
rect 78036 39058 78260 39060
rect 78036 39006 78206 39058
rect 78258 39006 78260 39058
rect 78036 39004 78260 39006
rect 77980 38994 78036 39004
rect 78204 38994 78260 39004
rect 78204 38836 78260 38846
rect 78092 38780 78204 38836
rect 77868 37214 77870 37266
rect 77922 37214 77924 37266
rect 77868 37202 77924 37214
rect 77980 38162 78036 38174
rect 77980 38110 77982 38162
rect 78034 38110 78036 38162
rect 77756 36642 77812 36652
rect 77868 36372 77924 36382
rect 77644 36370 77924 36372
rect 77644 36318 77870 36370
rect 77922 36318 77924 36370
rect 77644 36316 77924 36318
rect 77868 36306 77924 36316
rect 77532 36082 77588 36092
rect 77980 35922 78036 38110
rect 78092 36372 78148 38780
rect 78204 38770 78260 38780
rect 78428 37380 78484 37390
rect 78204 36372 78260 36382
rect 78092 36370 78372 36372
rect 78092 36318 78206 36370
rect 78258 36318 78372 36370
rect 78092 36316 78372 36318
rect 78204 36306 78260 36316
rect 77980 35870 77982 35922
rect 78034 35870 78036 35922
rect 77980 35858 78036 35870
rect 77532 35812 77588 35822
rect 77532 35718 77588 35756
rect 78092 35810 78148 35822
rect 78092 35758 78094 35810
rect 78146 35758 78148 35810
rect 77868 35474 77924 35486
rect 77868 35422 77870 35474
rect 77922 35422 77924 35474
rect 77868 35364 77924 35422
rect 77420 35308 77924 35364
rect 76524 34078 76526 34130
rect 76578 34078 76580 34130
rect 76524 34066 76580 34078
rect 76748 34300 77140 34356
rect 77196 35026 77252 35038
rect 77196 34974 77198 35026
rect 77250 34974 77252 35026
rect 76412 34020 76468 34030
rect 76412 33926 76468 33964
rect 76748 33572 76804 34300
rect 76860 34130 76916 34142
rect 77084 34132 77140 34142
rect 76860 34078 76862 34130
rect 76914 34078 76916 34130
rect 76860 33684 76916 34078
rect 76860 33618 76916 33628
rect 76972 34130 77140 34132
rect 76972 34078 77086 34130
rect 77138 34078 77140 34130
rect 76972 34076 77140 34078
rect 76748 33506 76804 33516
rect 76860 33460 76916 33470
rect 76860 33346 76916 33404
rect 76860 33294 76862 33346
rect 76914 33294 76916 33346
rect 76524 33236 76580 33246
rect 76300 33234 76580 33236
rect 76300 33182 76526 33234
rect 76578 33182 76580 33234
rect 76300 33180 76580 33182
rect 75964 32722 76020 32732
rect 76524 32676 76580 33180
rect 76636 33124 76692 33134
rect 76636 33030 76692 33068
rect 76860 33124 76916 33294
rect 76860 33058 76916 33068
rect 76748 32676 76804 32686
rect 76972 32676 77028 34076
rect 77084 34066 77140 34076
rect 77084 33684 77140 33694
rect 77084 33346 77140 33628
rect 77084 33294 77086 33346
rect 77138 33294 77140 33346
rect 77084 33282 77140 33294
rect 77196 32900 77252 34974
rect 77308 34018 77364 34030
rect 77308 33966 77310 34018
rect 77362 33966 77364 34018
rect 77308 33348 77364 33966
rect 77308 33282 77364 33292
rect 77420 33234 77476 35308
rect 77868 35140 77924 35150
rect 77868 34914 77924 35084
rect 77868 34862 77870 34914
rect 77922 34862 77924 34914
rect 77868 34850 77924 34862
rect 78092 34804 78148 35758
rect 78204 34804 78260 34814
rect 78092 34802 78260 34804
rect 78092 34750 78206 34802
rect 78258 34750 78260 34802
rect 78092 34748 78260 34750
rect 78204 34738 78260 34748
rect 77532 34580 77588 34590
rect 77532 34244 77588 34524
rect 78204 34580 78260 34590
rect 78204 34354 78260 34524
rect 78204 34302 78206 34354
rect 78258 34302 78260 34354
rect 78204 34290 78260 34302
rect 77532 34150 77588 34188
rect 77644 34130 77700 34142
rect 77644 34078 77646 34130
rect 77698 34078 77700 34130
rect 77644 33684 77700 34078
rect 77980 34132 78036 34142
rect 78036 34076 78148 34132
rect 77980 34066 78036 34076
rect 77868 33908 77924 33918
rect 77924 33852 78036 33908
rect 77868 33842 77924 33852
rect 77644 33618 77700 33628
rect 77756 33796 77812 33806
rect 77756 33346 77812 33740
rect 77756 33294 77758 33346
rect 77810 33294 77812 33346
rect 77756 33282 77812 33294
rect 77868 33572 77924 33582
rect 77420 33182 77422 33234
rect 77474 33182 77476 33234
rect 77420 33170 77476 33182
rect 77196 32844 77700 32900
rect 76524 32674 77028 32676
rect 76524 32622 76750 32674
rect 76802 32622 77028 32674
rect 76524 32620 77028 32622
rect 77532 32676 77588 32686
rect 76412 32562 76468 32574
rect 76412 32510 76414 32562
rect 76466 32510 76468 32562
rect 76412 32452 76468 32510
rect 76412 32386 76468 32396
rect 76524 31780 76580 31790
rect 76748 31780 76804 32620
rect 77308 32562 77364 32574
rect 77308 32510 77310 32562
rect 77362 32510 77364 32562
rect 77308 32452 77364 32510
rect 77420 32452 77476 32462
rect 77308 32396 77420 32452
rect 77420 32386 77476 32396
rect 77308 32116 77364 32126
rect 76524 31778 76804 31780
rect 76524 31726 76526 31778
rect 76578 31726 76804 31778
rect 76524 31724 76804 31726
rect 76860 31780 76916 31790
rect 76524 31714 76580 31724
rect 76860 31686 76916 31724
rect 77084 31666 77140 31678
rect 77084 31614 77086 31666
rect 77138 31614 77140 31666
rect 76636 31556 76692 31566
rect 76636 31462 76692 31500
rect 75852 31166 75854 31218
rect 75906 31166 75908 31218
rect 75852 31154 75908 31166
rect 76188 31164 76916 31220
rect 75516 31108 75572 31118
rect 75516 31014 75572 31052
rect 76188 31106 76244 31164
rect 76188 31054 76190 31106
rect 76242 31054 76244 31106
rect 76188 31042 76244 31054
rect 75404 30370 75460 30380
rect 76300 30882 76356 30894
rect 76300 30830 76302 30882
rect 76354 30830 76356 30882
rect 76300 30324 76356 30830
rect 76188 30268 76356 30324
rect 75180 30212 75236 30222
rect 76188 30212 76244 30268
rect 76412 30212 76468 31164
rect 75180 30210 75348 30212
rect 75180 30158 75182 30210
rect 75234 30158 75348 30210
rect 75180 30156 75348 30158
rect 75180 30146 75236 30156
rect 74844 29036 75124 29092
rect 74396 27570 74452 27580
rect 74508 28140 74676 28196
rect 74732 28644 74788 28654
rect 74284 26910 74286 26962
rect 74338 26910 74340 26962
rect 74284 26898 74340 26910
rect 74396 26740 74452 26750
rect 74060 26572 74340 26628
rect 73836 26292 73892 26302
rect 73836 26068 73892 26236
rect 74284 26290 74340 26572
rect 74284 26238 74286 26290
rect 74338 26238 74340 26290
rect 74284 26226 74340 26238
rect 73836 26002 73892 26012
rect 74060 26068 74116 26078
rect 74060 25974 74116 26012
rect 74172 25732 74228 25742
rect 73724 23774 73726 23826
rect 73778 23774 73780 23826
rect 73724 23762 73780 23774
rect 73836 25506 73892 25518
rect 73836 25454 73838 25506
rect 73890 25454 73892 25506
rect 73276 23548 73556 23604
rect 73276 22370 73332 23548
rect 73836 23380 73892 25454
rect 74172 25506 74228 25676
rect 74396 25730 74452 26684
rect 74396 25678 74398 25730
rect 74450 25678 74452 25730
rect 74396 25666 74452 25678
rect 74172 25454 74174 25506
rect 74226 25454 74228 25506
rect 74172 24946 74228 25454
rect 74172 24894 74174 24946
rect 74226 24894 74228 24946
rect 74172 24882 74228 24894
rect 74284 25620 74340 25630
rect 74284 24050 74340 25564
rect 74284 23998 74286 24050
rect 74338 23998 74340 24050
rect 73836 23314 73892 23324
rect 74172 23828 74228 23838
rect 73276 22318 73278 22370
rect 73330 22318 73332 22370
rect 73276 22306 73332 22318
rect 73500 23154 73556 23166
rect 73500 23102 73502 23154
rect 73554 23102 73556 23154
rect 73500 22148 73556 23102
rect 74172 22594 74228 23772
rect 74172 22542 74174 22594
rect 74226 22542 74228 22594
rect 74172 22530 74228 22542
rect 73500 22082 73556 22092
rect 73612 22370 73668 22382
rect 73612 22318 73614 22370
rect 73666 22318 73668 22370
rect 73612 22036 73668 22318
rect 73948 22372 74004 22382
rect 73948 22278 74004 22316
rect 73612 21970 73668 21980
rect 73276 21588 73332 21598
rect 73276 21494 73332 21532
rect 74060 21588 74116 21598
rect 74060 21494 74116 21532
rect 74284 21588 74340 23998
rect 74396 24276 74452 24286
rect 74396 23378 74452 24220
rect 74396 23326 74398 23378
rect 74450 23326 74452 23378
rect 74396 23314 74452 23326
rect 74508 23154 74564 28140
rect 74732 28084 74788 28588
rect 74620 28028 74788 28084
rect 74620 27524 74676 28028
rect 74732 27860 74788 27870
rect 74732 27766 74788 27804
rect 74844 27636 74900 29036
rect 75068 28530 75124 28542
rect 75068 28478 75070 28530
rect 75122 28478 75124 28530
rect 75068 28420 75124 28478
rect 75180 28532 75236 28542
rect 75180 28438 75236 28476
rect 74956 27972 75012 27982
rect 75068 27972 75124 28364
rect 75292 28420 75348 30156
rect 76188 30146 76244 30156
rect 76300 30156 76468 30212
rect 76524 30994 76580 31006
rect 76524 30942 76526 30994
rect 76578 30942 76580 30994
rect 76524 30884 76580 30942
rect 76636 30996 76692 31006
rect 76860 30996 76916 31164
rect 76972 30996 77028 31006
rect 76692 30940 76804 30996
rect 76860 30994 77028 30996
rect 76860 30942 76974 30994
rect 77026 30942 77028 30994
rect 76860 30940 77028 30942
rect 76636 30902 76692 30940
rect 76300 30098 76356 30156
rect 76300 30046 76302 30098
rect 76354 30046 76356 30098
rect 75516 29538 75572 29550
rect 75516 29486 75518 29538
rect 75570 29486 75572 29538
rect 75404 29316 75460 29326
rect 75404 29222 75460 29260
rect 75404 28980 75460 28990
rect 75404 28642 75460 28924
rect 75404 28590 75406 28642
rect 75458 28590 75460 28642
rect 75404 28578 75460 28590
rect 75292 28354 75348 28364
rect 75404 27972 75460 27982
rect 75068 27916 75404 27972
rect 74956 27878 75012 27916
rect 75292 27858 75348 27916
rect 75404 27906 75460 27916
rect 75292 27806 75294 27858
rect 75346 27806 75348 27858
rect 75292 27794 75348 27806
rect 75180 27746 75236 27758
rect 75180 27694 75182 27746
rect 75234 27694 75236 27746
rect 74844 27580 75124 27636
rect 74620 27468 75012 27524
rect 74620 26964 74676 26974
rect 74620 26870 74676 26908
rect 74844 26290 74900 26302
rect 74844 26238 74846 26290
rect 74898 26238 74900 26290
rect 74844 25396 74900 26238
rect 74956 25506 75012 27468
rect 75068 27188 75124 27580
rect 75068 27122 75124 27132
rect 75180 26908 75236 27694
rect 75404 27748 75460 27758
rect 75404 27186 75460 27692
rect 75516 27412 75572 29486
rect 76076 29540 76132 29550
rect 76300 29540 76356 30046
rect 76524 30100 76580 30828
rect 76748 30772 76804 30940
rect 76972 30930 77028 30940
rect 77084 30772 77140 31614
rect 76748 30716 77140 30772
rect 77196 30882 77252 30894
rect 77196 30830 77198 30882
rect 77250 30830 77252 30882
rect 76636 30212 76692 30222
rect 76636 30118 76692 30156
rect 76748 30210 76804 30716
rect 76748 30158 76750 30210
rect 76802 30158 76804 30210
rect 76748 30146 76804 30158
rect 76972 30212 77028 30222
rect 77028 30156 77140 30212
rect 76972 30146 77028 30156
rect 76524 30034 76580 30044
rect 76412 29986 76468 29998
rect 76412 29934 76414 29986
rect 76466 29934 76468 29986
rect 76412 29876 76468 29934
rect 76412 29810 76468 29820
rect 76132 29484 76356 29540
rect 76524 29540 76580 29550
rect 76076 29446 76132 29484
rect 76412 29428 76468 29438
rect 76524 29428 76580 29484
rect 76412 29426 76580 29428
rect 76412 29374 76414 29426
rect 76466 29374 76580 29426
rect 76412 29372 76580 29374
rect 76636 29426 76692 29438
rect 76636 29374 76638 29426
rect 76690 29374 76692 29426
rect 76412 29362 76468 29372
rect 76188 29316 76244 29326
rect 76188 29222 76244 29260
rect 75740 29204 75796 29214
rect 75740 29110 75796 29148
rect 76524 28980 76580 28990
rect 75628 28644 75684 28654
rect 75628 28550 75684 28588
rect 76524 28642 76580 28924
rect 76524 28590 76526 28642
rect 76578 28590 76580 28642
rect 76524 28578 76580 28590
rect 76636 28644 76692 29374
rect 76860 29204 76916 29214
rect 76692 28588 76804 28644
rect 76636 28550 76692 28588
rect 75852 28532 75908 28542
rect 75516 27346 75572 27356
rect 75628 28420 75684 28430
rect 75628 27300 75684 28364
rect 75852 27972 75908 28476
rect 76188 28532 76244 28542
rect 76188 28438 76244 28476
rect 76300 28418 76356 28430
rect 76300 28366 76302 28418
rect 76354 28366 76356 28418
rect 75964 28084 76020 28094
rect 75964 27990 76020 28028
rect 75852 27878 75908 27916
rect 76188 27972 76244 27982
rect 76188 27878 76244 27916
rect 75628 27234 75684 27244
rect 75964 27748 76020 27758
rect 75404 27134 75406 27186
rect 75458 27134 75460 27186
rect 75404 27122 75460 27134
rect 75516 27188 75572 27198
rect 74956 25454 74958 25506
rect 75010 25454 75012 25506
rect 74956 25442 75012 25454
rect 75068 26852 75236 26908
rect 75292 27074 75348 27086
rect 75292 27022 75294 27074
rect 75346 27022 75348 27074
rect 74844 25330 74900 25340
rect 75068 25172 75124 26852
rect 74844 25116 75124 25172
rect 74620 24722 74676 24734
rect 74620 24670 74622 24722
rect 74674 24670 74676 24722
rect 74620 24276 74676 24670
rect 74620 24210 74676 24220
rect 74732 24164 74788 24174
rect 74732 23940 74788 24108
rect 74844 24052 74900 25116
rect 74956 24948 75012 24958
rect 75292 24948 75348 27022
rect 75516 26908 75572 27132
rect 75404 26852 75572 26908
rect 75628 26962 75684 26974
rect 75628 26910 75630 26962
rect 75682 26910 75684 26962
rect 75404 26290 75460 26852
rect 75628 26740 75684 26910
rect 75964 26964 76020 27692
rect 76300 27636 76356 28366
rect 76748 28084 76804 28588
rect 76412 28082 76804 28084
rect 76412 28030 76750 28082
rect 76802 28030 76804 28082
rect 76412 28028 76804 28030
rect 76412 27970 76468 28028
rect 76748 28018 76804 28028
rect 76412 27918 76414 27970
rect 76466 27918 76468 27970
rect 76412 27906 76468 27918
rect 75964 26898 76020 26908
rect 76076 27580 76356 27636
rect 76636 27860 76692 27870
rect 75628 26674 75684 26684
rect 75628 26404 75684 26414
rect 75628 26402 75796 26404
rect 75628 26350 75630 26402
rect 75682 26350 75796 26402
rect 75628 26348 75796 26350
rect 75628 26338 75684 26348
rect 75404 26238 75406 26290
rect 75458 26238 75460 26290
rect 75404 26226 75460 26238
rect 75516 25508 75572 25518
rect 75516 25414 75572 25452
rect 74956 24946 75348 24948
rect 74956 24894 74958 24946
rect 75010 24894 75348 24946
rect 74956 24892 75348 24894
rect 75404 25396 75460 25406
rect 75404 24946 75460 25340
rect 75404 24894 75406 24946
rect 75458 24894 75460 24946
rect 74956 24882 75012 24892
rect 75404 24882 75460 24894
rect 75628 24722 75684 24734
rect 75628 24670 75630 24722
rect 75682 24670 75684 24722
rect 75292 24498 75348 24510
rect 75292 24446 75294 24498
rect 75346 24446 75348 24498
rect 75292 24164 75348 24446
rect 75292 24070 75348 24108
rect 74844 23996 75124 24052
rect 74732 23884 75012 23940
rect 74620 23828 74676 23838
rect 74620 23734 74676 23772
rect 74956 23826 75012 23884
rect 74956 23774 74958 23826
rect 75010 23774 75012 23826
rect 74956 23762 75012 23774
rect 74844 23716 74900 23726
rect 74844 23492 74900 23660
rect 75068 23604 75124 23996
rect 75404 23940 75460 23950
rect 75404 23846 75460 23884
rect 74508 23102 74510 23154
rect 74562 23102 74564 23154
rect 74508 23090 74564 23102
rect 74620 23436 74900 23492
rect 74956 23548 75124 23604
rect 75516 23714 75572 23726
rect 75516 23662 75518 23714
rect 75570 23662 75572 23714
rect 74620 21810 74676 23436
rect 74844 23154 74900 23166
rect 74844 23102 74846 23154
rect 74898 23102 74900 23154
rect 74844 23042 74900 23102
rect 74844 22990 74846 23042
rect 74898 22990 74900 23042
rect 74844 22148 74900 22990
rect 74956 22370 75012 23548
rect 75068 22932 75124 22942
rect 75068 22838 75124 22876
rect 74956 22318 74958 22370
rect 75010 22318 75012 22370
rect 74956 22306 75012 22318
rect 75068 22482 75124 22494
rect 75068 22430 75070 22482
rect 75122 22430 75124 22482
rect 74620 21758 74622 21810
rect 74674 21758 74676 21810
rect 74620 21746 74676 21758
rect 74732 22092 74900 22148
rect 74284 21028 74340 21532
rect 74284 20962 74340 20972
rect 73836 20914 73892 20926
rect 73836 20862 73838 20914
rect 73890 20862 73892 20914
rect 73500 20804 73556 20814
rect 73164 20802 73556 20804
rect 73164 20750 73502 20802
rect 73554 20750 73556 20802
rect 73164 20748 73556 20750
rect 73500 20738 73556 20748
rect 73836 20132 73892 20862
rect 74732 20914 74788 22092
rect 74956 21924 75012 21934
rect 74732 20862 74734 20914
rect 74786 20862 74788 20914
rect 74732 20850 74788 20862
rect 74844 21586 74900 21598
rect 74844 21534 74846 21586
rect 74898 21534 74900 21586
rect 74844 20916 74900 21534
rect 74844 20692 74900 20860
rect 74620 20636 74900 20692
rect 74620 20242 74676 20636
rect 74620 20190 74622 20242
rect 74674 20190 74676 20242
rect 74620 20178 74676 20190
rect 73836 20066 73892 20076
rect 73052 19394 73108 19404
rect 72268 17826 72324 17836
rect 74956 15148 75012 21868
rect 75068 20580 75124 22430
rect 75516 21924 75572 23662
rect 75628 22260 75684 24670
rect 75740 22372 75796 26348
rect 75964 26290 76020 26302
rect 75964 26238 75966 26290
rect 76018 26238 76020 26290
rect 75964 25620 76020 26238
rect 75964 25554 76020 25564
rect 76076 25060 76132 27580
rect 76188 27300 76244 27310
rect 76188 27206 76244 27244
rect 76524 26962 76580 26974
rect 76524 26910 76526 26962
rect 76578 26910 76580 26962
rect 76300 26852 76356 26862
rect 76300 26850 76468 26852
rect 76300 26798 76302 26850
rect 76354 26798 76468 26850
rect 76300 26796 76468 26798
rect 76300 26786 76356 26796
rect 76300 26404 76356 26414
rect 76300 26310 76356 26348
rect 75964 25004 76132 25060
rect 76188 25508 76244 25518
rect 75964 23154 76020 25004
rect 76188 24946 76244 25452
rect 76412 25394 76468 26796
rect 76524 26740 76580 26910
rect 76524 26674 76580 26684
rect 76412 25342 76414 25394
rect 76466 25342 76468 25394
rect 76412 25330 76468 25342
rect 76188 24894 76190 24946
rect 76242 24894 76244 24946
rect 76188 24882 76244 24894
rect 76076 24834 76132 24846
rect 76076 24782 76078 24834
rect 76130 24782 76132 24834
rect 76076 24612 76132 24782
rect 76076 23940 76132 24556
rect 76524 24724 76580 24734
rect 76300 24498 76356 24510
rect 76300 24446 76302 24498
rect 76354 24446 76356 24498
rect 76188 24164 76244 24174
rect 76300 24164 76356 24446
rect 76244 24108 76356 24164
rect 76524 24162 76580 24668
rect 76524 24110 76526 24162
rect 76578 24110 76580 24162
rect 76188 24070 76244 24108
rect 76524 24098 76580 24110
rect 76076 23874 76132 23884
rect 76524 23828 76580 23838
rect 76412 23716 76468 23726
rect 75964 23102 75966 23154
rect 76018 23102 76020 23154
rect 75964 23090 76020 23102
rect 76076 23714 76468 23716
rect 76076 23662 76414 23714
rect 76466 23662 76468 23714
rect 76076 23660 76468 23662
rect 75740 22306 75796 22316
rect 75628 22194 75684 22204
rect 75964 22260 76020 22270
rect 75852 21924 75908 21934
rect 75516 21868 75684 21924
rect 75180 21700 75236 21710
rect 75180 21606 75236 21644
rect 75516 21588 75572 21598
rect 75292 21476 75348 21486
rect 75292 21026 75348 21420
rect 75292 20974 75294 21026
rect 75346 20974 75348 21026
rect 75292 20962 75348 20974
rect 75516 20804 75572 21532
rect 75628 21252 75684 21868
rect 75852 21810 75908 21868
rect 75852 21758 75854 21810
rect 75906 21758 75908 21810
rect 75852 21746 75908 21758
rect 75628 21196 75908 21252
rect 75068 20514 75124 20524
rect 75180 20748 75572 20804
rect 75180 20130 75236 20748
rect 75628 20690 75684 20702
rect 75628 20638 75630 20690
rect 75682 20638 75684 20690
rect 75180 20078 75182 20130
rect 75234 20078 75236 20130
rect 75180 20066 75236 20078
rect 75404 20578 75460 20590
rect 75404 20526 75406 20578
rect 75458 20526 75460 20578
rect 75404 15988 75460 20526
rect 75628 20020 75684 20638
rect 75628 19954 75684 19964
rect 75852 19348 75908 21196
rect 75852 19282 75908 19292
rect 75964 20356 76020 22204
rect 76076 21924 76132 23660
rect 76412 23650 76468 23660
rect 76188 23154 76244 23166
rect 76188 23102 76190 23154
rect 76242 23102 76244 23154
rect 76188 22148 76244 23102
rect 76412 22930 76468 22942
rect 76412 22878 76414 22930
rect 76466 22878 76468 22930
rect 76412 22484 76468 22878
rect 76524 22708 76580 23772
rect 76636 22930 76692 27804
rect 76860 27300 76916 29148
rect 76860 27206 76916 27244
rect 76972 28196 77028 28206
rect 76972 27186 77028 28140
rect 77084 28084 77140 30156
rect 77196 29988 77252 30830
rect 77308 30772 77364 32060
rect 77532 32002 77588 32620
rect 77532 31950 77534 32002
rect 77586 31950 77588 32002
rect 77420 31892 77476 31902
rect 77420 31108 77476 31836
rect 77420 31014 77476 31052
rect 77308 30716 77476 30772
rect 77196 29922 77252 29932
rect 77308 30324 77364 30334
rect 77196 29204 77252 29214
rect 77196 28866 77252 29148
rect 77196 28814 77198 28866
rect 77250 28814 77252 28866
rect 77196 28802 77252 28814
rect 77308 28754 77364 30268
rect 77420 29314 77476 30716
rect 77532 30434 77588 31950
rect 77644 31890 77700 32844
rect 77756 32788 77812 32798
rect 77756 32694 77812 32732
rect 77644 31838 77646 31890
rect 77698 31838 77700 31890
rect 77644 31826 77700 31838
rect 77756 32564 77812 32574
rect 77644 30996 77700 31006
rect 77644 30902 77700 30940
rect 77532 30382 77534 30434
rect 77586 30382 77588 30434
rect 77532 30370 77588 30382
rect 77644 30436 77700 30446
rect 77644 30322 77700 30380
rect 77644 30270 77646 30322
rect 77698 30270 77700 30322
rect 77644 30258 77700 30270
rect 77756 29652 77812 32508
rect 77868 32450 77924 33516
rect 77868 32398 77870 32450
rect 77922 32398 77924 32450
rect 77868 32386 77924 32398
rect 77868 31780 77924 31790
rect 77980 31780 78036 33852
rect 77868 31778 78036 31780
rect 77868 31726 77870 31778
rect 77922 31726 78036 31778
rect 77868 31724 78036 31726
rect 77868 31714 77924 31724
rect 78092 31556 78148 34076
rect 78316 33458 78372 36316
rect 78316 33406 78318 33458
rect 78370 33406 78372 33458
rect 78316 33394 78372 33406
rect 78428 32452 78484 37324
rect 78540 37268 78596 37278
rect 78540 34580 78596 37212
rect 78652 37156 78708 40124
rect 78764 37380 78820 40236
rect 78764 37314 78820 37324
rect 78652 37100 78820 37156
rect 78540 34514 78596 34524
rect 78652 35700 78708 35710
rect 78428 32386 78484 32396
rect 77868 31500 78148 31556
rect 78204 32116 78260 32126
rect 77868 30210 77924 31500
rect 77868 30158 77870 30210
rect 77922 30158 77924 30210
rect 77868 30146 77924 30158
rect 77980 31332 78036 31342
rect 77868 29652 77924 29662
rect 77756 29650 77924 29652
rect 77756 29598 77870 29650
rect 77922 29598 77924 29650
rect 77756 29596 77924 29598
rect 77868 29586 77924 29596
rect 77532 29428 77588 29438
rect 77532 29426 77812 29428
rect 77532 29374 77534 29426
rect 77586 29374 77812 29426
rect 77532 29372 77812 29374
rect 77532 29362 77588 29372
rect 77420 29262 77422 29314
rect 77474 29262 77476 29314
rect 77420 29250 77476 29262
rect 77756 28980 77812 29372
rect 77756 28924 77924 28980
rect 77308 28702 77310 28754
rect 77362 28702 77364 28754
rect 77308 28690 77364 28702
rect 77532 28644 77588 28654
rect 77532 28642 77812 28644
rect 77532 28590 77534 28642
rect 77586 28590 77812 28642
rect 77532 28588 77812 28590
rect 77532 28578 77588 28588
rect 77756 28084 77812 28588
rect 77868 28530 77924 28924
rect 77868 28478 77870 28530
rect 77922 28478 77924 28530
rect 77868 28466 77924 28478
rect 77868 28084 77924 28094
rect 77084 28028 77252 28084
rect 77756 28082 77924 28084
rect 77756 28030 77870 28082
rect 77922 28030 77924 28082
rect 77756 28028 77924 28030
rect 77084 27858 77140 27870
rect 77084 27806 77086 27858
rect 77138 27806 77140 27858
rect 77084 27748 77140 27806
rect 77084 27682 77140 27692
rect 77196 27300 77252 28028
rect 77868 28018 77924 28028
rect 77644 27860 77700 27870
rect 77980 27860 78036 31276
rect 78092 31108 78148 31118
rect 78204 31108 78260 32060
rect 78148 31052 78260 31108
rect 78092 29540 78148 31052
rect 78204 30884 78260 30894
rect 78652 30884 78708 35644
rect 78764 34020 78820 37100
rect 78876 35364 78932 40348
rect 78876 35298 78932 35308
rect 78988 34244 79044 43652
rect 78988 34178 79044 34188
rect 78764 33964 78932 34020
rect 78204 30882 78708 30884
rect 78204 30830 78206 30882
rect 78258 30830 78708 30882
rect 78204 30828 78708 30830
rect 78764 33796 78820 33806
rect 78204 30818 78260 30828
rect 78316 30660 78372 30670
rect 78204 29540 78260 29550
rect 78092 29538 78260 29540
rect 78092 29486 78206 29538
rect 78258 29486 78260 29538
rect 78092 29484 78260 29486
rect 78204 29474 78260 29484
rect 78316 29092 78372 30604
rect 78204 28644 78260 28654
rect 78316 28644 78372 29036
rect 78540 29876 78596 29886
rect 78204 28642 78372 28644
rect 78204 28590 78206 28642
rect 78258 28590 78372 28642
rect 78204 28588 78372 28590
rect 78428 28756 78484 28766
rect 78204 28578 78260 28588
rect 78204 27972 78260 27982
rect 78204 27878 78260 27916
rect 77644 27858 78036 27860
rect 77644 27806 77646 27858
rect 77698 27806 78036 27858
rect 77644 27804 78036 27806
rect 77644 27794 77700 27804
rect 77756 27636 77812 27646
rect 76972 27134 76974 27186
rect 77026 27134 77028 27186
rect 76972 27122 77028 27134
rect 77084 27244 77252 27300
rect 77532 27300 77588 27310
rect 77084 26908 77140 27244
rect 76972 26852 77140 26908
rect 77196 27074 77252 27086
rect 77196 27022 77198 27074
rect 77250 27022 77252 27074
rect 76748 26516 76804 26526
rect 76748 25506 76804 26460
rect 76972 26514 77028 26852
rect 76972 26462 76974 26514
rect 77026 26462 77028 26514
rect 76972 26450 77028 26462
rect 77084 26740 77140 26750
rect 76748 25454 76750 25506
rect 76802 25454 76804 25506
rect 76748 25442 76804 25454
rect 77084 25732 77140 26684
rect 77196 26514 77252 27022
rect 77532 26962 77588 27244
rect 77532 26910 77534 26962
rect 77586 26910 77588 26962
rect 77532 26898 77588 26910
rect 77756 27076 77812 27580
rect 77196 26462 77198 26514
rect 77250 26462 77252 26514
rect 77196 26450 77252 26462
rect 77084 25394 77140 25676
rect 77420 26404 77476 26414
rect 77420 26180 77476 26348
rect 77532 26404 77588 26414
rect 77756 26404 77812 27020
rect 77868 26962 77924 26974
rect 77868 26910 77870 26962
rect 77922 26910 77924 26962
rect 77868 26908 77924 26910
rect 78428 26908 78484 28700
rect 78540 27972 78596 29820
rect 78540 27906 78596 27916
rect 78764 26908 78820 33740
rect 78876 31892 78932 33964
rect 78876 31826 78932 31836
rect 77868 26852 78148 26908
rect 77868 26740 77924 26750
rect 77868 26514 77924 26684
rect 77868 26462 77870 26514
rect 77922 26462 77924 26514
rect 77868 26450 77924 26462
rect 77532 26402 77812 26404
rect 77532 26350 77534 26402
rect 77586 26350 77812 26402
rect 77532 26348 77812 26350
rect 77532 26338 77588 26348
rect 77980 26180 78036 26852
rect 78092 26786 78148 26796
rect 78204 26852 78484 26908
rect 78540 26852 78820 26908
rect 77420 26124 78036 26180
rect 78092 26292 78148 26302
rect 77420 25506 77476 26124
rect 77756 25732 77812 25742
rect 77420 25454 77422 25506
rect 77474 25454 77476 25506
rect 77420 25442 77476 25454
rect 77532 25676 77756 25732
rect 77084 25342 77086 25394
rect 77138 25342 77140 25394
rect 77084 25330 77140 25342
rect 77196 25172 77252 25182
rect 77084 24836 77140 24846
rect 76636 22878 76638 22930
rect 76690 22878 76692 22930
rect 76636 22866 76692 22878
rect 76748 24834 77140 24836
rect 76748 24782 77086 24834
rect 77138 24782 77140 24834
rect 76748 24780 77140 24782
rect 76524 22652 76692 22708
rect 76524 22484 76580 22494
rect 76412 22482 76580 22484
rect 76412 22430 76526 22482
rect 76578 22430 76580 22482
rect 76412 22428 76580 22430
rect 76524 22418 76580 22428
rect 76636 22260 76692 22652
rect 76748 22484 76804 24780
rect 77084 24770 77140 24780
rect 77196 24610 77252 25116
rect 77532 24834 77588 25676
rect 77756 25638 77812 25676
rect 78092 25730 78148 26236
rect 78204 26290 78260 26852
rect 78540 26786 78596 26796
rect 78204 26238 78206 26290
rect 78258 26238 78260 26290
rect 78204 26180 78260 26238
rect 78204 26114 78260 26124
rect 78764 26516 78820 26526
rect 78092 25678 78094 25730
rect 78146 25678 78148 25730
rect 78092 25666 78148 25678
rect 78204 25396 78260 25406
rect 77644 25284 77700 25294
rect 77644 24946 77700 25228
rect 77644 24894 77646 24946
rect 77698 24894 77700 24946
rect 77644 24882 77700 24894
rect 77980 25282 78036 25294
rect 77980 25230 77982 25282
rect 78034 25230 78036 25282
rect 77532 24782 77534 24834
rect 77586 24782 77588 24834
rect 77532 24770 77588 24782
rect 77756 24834 77812 24846
rect 77756 24782 77758 24834
rect 77810 24782 77812 24834
rect 77196 24558 77198 24610
rect 77250 24558 77252 24610
rect 77196 24546 77252 24558
rect 76860 24500 76916 24510
rect 76860 24498 77140 24500
rect 76860 24446 76862 24498
rect 76914 24446 77140 24498
rect 76860 24444 77140 24446
rect 76860 24434 76916 24444
rect 76860 23828 76916 23838
rect 77084 23828 77140 24444
rect 77196 23828 77252 23838
rect 76860 23734 76916 23772
rect 76972 23826 77252 23828
rect 76972 23774 77198 23826
rect 77250 23774 77252 23826
rect 76972 23772 77252 23774
rect 77756 23828 77812 24782
rect 77868 23828 77924 23838
rect 77756 23826 77924 23828
rect 77756 23774 77870 23826
rect 77922 23774 77924 23826
rect 77756 23772 77924 23774
rect 76972 23380 77028 23772
rect 77196 23492 77252 23772
rect 77868 23762 77924 23772
rect 77196 23436 77588 23492
rect 76860 23324 77028 23380
rect 76860 23266 76916 23324
rect 76860 23214 76862 23266
rect 76914 23214 76916 23266
rect 76860 23202 76916 23214
rect 77084 23266 77140 23278
rect 77084 23214 77086 23266
rect 77138 23214 77140 23266
rect 76748 22418 76804 22428
rect 77084 22372 77140 23214
rect 77196 23268 77252 23278
rect 77196 23042 77252 23212
rect 77196 22990 77198 23042
rect 77250 22990 77252 23042
rect 77196 22978 77252 22990
rect 77532 23266 77588 23436
rect 77868 23380 77924 23390
rect 77756 23268 77812 23278
rect 77532 23214 77534 23266
rect 77586 23214 77588 23266
rect 77532 22594 77588 23214
rect 77532 22542 77534 22594
rect 77586 22542 77588 22594
rect 77532 22530 77588 22542
rect 77644 23266 77812 23268
rect 77644 23214 77758 23266
rect 77810 23214 77812 23266
rect 77644 23212 77812 23214
rect 77644 22372 77700 23212
rect 77756 23202 77812 23212
rect 77868 23042 77924 23324
rect 77868 22990 77870 23042
rect 77922 22990 77924 23042
rect 77868 22978 77924 22990
rect 77980 22820 78036 25230
rect 78204 23826 78260 25340
rect 78204 23774 78206 23826
rect 78258 23774 78260 23826
rect 78204 23716 78260 23774
rect 78204 23650 78260 23660
rect 78316 23940 78372 23950
rect 77084 22306 77140 22316
rect 77532 22316 77700 22372
rect 77756 22764 78036 22820
rect 78092 23604 78148 23614
rect 77756 22372 77812 22764
rect 77868 22596 77924 22606
rect 78092 22596 78148 23548
rect 77868 22594 78148 22596
rect 77868 22542 77870 22594
rect 77922 22542 78148 22594
rect 77868 22540 78148 22542
rect 78204 23156 78260 23166
rect 77868 22530 77924 22540
rect 77756 22316 77924 22372
rect 76748 22260 76804 22270
rect 76636 22258 76804 22260
rect 76636 22206 76750 22258
rect 76802 22206 76804 22258
rect 76636 22204 76804 22206
rect 76188 22092 76580 22148
rect 76412 21924 76468 21934
rect 76076 21868 76244 21924
rect 76188 20804 76244 21868
rect 76412 20916 76468 21868
rect 76524 21474 76580 22092
rect 76636 21924 76692 22204
rect 76748 22194 76804 22204
rect 77084 22148 77140 22158
rect 77420 22148 77476 22158
rect 77084 22146 77252 22148
rect 77084 22094 77086 22146
rect 77138 22094 77252 22146
rect 77084 22092 77252 22094
rect 77084 22082 77140 22092
rect 76636 21858 76692 21868
rect 76524 21422 76526 21474
rect 76578 21422 76580 21474
rect 76524 21410 76580 21422
rect 76636 21698 76692 21710
rect 76636 21646 76638 21698
rect 76690 21646 76692 21698
rect 76412 20860 76580 20916
rect 76188 20748 76468 20804
rect 76300 20578 76356 20590
rect 76300 20526 76302 20578
rect 76354 20526 76356 20578
rect 76300 20356 76356 20526
rect 75964 20300 76356 20356
rect 75404 15922 75460 15932
rect 74396 15092 74452 15102
rect 73052 12740 73108 12750
rect 71708 7588 71764 7598
rect 71708 7494 71764 7532
rect 72380 7588 72436 7598
rect 72380 7474 72436 7532
rect 72380 7422 72382 7474
rect 72434 7422 72436 7474
rect 72380 7410 72436 7422
rect 72268 6468 72324 6478
rect 72268 6374 72324 6412
rect 72268 5906 72324 5918
rect 72268 5854 72270 5906
rect 72322 5854 72324 5906
rect 71708 5796 71764 5806
rect 71708 5702 71764 5740
rect 72268 5796 72324 5854
rect 72268 5730 72324 5740
rect 72828 5236 72884 5246
rect 71036 5122 71428 5124
rect 71036 5070 71374 5122
rect 71426 5070 71428 5122
rect 71036 5068 71428 5070
rect 71036 4562 71092 5068
rect 71372 5058 71428 5068
rect 72156 5124 72212 5134
rect 71036 4510 71038 4562
rect 71090 4510 71092 4562
rect 71036 4498 71092 4510
rect 71708 4228 71764 4238
rect 71708 4134 71764 4172
rect 71260 3668 71316 3678
rect 71260 3574 71316 3612
rect 71484 3444 71540 3454
rect 71484 800 71540 3388
rect 72156 800 72212 5068
rect 72268 4900 72324 4910
rect 72268 4806 72324 4844
rect 72268 4338 72324 4350
rect 72268 4286 72270 4338
rect 72322 4286 72324 4338
rect 72268 4228 72324 4286
rect 72268 4162 72324 4172
rect 72828 800 72884 5180
rect 73052 4228 73108 12684
rect 73388 8818 73444 8830
rect 73388 8766 73390 8818
rect 73442 8766 73444 8818
rect 73276 5684 73332 5694
rect 73276 5590 73332 5628
rect 73388 5012 73444 8766
rect 73724 8372 73780 8382
rect 73724 6692 73780 8316
rect 74284 8370 74340 8382
rect 74284 8318 74286 8370
rect 74338 8318 74340 8370
rect 73724 6626 73780 6636
rect 73836 8148 73892 8158
rect 73836 5460 73892 8092
rect 73612 5404 73836 5460
rect 73388 4946 73444 4956
rect 73500 5348 73556 5358
rect 73052 4162 73108 4172
rect 73276 4116 73332 4126
rect 73276 4022 73332 4060
rect 73500 800 73556 5292
rect 73612 3666 73668 5404
rect 73836 5394 73892 5404
rect 73948 7362 74004 7374
rect 73948 7310 73950 7362
rect 74002 7310 74004 7362
rect 73948 5124 74004 7310
rect 73948 5058 74004 5068
rect 74172 4228 74228 4238
rect 73612 3614 73614 3666
rect 73666 3614 73668 3666
rect 73612 3602 73668 3614
rect 74060 4004 74116 4014
rect 74060 3554 74116 3948
rect 74060 3502 74062 3554
rect 74114 3502 74116 3554
rect 74060 3490 74116 3502
rect 74172 800 74228 4172
rect 74284 980 74340 8318
rect 74396 5908 74452 15036
rect 74732 15092 75012 15148
rect 74508 13076 74564 13086
rect 74732 13076 74788 15092
rect 74508 13074 74788 13076
rect 74508 13022 74510 13074
rect 74562 13022 74734 13074
rect 74786 13022 74788 13074
rect 74508 13020 74788 13022
rect 74508 13010 74564 13020
rect 74732 13010 74788 13020
rect 74956 13076 75012 13086
rect 74956 12982 75012 13020
rect 75628 13076 75684 13086
rect 75292 12740 75348 12750
rect 75292 12646 75348 12684
rect 75516 10052 75572 10062
rect 75292 9604 75348 9614
rect 75180 9602 75348 9604
rect 75180 9550 75294 9602
rect 75346 9550 75348 9602
rect 75180 9548 75348 9550
rect 74956 7588 75012 7598
rect 74508 6690 74564 6702
rect 74508 6638 74510 6690
rect 74562 6638 74564 6690
rect 74508 6356 74564 6638
rect 74732 6692 74788 6702
rect 74732 6690 74900 6692
rect 74732 6638 74734 6690
rect 74786 6638 74900 6690
rect 74732 6636 74900 6638
rect 74732 6626 74788 6636
rect 74508 6290 74564 6300
rect 74396 5234 74452 5852
rect 74396 5182 74398 5234
rect 74450 5182 74452 5234
rect 74396 5170 74452 5182
rect 74620 5460 74676 5470
rect 74620 5234 74676 5404
rect 74844 5348 74900 6636
rect 74956 6244 75012 7532
rect 75180 6804 75236 9548
rect 75292 9538 75348 9548
rect 75292 9042 75348 9054
rect 75292 8990 75294 9042
rect 75346 8990 75348 9042
rect 75292 7700 75348 8990
rect 75292 7634 75348 7644
rect 75404 8820 75460 8830
rect 75404 7588 75460 8764
rect 75516 8258 75572 9996
rect 75516 8206 75518 8258
rect 75570 8206 75572 8258
rect 75516 8194 75572 8206
rect 75404 7522 75460 7532
rect 75292 7476 75348 7486
rect 75292 7382 75348 7420
rect 75180 6738 75236 6748
rect 75404 7252 75460 7262
rect 75068 6468 75124 6478
rect 75068 6466 75348 6468
rect 75068 6414 75070 6466
rect 75122 6414 75348 6466
rect 75068 6412 75348 6414
rect 75068 6402 75124 6412
rect 74956 6188 75124 6244
rect 74956 5460 75012 5470
rect 74956 5348 75012 5404
rect 74844 5346 75012 5348
rect 74844 5294 74846 5346
rect 74898 5294 75012 5346
rect 74844 5292 75012 5294
rect 74844 5282 74900 5292
rect 74620 5182 74622 5234
rect 74674 5182 74676 5234
rect 74620 5170 74676 5182
rect 74956 5124 75012 5134
rect 74508 5012 74564 5022
rect 74508 2996 74564 4956
rect 74956 4900 75012 5068
rect 74508 2930 74564 2940
rect 74844 4844 75012 4900
rect 74284 914 74340 924
rect 74844 800 74900 4844
rect 75068 4116 75124 6188
rect 75180 5908 75236 5918
rect 75180 5814 75236 5852
rect 75180 4900 75236 4910
rect 75180 4806 75236 4844
rect 75180 4116 75236 4126
rect 75068 4060 75180 4116
rect 75180 4050 75236 4060
rect 75068 3780 75124 3790
rect 75068 3686 75124 3724
rect 75292 3556 75348 6412
rect 75404 6132 75460 7196
rect 75516 6466 75572 6478
rect 75516 6414 75518 6466
rect 75570 6414 75572 6466
rect 75516 6356 75572 6414
rect 75516 6290 75572 6300
rect 75404 6076 75572 6132
rect 75404 5572 75460 5582
rect 75404 4338 75460 5516
rect 75404 4286 75406 4338
rect 75458 4286 75460 4338
rect 75404 4274 75460 4286
rect 75292 3490 75348 3500
rect 75516 1876 75572 6076
rect 75628 5460 75684 13020
rect 75628 5122 75684 5404
rect 75628 5070 75630 5122
rect 75682 5070 75684 5122
rect 75628 4564 75684 5070
rect 75740 9602 75796 9614
rect 75740 9550 75742 9602
rect 75794 9550 75796 9602
rect 75740 5124 75796 9550
rect 75852 8820 75908 8830
rect 75852 8726 75908 8764
rect 75964 7924 76020 20300
rect 76188 20132 76244 20142
rect 76188 20038 76244 20076
rect 76300 20130 76356 20142
rect 76300 20078 76302 20130
rect 76354 20078 76356 20130
rect 76076 20020 76132 20030
rect 76076 19926 76132 19964
rect 76300 18564 76356 20078
rect 76300 18498 76356 18508
rect 76300 13076 76356 13086
rect 76300 12982 76356 13020
rect 76300 9602 76356 9614
rect 76300 9550 76302 9602
rect 76354 9550 76356 9602
rect 76300 8428 76356 9550
rect 76412 9380 76468 20748
rect 76524 20580 76580 20860
rect 76636 20804 76692 21646
rect 76636 20738 76692 20748
rect 76748 21700 76804 21710
rect 76748 20802 76804 21644
rect 77196 21698 77252 22092
rect 77308 22036 77364 22046
rect 77308 21810 77364 21980
rect 77308 21758 77310 21810
rect 77362 21758 77364 21810
rect 77308 21746 77364 21758
rect 77196 21646 77198 21698
rect 77250 21646 77252 21698
rect 76860 21586 76916 21598
rect 76860 21534 76862 21586
rect 76914 21534 76916 21586
rect 76860 21476 76916 21534
rect 77196 21476 77252 21646
rect 76860 21420 77252 21476
rect 77084 21028 77140 21038
rect 77196 21028 77252 21420
rect 77420 21364 77476 22092
rect 77532 21812 77588 22316
rect 77756 22148 77812 22158
rect 77756 22054 77812 22092
rect 77532 21756 77812 21812
rect 77532 21588 77588 21598
rect 77532 21586 77700 21588
rect 77532 21534 77534 21586
rect 77586 21534 77700 21586
rect 77532 21532 77700 21534
rect 77532 21522 77588 21532
rect 77420 21308 77588 21364
rect 77420 21028 77476 21038
rect 77084 21026 77476 21028
rect 77084 20974 77086 21026
rect 77138 20974 77422 21026
rect 77474 20974 77476 21026
rect 77084 20972 77476 20974
rect 77084 20962 77140 20972
rect 77420 20962 77476 20972
rect 77532 20914 77588 21308
rect 77532 20862 77534 20914
rect 77586 20862 77588 20914
rect 77532 20850 77588 20862
rect 76748 20750 76750 20802
rect 76802 20750 76804 20802
rect 76748 20738 76804 20750
rect 76972 20580 77028 20590
rect 76524 20524 76804 20580
rect 76748 20130 76804 20524
rect 76972 20486 77028 20524
rect 76748 20078 76750 20130
rect 76802 20078 76804 20130
rect 76748 20066 76804 20078
rect 77084 20130 77140 20142
rect 77644 20132 77700 21532
rect 77756 21028 77812 21756
rect 77868 21810 77924 22316
rect 77868 21758 77870 21810
rect 77922 21758 77924 21810
rect 77868 21746 77924 21758
rect 78092 22036 78148 22046
rect 77756 20972 78036 21028
rect 77084 20078 77086 20130
rect 77138 20078 77140 20130
rect 76636 20020 76692 20030
rect 76636 19460 76692 19964
rect 77084 20020 77140 20078
rect 77532 20076 77700 20132
rect 77756 20802 77812 20814
rect 77756 20750 77758 20802
rect 77810 20750 77812 20802
rect 77084 19954 77140 19964
rect 77420 20020 77476 20030
rect 76748 19460 76804 19470
rect 76636 19458 76804 19460
rect 76636 19406 76750 19458
rect 76802 19406 76804 19458
rect 76636 19404 76804 19406
rect 76748 19394 76804 19404
rect 77420 19458 77476 19964
rect 77420 19406 77422 19458
rect 77474 19406 77476 19458
rect 77420 19394 77476 19406
rect 76524 19348 76580 19358
rect 76580 19292 76692 19348
rect 76524 19282 76580 19292
rect 76524 19010 76580 19022
rect 76524 18958 76526 19010
rect 76578 18958 76580 19010
rect 76524 18900 76580 18958
rect 76524 18834 76580 18844
rect 76636 14196 76692 19292
rect 76860 19236 76916 19246
rect 77532 19236 77588 20076
rect 77644 19908 77700 19918
rect 77644 19814 77700 19852
rect 77756 19572 77812 20750
rect 77868 20804 77924 20814
rect 77868 20130 77924 20748
rect 77868 20078 77870 20130
rect 77922 20078 77924 20130
rect 77868 20066 77924 20078
rect 77756 19516 77924 19572
rect 77532 19180 77700 19236
rect 76860 19142 76916 19180
rect 76972 19010 77028 19022
rect 76972 18958 76974 19010
rect 77026 18958 77028 19010
rect 76972 18564 77028 18958
rect 77532 19012 77588 19022
rect 77532 18918 77588 18956
rect 76860 18508 77028 18564
rect 77308 18676 77364 18686
rect 76860 14420 76916 18508
rect 77308 18450 77364 18620
rect 77532 18676 77588 18686
rect 77644 18676 77700 19180
rect 77532 18674 77700 18676
rect 77532 18622 77534 18674
rect 77586 18622 77700 18674
rect 77532 18620 77700 18622
rect 77756 19234 77812 19246
rect 77756 19182 77758 19234
rect 77810 19182 77812 19234
rect 77532 18610 77588 18620
rect 77308 18398 77310 18450
rect 77362 18398 77364 18450
rect 76972 18340 77028 18350
rect 76972 18246 77028 18284
rect 77308 18340 77364 18398
rect 77308 18274 77364 18284
rect 77644 17556 77700 17566
rect 77644 17462 77700 17500
rect 77756 17108 77812 19182
rect 77868 18674 77924 19516
rect 77868 18622 77870 18674
rect 77922 18622 77924 18674
rect 77868 18610 77924 18622
rect 77868 18452 77924 18462
rect 77868 17554 77924 18396
rect 77868 17502 77870 17554
rect 77922 17502 77924 17554
rect 77868 17490 77924 17502
rect 77868 17108 77924 17118
rect 77756 17106 77924 17108
rect 77756 17054 77870 17106
rect 77922 17054 77924 17106
rect 77756 17052 77924 17054
rect 77868 17042 77924 17052
rect 77644 16884 77700 16894
rect 77644 16790 77700 16828
rect 77868 15988 77924 15998
rect 77868 15894 77924 15932
rect 77644 15876 77700 15886
rect 77644 15782 77700 15820
rect 77084 15204 77140 15214
rect 77140 15148 77252 15204
rect 77084 15138 77140 15148
rect 76860 14354 76916 14364
rect 76636 14140 77140 14196
rect 76524 11508 76580 11518
rect 76524 11414 76580 11452
rect 76972 11170 77028 11182
rect 76972 11118 76974 11170
rect 77026 11118 77028 11170
rect 76972 10836 77028 11118
rect 76972 10770 77028 10780
rect 76412 9314 76468 9324
rect 76524 10498 76580 10510
rect 76524 10446 76526 10498
rect 76578 10446 76580 10498
rect 75964 7858 76020 7868
rect 76188 8372 76356 8428
rect 76188 7252 76244 8372
rect 76300 8034 76356 8046
rect 76300 7982 76302 8034
rect 76354 7982 76356 8034
rect 76300 7476 76356 7982
rect 76300 7410 76356 7420
rect 75964 7196 76244 7252
rect 76300 7250 76356 7262
rect 76300 7198 76302 7250
rect 76354 7198 76356 7250
rect 75964 6692 76020 7196
rect 76188 6692 76244 6702
rect 75964 6690 76244 6692
rect 75964 6638 76190 6690
rect 76242 6638 76244 6690
rect 75964 6636 76244 6638
rect 76188 6580 76244 6636
rect 76188 6514 76244 6524
rect 76188 5682 76244 5694
rect 76188 5630 76190 5682
rect 76242 5630 76244 5682
rect 76188 5236 76244 5630
rect 76300 5348 76356 7198
rect 76524 7252 76580 10446
rect 76972 9602 77028 9614
rect 76972 9550 76974 9602
rect 77026 9550 77028 9602
rect 76860 8260 76916 8270
rect 76860 8166 76916 8204
rect 76972 8148 77028 9550
rect 77084 8428 77140 14140
rect 77196 11282 77252 15148
rect 77980 15148 78036 20972
rect 78092 20020 78148 21980
rect 78204 21698 78260 23100
rect 78316 21924 78372 23884
rect 78540 22148 78596 22158
rect 78596 22092 78708 22148
rect 78540 22082 78596 22092
rect 78316 21868 78596 21924
rect 78204 21646 78206 21698
rect 78258 21646 78260 21698
rect 78204 20244 78260 21646
rect 78428 21700 78484 21710
rect 78316 20916 78372 20926
rect 78428 20916 78484 21644
rect 78316 20914 78484 20916
rect 78316 20862 78318 20914
rect 78370 20862 78484 20914
rect 78316 20860 78484 20862
rect 78316 20850 78372 20860
rect 78540 20804 78596 21868
rect 78204 20178 78260 20188
rect 78428 20748 78596 20804
rect 78092 20018 78372 20020
rect 78092 19966 78094 20018
rect 78146 19966 78372 20018
rect 78092 19964 78372 19966
rect 78092 19954 78148 19964
rect 78204 19796 78260 19806
rect 78204 18900 78260 19740
rect 78316 19346 78372 19964
rect 78316 19294 78318 19346
rect 78370 19294 78372 19346
rect 78316 19282 78372 19294
rect 78204 18450 78260 18844
rect 78204 18398 78206 18450
rect 78258 18398 78260 18450
rect 78204 18386 78260 18398
rect 78204 17556 78260 17566
rect 78204 17462 78260 17500
rect 78204 16884 78260 16894
rect 78204 16436 78260 16828
rect 78204 16370 78260 16380
rect 78204 15986 78260 15998
rect 78204 15934 78206 15986
rect 78258 15934 78260 15986
rect 78204 15876 78260 15934
rect 78204 15316 78260 15820
rect 78204 15250 78260 15260
rect 78428 15148 78484 20748
rect 77980 15092 78148 15148
rect 77868 14420 77924 14430
rect 77868 14326 77924 14364
rect 77644 14306 77700 14318
rect 77644 14254 77646 14306
rect 77698 14254 77700 14306
rect 77644 14196 77700 14254
rect 77644 14130 77700 14140
rect 77868 13972 77924 13982
rect 77868 13878 77924 13916
rect 77644 13636 77700 13646
rect 77644 13542 77700 13580
rect 77756 12740 77812 12750
rect 77532 12292 77588 12302
rect 77196 11230 77198 11282
rect 77250 11230 77252 11282
rect 77196 11218 77252 11230
rect 77420 12290 77588 12292
rect 77420 12238 77534 12290
rect 77586 12238 77588 12290
rect 77420 12236 77588 12238
rect 77420 10052 77476 12236
rect 77532 12226 77588 12236
rect 77756 12178 77812 12684
rect 77756 12126 77758 12178
rect 77810 12126 77812 12178
rect 77756 12114 77812 12126
rect 77532 11282 77588 11294
rect 77532 11230 77534 11282
rect 77586 11230 77588 11282
rect 77532 10836 77588 11230
rect 77868 11284 77924 11294
rect 78092 11284 78148 15092
rect 78316 15092 78484 15148
rect 78204 14418 78260 14430
rect 78204 14366 78206 14418
rect 78258 14366 78260 14418
rect 78204 14196 78260 14366
rect 78204 14130 78260 14140
rect 78204 13746 78260 13758
rect 78204 13694 78206 13746
rect 78258 13694 78260 13746
rect 78204 13636 78260 13694
rect 78204 13076 78260 13580
rect 78204 13010 78260 13020
rect 78204 11956 78260 11966
rect 78204 11508 78260 11900
rect 78204 11394 78260 11452
rect 78204 11342 78206 11394
rect 78258 11342 78260 11394
rect 78204 11330 78260 11342
rect 77868 11282 78148 11284
rect 77868 11230 77870 11282
rect 77922 11230 78148 11282
rect 77868 11228 78148 11230
rect 77868 11218 77924 11228
rect 78316 11172 78372 15092
rect 77532 10770 77588 10780
rect 77980 11116 78372 11172
rect 77420 9986 77476 9996
rect 77644 9716 77700 9726
rect 77644 9622 77700 9660
rect 77868 9604 77924 9614
rect 77868 9510 77924 9548
rect 77868 9380 77924 9390
rect 77756 9042 77812 9054
rect 77756 8990 77758 9042
rect 77810 8990 77812 9042
rect 77756 8428 77812 8990
rect 77084 8372 77252 8428
rect 76972 8082 77028 8092
rect 77196 8146 77252 8372
rect 77196 8094 77198 8146
rect 77250 8094 77252 8146
rect 77196 8082 77252 8094
rect 77308 8372 77812 8428
rect 76860 7924 76916 7934
rect 76916 7868 77252 7924
rect 76860 7858 76916 7868
rect 76524 7186 76580 7196
rect 76300 5282 76356 5292
rect 76412 6690 76468 6702
rect 76412 6638 76414 6690
rect 76466 6638 76468 6690
rect 76188 5170 76244 5180
rect 75740 5058 75796 5068
rect 76300 5124 76356 5134
rect 76300 5030 76356 5068
rect 75628 4498 75684 4508
rect 76412 4564 76468 6638
rect 76636 6692 76692 6702
rect 76636 5234 76692 6636
rect 77196 6578 77252 7868
rect 77196 6526 77198 6578
rect 77250 6526 77252 6578
rect 77196 6514 77252 6526
rect 76748 6468 76804 6478
rect 76748 6374 76804 6412
rect 76636 5182 76638 5234
rect 76690 5182 76692 5234
rect 76636 5170 76692 5182
rect 77196 5122 77252 5134
rect 77196 5070 77198 5122
rect 77250 5070 77252 5122
rect 76412 4498 76468 4508
rect 76972 4900 77028 4910
rect 76188 4114 76244 4126
rect 76188 4062 76190 4114
rect 76242 4062 76244 4114
rect 76188 3444 76244 4062
rect 76972 3554 77028 4844
rect 77196 4564 77252 5070
rect 77196 4498 77252 4508
rect 76972 3502 76974 3554
rect 77026 3502 77028 3554
rect 76972 3490 77028 3502
rect 76188 3378 76244 3388
rect 77308 3442 77364 8372
rect 77532 8148 77588 8158
rect 77420 7700 77476 7710
rect 77420 6356 77476 7644
rect 77532 7476 77588 8092
rect 77868 8146 77924 9324
rect 77868 8094 77870 8146
rect 77922 8094 77924 8146
rect 77868 8082 77924 8094
rect 77532 7410 77588 7420
rect 77980 7028 78036 11116
rect 78204 10612 78260 10622
rect 78204 10610 78484 10612
rect 78204 10558 78206 10610
rect 78258 10558 78484 10610
rect 78204 10556 78484 10558
rect 78204 10546 78260 10556
rect 78204 9716 78260 9726
rect 78204 9622 78260 9660
rect 78204 8596 78260 8606
rect 78092 8260 78148 8270
rect 78204 8260 78260 8540
rect 78148 8204 78260 8260
rect 78092 8166 78148 8204
rect 77868 6972 78036 7028
rect 77532 6804 77588 6814
rect 77532 6580 77588 6748
rect 77532 6578 77700 6580
rect 77532 6526 77534 6578
rect 77586 6526 77700 6578
rect 77532 6524 77700 6526
rect 77532 6514 77588 6524
rect 77420 6300 77588 6356
rect 77532 5010 77588 6300
rect 77644 5236 77700 6524
rect 77868 6578 77924 6972
rect 77868 6526 77870 6578
rect 77922 6526 77924 6578
rect 77868 6514 77924 6526
rect 78204 6578 78260 6590
rect 78204 6526 78206 6578
rect 78258 6526 78260 6578
rect 77644 5170 77700 5180
rect 77756 6468 77812 6478
rect 77756 5122 77812 6412
rect 78204 6356 78260 6526
rect 78316 6356 78372 6366
rect 78204 6300 78316 6356
rect 78316 6130 78372 6300
rect 78316 6078 78318 6130
rect 78370 6078 78372 6130
rect 78316 6066 78372 6078
rect 77756 5070 77758 5122
rect 77810 5070 77812 5122
rect 77756 5058 77812 5070
rect 77532 4958 77534 5010
rect 77586 4958 77588 5010
rect 77532 4946 77588 4958
rect 78204 4564 78260 4574
rect 78204 4470 78260 4508
rect 77868 3556 77924 3566
rect 77868 3462 77924 3500
rect 77308 3390 77310 3442
rect 77362 3390 77364 3442
rect 77308 3378 77364 3390
rect 78204 3444 78260 3454
rect 78428 3444 78484 10556
rect 78652 9604 78708 22092
rect 78764 21700 78820 26460
rect 78764 21634 78820 21644
rect 78652 9538 78708 9548
rect 78204 3442 78484 3444
rect 78204 3390 78206 3442
rect 78258 3390 78484 3442
rect 78204 3388 78484 3390
rect 78204 3378 78260 3388
rect 75516 1810 75572 1820
rect 4060 700 4788 756
rect 4928 0 5040 800
rect 5600 0 5712 800
rect 6272 0 6384 800
rect 6944 0 7056 800
rect 7616 0 7728 800
rect 8288 0 8400 800
rect 8960 0 9072 800
rect 9632 0 9744 800
rect 10304 0 10416 800
rect 10976 0 11088 800
rect 11648 0 11760 800
rect 12320 0 12432 800
rect 12992 0 13104 800
rect 13664 0 13776 800
rect 14336 0 14448 800
rect 15008 0 15120 800
rect 15680 0 15792 800
rect 16352 0 16464 800
rect 17024 0 17136 800
rect 17696 0 17808 800
rect 18368 0 18480 800
rect 19040 0 19152 800
rect 19712 0 19824 800
rect 20384 0 20496 800
rect 21056 0 21168 800
rect 21728 0 21840 800
rect 22400 0 22512 800
rect 23072 0 23184 800
rect 23744 0 23856 800
rect 24416 0 24528 800
rect 25088 0 25200 800
rect 25760 0 25872 800
rect 26432 0 26544 800
rect 27104 0 27216 800
rect 27776 0 27888 800
rect 28448 0 28560 800
rect 29120 0 29232 800
rect 29792 0 29904 800
rect 30464 0 30576 800
rect 31136 0 31248 800
rect 31808 0 31920 800
rect 32480 0 32592 800
rect 33152 0 33264 800
rect 33824 0 33936 800
rect 34496 0 34608 800
rect 35168 0 35280 800
rect 35840 0 35952 800
rect 36512 0 36624 800
rect 37184 0 37296 800
rect 37856 0 37968 800
rect 38528 0 38640 800
rect 39200 0 39312 800
rect 39872 0 39984 800
rect 40544 0 40656 800
rect 41216 0 41328 800
rect 41888 0 42000 800
rect 42560 0 42672 800
rect 43232 0 43344 800
rect 43904 0 44016 800
rect 44576 0 44688 800
rect 45248 0 45360 800
rect 45920 0 46032 800
rect 46592 0 46704 800
rect 47264 0 47376 800
rect 47936 0 48048 800
rect 48608 0 48720 800
rect 49280 0 49392 800
rect 49952 0 50064 800
rect 50624 0 50736 800
rect 51296 0 51408 800
rect 51968 0 52080 800
rect 52640 0 52752 800
rect 53312 0 53424 800
rect 53984 0 54096 800
rect 54656 0 54768 800
rect 55328 0 55440 800
rect 56000 0 56112 800
rect 56672 0 56784 800
rect 57344 0 57456 800
rect 58016 0 58128 800
rect 58688 0 58800 800
rect 59360 0 59472 800
rect 60032 0 60144 800
rect 60704 0 60816 800
rect 61376 0 61488 800
rect 62048 0 62160 800
rect 62720 0 62832 800
rect 63392 0 63504 800
rect 64064 0 64176 800
rect 64736 0 64848 800
rect 65408 0 65520 800
rect 66080 0 66192 800
rect 66752 0 66864 800
rect 67424 0 67536 800
rect 68096 0 68208 800
rect 68768 0 68880 800
rect 69440 0 69552 800
rect 70112 0 70224 800
rect 70784 0 70896 800
rect 71456 0 71568 800
rect 72128 0 72240 800
rect 72800 0 72912 800
rect 73472 0 73584 800
rect 74144 0 74256 800
rect 74816 0 74928 800
<< via2 >>
rect 2156 77308 2212 77364
rect 1932 76242 1988 76244
rect 1932 76190 1934 76242
rect 1934 76190 1986 76242
rect 1986 76190 1988 76242
rect 1932 76188 1988 76190
rect 1932 75292 1988 75348
rect 4476 76074 4532 76076
rect 4476 76022 4478 76074
rect 4478 76022 4530 76074
rect 4530 76022 4532 76074
rect 4476 76020 4532 76022
rect 4580 76074 4636 76076
rect 4580 76022 4582 76074
rect 4582 76022 4634 76074
rect 4634 76022 4636 76074
rect 4580 76020 4636 76022
rect 4684 76074 4740 76076
rect 4684 76022 4686 76074
rect 4686 76022 4738 76074
rect 4738 76022 4740 76074
rect 4684 76020 4740 76022
rect 4476 74506 4532 74508
rect 4476 74454 4478 74506
rect 4478 74454 4530 74506
rect 4530 74454 4532 74506
rect 4476 74452 4532 74454
rect 4580 74506 4636 74508
rect 4580 74454 4582 74506
rect 4582 74454 4634 74506
rect 4634 74454 4636 74506
rect 4580 74452 4636 74454
rect 4684 74506 4740 74508
rect 4684 74454 4686 74506
rect 4686 74454 4738 74506
rect 4738 74454 4740 74506
rect 4684 74452 4740 74454
rect 1932 74226 1988 74228
rect 1932 74174 1934 74226
rect 1934 74174 1986 74226
rect 1986 74174 1988 74226
rect 1932 74172 1988 74174
rect 1932 73106 1988 73108
rect 1932 73054 1934 73106
rect 1934 73054 1986 73106
rect 1986 73054 1988 73106
rect 1932 73052 1988 73054
rect 4476 72938 4532 72940
rect 4476 72886 4478 72938
rect 4478 72886 4530 72938
rect 4530 72886 4532 72938
rect 4476 72884 4532 72886
rect 4580 72938 4636 72940
rect 4580 72886 4582 72938
rect 4582 72886 4634 72938
rect 4634 72886 4636 72938
rect 4580 72884 4636 72886
rect 4684 72938 4740 72940
rect 4684 72886 4686 72938
rect 4686 72886 4738 72938
rect 4738 72886 4740 72938
rect 4684 72884 4740 72886
rect 1932 71932 1988 71988
rect 3164 71986 3220 71988
rect 3164 71934 3166 71986
rect 3166 71934 3218 71986
rect 3218 71934 3220 71986
rect 3164 71932 3220 71934
rect 2492 71874 2548 71876
rect 2492 71822 2494 71874
rect 2494 71822 2546 71874
rect 2546 71822 2548 71874
rect 2492 71820 2548 71822
rect 2940 71820 2996 71876
rect 3948 71932 4004 71988
rect 1932 70588 1988 70644
rect 2716 70140 2772 70196
rect 1932 69468 1988 69524
rect 1932 67228 1988 67284
rect 4508 71874 4564 71876
rect 4508 71822 4510 71874
rect 4510 71822 4562 71874
rect 4562 71822 4564 71874
rect 4508 71820 4564 71822
rect 12460 76300 12516 76356
rect 11900 75906 11956 75908
rect 11900 75854 11902 75906
rect 11902 75854 11954 75906
rect 11954 75854 11956 75906
rect 11900 75852 11956 75854
rect 11564 75516 11620 75572
rect 11676 74844 11732 74900
rect 5740 71820 5796 71876
rect 4476 71370 4532 71372
rect 4476 71318 4478 71370
rect 4478 71318 4530 71370
rect 4530 71318 4532 71370
rect 4476 71316 4532 71318
rect 4580 71370 4636 71372
rect 4580 71318 4582 71370
rect 4582 71318 4634 71370
rect 4634 71318 4636 71370
rect 4580 71316 4636 71318
rect 4684 71370 4740 71372
rect 4684 71318 4686 71370
rect 4686 71318 4738 71370
rect 4738 71318 4740 71370
rect 4684 71316 4740 71318
rect 3836 70194 3892 70196
rect 3836 70142 3838 70194
rect 3838 70142 3890 70194
rect 3890 70142 3892 70194
rect 3836 70140 3892 70142
rect 4476 69802 4532 69804
rect 4476 69750 4478 69802
rect 4478 69750 4530 69802
rect 4530 69750 4532 69802
rect 4476 69748 4532 69750
rect 4580 69802 4636 69804
rect 4580 69750 4582 69802
rect 4582 69750 4634 69802
rect 4634 69750 4636 69802
rect 4580 69748 4636 69750
rect 4684 69802 4740 69804
rect 4684 69750 4686 69802
rect 4686 69750 4738 69802
rect 4738 69750 4740 69802
rect 4684 69748 4740 69750
rect 2716 68402 2772 68404
rect 2716 68350 2718 68402
rect 2718 68350 2770 68402
rect 2770 68350 2772 68402
rect 2716 68348 2772 68350
rect 4476 68234 4532 68236
rect 4476 68182 4478 68234
rect 4478 68182 4530 68234
rect 4530 68182 4532 68234
rect 4476 68180 4532 68182
rect 4580 68234 4636 68236
rect 4580 68182 4582 68234
rect 4582 68182 4634 68234
rect 4634 68182 4636 68234
rect 4580 68180 4636 68182
rect 4684 68234 4740 68236
rect 4684 68182 4686 68234
rect 4686 68182 4738 68234
rect 4738 68182 4740 68234
rect 4684 68180 4740 68182
rect 2380 67170 2436 67172
rect 2380 67118 2382 67170
rect 2382 67118 2434 67170
rect 2434 67118 2436 67170
rect 2380 67116 2436 67118
rect 3052 67170 3108 67172
rect 3052 67118 3054 67170
rect 3054 67118 3106 67170
rect 3106 67118 3108 67170
rect 3052 67116 3108 67118
rect 1932 65266 1988 65268
rect 1932 65214 1934 65266
rect 1934 65214 1986 65266
rect 1986 65214 1988 65266
rect 1932 65212 1988 65214
rect 4476 66666 4532 66668
rect 4476 66614 4478 66666
rect 4478 66614 4530 66666
rect 4530 66614 4532 66666
rect 4476 66612 4532 66614
rect 4580 66666 4636 66668
rect 4580 66614 4582 66666
rect 4582 66614 4634 66666
rect 4634 66614 4636 66666
rect 4580 66612 4636 66614
rect 4684 66666 4740 66668
rect 4684 66614 4686 66666
rect 4686 66614 4738 66666
rect 4738 66614 4740 66666
rect 4684 66612 4740 66614
rect 2716 66050 2772 66052
rect 2716 65998 2718 66050
rect 2718 65998 2770 66050
rect 2770 65998 2772 66050
rect 2716 65996 2772 65998
rect 4476 65098 4532 65100
rect 4476 65046 4478 65098
rect 4478 65046 4530 65098
rect 4530 65046 4532 65098
rect 4476 65044 4532 65046
rect 4580 65098 4636 65100
rect 4580 65046 4582 65098
rect 4582 65046 4634 65098
rect 4634 65046 4636 65098
rect 4580 65044 4636 65046
rect 4684 65098 4740 65100
rect 4684 65046 4686 65098
rect 4686 65046 4738 65098
rect 4738 65046 4740 65098
rect 4684 65044 4740 65046
rect 1932 63868 1988 63924
rect 3612 64540 3668 64596
rect 1932 62748 1988 62804
rect 1932 61628 1988 61684
rect 2492 63868 2548 63924
rect 2940 63922 2996 63924
rect 2940 63870 2942 63922
rect 2942 63870 2994 63922
rect 2994 63870 2996 63922
rect 2940 63868 2996 63870
rect 4956 64594 5012 64596
rect 4956 64542 4958 64594
rect 4958 64542 5010 64594
rect 5010 64542 5012 64594
rect 4956 64540 5012 64542
rect 3612 63922 3668 63924
rect 3612 63870 3614 63922
rect 3614 63870 3666 63922
rect 3666 63870 3668 63922
rect 3612 63868 3668 63870
rect 4476 63530 4532 63532
rect 4476 63478 4478 63530
rect 4478 63478 4530 63530
rect 4530 63478 4532 63530
rect 4476 63476 4532 63478
rect 4580 63530 4636 63532
rect 4580 63478 4582 63530
rect 4582 63478 4634 63530
rect 4634 63478 4636 63530
rect 4580 63476 4636 63478
rect 4684 63530 4740 63532
rect 4684 63478 4686 63530
rect 4686 63478 4738 63530
rect 4738 63478 4740 63530
rect 4684 63476 4740 63478
rect 2940 61516 2996 61572
rect 4476 61962 4532 61964
rect 4476 61910 4478 61962
rect 4478 61910 4530 61962
rect 4530 61910 4532 61962
rect 4476 61908 4532 61910
rect 4580 61962 4636 61964
rect 4580 61910 4582 61962
rect 4582 61910 4634 61962
rect 4634 61910 4636 61962
rect 4580 61908 4636 61910
rect 4684 61962 4740 61964
rect 4684 61910 4686 61962
rect 4686 61910 4738 61962
rect 4738 61910 4740 61962
rect 4684 61908 4740 61910
rect 3612 61570 3668 61572
rect 3612 61518 3614 61570
rect 3614 61518 3666 61570
rect 3666 61518 3668 61570
rect 3612 61516 3668 61518
rect 3052 61292 3108 61348
rect 4172 61292 4228 61348
rect 2716 60562 2772 60564
rect 2716 60510 2718 60562
rect 2718 60510 2770 60562
rect 2770 60510 2772 60562
rect 2716 60508 2772 60510
rect 1932 59388 1988 59444
rect 2716 59948 2772 60004
rect 3836 60002 3892 60004
rect 3836 59950 3838 60002
rect 3838 59950 3890 60002
rect 3890 59950 3892 60002
rect 3836 59948 3892 59950
rect 2156 59164 2212 59220
rect 1932 57426 1988 57428
rect 1932 57374 1934 57426
rect 1934 57374 1986 57426
rect 1986 57374 1988 57426
rect 1932 57372 1988 57374
rect 1932 56028 1988 56084
rect 1932 53788 1988 53844
rect 2940 59218 2996 59220
rect 2940 59166 2942 59218
rect 2942 59166 2994 59218
rect 2994 59166 2996 59218
rect 2940 59164 2996 59166
rect 3500 59218 3556 59220
rect 3500 59166 3502 59218
rect 3502 59166 3554 59218
rect 3554 59166 3556 59218
rect 3500 59164 3556 59166
rect 2716 58210 2772 58212
rect 2716 58158 2718 58210
rect 2718 58158 2770 58210
rect 2770 58158 2772 58210
rect 2716 58156 2772 58158
rect 2716 56140 2772 56196
rect 3388 56194 3444 56196
rect 3388 56142 3390 56194
rect 3390 56142 3442 56194
rect 3442 56142 3444 56194
rect 3388 56140 3444 56142
rect 2716 55074 2772 55076
rect 2716 55022 2718 55074
rect 2718 55022 2770 55074
rect 2770 55022 2772 55074
rect 2716 55020 2772 55022
rect 4476 60394 4532 60396
rect 4476 60342 4478 60394
rect 4478 60342 4530 60394
rect 4530 60342 4532 60394
rect 4476 60340 4532 60342
rect 4580 60394 4636 60396
rect 4580 60342 4582 60394
rect 4582 60342 4634 60394
rect 4634 60342 4636 60394
rect 4580 60340 4636 60342
rect 4684 60394 4740 60396
rect 4684 60342 4686 60394
rect 4686 60342 4738 60394
rect 4738 60342 4740 60394
rect 4684 60340 4740 60342
rect 4476 58826 4532 58828
rect 4476 58774 4478 58826
rect 4478 58774 4530 58826
rect 4530 58774 4532 58826
rect 4476 58772 4532 58774
rect 4580 58826 4636 58828
rect 4580 58774 4582 58826
rect 4582 58774 4634 58826
rect 4634 58774 4636 58826
rect 4580 58772 4636 58774
rect 4684 58826 4740 58828
rect 4684 58774 4686 58826
rect 4686 58774 4738 58826
rect 4738 58774 4740 58826
rect 4684 58772 4740 58774
rect 4476 57258 4532 57260
rect 4476 57206 4478 57258
rect 4478 57206 4530 57258
rect 4530 57206 4532 57258
rect 4476 57204 4532 57206
rect 4580 57258 4636 57260
rect 4580 57206 4582 57258
rect 4582 57206 4634 57258
rect 4634 57206 4636 57258
rect 4580 57204 4636 57206
rect 4684 57258 4740 57260
rect 4684 57206 4686 57258
rect 4686 57206 4738 57258
rect 4738 57206 4740 57258
rect 4684 57204 4740 57206
rect 4844 56140 4900 56196
rect 4476 55690 4532 55692
rect 4476 55638 4478 55690
rect 4478 55638 4530 55690
rect 4530 55638 4532 55690
rect 4476 55636 4532 55638
rect 4580 55690 4636 55692
rect 4580 55638 4582 55690
rect 4582 55638 4634 55690
rect 4634 55638 4636 55690
rect 4580 55636 4636 55638
rect 4684 55690 4740 55692
rect 4684 55638 4686 55690
rect 4686 55638 4738 55690
rect 4738 55638 4740 55690
rect 4684 55636 4740 55638
rect 1932 52722 1988 52724
rect 1932 52670 1934 52722
rect 1934 52670 1986 52722
rect 1986 52670 1988 52722
rect 1932 52668 1988 52670
rect 1932 51548 1988 51604
rect 1932 50706 1988 50708
rect 1932 50654 1934 50706
rect 1934 50654 1986 50706
rect 1986 50654 1988 50706
rect 1932 50652 1988 50654
rect 1932 49586 1988 49588
rect 1932 49534 1934 49586
rect 1934 49534 1986 49586
rect 1986 49534 1988 49586
rect 1932 49532 1988 49534
rect 1932 48188 1988 48244
rect 1932 45948 1988 46004
rect 2492 53506 2548 53508
rect 2492 53454 2494 53506
rect 2494 53454 2546 53506
rect 2546 53454 2548 53506
rect 2492 53452 2548 53454
rect 3164 53618 3220 53620
rect 3164 53566 3166 53618
rect 3166 53566 3218 53618
rect 3218 53566 3220 53618
rect 3164 53564 3220 53566
rect 2940 53452 2996 53508
rect 3836 53452 3892 53508
rect 3948 53564 4004 53620
rect 2828 50540 2884 50596
rect 3836 50594 3892 50596
rect 3836 50542 3838 50594
rect 3838 50542 3890 50594
rect 3890 50542 3892 50594
rect 3836 50540 3892 50542
rect 3164 49532 3220 49588
rect 2716 48972 2772 49028
rect 3612 49532 3668 49588
rect 3836 49026 3892 49028
rect 3836 48974 3838 49026
rect 3838 48974 3890 49026
rect 3890 48974 3892 49026
rect 3836 48972 3892 48974
rect 2716 47234 2772 47236
rect 2716 47182 2718 47234
rect 2718 47182 2770 47234
rect 2770 47182 2772 47234
rect 2716 47180 2772 47182
rect 2380 45890 2436 45892
rect 2380 45838 2382 45890
rect 2382 45838 2434 45890
rect 2434 45838 2436 45890
rect 2380 45836 2436 45838
rect 2828 45724 2884 45780
rect 3052 45836 3108 45892
rect 3276 45724 3332 45780
rect 2716 44882 2772 44884
rect 2716 44830 2718 44882
rect 2718 44830 2770 44882
rect 2770 44830 2772 44882
rect 2716 44828 2772 44830
rect 2716 44098 2772 44100
rect 2716 44046 2718 44098
rect 2718 44046 2770 44098
rect 2770 44046 2772 44098
rect 2716 44044 2772 44046
rect 2268 43538 2324 43540
rect 2268 43486 2270 43538
rect 2270 43486 2322 43538
rect 2322 43486 2324 43538
rect 2268 43484 2324 43486
rect 1932 42866 1988 42868
rect 1932 42814 1934 42866
rect 1934 42814 1986 42866
rect 1986 42814 1988 42866
rect 1932 42812 1988 42814
rect 1708 41916 1764 41972
rect 1932 41746 1988 41748
rect 1932 41694 1934 41746
rect 1934 41694 1986 41746
rect 1986 41694 1988 41746
rect 1932 41692 1988 41694
rect 1932 40348 1988 40404
rect 1932 39228 1988 39284
rect 2268 40626 2324 40628
rect 2268 40574 2270 40626
rect 2270 40574 2322 40626
rect 2322 40574 2324 40626
rect 2268 40572 2324 40574
rect 2828 43484 2884 43540
rect 2716 42700 2772 42756
rect 3164 40402 3220 40404
rect 3164 40350 3166 40402
rect 3166 40350 3218 40402
rect 3218 40350 3220 40402
rect 3164 40348 3220 40350
rect 2604 39564 2660 39620
rect 2940 38668 2996 38724
rect 3612 45890 3668 45892
rect 3612 45838 3614 45890
rect 3614 45838 3666 45890
rect 3666 45838 3668 45890
rect 3612 45836 3668 45838
rect 3836 42754 3892 42756
rect 3836 42702 3838 42754
rect 3838 42702 3890 42754
rect 3890 42702 3892 42754
rect 3836 42700 3892 42702
rect 3836 41970 3892 41972
rect 3836 41918 3838 41970
rect 3838 41918 3890 41970
rect 3890 41918 3892 41970
rect 3836 41916 3892 41918
rect 4476 54122 4532 54124
rect 4476 54070 4478 54122
rect 4478 54070 4530 54122
rect 4530 54070 4532 54122
rect 4476 54068 4532 54070
rect 4580 54122 4636 54124
rect 4580 54070 4582 54122
rect 4582 54070 4634 54122
rect 4634 54070 4636 54122
rect 4580 54068 4636 54070
rect 4684 54122 4740 54124
rect 4684 54070 4686 54122
rect 4686 54070 4738 54122
rect 4738 54070 4740 54122
rect 4684 54068 4740 54070
rect 4476 52554 4532 52556
rect 4476 52502 4478 52554
rect 4478 52502 4530 52554
rect 4530 52502 4532 52554
rect 4476 52500 4532 52502
rect 4580 52554 4636 52556
rect 4580 52502 4582 52554
rect 4582 52502 4634 52554
rect 4634 52502 4636 52554
rect 4580 52500 4636 52502
rect 4684 52554 4740 52556
rect 4684 52502 4686 52554
rect 4686 52502 4738 52554
rect 4738 52502 4740 52554
rect 4684 52500 4740 52502
rect 4476 50986 4532 50988
rect 4476 50934 4478 50986
rect 4478 50934 4530 50986
rect 4530 50934 4532 50986
rect 4476 50932 4532 50934
rect 4580 50986 4636 50988
rect 4580 50934 4582 50986
rect 4582 50934 4634 50986
rect 4634 50934 4636 50986
rect 4580 50932 4636 50934
rect 4684 50986 4740 50988
rect 4684 50934 4686 50986
rect 4686 50934 4738 50986
rect 4738 50934 4740 50986
rect 4684 50932 4740 50934
rect 4476 49418 4532 49420
rect 4476 49366 4478 49418
rect 4478 49366 4530 49418
rect 4530 49366 4532 49418
rect 4476 49364 4532 49366
rect 4580 49418 4636 49420
rect 4580 49366 4582 49418
rect 4582 49366 4634 49418
rect 4634 49366 4636 49418
rect 4580 49364 4636 49366
rect 4684 49418 4740 49420
rect 4684 49366 4686 49418
rect 4686 49366 4738 49418
rect 4738 49366 4740 49418
rect 4684 49364 4740 49366
rect 4476 47850 4532 47852
rect 4476 47798 4478 47850
rect 4478 47798 4530 47850
rect 4530 47798 4532 47850
rect 4476 47796 4532 47798
rect 4580 47850 4636 47852
rect 4580 47798 4582 47850
rect 4582 47798 4634 47850
rect 4634 47798 4636 47850
rect 4580 47796 4636 47798
rect 4684 47850 4740 47852
rect 4684 47798 4686 47850
rect 4686 47798 4738 47850
rect 4738 47798 4740 47850
rect 4684 47796 4740 47798
rect 4476 46282 4532 46284
rect 4476 46230 4478 46282
rect 4478 46230 4530 46282
rect 4530 46230 4532 46282
rect 4476 46228 4532 46230
rect 4580 46282 4636 46284
rect 4580 46230 4582 46282
rect 4582 46230 4634 46282
rect 4634 46230 4636 46282
rect 4580 46228 4636 46230
rect 4684 46282 4740 46284
rect 4684 46230 4686 46282
rect 4686 46230 4738 46282
rect 4738 46230 4740 46282
rect 4684 46228 4740 46230
rect 4284 45778 4340 45780
rect 4284 45726 4286 45778
rect 4286 45726 4338 45778
rect 4338 45726 4340 45778
rect 4284 45724 4340 45726
rect 4476 44714 4532 44716
rect 4476 44662 4478 44714
rect 4478 44662 4530 44714
rect 4530 44662 4532 44714
rect 4476 44660 4532 44662
rect 4580 44714 4636 44716
rect 4580 44662 4582 44714
rect 4582 44662 4634 44714
rect 4634 44662 4636 44714
rect 4580 44660 4636 44662
rect 4684 44714 4740 44716
rect 4684 44662 4686 44714
rect 4686 44662 4738 44714
rect 4738 44662 4740 44714
rect 4684 44660 4740 44662
rect 4476 43146 4532 43148
rect 4476 43094 4478 43146
rect 4478 43094 4530 43146
rect 4530 43094 4532 43146
rect 4476 43092 4532 43094
rect 4580 43146 4636 43148
rect 4580 43094 4582 43146
rect 4582 43094 4634 43146
rect 4634 43094 4636 43146
rect 4580 43092 4636 43094
rect 4684 43146 4740 43148
rect 4684 43094 4686 43146
rect 4686 43094 4738 43146
rect 4738 43094 4740 43146
rect 4684 43092 4740 43094
rect 4732 41970 4788 41972
rect 4732 41918 4734 41970
rect 4734 41918 4786 41970
rect 4786 41918 4788 41970
rect 4732 41916 4788 41918
rect 4476 41578 4532 41580
rect 4476 41526 4478 41578
rect 4478 41526 4530 41578
rect 4530 41526 4532 41578
rect 4476 41524 4532 41526
rect 4580 41578 4636 41580
rect 4580 41526 4582 41578
rect 4582 41526 4634 41578
rect 4634 41526 4636 41578
rect 4580 41524 4636 41526
rect 4684 41578 4740 41580
rect 4684 41526 4686 41578
rect 4686 41526 4738 41578
rect 4738 41526 4740 41578
rect 4684 41524 4740 41526
rect 5404 40572 5460 40628
rect 4060 40514 4116 40516
rect 4060 40462 4062 40514
rect 4062 40462 4114 40514
rect 4114 40462 4116 40514
rect 4060 40460 4116 40462
rect 4508 40514 4564 40516
rect 4508 40462 4510 40514
rect 4510 40462 4562 40514
rect 4562 40462 4564 40514
rect 4508 40460 4564 40462
rect 5180 40460 5236 40516
rect 4956 40402 5012 40404
rect 4956 40350 4958 40402
rect 4958 40350 5010 40402
rect 5010 40350 5012 40402
rect 4956 40348 5012 40350
rect 4476 40010 4532 40012
rect 4476 39958 4478 40010
rect 4478 39958 4530 40010
rect 4530 39958 4532 40010
rect 4476 39956 4532 39958
rect 4580 40010 4636 40012
rect 4580 39958 4582 40010
rect 4582 39958 4634 40010
rect 4634 39958 4636 40010
rect 4580 39956 4636 39958
rect 4684 40010 4740 40012
rect 4684 39958 4686 40010
rect 4686 39958 4738 40010
rect 4738 39958 4740 40010
rect 4684 39956 4740 39958
rect 3836 39618 3892 39620
rect 3836 39566 3838 39618
rect 3838 39566 3890 39618
rect 3890 39566 3892 39618
rect 3836 39564 3892 39566
rect 4732 39618 4788 39620
rect 4732 39566 4734 39618
rect 4734 39566 4786 39618
rect 4786 39566 4788 39618
rect 4732 39564 4788 39566
rect 5180 39340 5236 39396
rect 3276 38668 3332 38724
rect 4476 38442 4532 38444
rect 4476 38390 4478 38442
rect 4478 38390 4530 38442
rect 4530 38390 4532 38442
rect 4476 38388 4532 38390
rect 4580 38442 4636 38444
rect 4580 38390 4582 38442
rect 4582 38390 4634 38442
rect 4634 38390 4636 38442
rect 4580 38388 4636 38390
rect 4684 38442 4740 38444
rect 4684 38390 4686 38442
rect 4686 38390 4738 38442
rect 4738 38390 4740 38442
rect 4684 38388 4740 38390
rect 3388 38108 3444 38164
rect 2044 37378 2100 37380
rect 2044 37326 2046 37378
rect 2046 37326 2098 37378
rect 2098 37326 2100 37378
rect 2044 37324 2100 37326
rect 1708 36988 1764 37044
rect 2492 36988 2548 37044
rect 4476 36874 4532 36876
rect 4476 36822 4478 36874
rect 4478 36822 4530 36874
rect 4530 36822 4532 36874
rect 4476 36820 4532 36822
rect 4580 36874 4636 36876
rect 4580 36822 4582 36874
rect 4582 36822 4634 36874
rect 4634 36822 4636 36874
rect 4580 36820 4636 36822
rect 4684 36874 4740 36876
rect 4684 36822 4686 36874
rect 4686 36822 4738 36874
rect 4738 36822 4740 36874
rect 4684 36820 4740 36822
rect 2044 36258 2100 36260
rect 2044 36206 2046 36258
rect 2046 36206 2098 36258
rect 2098 36206 2100 36258
rect 2044 36204 2100 36206
rect 1708 35868 1764 35924
rect 2492 35868 2548 35924
rect 4476 35306 4532 35308
rect 4476 35254 4478 35306
rect 4478 35254 4530 35306
rect 4530 35254 4532 35306
rect 4476 35252 4532 35254
rect 4580 35306 4636 35308
rect 4580 35254 4582 35306
rect 4582 35254 4634 35306
rect 4634 35254 4636 35306
rect 4580 35252 4636 35254
rect 4684 35306 4740 35308
rect 4684 35254 4686 35306
rect 4686 35254 4738 35306
rect 4738 35254 4740 35306
rect 4684 35252 4740 35254
rect 1708 34802 1764 34804
rect 1708 34750 1710 34802
rect 1710 34750 1762 34802
rect 1762 34750 1764 34802
rect 1708 34748 1764 34750
rect 2492 34802 2548 34804
rect 2492 34750 2494 34802
rect 2494 34750 2546 34802
rect 2546 34750 2548 34802
rect 2492 34748 2548 34750
rect 2044 34690 2100 34692
rect 2044 34638 2046 34690
rect 2046 34638 2098 34690
rect 2098 34638 2100 34690
rect 2044 34636 2100 34638
rect 1708 33628 1764 33684
rect 2492 33628 2548 33684
rect 4476 33738 4532 33740
rect 4476 33686 4478 33738
rect 4478 33686 4530 33738
rect 4530 33686 4532 33738
rect 4476 33684 4532 33686
rect 4580 33738 4636 33740
rect 4580 33686 4582 33738
rect 4582 33686 4634 33738
rect 4634 33686 4636 33738
rect 4580 33684 4636 33686
rect 4684 33738 4740 33740
rect 4684 33686 4686 33738
rect 4686 33686 4738 33738
rect 4738 33686 4740 33738
rect 4684 33684 4740 33686
rect 2044 33292 2100 33348
rect 2044 33122 2100 33124
rect 2044 33070 2046 33122
rect 2046 33070 2098 33122
rect 2098 33070 2100 33122
rect 2044 33068 2100 33070
rect 1708 32508 1764 32564
rect 2492 32508 2548 32564
rect 4476 32170 4532 32172
rect 4476 32118 4478 32170
rect 4478 32118 4530 32170
rect 4530 32118 4532 32170
rect 4476 32116 4532 32118
rect 4580 32170 4636 32172
rect 4580 32118 4582 32170
rect 4582 32118 4634 32170
rect 4634 32118 4636 32170
rect 4580 32116 4636 32118
rect 4684 32170 4740 32172
rect 4684 32118 4686 32170
rect 4686 32118 4738 32170
rect 4738 32118 4740 32170
rect 4684 32116 4740 32118
rect 2044 31554 2100 31556
rect 2044 31502 2046 31554
rect 2046 31502 2098 31554
rect 2098 31502 2100 31554
rect 2044 31500 2100 31502
rect 1708 31388 1764 31444
rect 2492 31388 2548 31444
rect 2044 31106 2100 31108
rect 2044 31054 2046 31106
rect 2046 31054 2098 31106
rect 2098 31054 2100 31106
rect 2044 31052 2100 31054
rect 1708 30828 1764 30884
rect 2492 30882 2548 30884
rect 2492 30830 2494 30882
rect 2494 30830 2546 30882
rect 2546 30830 2548 30882
rect 2492 30828 2548 30830
rect 4476 30602 4532 30604
rect 4476 30550 4478 30602
rect 4478 30550 4530 30602
rect 4530 30550 4532 30602
rect 4476 30548 4532 30550
rect 4580 30602 4636 30604
rect 4580 30550 4582 30602
rect 4582 30550 4634 30602
rect 4634 30550 4636 30602
rect 4580 30548 4636 30550
rect 4684 30602 4740 30604
rect 4684 30550 4686 30602
rect 4686 30550 4738 30602
rect 4738 30550 4740 30602
rect 4684 30548 4740 30550
rect 1708 30268 1764 30324
rect 2044 29538 2100 29540
rect 2044 29486 2046 29538
rect 2046 29486 2098 29538
rect 2098 29486 2100 29538
rect 2044 29484 2100 29486
rect 1708 29148 1764 29204
rect 2492 29148 2548 29204
rect 4476 29034 4532 29036
rect 4476 28982 4478 29034
rect 4478 28982 4530 29034
rect 4530 28982 4532 29034
rect 4476 28980 4532 28982
rect 4580 29034 4636 29036
rect 4580 28982 4582 29034
rect 4582 28982 4634 29034
rect 4634 28982 4636 29034
rect 4580 28980 4636 28982
rect 4684 29034 4740 29036
rect 4684 28982 4686 29034
rect 4686 28982 4738 29034
rect 4738 28982 4740 29034
rect 4684 28980 4740 28982
rect 2044 28588 2100 28644
rect 1708 28028 1764 28084
rect 2492 28028 2548 28084
rect 5404 27692 5460 27748
rect 2044 27580 2100 27636
rect 1708 26962 1764 26964
rect 1708 26910 1710 26962
rect 1710 26910 1762 26962
rect 1762 26910 1764 26962
rect 1708 26908 1764 26910
rect 4476 27466 4532 27468
rect 4476 27414 4478 27466
rect 4478 27414 4530 27466
rect 4530 27414 4532 27466
rect 4476 27412 4532 27414
rect 4580 27466 4636 27468
rect 4580 27414 4582 27466
rect 4582 27414 4634 27466
rect 4634 27414 4636 27466
rect 4580 27412 4636 27414
rect 4684 27466 4740 27468
rect 4684 27414 4686 27466
rect 4686 27414 4738 27466
rect 4738 27414 4740 27466
rect 4684 27412 4740 27414
rect 2492 26962 2548 26964
rect 2492 26910 2494 26962
rect 2494 26910 2546 26962
rect 2546 26910 2548 26962
rect 2492 26908 2548 26910
rect 2156 26460 2212 26516
rect 2044 26402 2100 26404
rect 2044 26350 2046 26402
rect 2046 26350 2098 26402
rect 2098 26350 2100 26402
rect 2044 26348 2100 26350
rect 1708 25788 1764 25844
rect 2492 25788 2548 25844
rect 4476 25898 4532 25900
rect 4476 25846 4478 25898
rect 4478 25846 4530 25898
rect 4530 25846 4532 25898
rect 4476 25844 4532 25846
rect 4580 25898 4636 25900
rect 4580 25846 4582 25898
rect 4582 25846 4634 25898
rect 4634 25846 4636 25898
rect 4580 25844 4636 25846
rect 4684 25898 4740 25900
rect 4684 25846 4686 25898
rect 4686 25846 4738 25898
rect 4738 25846 4740 25898
rect 4684 25844 4740 25846
rect 1708 24668 1764 24724
rect 2492 24668 2548 24724
rect 4476 24330 4532 24332
rect 4476 24278 4478 24330
rect 4478 24278 4530 24330
rect 4530 24278 4532 24330
rect 4476 24276 4532 24278
rect 4580 24330 4636 24332
rect 4580 24278 4582 24330
rect 4582 24278 4634 24330
rect 4634 24278 4636 24330
rect 4580 24276 4636 24278
rect 4684 24330 4740 24332
rect 4684 24278 4686 24330
rect 4686 24278 4738 24330
rect 4738 24278 4740 24330
rect 4684 24276 4740 24278
rect 2044 23996 2100 24052
rect 1708 23548 1764 23604
rect 2492 23548 2548 23604
rect 11564 23548 11620 23604
rect 2156 23436 2212 23492
rect 1708 22988 1764 23044
rect 2044 22876 2100 22932
rect 2492 23042 2548 23044
rect 2492 22990 2494 23042
rect 2494 22990 2546 23042
rect 2546 22990 2548 23042
rect 2492 22988 2548 22990
rect 4476 22762 4532 22764
rect 4476 22710 4478 22762
rect 4478 22710 4530 22762
rect 4530 22710 4532 22762
rect 4476 22708 4532 22710
rect 4580 22762 4636 22764
rect 4580 22710 4582 22762
rect 4582 22710 4634 22762
rect 4634 22710 4636 22762
rect 4580 22708 4636 22710
rect 4684 22762 4740 22764
rect 4684 22710 4686 22762
rect 4686 22710 4738 22762
rect 4738 22710 4740 22762
rect 4684 22708 4740 22710
rect 1708 22428 1764 22484
rect 2156 21756 2212 21812
rect 1708 21308 1764 21364
rect 2492 21308 2548 21364
rect 4476 21194 4532 21196
rect 4476 21142 4478 21194
rect 4478 21142 4530 21194
rect 4530 21142 4532 21194
rect 4476 21140 4532 21142
rect 4580 21194 4636 21196
rect 4580 21142 4582 21194
rect 4582 21142 4634 21194
rect 4634 21142 4636 21194
rect 4580 21140 4636 21142
rect 4684 21194 4740 21196
rect 4684 21142 4686 21194
rect 4686 21142 4738 21194
rect 4738 21142 4740 21194
rect 4684 21140 4740 21142
rect 1708 20188 1764 20244
rect 2044 20300 2100 20356
rect 1708 19122 1764 19124
rect 1708 19070 1710 19122
rect 1710 19070 1762 19122
rect 1762 19070 1764 19122
rect 1708 19068 1764 19070
rect 2492 20188 2548 20244
rect 7532 19740 7588 19796
rect 4476 19626 4532 19628
rect 4476 19574 4478 19626
rect 4478 19574 4530 19626
rect 4530 19574 4532 19626
rect 4476 19572 4532 19574
rect 4580 19626 4636 19628
rect 4580 19574 4582 19626
rect 4582 19574 4634 19626
rect 4634 19574 4636 19626
rect 4580 19572 4636 19574
rect 4684 19626 4740 19628
rect 4684 19574 4686 19626
rect 4686 19574 4738 19626
rect 4738 19574 4740 19626
rect 4684 19572 4740 19574
rect 2492 19122 2548 19124
rect 2492 19070 2494 19122
rect 2494 19070 2546 19122
rect 2546 19070 2548 19122
rect 2492 19068 2548 19070
rect 1708 17948 1764 18004
rect 2492 17948 2548 18004
rect 4476 18058 4532 18060
rect 4476 18006 4478 18058
rect 4478 18006 4530 18058
rect 4530 18006 4532 18058
rect 4476 18004 4532 18006
rect 4580 18058 4636 18060
rect 4580 18006 4582 18058
rect 4582 18006 4634 18058
rect 4634 18006 4636 18058
rect 4580 18004 4636 18006
rect 4684 18058 4740 18060
rect 4684 18006 4686 18058
rect 4686 18006 4738 18058
rect 4738 18006 4740 18058
rect 4684 18004 4740 18006
rect 2044 17836 2100 17892
rect 1708 17388 1764 17444
rect 2492 17442 2548 17444
rect 2492 17390 2494 17442
rect 2494 17390 2546 17442
rect 2546 17390 2548 17442
rect 2492 17388 2548 17390
rect 2044 17052 2100 17108
rect 1708 16828 1764 16884
rect 4476 16490 4532 16492
rect 4476 16438 4478 16490
rect 4478 16438 4530 16490
rect 4530 16438 4532 16490
rect 4476 16436 4532 16438
rect 4580 16490 4636 16492
rect 4580 16438 4582 16490
rect 4582 16438 4634 16490
rect 4634 16438 4636 16490
rect 4580 16436 4636 16438
rect 4684 16490 4740 16492
rect 4684 16438 4686 16490
rect 4686 16438 4738 16490
rect 4738 16438 4740 16490
rect 4684 16436 4740 16438
rect 2044 16268 2100 16324
rect 1932 16044 1988 16100
rect 1708 15708 1764 15764
rect 1708 14588 1764 14644
rect 1708 13468 1764 13524
rect 1708 12348 1764 12404
rect 1708 11282 1764 11284
rect 1708 11230 1710 11282
rect 1710 11230 1762 11282
rect 1762 11230 1764 11282
rect 1708 11228 1764 11230
rect 1708 10108 1764 10164
rect 1708 9548 1764 9604
rect 1708 8988 1764 9044
rect 1708 7868 1764 7924
rect 1708 7308 1764 7364
rect 1708 6748 1764 6804
rect 5964 15932 6020 15988
rect 2492 15708 2548 15764
rect 2044 15426 2100 15428
rect 2044 15374 2046 15426
rect 2046 15374 2098 15426
rect 2098 15374 2100 15426
rect 2044 15372 2100 15374
rect 2156 14700 2212 14756
rect 2044 13970 2100 13972
rect 2044 13918 2046 13970
rect 2046 13918 2098 13970
rect 2098 13918 2100 13970
rect 2044 13916 2100 13918
rect 4476 14922 4532 14924
rect 4476 14870 4478 14922
rect 4478 14870 4530 14922
rect 4530 14870 4532 14922
rect 4476 14868 4532 14870
rect 4580 14922 4636 14924
rect 4580 14870 4582 14922
rect 4582 14870 4634 14922
rect 4634 14870 4636 14922
rect 4580 14868 4636 14870
rect 4684 14922 4740 14924
rect 4684 14870 4686 14922
rect 4686 14870 4738 14922
rect 4738 14870 4740 14922
rect 4684 14868 4740 14870
rect 2492 14588 2548 14644
rect 2492 13468 2548 13524
rect 4476 13354 4532 13356
rect 4476 13302 4478 13354
rect 4478 13302 4530 13354
rect 4530 13302 4532 13354
rect 4476 13300 4532 13302
rect 4580 13354 4636 13356
rect 4580 13302 4582 13354
rect 4582 13302 4634 13354
rect 4634 13302 4636 13354
rect 4580 13300 4636 13302
rect 4684 13354 4740 13356
rect 4684 13302 4686 13354
rect 4686 13302 4738 13354
rect 4738 13302 4740 13354
rect 4684 13300 4740 13302
rect 2492 12348 2548 12404
rect 2156 12236 2212 12292
rect 2044 11170 2100 11172
rect 2044 11118 2046 11170
rect 2046 11118 2098 11170
rect 2098 11118 2100 11170
rect 2044 11116 2100 11118
rect 4476 11786 4532 11788
rect 4476 11734 4478 11786
rect 4478 11734 4530 11786
rect 4530 11734 4532 11786
rect 4476 11732 4532 11734
rect 4580 11786 4636 11788
rect 4580 11734 4582 11786
rect 4582 11734 4634 11786
rect 4634 11734 4636 11786
rect 4580 11732 4636 11734
rect 4684 11786 4740 11788
rect 4684 11734 4686 11786
rect 4686 11734 4738 11786
rect 4738 11734 4740 11786
rect 4684 11732 4740 11734
rect 2492 11282 2548 11284
rect 2492 11230 2494 11282
rect 2494 11230 2546 11282
rect 2546 11230 2548 11282
rect 2492 11228 2548 11230
rect 2380 10892 2436 10948
rect 2044 9996 2100 10052
rect 2492 10108 2548 10164
rect 4476 10218 4532 10220
rect 4476 10166 4478 10218
rect 4478 10166 4530 10218
rect 4530 10166 4532 10218
rect 4476 10164 4532 10166
rect 4580 10218 4636 10220
rect 4580 10166 4582 10218
rect 4582 10166 4634 10218
rect 4634 10166 4636 10218
rect 4580 10164 4636 10166
rect 4684 10218 4740 10220
rect 4684 10166 4686 10218
rect 4686 10166 4738 10218
rect 4738 10166 4740 10218
rect 4684 10164 4740 10166
rect 2492 9602 2548 9604
rect 2492 9550 2494 9602
rect 2494 9550 2546 9602
rect 2546 9550 2548 9602
rect 2492 9548 2548 9550
rect 4476 8650 4532 8652
rect 4476 8598 4478 8650
rect 4478 8598 4530 8650
rect 4530 8598 4532 8650
rect 4476 8596 4532 8598
rect 4580 8650 4636 8652
rect 4580 8598 4582 8650
rect 4582 8598 4634 8650
rect 4634 8598 4636 8650
rect 4580 8596 4636 8598
rect 4684 8650 4740 8652
rect 4684 8598 4686 8650
rect 4686 8598 4738 8650
rect 4738 8598 4740 8650
rect 4684 8596 4740 8598
rect 2492 7868 2548 7924
rect 2044 7698 2100 7700
rect 2044 7646 2046 7698
rect 2046 7646 2098 7698
rect 2098 7646 2100 7698
rect 2044 7644 2100 7646
rect 2492 7362 2548 7364
rect 2492 7310 2494 7362
rect 2494 7310 2546 7362
rect 2546 7310 2548 7362
rect 2492 7308 2548 7310
rect 4476 7082 4532 7084
rect 4476 7030 4478 7082
rect 4478 7030 4530 7082
rect 4530 7030 4532 7082
rect 4476 7028 4532 7030
rect 4580 7082 4636 7084
rect 4580 7030 4582 7082
rect 4582 7030 4634 7082
rect 4634 7030 4636 7082
rect 4580 7028 4636 7030
rect 4684 7082 4740 7084
rect 4684 7030 4686 7082
rect 4686 7030 4738 7082
rect 4738 7030 4740 7082
rect 4684 7028 4740 7030
rect 2716 6748 2772 6804
rect 1708 5628 1764 5684
rect 2044 5740 2100 5796
rect 2492 5628 2548 5684
rect 1708 4508 1764 4564
rect 2044 4732 2100 4788
rect 1708 3442 1764 3444
rect 1708 3390 1710 3442
rect 1710 3390 1762 3442
rect 1762 3390 1764 3442
rect 1708 3388 1764 3390
rect 2492 4508 2548 4564
rect 4284 5628 4340 5684
rect 3164 3442 3220 3444
rect 3164 3390 3166 3442
rect 3166 3390 3218 3442
rect 3218 3390 3220 3442
rect 3164 3388 3220 3390
rect 4476 5514 4532 5516
rect 4476 5462 4478 5514
rect 4478 5462 4530 5514
rect 4530 5462 4532 5514
rect 4476 5460 4532 5462
rect 4580 5514 4636 5516
rect 4580 5462 4582 5514
rect 4582 5462 4634 5514
rect 4634 5462 4636 5514
rect 4580 5460 4636 5462
rect 4684 5514 4740 5516
rect 4684 5462 4686 5514
rect 4686 5462 4738 5514
rect 4738 5462 4740 5514
rect 4684 5460 4740 5462
rect 4956 5292 5012 5348
rect 4476 3946 4532 3948
rect 4476 3894 4478 3946
rect 4478 3894 4530 3946
rect 4530 3894 4532 3946
rect 4476 3892 4532 3894
rect 4580 3946 4636 3948
rect 4580 3894 4582 3946
rect 4582 3894 4634 3946
rect 4634 3894 4636 3946
rect 4580 3892 4636 3894
rect 4684 3946 4740 3948
rect 4684 3894 4686 3946
rect 4686 3894 4738 3946
rect 4738 3894 4740 3946
rect 4684 3892 4740 3894
rect 4732 3388 4788 3444
rect 5180 4898 5236 4900
rect 5180 4846 5182 4898
rect 5182 4846 5234 4898
rect 5234 4846 5236 4898
rect 5180 4844 5236 4846
rect 6972 14476 7028 14532
rect 6636 13020 6692 13076
rect 6636 7644 6692 7700
rect 6300 6412 6356 6468
rect 5964 4732 6020 4788
rect 6188 4732 6244 4788
rect 6748 5852 6804 5908
rect 6412 4844 6468 4900
rect 5628 3836 5684 3892
rect 5740 3612 5796 3668
rect 2380 2268 2436 2324
rect 5964 3612 6020 3668
rect 6076 4284 6132 4340
rect 6412 3724 6468 3780
rect 6300 3388 6356 3444
rect 7420 6860 7476 6916
rect 6972 5740 7028 5796
rect 6860 4844 6916 4900
rect 6748 3836 6804 3892
rect 7196 5740 7252 5796
rect 7084 4620 7140 4676
rect 9996 17948 10052 18004
rect 7532 6748 7588 6804
rect 8316 9548 8372 9604
rect 8876 8428 8932 8484
rect 8428 6802 8484 6804
rect 8428 6750 8430 6802
rect 8430 6750 8482 6802
rect 8482 6750 8484 6802
rect 8428 6748 8484 6750
rect 7420 5404 7476 5460
rect 7644 4450 7700 4452
rect 7644 4398 7646 4450
rect 7646 4398 7698 4450
rect 7698 4398 7700 4450
rect 7644 4396 7700 4398
rect 7420 4060 7476 4116
rect 7196 3554 7252 3556
rect 7196 3502 7198 3554
rect 7198 3502 7250 3554
rect 7250 3502 7252 3554
rect 7196 3500 7252 3502
rect 7644 3836 7700 3892
rect 8204 6466 8260 6468
rect 8204 6414 8206 6466
rect 8206 6414 8258 6466
rect 8258 6414 8260 6466
rect 8204 6412 8260 6414
rect 8316 6076 8372 6132
rect 7868 5516 7924 5572
rect 7980 4508 8036 4564
rect 7980 4338 8036 4340
rect 7980 4286 7982 4338
rect 7982 4286 8034 4338
rect 8034 4286 8036 4338
rect 7980 4284 8036 4286
rect 8204 5180 8260 5236
rect 8652 5906 8708 5908
rect 8652 5854 8654 5906
rect 8654 5854 8706 5906
rect 8706 5854 8708 5906
rect 8652 5852 8708 5854
rect 9884 12066 9940 12068
rect 9884 12014 9886 12066
rect 9886 12014 9938 12066
rect 9938 12014 9940 12066
rect 9884 12012 9940 12014
rect 9996 10892 10052 10948
rect 10108 14588 10164 14644
rect 9436 10444 9492 10500
rect 9548 9714 9604 9716
rect 9548 9662 9550 9714
rect 9550 9662 9602 9714
rect 9602 9662 9604 9714
rect 9548 9660 9604 9662
rect 9324 9602 9380 9604
rect 9324 9550 9326 9602
rect 9326 9550 9378 9602
rect 9378 9550 9380 9602
rect 9324 9548 9380 9550
rect 13356 76354 13412 76356
rect 13356 76302 13358 76354
rect 13358 76302 13410 76354
rect 13410 76302 13412 76354
rect 13356 76300 13412 76302
rect 12572 75852 12628 75908
rect 12572 75682 12628 75684
rect 12572 75630 12574 75682
rect 12574 75630 12626 75682
rect 12626 75630 12628 75682
rect 12572 75628 12628 75630
rect 13580 75682 13636 75684
rect 13580 75630 13582 75682
rect 13582 75630 13634 75682
rect 13634 75630 13636 75682
rect 13580 75628 13636 75630
rect 13916 75516 13972 75572
rect 14140 76300 14196 76356
rect 13468 74898 13524 74900
rect 13468 74846 13470 74898
rect 13470 74846 13522 74898
rect 13522 74846 13524 74898
rect 13468 74844 13524 74846
rect 14252 74844 14308 74900
rect 12684 73948 12740 74004
rect 14028 73276 14084 73332
rect 12460 24444 12516 24500
rect 11676 21644 11732 21700
rect 13468 25228 13524 25284
rect 14364 74002 14420 74004
rect 14364 73950 14366 74002
rect 14366 73950 14418 74002
rect 14418 73950 14420 74002
rect 14364 73948 14420 73950
rect 14700 75682 14756 75684
rect 14700 75630 14702 75682
rect 14702 75630 14754 75682
rect 14754 75630 14756 75682
rect 14700 75628 14756 75630
rect 15372 76690 15428 76692
rect 15372 76638 15374 76690
rect 15374 76638 15426 76690
rect 15426 76638 15428 76690
rect 15372 76636 15428 76638
rect 16604 76636 16660 76692
rect 16380 76300 16436 76356
rect 17164 76354 17220 76356
rect 17164 76302 17166 76354
rect 17166 76302 17218 76354
rect 17218 76302 17220 76354
rect 17164 76300 17220 76302
rect 16492 75628 16548 75684
rect 18060 76466 18116 76468
rect 18060 76414 18062 76466
rect 18062 76414 18114 76466
rect 18114 76414 18116 76466
rect 18060 76412 18116 76414
rect 19836 76858 19892 76860
rect 19836 76806 19838 76858
rect 19838 76806 19890 76858
rect 19890 76806 19892 76858
rect 19836 76804 19892 76806
rect 19940 76858 19996 76860
rect 19940 76806 19942 76858
rect 19942 76806 19994 76858
rect 19994 76806 19996 76858
rect 19940 76804 19996 76806
rect 20044 76858 20100 76860
rect 20044 76806 20046 76858
rect 20046 76806 20098 76858
rect 20098 76806 20100 76858
rect 20044 76804 20100 76806
rect 19404 76412 19460 76468
rect 17948 75516 18004 75572
rect 19180 75516 19236 75572
rect 16268 73276 16324 73332
rect 14252 24780 14308 24836
rect 14812 24780 14868 24836
rect 13468 23548 13524 23604
rect 13804 23548 13860 23604
rect 12796 23100 12852 23156
rect 14028 18508 14084 18564
rect 11564 11116 11620 11172
rect 10332 10498 10388 10500
rect 10332 10446 10334 10498
rect 10334 10446 10386 10498
rect 10386 10446 10388 10498
rect 10332 10444 10388 10446
rect 11788 12066 11844 12068
rect 11788 12014 11790 12066
rect 11790 12014 11842 12066
rect 11842 12014 11844 12066
rect 11788 12012 11844 12014
rect 12012 11116 12068 11172
rect 11788 10108 11844 10164
rect 10108 9996 10164 10052
rect 9324 8876 9380 8932
rect 9436 8146 9492 8148
rect 9436 8094 9438 8146
rect 9438 8094 9490 8146
rect 9490 8094 9492 8146
rect 9436 8092 9492 8094
rect 11116 9548 11172 9604
rect 10332 8930 10388 8932
rect 10332 8878 10334 8930
rect 10334 8878 10386 8930
rect 10386 8878 10388 8930
rect 10332 8876 10388 8878
rect 11004 8258 11060 8260
rect 11004 8206 11006 8258
rect 11006 8206 11058 8258
rect 11058 8206 11060 8258
rect 11004 8204 11060 8206
rect 9660 7756 9716 7812
rect 10556 7756 10612 7812
rect 9100 6802 9156 6804
rect 9100 6750 9102 6802
rect 9102 6750 9154 6802
rect 9154 6750 9156 6802
rect 9100 6748 9156 6750
rect 9772 6802 9828 6804
rect 9772 6750 9774 6802
rect 9774 6750 9826 6802
rect 9826 6750 9828 6802
rect 9772 6748 9828 6750
rect 9884 6524 9940 6580
rect 10444 6188 10500 6244
rect 9884 5906 9940 5908
rect 9884 5854 9886 5906
rect 9886 5854 9938 5906
rect 9938 5854 9940 5906
rect 9884 5852 9940 5854
rect 9548 5628 9604 5684
rect 9436 5516 9492 5572
rect 8876 5292 8932 5348
rect 9324 5404 9380 5460
rect 8764 5122 8820 5124
rect 8764 5070 8766 5122
rect 8766 5070 8818 5122
rect 8818 5070 8820 5122
rect 8764 5068 8820 5070
rect 8428 4956 8484 5012
rect 9212 5010 9268 5012
rect 9212 4958 9214 5010
rect 9214 4958 9266 5010
rect 9266 4958 9268 5010
rect 9212 4956 9268 4958
rect 8652 4898 8708 4900
rect 8652 4846 8654 4898
rect 8654 4846 8706 4898
rect 8706 4846 8708 4898
rect 8652 4844 8708 4846
rect 9548 5292 9604 5348
rect 9884 5010 9940 5012
rect 9884 4958 9886 5010
rect 9886 4958 9938 5010
rect 9938 4958 9940 5010
rect 9884 4956 9940 4958
rect 9436 4508 9492 4564
rect 8316 4450 8372 4452
rect 8316 4398 8318 4450
rect 8318 4398 8370 4450
rect 8370 4398 8372 4450
rect 8316 4396 8372 4398
rect 8764 4396 8820 4452
rect 7868 3836 7924 3892
rect 8316 3612 8372 3668
rect 8092 3442 8148 3444
rect 8092 3390 8094 3442
rect 8094 3390 8146 3442
rect 8146 3390 8148 3442
rect 8092 3388 8148 3390
rect 8764 3948 8820 4004
rect 8988 3724 9044 3780
rect 8540 3612 8596 3668
rect 8764 3164 8820 3220
rect 9772 4732 9828 4788
rect 10108 5292 10164 5348
rect 9772 4396 9828 4452
rect 9884 4284 9940 4340
rect 10332 4844 10388 4900
rect 12460 11116 12516 11172
rect 12348 9826 12404 9828
rect 12348 9774 12350 9826
rect 12350 9774 12402 9826
rect 12402 9774 12404 9826
rect 12348 9772 12404 9774
rect 11900 9714 11956 9716
rect 11900 9662 11902 9714
rect 11902 9662 11954 9714
rect 11954 9662 11956 9714
rect 11900 9660 11956 9662
rect 12012 8258 12068 8260
rect 12012 8206 12014 8258
rect 12014 8206 12066 8258
rect 12066 8206 12068 8258
rect 12012 8204 12068 8206
rect 12684 11788 12740 11844
rect 13020 11116 13076 11172
rect 13692 11452 13748 11508
rect 13468 11170 13524 11172
rect 13468 11118 13470 11170
rect 13470 11118 13522 11170
rect 13522 11118 13524 11170
rect 13468 11116 13524 11118
rect 13020 10108 13076 10164
rect 13804 10444 13860 10500
rect 13356 10108 13412 10164
rect 13468 9772 13524 9828
rect 13132 8428 13188 8484
rect 12572 8204 12628 8260
rect 11900 8146 11956 8148
rect 11900 8094 11902 8146
rect 11902 8094 11954 8146
rect 11954 8094 11956 8146
rect 11900 8092 11956 8094
rect 13020 8146 13076 8148
rect 13020 8094 13022 8146
rect 13022 8094 13074 8146
rect 13074 8094 13076 8146
rect 13020 8092 13076 8094
rect 11452 7420 11508 7476
rect 10892 6860 10948 6916
rect 10668 5964 10724 6020
rect 13468 7420 13524 7476
rect 11676 7308 11732 7364
rect 11228 6914 11284 6916
rect 11228 6862 11230 6914
rect 11230 6862 11282 6914
rect 11282 6862 11284 6914
rect 11228 6860 11284 6862
rect 10668 5180 10724 5236
rect 10892 5234 10948 5236
rect 10892 5182 10894 5234
rect 10894 5182 10946 5234
rect 10946 5182 10948 5234
rect 10892 5180 10948 5182
rect 10220 4172 10276 4228
rect 10108 4060 10164 4116
rect 10892 4060 10948 4116
rect 10332 3948 10388 4004
rect 10220 3724 10276 3780
rect 10780 3948 10836 4004
rect 10780 3724 10836 3780
rect 11004 3724 11060 3780
rect 10556 3612 10612 3668
rect 10892 3388 10948 3444
rect 11228 5964 11284 6020
rect 11228 3948 11284 4004
rect 13244 6636 13300 6692
rect 12124 6466 12180 6468
rect 12124 6414 12126 6466
rect 12126 6414 12178 6466
rect 12178 6414 12180 6466
rect 12124 6412 12180 6414
rect 11340 5292 11396 5348
rect 11228 3442 11284 3444
rect 11228 3390 11230 3442
rect 11230 3390 11282 3442
rect 11282 3390 11284 3442
rect 11228 3388 11284 3390
rect 12236 6188 12292 6244
rect 11564 5122 11620 5124
rect 11564 5070 11566 5122
rect 11566 5070 11618 5122
rect 11618 5070 11620 5122
rect 11564 5068 11620 5070
rect 11900 5122 11956 5124
rect 11900 5070 11902 5122
rect 11902 5070 11954 5122
rect 11954 5070 11956 5122
rect 11900 5068 11956 5070
rect 11452 4060 11508 4116
rect 11676 4844 11732 4900
rect 11340 2380 11396 2436
rect 11900 3442 11956 3444
rect 11900 3390 11902 3442
rect 11902 3390 11954 3442
rect 11954 3390 11956 3442
rect 11900 3388 11956 3390
rect 11900 3276 11956 3332
rect 12460 5740 12516 5796
rect 12572 5628 12628 5684
rect 13020 5964 13076 6020
rect 12460 5122 12516 5124
rect 12460 5070 12462 5122
rect 12462 5070 12514 5122
rect 12514 5070 12516 5122
rect 12460 5068 12516 5070
rect 12572 5010 12628 5012
rect 12572 4958 12574 5010
rect 12574 4958 12626 5010
rect 12626 4958 12628 5010
rect 12572 4956 12628 4958
rect 12348 4898 12404 4900
rect 12348 4846 12350 4898
rect 12350 4846 12402 4898
rect 12402 4846 12404 4898
rect 12348 4844 12404 4846
rect 12572 3948 12628 4004
rect 12348 3500 12404 3556
rect 13132 5740 13188 5796
rect 13244 6076 13300 6132
rect 13244 5292 13300 5348
rect 13468 6466 13524 6468
rect 13468 6414 13470 6466
rect 13470 6414 13522 6466
rect 13522 6414 13524 6466
rect 13468 6412 13524 6414
rect 13020 5122 13076 5124
rect 13020 5070 13022 5122
rect 13022 5070 13074 5122
rect 13074 5070 13076 5122
rect 13020 5068 13076 5070
rect 13804 9884 13860 9940
rect 13916 9772 13972 9828
rect 14028 10108 14084 10164
rect 13580 6018 13636 6020
rect 13580 5966 13582 6018
rect 13582 5966 13634 6018
rect 13634 5966 13636 6018
rect 13580 5964 13636 5966
rect 13804 8876 13860 8932
rect 14140 9884 14196 9940
rect 13692 7756 13748 7812
rect 14252 8146 14308 8148
rect 14252 8094 14254 8146
rect 14254 8094 14306 8146
rect 14306 8094 14308 8146
rect 14252 8092 14308 8094
rect 14476 11506 14532 11508
rect 14476 11454 14478 11506
rect 14478 11454 14530 11506
rect 14530 11454 14532 11506
rect 14476 11452 14532 11454
rect 14476 10498 14532 10500
rect 14476 10446 14478 10498
rect 14478 10446 14530 10498
rect 14530 10446 14532 10498
rect 14476 10444 14532 10446
rect 14700 9714 14756 9716
rect 14700 9662 14702 9714
rect 14702 9662 14754 9714
rect 14754 9662 14756 9714
rect 14700 9660 14756 9662
rect 14476 9602 14532 9604
rect 14476 9550 14478 9602
rect 14478 9550 14530 9602
rect 14530 9550 14532 9602
rect 14476 9548 14532 9550
rect 14588 8876 14644 8932
rect 14364 7868 14420 7924
rect 13916 6636 13972 6692
rect 14252 7474 14308 7476
rect 14252 7422 14254 7474
rect 14254 7422 14306 7474
rect 14306 7422 14308 7474
rect 14252 7420 14308 7422
rect 14140 6860 14196 6916
rect 14028 6412 14084 6468
rect 14476 6466 14532 6468
rect 14476 6414 14478 6466
rect 14478 6414 14530 6466
rect 14530 6414 14532 6466
rect 14476 6412 14532 6414
rect 17612 73164 17668 73220
rect 17836 73388 17892 73444
rect 16268 23548 16324 23604
rect 16604 24668 16660 24724
rect 18284 73948 18340 74004
rect 18844 74732 18900 74788
rect 18172 73388 18228 73444
rect 18060 73218 18116 73220
rect 18060 73166 18062 73218
rect 18062 73166 18114 73218
rect 18114 73166 18116 73218
rect 18060 73164 18116 73166
rect 18060 29372 18116 29428
rect 17164 24780 17220 24836
rect 17500 24722 17556 24724
rect 17500 24670 17502 24722
rect 17502 24670 17554 24722
rect 17554 24670 17556 24722
rect 17500 24668 17556 24670
rect 17612 24556 17668 24612
rect 18172 24610 18228 24612
rect 18172 24558 18174 24610
rect 18174 24558 18226 24610
rect 18226 24558 18228 24610
rect 18172 24556 18228 24558
rect 18396 24556 18452 24612
rect 17724 24220 17780 24276
rect 18396 24220 18452 24276
rect 18060 23884 18116 23940
rect 17164 23772 17220 23828
rect 16828 23212 16884 23268
rect 15596 21644 15652 21700
rect 15596 21420 15652 21476
rect 17948 23660 18004 23716
rect 17612 23436 17668 23492
rect 17500 23266 17556 23268
rect 17500 23214 17502 23266
rect 17502 23214 17554 23266
rect 17554 23214 17556 23266
rect 17500 23212 17556 23214
rect 17164 21532 17220 21588
rect 17276 21980 17332 22036
rect 16716 18508 16772 18564
rect 15372 11788 15428 11844
rect 16604 11788 16660 11844
rect 15596 11452 15652 11508
rect 14812 7420 14868 7476
rect 14924 8540 14980 8596
rect 14924 7756 14980 7812
rect 14924 6636 14980 6692
rect 15036 8092 15092 8148
rect 14700 6466 14756 6468
rect 14700 6414 14702 6466
rect 14702 6414 14754 6466
rect 14754 6414 14756 6466
rect 14700 6412 14756 6414
rect 15372 8540 15428 8596
rect 15596 8988 15652 9044
rect 15484 7474 15540 7476
rect 15484 7422 15486 7474
rect 15486 7422 15538 7474
rect 15538 7422 15540 7474
rect 15484 7420 15540 7422
rect 15260 7362 15316 7364
rect 15260 7310 15262 7362
rect 15262 7310 15314 7362
rect 15314 7310 15316 7362
rect 15260 7308 15316 7310
rect 13916 6018 13972 6020
rect 13916 5966 13918 6018
rect 13918 5966 13970 6018
rect 13970 5966 13972 6018
rect 13916 5964 13972 5966
rect 14476 5906 14532 5908
rect 14476 5854 14478 5906
rect 14478 5854 14530 5906
rect 14530 5854 14532 5906
rect 14476 5852 14532 5854
rect 13692 5516 13748 5572
rect 13692 5292 13748 5348
rect 13580 5234 13636 5236
rect 13580 5182 13582 5234
rect 13582 5182 13634 5234
rect 13634 5182 13636 5234
rect 13580 5180 13636 5182
rect 13468 4844 13524 4900
rect 13468 4396 13524 4452
rect 13356 4172 13412 4228
rect 14364 5516 14420 5572
rect 14028 5292 14084 5348
rect 13916 5180 13972 5236
rect 13916 4956 13972 5012
rect 14140 5122 14196 5124
rect 14140 5070 14142 5122
rect 14142 5070 14194 5122
rect 14194 5070 14196 5122
rect 14140 5068 14196 5070
rect 14812 5964 14868 6020
rect 14812 5516 14868 5572
rect 15260 5404 15316 5460
rect 15372 5628 15428 5684
rect 15148 5292 15204 5348
rect 14700 5068 14756 5124
rect 14252 4508 14308 4564
rect 14140 3554 14196 3556
rect 14140 3502 14142 3554
rect 14142 3502 14194 3554
rect 14194 3502 14196 3554
rect 14140 3500 14196 3502
rect 14588 3724 14644 3780
rect 14812 4450 14868 4452
rect 14812 4398 14814 4450
rect 14814 4398 14866 4450
rect 14866 4398 14868 4450
rect 14812 4396 14868 4398
rect 14700 3388 14756 3444
rect 14812 3836 14868 3892
rect 15036 3836 15092 3892
rect 15372 4956 15428 5012
rect 15820 7980 15876 8036
rect 15708 6466 15764 6468
rect 15708 6414 15710 6466
rect 15710 6414 15762 6466
rect 15762 6414 15764 6466
rect 15708 6412 15764 6414
rect 15484 4732 15540 4788
rect 15372 3554 15428 3556
rect 15372 3502 15374 3554
rect 15374 3502 15426 3554
rect 15426 3502 15428 3554
rect 15372 3500 15428 3502
rect 16156 9212 16212 9268
rect 16716 9324 16772 9380
rect 16044 8092 16100 8148
rect 16380 8540 16436 8596
rect 16156 6578 16212 6580
rect 16156 6526 16158 6578
rect 16158 6526 16210 6578
rect 16210 6526 16212 6578
rect 16156 6524 16212 6526
rect 15484 3276 15540 3332
rect 16156 6076 16212 6132
rect 15596 3724 15652 3780
rect 14364 2268 14420 2324
rect 15148 3164 15204 3220
rect 16716 8428 16772 8484
rect 16492 8316 16548 8372
rect 16380 6690 16436 6692
rect 16380 6638 16382 6690
rect 16382 6638 16434 6690
rect 16434 6638 16436 6690
rect 16380 6636 16436 6638
rect 16492 4508 16548 4564
rect 17052 7308 17108 7364
rect 16828 5740 16884 5796
rect 16492 4338 16548 4340
rect 16492 4286 16494 4338
rect 16494 4286 16546 4338
rect 16546 4286 16548 4338
rect 16492 4284 16548 4286
rect 16828 4284 16884 4340
rect 16828 4114 16884 4116
rect 16828 4062 16830 4114
rect 16830 4062 16882 4114
rect 16882 4062 16884 4114
rect 16828 4060 16884 4062
rect 17164 6690 17220 6692
rect 17164 6638 17166 6690
rect 17166 6638 17218 6690
rect 17218 6638 17220 6690
rect 17164 6636 17220 6638
rect 17052 4732 17108 4788
rect 17164 6300 17220 6356
rect 16940 3724 16996 3780
rect 17052 4172 17108 4228
rect 17948 21980 18004 22036
rect 17948 21586 18004 21588
rect 17948 21534 17950 21586
rect 17950 21534 18002 21586
rect 18002 21534 18004 21586
rect 17948 21532 18004 21534
rect 17724 21308 17780 21364
rect 18508 23826 18564 23828
rect 18508 23774 18510 23826
rect 18510 23774 18562 23826
rect 18562 23774 18564 23826
rect 18508 23772 18564 23774
rect 18732 23772 18788 23828
rect 18620 23436 18676 23492
rect 18732 22092 18788 22148
rect 18396 21308 18452 21364
rect 18620 20802 18676 20804
rect 18620 20750 18622 20802
rect 18622 20750 18674 20802
rect 18674 20750 18676 20802
rect 18620 20748 18676 20750
rect 18396 20130 18452 20132
rect 18396 20078 18398 20130
rect 18398 20078 18450 20130
rect 18450 20078 18452 20130
rect 18396 20076 18452 20078
rect 18172 18620 18228 18676
rect 18060 18226 18116 18228
rect 18060 18174 18062 18226
rect 18062 18174 18114 18226
rect 18114 18174 18116 18226
rect 18060 18172 18116 18174
rect 17388 9042 17444 9044
rect 17388 8990 17390 9042
rect 17390 8990 17442 9042
rect 17442 8990 17444 9042
rect 17388 8988 17444 8990
rect 18060 13580 18116 13636
rect 21084 76690 21140 76692
rect 21084 76638 21086 76690
rect 21086 76638 21138 76690
rect 21138 76638 21140 76690
rect 21084 76636 21140 76638
rect 20636 75852 20692 75908
rect 20748 76300 20804 76356
rect 21980 76636 22036 76692
rect 19836 75290 19892 75292
rect 19836 75238 19838 75290
rect 19838 75238 19890 75290
rect 19890 75238 19892 75290
rect 19836 75236 19892 75238
rect 19940 75290 19996 75292
rect 19940 75238 19942 75290
rect 19942 75238 19994 75290
rect 19994 75238 19996 75290
rect 19940 75236 19996 75238
rect 20044 75290 20100 75292
rect 20044 75238 20046 75290
rect 20046 75238 20098 75290
rect 20098 75238 20100 75290
rect 20044 75236 20100 75238
rect 19852 74786 19908 74788
rect 19852 74734 19854 74786
rect 19854 74734 19906 74786
rect 19906 74734 19908 74786
rect 19852 74732 19908 74734
rect 20300 74732 20356 74788
rect 19836 73722 19892 73724
rect 19836 73670 19838 73722
rect 19838 73670 19890 73722
rect 19890 73670 19892 73722
rect 19836 73668 19892 73670
rect 19940 73722 19996 73724
rect 19940 73670 19942 73722
rect 19942 73670 19994 73722
rect 19994 73670 19996 73722
rect 19940 73668 19996 73670
rect 20044 73722 20100 73724
rect 20044 73670 20046 73722
rect 20046 73670 20098 73722
rect 20098 73670 20100 73722
rect 20044 73668 20100 73670
rect 19836 72154 19892 72156
rect 19836 72102 19838 72154
rect 19838 72102 19890 72154
rect 19890 72102 19892 72154
rect 19836 72100 19892 72102
rect 19940 72154 19996 72156
rect 19940 72102 19942 72154
rect 19942 72102 19994 72154
rect 19994 72102 19996 72154
rect 19940 72100 19996 72102
rect 20044 72154 20100 72156
rect 20044 72102 20046 72154
rect 20046 72102 20098 72154
rect 20098 72102 20100 72154
rect 20044 72100 20100 72102
rect 19836 70586 19892 70588
rect 19836 70534 19838 70586
rect 19838 70534 19890 70586
rect 19890 70534 19892 70586
rect 19836 70532 19892 70534
rect 19940 70586 19996 70588
rect 19940 70534 19942 70586
rect 19942 70534 19994 70586
rect 19994 70534 19996 70586
rect 19940 70532 19996 70534
rect 20044 70586 20100 70588
rect 20044 70534 20046 70586
rect 20046 70534 20098 70586
rect 20098 70534 20100 70586
rect 20044 70532 20100 70534
rect 19836 69018 19892 69020
rect 19836 68966 19838 69018
rect 19838 68966 19890 69018
rect 19890 68966 19892 69018
rect 19836 68964 19892 68966
rect 19940 69018 19996 69020
rect 19940 68966 19942 69018
rect 19942 68966 19994 69018
rect 19994 68966 19996 69018
rect 19940 68964 19996 68966
rect 20044 69018 20100 69020
rect 20044 68966 20046 69018
rect 20046 68966 20098 69018
rect 20098 68966 20100 69018
rect 20044 68964 20100 68966
rect 19836 67450 19892 67452
rect 19836 67398 19838 67450
rect 19838 67398 19890 67450
rect 19890 67398 19892 67450
rect 19836 67396 19892 67398
rect 19940 67450 19996 67452
rect 19940 67398 19942 67450
rect 19942 67398 19994 67450
rect 19994 67398 19996 67450
rect 19940 67396 19996 67398
rect 20044 67450 20100 67452
rect 20044 67398 20046 67450
rect 20046 67398 20098 67450
rect 20098 67398 20100 67450
rect 20044 67396 20100 67398
rect 19836 65882 19892 65884
rect 19836 65830 19838 65882
rect 19838 65830 19890 65882
rect 19890 65830 19892 65882
rect 19836 65828 19892 65830
rect 19940 65882 19996 65884
rect 19940 65830 19942 65882
rect 19942 65830 19994 65882
rect 19994 65830 19996 65882
rect 19940 65828 19996 65830
rect 20044 65882 20100 65884
rect 20044 65830 20046 65882
rect 20046 65830 20098 65882
rect 20098 65830 20100 65882
rect 20044 65828 20100 65830
rect 19836 64314 19892 64316
rect 19836 64262 19838 64314
rect 19838 64262 19890 64314
rect 19890 64262 19892 64314
rect 19836 64260 19892 64262
rect 19940 64314 19996 64316
rect 19940 64262 19942 64314
rect 19942 64262 19994 64314
rect 19994 64262 19996 64314
rect 19940 64260 19996 64262
rect 20044 64314 20100 64316
rect 20044 64262 20046 64314
rect 20046 64262 20098 64314
rect 20098 64262 20100 64314
rect 20044 64260 20100 64262
rect 19836 62746 19892 62748
rect 19836 62694 19838 62746
rect 19838 62694 19890 62746
rect 19890 62694 19892 62746
rect 19836 62692 19892 62694
rect 19940 62746 19996 62748
rect 19940 62694 19942 62746
rect 19942 62694 19994 62746
rect 19994 62694 19996 62746
rect 19940 62692 19996 62694
rect 20044 62746 20100 62748
rect 20044 62694 20046 62746
rect 20046 62694 20098 62746
rect 20098 62694 20100 62746
rect 20044 62692 20100 62694
rect 19836 61178 19892 61180
rect 19836 61126 19838 61178
rect 19838 61126 19890 61178
rect 19890 61126 19892 61178
rect 19836 61124 19892 61126
rect 19940 61178 19996 61180
rect 19940 61126 19942 61178
rect 19942 61126 19994 61178
rect 19994 61126 19996 61178
rect 19940 61124 19996 61126
rect 20044 61178 20100 61180
rect 20044 61126 20046 61178
rect 20046 61126 20098 61178
rect 20098 61126 20100 61178
rect 20044 61124 20100 61126
rect 19836 59610 19892 59612
rect 19836 59558 19838 59610
rect 19838 59558 19890 59610
rect 19890 59558 19892 59610
rect 19836 59556 19892 59558
rect 19940 59610 19996 59612
rect 19940 59558 19942 59610
rect 19942 59558 19994 59610
rect 19994 59558 19996 59610
rect 19940 59556 19996 59558
rect 20044 59610 20100 59612
rect 20044 59558 20046 59610
rect 20046 59558 20098 59610
rect 20098 59558 20100 59610
rect 20044 59556 20100 59558
rect 19836 58042 19892 58044
rect 19836 57990 19838 58042
rect 19838 57990 19890 58042
rect 19890 57990 19892 58042
rect 19836 57988 19892 57990
rect 19940 58042 19996 58044
rect 19940 57990 19942 58042
rect 19942 57990 19994 58042
rect 19994 57990 19996 58042
rect 19940 57988 19996 57990
rect 20044 58042 20100 58044
rect 20044 57990 20046 58042
rect 20046 57990 20098 58042
rect 20098 57990 20100 58042
rect 20044 57988 20100 57990
rect 19836 56474 19892 56476
rect 19836 56422 19838 56474
rect 19838 56422 19890 56474
rect 19890 56422 19892 56474
rect 19836 56420 19892 56422
rect 19940 56474 19996 56476
rect 19940 56422 19942 56474
rect 19942 56422 19994 56474
rect 19994 56422 19996 56474
rect 19940 56420 19996 56422
rect 20044 56474 20100 56476
rect 20044 56422 20046 56474
rect 20046 56422 20098 56474
rect 20098 56422 20100 56474
rect 20044 56420 20100 56422
rect 19180 23042 19236 23044
rect 19180 22990 19182 23042
rect 19182 22990 19234 23042
rect 19234 22990 19236 23042
rect 19180 22988 19236 22990
rect 19180 21980 19236 22036
rect 19836 54906 19892 54908
rect 19836 54854 19838 54906
rect 19838 54854 19890 54906
rect 19890 54854 19892 54906
rect 19836 54852 19892 54854
rect 19940 54906 19996 54908
rect 19940 54854 19942 54906
rect 19942 54854 19994 54906
rect 19994 54854 19996 54906
rect 19940 54852 19996 54854
rect 20044 54906 20100 54908
rect 20044 54854 20046 54906
rect 20046 54854 20098 54906
rect 20098 54854 20100 54906
rect 20044 54852 20100 54854
rect 19836 53338 19892 53340
rect 19836 53286 19838 53338
rect 19838 53286 19890 53338
rect 19890 53286 19892 53338
rect 19836 53284 19892 53286
rect 19940 53338 19996 53340
rect 19940 53286 19942 53338
rect 19942 53286 19994 53338
rect 19994 53286 19996 53338
rect 19940 53284 19996 53286
rect 20044 53338 20100 53340
rect 20044 53286 20046 53338
rect 20046 53286 20098 53338
rect 20098 53286 20100 53338
rect 20044 53284 20100 53286
rect 19836 51770 19892 51772
rect 19836 51718 19838 51770
rect 19838 51718 19890 51770
rect 19890 51718 19892 51770
rect 19836 51716 19892 51718
rect 19940 51770 19996 51772
rect 19940 51718 19942 51770
rect 19942 51718 19994 51770
rect 19994 51718 19996 51770
rect 19940 51716 19996 51718
rect 20044 51770 20100 51772
rect 20044 51718 20046 51770
rect 20046 51718 20098 51770
rect 20098 51718 20100 51770
rect 20044 51716 20100 51718
rect 19836 50202 19892 50204
rect 19836 50150 19838 50202
rect 19838 50150 19890 50202
rect 19890 50150 19892 50202
rect 19836 50148 19892 50150
rect 19940 50202 19996 50204
rect 19940 50150 19942 50202
rect 19942 50150 19994 50202
rect 19994 50150 19996 50202
rect 19940 50148 19996 50150
rect 20044 50202 20100 50204
rect 20044 50150 20046 50202
rect 20046 50150 20098 50202
rect 20098 50150 20100 50202
rect 20044 50148 20100 50150
rect 19836 48634 19892 48636
rect 19836 48582 19838 48634
rect 19838 48582 19890 48634
rect 19890 48582 19892 48634
rect 19836 48580 19892 48582
rect 19940 48634 19996 48636
rect 19940 48582 19942 48634
rect 19942 48582 19994 48634
rect 19994 48582 19996 48634
rect 19940 48580 19996 48582
rect 20044 48634 20100 48636
rect 20044 48582 20046 48634
rect 20046 48582 20098 48634
rect 20098 48582 20100 48634
rect 20044 48580 20100 48582
rect 19836 47066 19892 47068
rect 19836 47014 19838 47066
rect 19838 47014 19890 47066
rect 19890 47014 19892 47066
rect 19836 47012 19892 47014
rect 19940 47066 19996 47068
rect 19940 47014 19942 47066
rect 19942 47014 19994 47066
rect 19994 47014 19996 47066
rect 19940 47012 19996 47014
rect 20044 47066 20100 47068
rect 20044 47014 20046 47066
rect 20046 47014 20098 47066
rect 20098 47014 20100 47066
rect 20044 47012 20100 47014
rect 19836 45498 19892 45500
rect 19836 45446 19838 45498
rect 19838 45446 19890 45498
rect 19890 45446 19892 45498
rect 19836 45444 19892 45446
rect 19940 45498 19996 45500
rect 19940 45446 19942 45498
rect 19942 45446 19994 45498
rect 19994 45446 19996 45498
rect 19940 45444 19996 45446
rect 20044 45498 20100 45500
rect 20044 45446 20046 45498
rect 20046 45446 20098 45498
rect 20098 45446 20100 45498
rect 20044 45444 20100 45446
rect 19836 43930 19892 43932
rect 19836 43878 19838 43930
rect 19838 43878 19890 43930
rect 19890 43878 19892 43930
rect 19836 43876 19892 43878
rect 19940 43930 19996 43932
rect 19940 43878 19942 43930
rect 19942 43878 19994 43930
rect 19994 43878 19996 43930
rect 19940 43876 19996 43878
rect 20044 43930 20100 43932
rect 20044 43878 20046 43930
rect 20046 43878 20098 43930
rect 20098 43878 20100 43930
rect 20044 43876 20100 43878
rect 19836 42362 19892 42364
rect 19836 42310 19838 42362
rect 19838 42310 19890 42362
rect 19890 42310 19892 42362
rect 19836 42308 19892 42310
rect 19940 42362 19996 42364
rect 19940 42310 19942 42362
rect 19942 42310 19994 42362
rect 19994 42310 19996 42362
rect 19940 42308 19996 42310
rect 20044 42362 20100 42364
rect 20044 42310 20046 42362
rect 20046 42310 20098 42362
rect 20098 42310 20100 42362
rect 20044 42308 20100 42310
rect 19836 40794 19892 40796
rect 19836 40742 19838 40794
rect 19838 40742 19890 40794
rect 19890 40742 19892 40794
rect 19836 40740 19892 40742
rect 19940 40794 19996 40796
rect 19940 40742 19942 40794
rect 19942 40742 19994 40794
rect 19994 40742 19996 40794
rect 19940 40740 19996 40742
rect 20044 40794 20100 40796
rect 20044 40742 20046 40794
rect 20046 40742 20098 40794
rect 20098 40742 20100 40794
rect 20044 40740 20100 40742
rect 19836 39226 19892 39228
rect 19836 39174 19838 39226
rect 19838 39174 19890 39226
rect 19890 39174 19892 39226
rect 19836 39172 19892 39174
rect 19940 39226 19996 39228
rect 19940 39174 19942 39226
rect 19942 39174 19994 39226
rect 19994 39174 19996 39226
rect 19940 39172 19996 39174
rect 20044 39226 20100 39228
rect 20044 39174 20046 39226
rect 20046 39174 20098 39226
rect 20098 39174 20100 39226
rect 20044 39172 20100 39174
rect 19836 37658 19892 37660
rect 19836 37606 19838 37658
rect 19838 37606 19890 37658
rect 19890 37606 19892 37658
rect 19836 37604 19892 37606
rect 19940 37658 19996 37660
rect 19940 37606 19942 37658
rect 19942 37606 19994 37658
rect 19994 37606 19996 37658
rect 19940 37604 19996 37606
rect 20044 37658 20100 37660
rect 20044 37606 20046 37658
rect 20046 37606 20098 37658
rect 20098 37606 20100 37658
rect 20044 37604 20100 37606
rect 19836 36090 19892 36092
rect 19836 36038 19838 36090
rect 19838 36038 19890 36090
rect 19890 36038 19892 36090
rect 19836 36036 19892 36038
rect 19940 36090 19996 36092
rect 19940 36038 19942 36090
rect 19942 36038 19994 36090
rect 19994 36038 19996 36090
rect 19940 36036 19996 36038
rect 20044 36090 20100 36092
rect 20044 36038 20046 36090
rect 20046 36038 20098 36090
rect 20098 36038 20100 36090
rect 20044 36036 20100 36038
rect 19836 34522 19892 34524
rect 19836 34470 19838 34522
rect 19838 34470 19890 34522
rect 19890 34470 19892 34522
rect 19836 34468 19892 34470
rect 19940 34522 19996 34524
rect 19940 34470 19942 34522
rect 19942 34470 19994 34522
rect 19994 34470 19996 34522
rect 19940 34468 19996 34470
rect 20044 34522 20100 34524
rect 20044 34470 20046 34522
rect 20046 34470 20098 34522
rect 20098 34470 20100 34522
rect 20044 34468 20100 34470
rect 19836 32954 19892 32956
rect 19836 32902 19838 32954
rect 19838 32902 19890 32954
rect 19890 32902 19892 32954
rect 19836 32900 19892 32902
rect 19940 32954 19996 32956
rect 19940 32902 19942 32954
rect 19942 32902 19994 32954
rect 19994 32902 19996 32954
rect 19940 32900 19996 32902
rect 20044 32954 20100 32956
rect 20044 32902 20046 32954
rect 20046 32902 20098 32954
rect 20098 32902 20100 32954
rect 20044 32900 20100 32902
rect 21980 75906 22036 75908
rect 21980 75854 21982 75906
rect 21982 75854 22034 75906
rect 22034 75854 22036 75906
rect 21980 75852 22036 75854
rect 23772 75628 23828 75684
rect 25228 75682 25284 75684
rect 25228 75630 25230 75682
rect 25230 75630 25282 75682
rect 25282 75630 25284 75682
rect 25228 75628 25284 75630
rect 25900 75628 25956 75684
rect 20860 73948 20916 74004
rect 19836 31386 19892 31388
rect 19836 31334 19838 31386
rect 19838 31334 19890 31386
rect 19890 31334 19892 31386
rect 19836 31332 19892 31334
rect 19940 31386 19996 31388
rect 19940 31334 19942 31386
rect 19942 31334 19994 31386
rect 19994 31334 19996 31386
rect 19940 31332 19996 31334
rect 20044 31386 20100 31388
rect 20044 31334 20046 31386
rect 20046 31334 20098 31386
rect 20098 31334 20100 31386
rect 20044 31332 20100 31334
rect 19836 29818 19892 29820
rect 19836 29766 19838 29818
rect 19838 29766 19890 29818
rect 19890 29766 19892 29818
rect 19836 29764 19892 29766
rect 19940 29818 19996 29820
rect 19940 29766 19942 29818
rect 19942 29766 19994 29818
rect 19994 29766 19996 29818
rect 19940 29764 19996 29766
rect 20044 29818 20100 29820
rect 20044 29766 20046 29818
rect 20046 29766 20098 29818
rect 20098 29766 20100 29818
rect 20044 29764 20100 29766
rect 19836 28250 19892 28252
rect 19836 28198 19838 28250
rect 19838 28198 19890 28250
rect 19890 28198 19892 28250
rect 19836 28196 19892 28198
rect 19940 28250 19996 28252
rect 19940 28198 19942 28250
rect 19942 28198 19994 28250
rect 19994 28198 19996 28250
rect 19940 28196 19996 28198
rect 20044 28250 20100 28252
rect 20044 28198 20046 28250
rect 20046 28198 20098 28250
rect 20098 28198 20100 28250
rect 20044 28196 20100 28198
rect 19836 26682 19892 26684
rect 19836 26630 19838 26682
rect 19838 26630 19890 26682
rect 19890 26630 19892 26682
rect 19836 26628 19892 26630
rect 19940 26682 19996 26684
rect 19940 26630 19942 26682
rect 19942 26630 19994 26682
rect 19994 26630 19996 26682
rect 19940 26628 19996 26630
rect 20044 26682 20100 26684
rect 20044 26630 20046 26682
rect 20046 26630 20098 26682
rect 20098 26630 20100 26682
rect 20044 26628 20100 26630
rect 19836 25114 19892 25116
rect 19836 25062 19838 25114
rect 19838 25062 19890 25114
rect 19890 25062 19892 25114
rect 19836 25060 19892 25062
rect 19940 25114 19996 25116
rect 19940 25062 19942 25114
rect 19942 25062 19994 25114
rect 19994 25062 19996 25114
rect 19940 25060 19996 25062
rect 20044 25114 20100 25116
rect 20044 25062 20046 25114
rect 20046 25062 20098 25114
rect 20098 25062 20100 25114
rect 20044 25060 20100 25062
rect 19740 24220 19796 24276
rect 20636 24722 20692 24724
rect 20636 24670 20638 24722
rect 20638 24670 20690 24722
rect 20690 24670 20692 24722
rect 20636 24668 20692 24670
rect 19516 23772 19572 23828
rect 19404 23548 19460 23604
rect 19836 23546 19892 23548
rect 19836 23494 19838 23546
rect 19838 23494 19890 23546
rect 19890 23494 19892 23546
rect 19836 23492 19892 23494
rect 19940 23546 19996 23548
rect 19940 23494 19942 23546
rect 19942 23494 19994 23546
rect 19994 23494 19996 23546
rect 19940 23492 19996 23494
rect 20044 23546 20100 23548
rect 20044 23494 20046 23546
rect 20046 23494 20098 23546
rect 20098 23494 20100 23546
rect 20044 23492 20100 23494
rect 19404 22482 19460 22484
rect 19404 22430 19406 22482
rect 19406 22430 19458 22482
rect 19458 22430 19460 22482
rect 19404 22428 19460 22430
rect 19628 22988 19684 23044
rect 19852 22316 19908 22372
rect 19852 22092 19908 22148
rect 19836 21978 19892 21980
rect 19836 21926 19838 21978
rect 19838 21926 19890 21978
rect 19890 21926 19892 21978
rect 19836 21924 19892 21926
rect 19940 21978 19996 21980
rect 19940 21926 19942 21978
rect 19942 21926 19994 21978
rect 19994 21926 19996 21978
rect 19940 21924 19996 21926
rect 20044 21978 20100 21980
rect 20044 21926 20046 21978
rect 20046 21926 20098 21978
rect 20098 21926 20100 21978
rect 20044 21924 20100 21926
rect 19068 20748 19124 20804
rect 18956 20076 19012 20132
rect 19068 20412 19124 20468
rect 20412 23826 20468 23828
rect 20412 23774 20414 23826
rect 20414 23774 20466 23826
rect 20466 23774 20468 23826
rect 20412 23772 20468 23774
rect 20524 23714 20580 23716
rect 20524 23662 20526 23714
rect 20526 23662 20578 23714
rect 20578 23662 20580 23714
rect 20524 23660 20580 23662
rect 20188 20748 20244 20804
rect 20748 23938 20804 23940
rect 20748 23886 20750 23938
rect 20750 23886 20802 23938
rect 20802 23886 20804 23938
rect 20748 23884 20804 23886
rect 19404 20412 19460 20468
rect 19836 20410 19892 20412
rect 19836 20358 19838 20410
rect 19838 20358 19890 20410
rect 19890 20358 19892 20410
rect 19836 20356 19892 20358
rect 19940 20410 19996 20412
rect 19940 20358 19942 20410
rect 19942 20358 19994 20410
rect 19994 20358 19996 20410
rect 19940 20356 19996 20358
rect 20044 20410 20100 20412
rect 20044 20358 20046 20410
rect 20046 20358 20098 20410
rect 20098 20358 20100 20410
rect 20044 20356 20100 20358
rect 19180 19852 19236 19908
rect 19628 19906 19684 19908
rect 19628 19854 19630 19906
rect 19630 19854 19682 19906
rect 19682 19854 19684 19906
rect 19628 19852 19684 19854
rect 19404 19516 19460 19572
rect 18620 18508 18676 18564
rect 18732 17554 18788 17556
rect 18732 17502 18734 17554
rect 18734 17502 18786 17554
rect 18786 17502 18788 17554
rect 18732 17500 18788 17502
rect 18620 13858 18676 13860
rect 18620 13806 18622 13858
rect 18622 13806 18674 13858
rect 18674 13806 18676 13858
rect 18620 13804 18676 13806
rect 17836 10892 17892 10948
rect 17724 10610 17780 10612
rect 17724 10558 17726 10610
rect 17726 10558 17778 10610
rect 17778 10558 17780 10610
rect 17724 10556 17780 10558
rect 17612 9266 17668 9268
rect 17612 9214 17614 9266
rect 17614 9214 17666 9266
rect 17666 9214 17668 9266
rect 17612 9212 17668 9214
rect 18284 10556 18340 10612
rect 18396 9212 18452 9268
rect 18508 9660 18564 9716
rect 18620 9324 18676 9380
rect 17836 8370 17892 8372
rect 17836 8318 17838 8370
rect 17838 8318 17890 8370
rect 17890 8318 17892 8370
rect 17836 8316 17892 8318
rect 19180 18620 19236 18676
rect 19292 18338 19348 18340
rect 19292 18286 19294 18338
rect 19294 18286 19346 18338
rect 19346 18286 19348 18338
rect 19292 18284 19348 18286
rect 19516 19010 19572 19012
rect 19516 18958 19518 19010
rect 19518 18958 19570 19010
rect 19570 18958 19572 19010
rect 19516 18956 19572 18958
rect 20412 22482 20468 22484
rect 20412 22430 20414 22482
rect 20414 22430 20466 22482
rect 20466 22430 20468 22482
rect 20412 22428 20468 22430
rect 20748 21308 20804 21364
rect 20300 19852 20356 19908
rect 20412 19234 20468 19236
rect 20412 19182 20414 19234
rect 20414 19182 20466 19234
rect 20466 19182 20468 19234
rect 20412 19180 20468 19182
rect 19836 18842 19892 18844
rect 19836 18790 19838 18842
rect 19838 18790 19890 18842
rect 19890 18790 19892 18842
rect 19836 18788 19892 18790
rect 19940 18842 19996 18844
rect 19940 18790 19942 18842
rect 19942 18790 19994 18842
rect 19994 18790 19996 18842
rect 19940 18788 19996 18790
rect 20044 18842 20100 18844
rect 20044 18790 20046 18842
rect 20046 18790 20098 18842
rect 20098 18790 20100 18842
rect 20044 18788 20100 18790
rect 20188 18620 20244 18676
rect 20524 18844 20580 18900
rect 19628 18508 19684 18564
rect 19404 17666 19460 17668
rect 19404 17614 19406 17666
rect 19406 17614 19458 17666
rect 19458 17614 19460 17666
rect 19404 17612 19460 17614
rect 19292 17500 19348 17556
rect 18956 14252 19012 14308
rect 19180 13804 19236 13860
rect 19068 13634 19124 13636
rect 19068 13582 19070 13634
rect 19070 13582 19122 13634
rect 19122 13582 19124 13634
rect 19068 13580 19124 13582
rect 19516 13746 19572 13748
rect 19516 13694 19518 13746
rect 19518 13694 19570 13746
rect 19570 13694 19572 13746
rect 19516 13692 19572 13694
rect 20188 17666 20244 17668
rect 20188 17614 20190 17666
rect 20190 17614 20242 17666
rect 20242 17614 20244 17666
rect 20188 17612 20244 17614
rect 20636 18620 20692 18676
rect 20748 19180 20804 19236
rect 20636 18284 20692 18340
rect 21196 23938 21252 23940
rect 21196 23886 21198 23938
rect 21198 23886 21250 23938
rect 21250 23886 21252 23938
rect 21196 23884 21252 23886
rect 21644 23714 21700 23716
rect 21644 23662 21646 23714
rect 21646 23662 21698 23714
rect 21698 23662 21700 23714
rect 21644 23660 21700 23662
rect 21196 22370 21252 22372
rect 21196 22318 21198 22370
rect 21198 22318 21250 22370
rect 21250 22318 21252 22370
rect 21196 22316 21252 22318
rect 21644 21980 21700 22036
rect 22316 23714 22372 23716
rect 22316 23662 22318 23714
rect 22318 23662 22370 23714
rect 22370 23662 22372 23714
rect 22316 23660 22372 23662
rect 21868 21644 21924 21700
rect 22092 21868 22148 21924
rect 22316 21698 22372 21700
rect 22316 21646 22318 21698
rect 22318 21646 22370 21698
rect 22370 21646 22372 21698
rect 22316 21644 22372 21646
rect 21420 19068 21476 19124
rect 21532 18844 21588 18900
rect 21756 19404 21812 19460
rect 21644 18620 21700 18676
rect 23660 25282 23716 25284
rect 23660 25230 23662 25282
rect 23662 25230 23714 25282
rect 23714 25230 23716 25282
rect 23660 25228 23716 25230
rect 23324 24444 23380 24500
rect 24108 25282 24164 25284
rect 24108 25230 24110 25282
rect 24110 25230 24162 25282
rect 24162 25230 24164 25282
rect 24108 25228 24164 25230
rect 24332 25004 24388 25060
rect 23996 23938 24052 23940
rect 23996 23886 23998 23938
rect 23998 23886 24050 23938
rect 24050 23886 24052 23938
rect 23996 23884 24052 23886
rect 24220 23660 24276 23716
rect 24108 23212 24164 23268
rect 23996 23100 24052 23156
rect 24220 23100 24276 23156
rect 23548 22092 23604 22148
rect 22988 21980 23044 22036
rect 23548 21474 23604 21476
rect 23548 21422 23550 21474
rect 23550 21422 23602 21474
rect 23602 21422 23604 21474
rect 23548 21420 23604 21422
rect 24332 21868 24388 21924
rect 30156 75628 30212 75684
rect 26908 40348 26964 40404
rect 26908 38892 26964 38948
rect 26908 37324 26964 37380
rect 26908 36316 26964 36372
rect 28476 33068 28532 33124
rect 33628 75740 33684 75796
rect 33516 75682 33572 75684
rect 33516 75630 33518 75682
rect 33518 75630 33570 75682
rect 33570 75630 33572 75682
rect 33516 75628 33572 75630
rect 28476 31612 28532 31668
rect 31052 74732 31108 74788
rect 26908 31052 26964 31108
rect 26908 30044 26964 30100
rect 25228 25004 25284 25060
rect 25564 24722 25620 24724
rect 25564 24670 25566 24722
rect 25566 24670 25618 24722
rect 25618 24670 25620 24722
rect 25564 24668 25620 24670
rect 25004 24556 25060 24612
rect 25676 24610 25732 24612
rect 25676 24558 25678 24610
rect 25678 24558 25730 24610
rect 25730 24558 25732 24610
rect 25676 24556 25732 24558
rect 26012 23212 26068 23268
rect 25116 23154 25172 23156
rect 25116 23102 25118 23154
rect 25118 23102 25170 23154
rect 25170 23102 25172 23154
rect 25116 23100 25172 23102
rect 25564 23154 25620 23156
rect 25564 23102 25566 23154
rect 25566 23102 25618 23154
rect 25618 23102 25620 23154
rect 25564 23100 25620 23102
rect 24556 23042 24612 23044
rect 24556 22990 24558 23042
rect 24558 22990 24610 23042
rect 24610 22990 24612 23042
rect 24556 22988 24612 22990
rect 24444 21644 24500 21700
rect 25676 21698 25732 21700
rect 25676 21646 25678 21698
rect 25678 21646 25730 21698
rect 25730 21646 25732 21698
rect 25676 21644 25732 21646
rect 23996 21420 24052 21476
rect 23660 20748 23716 20804
rect 24780 20748 24836 20804
rect 22652 20076 22708 20132
rect 22540 19292 22596 19348
rect 21980 19180 22036 19236
rect 23212 20076 23268 20132
rect 22988 19404 23044 19460
rect 22652 19234 22708 19236
rect 22652 19182 22654 19234
rect 22654 19182 22706 19234
rect 22706 19182 22708 19234
rect 22652 19180 22708 19182
rect 20860 17500 20916 17556
rect 21980 18172 22036 18228
rect 22316 18172 22372 18228
rect 21868 17500 21924 17556
rect 23100 19010 23156 19012
rect 23100 18958 23102 19010
rect 23102 18958 23154 19010
rect 23154 18958 23156 19010
rect 23100 18956 23156 18958
rect 19836 17274 19892 17276
rect 19836 17222 19838 17274
rect 19838 17222 19890 17274
rect 19890 17222 19892 17274
rect 19836 17220 19892 17222
rect 19940 17274 19996 17276
rect 19940 17222 19942 17274
rect 19942 17222 19994 17274
rect 19994 17222 19996 17274
rect 19940 17220 19996 17222
rect 20044 17274 20100 17276
rect 20044 17222 20046 17274
rect 20046 17222 20098 17274
rect 20098 17222 20100 17274
rect 20044 17220 20100 17222
rect 19836 15706 19892 15708
rect 19836 15654 19838 15706
rect 19838 15654 19890 15706
rect 19890 15654 19892 15706
rect 19836 15652 19892 15654
rect 19940 15706 19996 15708
rect 19940 15654 19942 15706
rect 19942 15654 19994 15706
rect 19994 15654 19996 15706
rect 19940 15652 19996 15654
rect 20044 15706 20100 15708
rect 20044 15654 20046 15706
rect 20046 15654 20098 15706
rect 20098 15654 20100 15706
rect 20044 15652 20100 15654
rect 24668 19852 24724 19908
rect 24444 19516 24500 19572
rect 23548 19122 23604 19124
rect 23548 19070 23550 19122
rect 23550 19070 23602 19122
rect 23602 19070 23604 19122
rect 23548 19068 23604 19070
rect 24892 20524 24948 20580
rect 24444 18956 24500 19012
rect 23884 18844 23940 18900
rect 24668 18338 24724 18340
rect 24668 18286 24670 18338
rect 24670 18286 24722 18338
rect 24722 18286 24724 18338
rect 24668 18284 24724 18286
rect 21868 14812 21924 14868
rect 19740 14252 19796 14308
rect 20076 14306 20132 14308
rect 20076 14254 20078 14306
rect 20078 14254 20130 14306
rect 20130 14254 20132 14306
rect 20076 14252 20132 14254
rect 19836 14138 19892 14140
rect 19836 14086 19838 14138
rect 19838 14086 19890 14138
rect 19890 14086 19892 14138
rect 19836 14084 19892 14086
rect 19940 14138 19996 14140
rect 19940 14086 19942 14138
rect 19942 14086 19994 14138
rect 19994 14086 19996 14138
rect 19940 14084 19996 14086
rect 20044 14138 20100 14140
rect 20044 14086 20046 14138
rect 20046 14086 20098 14138
rect 20098 14086 20100 14138
rect 20044 14084 20100 14086
rect 21420 14306 21476 14308
rect 21420 14254 21422 14306
rect 21422 14254 21474 14306
rect 21474 14254 21476 14306
rect 21420 14252 21476 14254
rect 20300 13692 20356 13748
rect 19836 12570 19892 12572
rect 19836 12518 19838 12570
rect 19838 12518 19890 12570
rect 19890 12518 19892 12570
rect 19836 12516 19892 12518
rect 19940 12570 19996 12572
rect 19940 12518 19942 12570
rect 19942 12518 19994 12570
rect 19994 12518 19996 12570
rect 19940 12516 19996 12518
rect 20044 12570 20100 12572
rect 20044 12518 20046 12570
rect 20046 12518 20098 12570
rect 20098 12518 20100 12570
rect 20044 12516 20100 12518
rect 19964 11452 20020 11508
rect 18956 11116 19012 11172
rect 18732 8988 18788 9044
rect 18844 9266 18900 9268
rect 18844 9214 18846 9266
rect 18846 9214 18898 9266
rect 18898 9214 18900 9266
rect 18844 9212 18900 9214
rect 18732 8764 18788 8820
rect 18620 8316 18676 8372
rect 18508 8034 18564 8036
rect 18508 7982 18510 8034
rect 18510 7982 18562 8034
rect 18562 7982 18564 8034
rect 18508 7980 18564 7982
rect 17948 7868 18004 7924
rect 17836 7756 17892 7812
rect 17612 7532 17668 7588
rect 17276 5852 17332 5908
rect 17388 5964 17444 6020
rect 17388 5180 17444 5236
rect 17276 4172 17332 4228
rect 17500 5068 17556 5124
rect 17836 5516 17892 5572
rect 18396 7756 18452 7812
rect 18172 6636 18228 6692
rect 18396 7196 18452 7252
rect 18396 5292 18452 5348
rect 18844 7644 18900 7700
rect 19740 11170 19796 11172
rect 19740 11118 19742 11170
rect 19742 11118 19794 11170
rect 19794 11118 19796 11170
rect 19740 11116 19796 11118
rect 19404 9042 19460 9044
rect 19404 8990 19406 9042
rect 19406 8990 19458 9042
rect 19458 8990 19460 9042
rect 19404 8988 19460 8990
rect 19180 8428 19236 8484
rect 19516 8876 19572 8932
rect 19404 8204 19460 8260
rect 18956 7756 19012 7812
rect 17948 4956 18004 5012
rect 17836 4284 17892 4340
rect 17500 3612 17556 3668
rect 17948 4114 18004 4116
rect 17948 4062 17950 4114
rect 17950 4062 18002 4114
rect 18002 4062 18004 4114
rect 17948 4060 18004 4062
rect 17724 3388 17780 3444
rect 17948 3388 18004 3444
rect 18732 6748 18788 6804
rect 19836 11002 19892 11004
rect 19836 10950 19838 11002
rect 19838 10950 19890 11002
rect 19890 10950 19892 11002
rect 19836 10948 19892 10950
rect 19940 11002 19996 11004
rect 19940 10950 19942 11002
rect 19942 10950 19994 11002
rect 19994 10950 19996 11002
rect 19940 10948 19996 10950
rect 20044 11002 20100 11004
rect 20044 10950 20046 11002
rect 20046 10950 20098 11002
rect 20098 10950 20100 11002
rect 20044 10948 20100 10950
rect 19836 9434 19892 9436
rect 19836 9382 19838 9434
rect 19838 9382 19890 9434
rect 19890 9382 19892 9434
rect 19836 9380 19892 9382
rect 19940 9434 19996 9436
rect 19940 9382 19942 9434
rect 19942 9382 19994 9434
rect 19994 9382 19996 9434
rect 19940 9380 19996 9382
rect 20044 9434 20100 9436
rect 20044 9382 20046 9434
rect 20046 9382 20098 9434
rect 20098 9382 20100 9434
rect 20044 9380 20100 9382
rect 20076 8930 20132 8932
rect 20076 8878 20078 8930
rect 20078 8878 20130 8930
rect 20130 8878 20132 8930
rect 20076 8876 20132 8878
rect 25340 20802 25396 20804
rect 25340 20750 25342 20802
rect 25342 20750 25394 20802
rect 25394 20750 25396 20802
rect 25340 20748 25396 20750
rect 26012 20802 26068 20804
rect 26012 20750 26014 20802
rect 26014 20750 26066 20802
rect 26066 20750 26068 20802
rect 26012 20748 26068 20750
rect 25564 20524 25620 20580
rect 26124 20578 26180 20580
rect 26124 20526 26126 20578
rect 26126 20526 26178 20578
rect 26178 20526 26180 20578
rect 26124 20524 26180 20526
rect 25900 20412 25956 20468
rect 25564 19404 25620 19460
rect 25452 19292 25508 19348
rect 25116 19122 25172 19124
rect 25116 19070 25118 19122
rect 25118 19070 25170 19122
rect 25170 19070 25172 19122
rect 25116 19068 25172 19070
rect 25788 19122 25844 19124
rect 25788 19070 25790 19122
rect 25790 19070 25842 19122
rect 25842 19070 25844 19122
rect 25788 19068 25844 19070
rect 25340 18338 25396 18340
rect 25340 18286 25342 18338
rect 25342 18286 25394 18338
rect 25394 18286 25396 18338
rect 25340 18284 25396 18286
rect 25676 18172 25732 18228
rect 24892 14812 24948 14868
rect 25116 17554 25172 17556
rect 25116 17502 25118 17554
rect 25118 17502 25170 17554
rect 25170 17502 25172 17554
rect 25116 17500 25172 17502
rect 22876 14252 22932 14308
rect 25564 16380 25620 16436
rect 25676 15820 25732 15876
rect 23548 13804 23604 13860
rect 22540 13692 22596 13748
rect 20748 11506 20804 11508
rect 20748 11454 20750 11506
rect 20750 11454 20802 11506
rect 20802 11454 20804 11506
rect 20748 11452 20804 11454
rect 21756 11452 21812 11508
rect 20300 9826 20356 9828
rect 20300 9774 20302 9826
rect 20302 9774 20354 9826
rect 20354 9774 20356 9826
rect 20300 9772 20356 9774
rect 20188 8764 20244 8820
rect 20412 8652 20468 8708
rect 19628 8316 19684 8372
rect 19964 8370 20020 8372
rect 19964 8318 19966 8370
rect 19966 8318 20018 8370
rect 20018 8318 20020 8370
rect 19964 8316 20020 8318
rect 20076 8258 20132 8260
rect 20076 8206 20078 8258
rect 20078 8206 20130 8258
rect 20130 8206 20132 8258
rect 20076 8204 20132 8206
rect 20188 8092 20244 8148
rect 19628 8034 19684 8036
rect 19628 7982 19630 8034
rect 19630 7982 19682 8034
rect 19682 7982 19684 8034
rect 19628 7980 19684 7982
rect 19836 7866 19892 7868
rect 19836 7814 19838 7866
rect 19838 7814 19890 7866
rect 19890 7814 19892 7866
rect 19836 7812 19892 7814
rect 19940 7866 19996 7868
rect 19940 7814 19942 7866
rect 19942 7814 19994 7866
rect 19994 7814 19996 7866
rect 19940 7812 19996 7814
rect 20044 7866 20100 7868
rect 20044 7814 20046 7866
rect 20046 7814 20098 7866
rect 20098 7814 20100 7866
rect 20044 7812 20100 7814
rect 19740 7586 19796 7588
rect 19740 7534 19742 7586
rect 19742 7534 19794 7586
rect 19794 7534 19796 7586
rect 19740 7532 19796 7534
rect 19852 7420 19908 7476
rect 20300 7698 20356 7700
rect 20300 7646 20302 7698
rect 20302 7646 20354 7698
rect 20354 7646 20356 7698
rect 20300 7644 20356 7646
rect 20188 7532 20244 7588
rect 20076 7420 20132 7476
rect 19628 6636 19684 6692
rect 19516 6412 19572 6468
rect 19068 6188 19124 6244
rect 18956 5852 19012 5908
rect 18172 5010 18228 5012
rect 18172 4958 18174 5010
rect 18174 4958 18226 5010
rect 18226 4958 18228 5010
rect 18172 4956 18228 4958
rect 18284 4956 18340 5012
rect 18284 4732 18340 4788
rect 20076 6412 20132 6468
rect 19836 6298 19892 6300
rect 19836 6246 19838 6298
rect 19838 6246 19890 6298
rect 19890 6246 19892 6298
rect 19836 6244 19892 6246
rect 19940 6298 19996 6300
rect 19940 6246 19942 6298
rect 19942 6246 19994 6298
rect 19994 6246 19996 6298
rect 19940 6244 19996 6246
rect 20044 6298 20100 6300
rect 20044 6246 20046 6298
rect 20046 6246 20098 6298
rect 20098 6246 20100 6298
rect 20044 6244 20100 6246
rect 19068 4732 19124 4788
rect 19068 4508 19124 4564
rect 18284 3612 18340 3668
rect 18620 4060 18676 4116
rect 19516 5740 19572 5796
rect 19404 5628 19460 5684
rect 23436 12012 23492 12068
rect 20860 9826 20916 9828
rect 20860 9774 20862 9826
rect 20862 9774 20914 9826
rect 20914 9774 20916 9826
rect 20860 9772 20916 9774
rect 21420 8876 21476 8932
rect 22652 11282 22708 11284
rect 22652 11230 22654 11282
rect 22654 11230 22706 11282
rect 22706 11230 22708 11282
rect 22652 11228 22708 11230
rect 22092 8988 22148 9044
rect 20972 7868 21028 7924
rect 20636 7756 20692 7812
rect 20748 7532 20804 7588
rect 20636 6524 20692 6580
rect 19964 5404 20020 5460
rect 19836 4730 19892 4732
rect 19836 4678 19838 4730
rect 19838 4678 19890 4730
rect 19890 4678 19892 4730
rect 19836 4676 19892 4678
rect 19940 4730 19996 4732
rect 19940 4678 19942 4730
rect 19942 4678 19994 4730
rect 19994 4678 19996 4730
rect 19940 4676 19996 4678
rect 20044 4730 20100 4732
rect 20044 4678 20046 4730
rect 20046 4678 20098 4730
rect 20098 4678 20100 4730
rect 20044 4676 20100 4678
rect 19404 4172 19460 4228
rect 19292 4060 19348 4116
rect 18396 3500 18452 3556
rect 19068 3612 19124 3668
rect 18844 1260 18900 1316
rect 19292 3612 19348 3668
rect 19628 4172 19684 4228
rect 19628 3612 19684 3668
rect 19516 3500 19572 3556
rect 20412 5010 20468 5012
rect 20412 4958 20414 5010
rect 20414 4958 20466 5010
rect 20466 4958 20468 5010
rect 20412 4956 20468 4958
rect 20412 4508 20468 4564
rect 21196 7532 21252 7588
rect 21196 5906 21252 5908
rect 21196 5854 21198 5906
rect 21198 5854 21250 5906
rect 21250 5854 21252 5906
rect 21196 5852 21252 5854
rect 21644 7756 21700 7812
rect 21532 6188 21588 6244
rect 21532 5906 21588 5908
rect 21532 5854 21534 5906
rect 21534 5854 21586 5906
rect 21586 5854 21588 5906
rect 21532 5852 21588 5854
rect 21532 5516 21588 5572
rect 22316 9266 22372 9268
rect 22316 9214 22318 9266
rect 22318 9214 22370 9266
rect 22370 9214 22372 9266
rect 22316 9212 22372 9214
rect 22316 8204 22372 8260
rect 21980 6300 22036 6356
rect 22428 7084 22484 7140
rect 22540 6748 22596 6804
rect 22764 9826 22820 9828
rect 22764 9774 22766 9826
rect 22766 9774 22818 9826
rect 22818 9774 22820 9826
rect 22764 9772 22820 9774
rect 22988 10498 23044 10500
rect 22988 10446 22990 10498
rect 22990 10446 23042 10498
rect 23042 10446 23044 10498
rect 22988 10444 23044 10446
rect 23436 9548 23492 9604
rect 23212 8988 23268 9044
rect 22876 7084 22932 7140
rect 21868 5628 21924 5684
rect 22764 6018 22820 6020
rect 22764 5966 22766 6018
rect 22766 5966 22818 6018
rect 22818 5966 22820 6018
rect 22764 5964 22820 5966
rect 22204 5852 22260 5908
rect 22428 5292 22484 5348
rect 21644 5180 21700 5236
rect 20300 4396 20356 4452
rect 20300 3724 20356 3780
rect 20076 3276 20132 3332
rect 19836 3162 19892 3164
rect 19836 3110 19838 3162
rect 19838 3110 19890 3162
rect 19890 3110 19892 3162
rect 19836 3108 19892 3110
rect 19940 3162 19996 3164
rect 19940 3110 19942 3162
rect 19942 3110 19994 3162
rect 19994 3110 19996 3162
rect 19940 3108 19996 3110
rect 20044 3162 20100 3164
rect 20044 3110 20046 3162
rect 20046 3110 20098 3162
rect 20098 3110 20100 3162
rect 20044 3108 20100 3110
rect 19628 1708 19684 1764
rect 20636 3724 20692 3780
rect 20860 3836 20916 3892
rect 20972 3724 21028 3780
rect 21084 3388 21140 3444
rect 21308 4450 21364 4452
rect 21308 4398 21310 4450
rect 21310 4398 21362 4450
rect 21362 4398 21364 4450
rect 21308 4396 21364 4398
rect 21196 3052 21252 3108
rect 21532 4172 21588 4228
rect 22092 4956 22148 5012
rect 21868 4898 21924 4900
rect 21868 4846 21870 4898
rect 21870 4846 21922 4898
rect 21922 4846 21924 4898
rect 21868 4844 21924 4846
rect 22540 5010 22596 5012
rect 22540 4958 22542 5010
rect 22542 4958 22594 5010
rect 22594 4958 22596 5010
rect 22540 4956 22596 4958
rect 21980 4450 22036 4452
rect 21980 4398 21982 4450
rect 21982 4398 22034 4450
rect 22034 4398 22036 4450
rect 21980 4396 22036 4398
rect 22652 4732 22708 4788
rect 21756 3948 21812 4004
rect 21756 3612 21812 3668
rect 22428 4508 22484 4564
rect 22876 4620 22932 4676
rect 22316 4172 22372 4228
rect 22428 4060 22484 4116
rect 21532 2492 21588 2548
rect 21308 1484 21364 1540
rect 22652 1372 22708 1428
rect 24892 13692 24948 13748
rect 24668 13580 24724 13636
rect 25452 13468 25508 13524
rect 26348 20690 26404 20692
rect 26348 20638 26350 20690
rect 26350 20638 26402 20690
rect 26402 20638 26404 20690
rect 26348 20636 26404 20638
rect 26348 20130 26404 20132
rect 26348 20078 26350 20130
rect 26350 20078 26402 20130
rect 26402 20078 26404 20130
rect 26348 20076 26404 20078
rect 27020 24668 27076 24724
rect 27468 23938 27524 23940
rect 27468 23886 27470 23938
rect 27470 23886 27522 23938
rect 27522 23886 27524 23938
rect 27468 23884 27524 23886
rect 27580 23378 27636 23380
rect 27580 23326 27582 23378
rect 27582 23326 27634 23378
rect 27634 23326 27636 23378
rect 27580 23324 27636 23326
rect 26908 23154 26964 23156
rect 26908 23102 26910 23154
rect 26910 23102 26962 23154
rect 26962 23102 26964 23154
rect 26908 23100 26964 23102
rect 27132 22876 27188 22932
rect 28476 24668 28532 24724
rect 27916 23826 27972 23828
rect 27916 23774 27918 23826
rect 27918 23774 27970 23826
rect 27970 23774 27972 23826
rect 27916 23772 27972 23774
rect 28140 23324 28196 23380
rect 28476 23324 28532 23380
rect 30492 24722 30548 24724
rect 30492 24670 30494 24722
rect 30494 24670 30546 24722
rect 30546 24670 30548 24722
rect 30492 24668 30548 24670
rect 30492 23772 30548 23828
rect 29932 23212 29988 23268
rect 27468 23042 27524 23044
rect 27468 22990 27470 23042
rect 27470 22990 27522 23042
rect 27522 22990 27524 23042
rect 27468 22988 27524 22990
rect 27692 22316 27748 22372
rect 27132 22092 27188 22148
rect 27692 22146 27748 22148
rect 27692 22094 27694 22146
rect 27694 22094 27746 22146
rect 27746 22094 27748 22146
rect 27692 22092 27748 22094
rect 27244 20802 27300 20804
rect 27244 20750 27246 20802
rect 27246 20750 27298 20802
rect 27298 20750 27300 20802
rect 27244 20748 27300 20750
rect 26684 20524 26740 20580
rect 26908 20130 26964 20132
rect 26908 20078 26910 20130
rect 26910 20078 26962 20130
rect 26962 20078 26964 20130
rect 26908 20076 26964 20078
rect 26460 19292 26516 19348
rect 26460 19010 26516 19012
rect 26460 18958 26462 19010
rect 26462 18958 26514 19010
rect 26514 18958 26516 19010
rect 26460 18956 26516 18958
rect 26460 18450 26516 18452
rect 26460 18398 26462 18450
rect 26462 18398 26514 18450
rect 26514 18398 26516 18450
rect 26460 18396 26516 18398
rect 27356 20578 27412 20580
rect 27356 20526 27358 20578
rect 27358 20526 27410 20578
rect 27410 20526 27412 20578
rect 27356 20524 27412 20526
rect 27580 20076 27636 20132
rect 27132 19964 27188 20020
rect 27692 19964 27748 20020
rect 27468 19906 27524 19908
rect 27468 19854 27470 19906
rect 27470 19854 27522 19906
rect 27522 19854 27524 19906
rect 27468 19852 27524 19854
rect 27468 19180 27524 19236
rect 28700 23042 28756 23044
rect 28700 22990 28702 23042
rect 28702 22990 28754 23042
rect 28754 22990 28756 23042
rect 28700 22988 28756 22990
rect 30156 22540 30212 22596
rect 28252 22092 28308 22148
rect 27916 20578 27972 20580
rect 27916 20526 27918 20578
rect 27918 20526 27970 20578
rect 27970 20526 27972 20578
rect 27916 20524 27972 20526
rect 30940 22370 30996 22372
rect 30940 22318 30942 22370
rect 30942 22318 30994 22370
rect 30994 22318 30996 22370
rect 30940 22316 30996 22318
rect 29036 20636 29092 20692
rect 28476 20524 28532 20580
rect 29596 20578 29652 20580
rect 29596 20526 29598 20578
rect 29598 20526 29650 20578
rect 29650 20526 29652 20578
rect 29596 20524 29652 20526
rect 29708 19964 29764 20020
rect 28252 19516 28308 19572
rect 27804 19068 27860 19124
rect 27468 19010 27524 19012
rect 27468 18958 27470 19010
rect 27470 18958 27522 19010
rect 27522 18958 27524 19010
rect 27468 18956 27524 18958
rect 28476 19180 28532 19236
rect 28140 19010 28196 19012
rect 28140 18958 28142 19010
rect 28142 18958 28194 19010
rect 28194 18958 28196 19010
rect 28140 18956 28196 18958
rect 28700 19068 28756 19124
rect 27804 18620 27860 18676
rect 26572 18060 26628 18116
rect 27132 18284 27188 18340
rect 26572 16380 26628 16436
rect 28476 17836 28532 17892
rect 28140 17724 28196 17780
rect 27804 16380 27860 16436
rect 27132 15932 27188 15988
rect 26012 15484 26068 15540
rect 26796 15708 26852 15764
rect 27356 15820 27412 15876
rect 27692 15596 27748 15652
rect 27468 15484 27524 15540
rect 27804 15260 27860 15316
rect 28140 16828 28196 16884
rect 28252 16492 28308 16548
rect 28028 15596 28084 15652
rect 25900 13804 25956 13860
rect 25788 12796 25844 12852
rect 27020 13858 27076 13860
rect 27020 13806 27022 13858
rect 27022 13806 27074 13858
rect 27074 13806 27076 13858
rect 27020 13804 27076 13806
rect 27132 13692 27188 13748
rect 27692 13580 27748 13636
rect 24892 11282 24948 11284
rect 24892 11230 24894 11282
rect 24894 11230 24946 11282
rect 24946 11230 24948 11282
rect 24892 11228 24948 11230
rect 25340 12066 25396 12068
rect 25340 12014 25342 12066
rect 25342 12014 25394 12066
rect 25394 12014 25396 12066
rect 25340 12012 25396 12014
rect 25228 10892 25284 10948
rect 25340 10498 25396 10500
rect 25340 10446 25342 10498
rect 25342 10446 25394 10498
rect 25394 10446 25396 10498
rect 25340 10444 25396 10446
rect 24668 9884 24724 9940
rect 23548 9212 23604 9268
rect 24668 9266 24724 9268
rect 24668 9214 24670 9266
rect 24670 9214 24722 9266
rect 24722 9214 24724 9266
rect 24668 9212 24724 9214
rect 23660 8988 23716 9044
rect 23436 6972 23492 7028
rect 24108 6860 24164 6916
rect 23324 6578 23380 6580
rect 23324 6526 23326 6578
rect 23326 6526 23378 6578
rect 23378 6526 23380 6578
rect 23324 6524 23380 6526
rect 23660 6524 23716 6580
rect 23548 6300 23604 6356
rect 23436 5628 23492 5684
rect 23324 5068 23380 5124
rect 22988 4508 23044 4564
rect 23212 4844 23268 4900
rect 22988 4338 23044 4340
rect 22988 4286 22990 4338
rect 22990 4286 23042 4338
rect 23042 4286 23044 4338
rect 22988 4284 23044 4286
rect 23212 4226 23268 4228
rect 23212 4174 23214 4226
rect 23214 4174 23266 4226
rect 23266 4174 23268 4226
rect 23212 4172 23268 4174
rect 23548 4956 23604 5012
rect 23660 5404 23716 5460
rect 22988 3554 23044 3556
rect 22988 3502 22990 3554
rect 22990 3502 23042 3554
rect 23042 3502 23044 3554
rect 22988 3500 23044 3502
rect 23548 3388 23604 3444
rect 23884 5180 23940 5236
rect 24220 5740 24276 5796
rect 23996 3836 24052 3892
rect 23660 3276 23716 3332
rect 23884 2268 23940 2324
rect 25228 9266 25284 9268
rect 25228 9214 25230 9266
rect 25230 9214 25282 9266
rect 25282 9214 25284 9266
rect 25228 9212 25284 9214
rect 25788 10220 25844 10276
rect 25340 8988 25396 9044
rect 24668 8092 24724 8148
rect 24780 6972 24836 7028
rect 24668 6466 24724 6468
rect 24668 6414 24670 6466
rect 24670 6414 24722 6466
rect 24722 6414 24724 6466
rect 24668 6412 24724 6414
rect 24332 4060 24388 4116
rect 24444 4508 24500 4564
rect 24220 3276 24276 3332
rect 24220 2716 24276 2772
rect 24108 2156 24164 2212
rect 23772 1708 23828 1764
rect 24668 4450 24724 4452
rect 24668 4398 24670 4450
rect 24670 4398 24722 4450
rect 24722 4398 24724 4450
rect 24668 4396 24724 4398
rect 24556 3724 24612 3780
rect 24556 3500 24612 3556
rect 24780 3724 24836 3780
rect 25564 8258 25620 8260
rect 25564 8206 25566 8258
rect 25566 8206 25618 8258
rect 25618 8206 25620 8258
rect 25564 8204 25620 8206
rect 26236 11564 26292 11620
rect 27132 11116 27188 11172
rect 26684 10892 26740 10948
rect 25900 9042 25956 9044
rect 25900 8990 25902 9042
rect 25902 8990 25954 9042
rect 25954 8990 25956 9042
rect 25900 8988 25956 8990
rect 26236 10332 26292 10388
rect 25788 8092 25844 8148
rect 25900 8428 25956 8484
rect 25340 7756 25396 7812
rect 25564 7308 25620 7364
rect 25452 7196 25508 7252
rect 25340 6412 25396 6468
rect 25788 7420 25844 7476
rect 25788 6972 25844 7028
rect 25676 6748 25732 6804
rect 25788 6076 25844 6132
rect 25452 5794 25508 5796
rect 25452 5742 25454 5794
rect 25454 5742 25506 5794
rect 25506 5742 25508 5794
rect 25452 5740 25508 5742
rect 25452 5404 25508 5460
rect 26012 8204 26068 8260
rect 26796 8988 26852 9044
rect 26348 8876 26404 8932
rect 26684 8930 26740 8932
rect 26684 8878 26686 8930
rect 26686 8878 26738 8930
rect 26738 8878 26740 8930
rect 26684 8876 26740 8878
rect 26572 8764 26628 8820
rect 26236 8092 26292 8148
rect 26908 8370 26964 8372
rect 26908 8318 26910 8370
rect 26910 8318 26962 8370
rect 26962 8318 26964 8370
rect 26908 8316 26964 8318
rect 27020 8204 27076 8260
rect 26572 8146 26628 8148
rect 26572 8094 26574 8146
rect 26574 8094 26626 8146
rect 26626 8094 26628 8146
rect 26572 8092 26628 8094
rect 26460 7756 26516 7812
rect 26348 7698 26404 7700
rect 26348 7646 26350 7698
rect 26350 7646 26402 7698
rect 26402 7646 26404 7698
rect 26348 7644 26404 7646
rect 26012 6748 26068 6804
rect 26124 6860 26180 6916
rect 26012 5682 26068 5684
rect 26012 5630 26014 5682
rect 26014 5630 26066 5682
rect 26066 5630 26068 5682
rect 26012 5628 26068 5630
rect 26012 5180 26068 5236
rect 26348 6748 26404 6804
rect 26572 5906 26628 5908
rect 26572 5854 26574 5906
rect 26574 5854 26626 5906
rect 26626 5854 26628 5906
rect 26572 5852 26628 5854
rect 26348 5404 26404 5460
rect 26012 4226 26068 4228
rect 26012 4174 26014 4226
rect 26014 4174 26066 4226
rect 26066 4174 26068 4226
rect 26012 4172 26068 4174
rect 26236 3724 26292 3780
rect 25788 3612 25844 3668
rect 25004 3276 25060 3332
rect 25116 3500 25172 3556
rect 25340 2044 25396 2100
rect 26684 5404 26740 5460
rect 28140 15484 28196 15540
rect 28588 17778 28644 17780
rect 28588 17726 28590 17778
rect 28590 17726 28642 17778
rect 28642 17726 28644 17778
rect 28588 17724 28644 17726
rect 30268 19122 30324 19124
rect 30268 19070 30270 19122
rect 30270 19070 30322 19122
rect 30322 19070 30324 19122
rect 30268 19068 30324 19070
rect 30940 20076 30996 20132
rect 30828 19068 30884 19124
rect 29484 18956 29540 19012
rect 29484 18732 29540 18788
rect 29260 17276 29316 17332
rect 28476 16044 28532 16100
rect 28588 15932 28644 15988
rect 28476 15260 28532 15316
rect 30716 18060 30772 18116
rect 30380 17500 30436 17556
rect 34748 75682 34804 75684
rect 34748 75630 34750 75682
rect 34750 75630 34802 75682
rect 34802 75630 34804 75682
rect 34748 75628 34804 75630
rect 34972 75852 35028 75908
rect 35196 76074 35252 76076
rect 35196 76022 35198 76074
rect 35198 76022 35250 76074
rect 35250 76022 35252 76074
rect 35196 76020 35252 76022
rect 35300 76074 35356 76076
rect 35300 76022 35302 76074
rect 35302 76022 35354 76074
rect 35354 76022 35356 76074
rect 35300 76020 35356 76022
rect 35404 76074 35460 76076
rect 35404 76022 35406 76074
rect 35406 76022 35458 76074
rect 35458 76022 35460 76074
rect 35404 76020 35460 76022
rect 35196 75794 35252 75796
rect 35196 75742 35198 75794
rect 35198 75742 35250 75794
rect 35250 75742 35252 75794
rect 35196 75740 35252 75742
rect 35532 75628 35588 75684
rect 35084 74786 35140 74788
rect 35084 74734 35086 74786
rect 35086 74734 35138 74786
rect 35138 74734 35140 74786
rect 35084 74732 35140 74734
rect 35196 74506 35252 74508
rect 35196 74454 35198 74506
rect 35198 74454 35250 74506
rect 35250 74454 35252 74506
rect 35196 74452 35252 74454
rect 35300 74506 35356 74508
rect 35300 74454 35302 74506
rect 35302 74454 35354 74506
rect 35354 74454 35356 74506
rect 35300 74452 35356 74454
rect 35404 74506 35460 74508
rect 35404 74454 35406 74506
rect 35406 74454 35458 74506
rect 35458 74454 35460 74506
rect 35404 74452 35460 74454
rect 35196 72938 35252 72940
rect 35196 72886 35198 72938
rect 35198 72886 35250 72938
rect 35250 72886 35252 72938
rect 35196 72884 35252 72886
rect 35300 72938 35356 72940
rect 35300 72886 35302 72938
rect 35302 72886 35354 72938
rect 35354 72886 35356 72938
rect 35300 72884 35356 72886
rect 35404 72938 35460 72940
rect 35404 72886 35406 72938
rect 35406 72886 35458 72938
rect 35458 72886 35460 72938
rect 35404 72884 35460 72886
rect 35196 71370 35252 71372
rect 35196 71318 35198 71370
rect 35198 71318 35250 71370
rect 35250 71318 35252 71370
rect 35196 71316 35252 71318
rect 35300 71370 35356 71372
rect 35300 71318 35302 71370
rect 35302 71318 35354 71370
rect 35354 71318 35356 71370
rect 35300 71316 35356 71318
rect 35404 71370 35460 71372
rect 35404 71318 35406 71370
rect 35406 71318 35458 71370
rect 35458 71318 35460 71370
rect 35404 71316 35460 71318
rect 35196 69802 35252 69804
rect 35196 69750 35198 69802
rect 35198 69750 35250 69802
rect 35250 69750 35252 69802
rect 35196 69748 35252 69750
rect 35300 69802 35356 69804
rect 35300 69750 35302 69802
rect 35302 69750 35354 69802
rect 35354 69750 35356 69802
rect 35300 69748 35356 69750
rect 35404 69802 35460 69804
rect 35404 69750 35406 69802
rect 35406 69750 35458 69802
rect 35458 69750 35460 69802
rect 35404 69748 35460 69750
rect 35196 68234 35252 68236
rect 35196 68182 35198 68234
rect 35198 68182 35250 68234
rect 35250 68182 35252 68234
rect 35196 68180 35252 68182
rect 35300 68234 35356 68236
rect 35300 68182 35302 68234
rect 35302 68182 35354 68234
rect 35354 68182 35356 68234
rect 35300 68180 35356 68182
rect 35404 68234 35460 68236
rect 35404 68182 35406 68234
rect 35406 68182 35458 68234
rect 35458 68182 35460 68234
rect 35404 68180 35460 68182
rect 35196 66666 35252 66668
rect 35196 66614 35198 66666
rect 35198 66614 35250 66666
rect 35250 66614 35252 66666
rect 35196 66612 35252 66614
rect 35300 66666 35356 66668
rect 35300 66614 35302 66666
rect 35302 66614 35354 66666
rect 35354 66614 35356 66666
rect 35300 66612 35356 66614
rect 35404 66666 35460 66668
rect 35404 66614 35406 66666
rect 35406 66614 35458 66666
rect 35458 66614 35460 66666
rect 35404 66612 35460 66614
rect 35196 65098 35252 65100
rect 35196 65046 35198 65098
rect 35198 65046 35250 65098
rect 35250 65046 35252 65098
rect 35196 65044 35252 65046
rect 35300 65098 35356 65100
rect 35300 65046 35302 65098
rect 35302 65046 35354 65098
rect 35354 65046 35356 65098
rect 35300 65044 35356 65046
rect 35404 65098 35460 65100
rect 35404 65046 35406 65098
rect 35406 65046 35458 65098
rect 35458 65046 35460 65098
rect 35404 65044 35460 65046
rect 35196 63530 35252 63532
rect 35196 63478 35198 63530
rect 35198 63478 35250 63530
rect 35250 63478 35252 63530
rect 35196 63476 35252 63478
rect 35300 63530 35356 63532
rect 35300 63478 35302 63530
rect 35302 63478 35354 63530
rect 35354 63478 35356 63530
rect 35300 63476 35356 63478
rect 35404 63530 35460 63532
rect 35404 63478 35406 63530
rect 35406 63478 35458 63530
rect 35458 63478 35460 63530
rect 35404 63476 35460 63478
rect 35196 61962 35252 61964
rect 35196 61910 35198 61962
rect 35198 61910 35250 61962
rect 35250 61910 35252 61962
rect 35196 61908 35252 61910
rect 35300 61962 35356 61964
rect 35300 61910 35302 61962
rect 35302 61910 35354 61962
rect 35354 61910 35356 61962
rect 35300 61908 35356 61910
rect 35404 61962 35460 61964
rect 35404 61910 35406 61962
rect 35406 61910 35458 61962
rect 35458 61910 35460 61962
rect 35404 61908 35460 61910
rect 35196 60394 35252 60396
rect 35196 60342 35198 60394
rect 35198 60342 35250 60394
rect 35250 60342 35252 60394
rect 35196 60340 35252 60342
rect 35300 60394 35356 60396
rect 35300 60342 35302 60394
rect 35302 60342 35354 60394
rect 35354 60342 35356 60394
rect 35300 60340 35356 60342
rect 35404 60394 35460 60396
rect 35404 60342 35406 60394
rect 35406 60342 35458 60394
rect 35458 60342 35460 60394
rect 35404 60340 35460 60342
rect 35196 58826 35252 58828
rect 35196 58774 35198 58826
rect 35198 58774 35250 58826
rect 35250 58774 35252 58826
rect 35196 58772 35252 58774
rect 35300 58826 35356 58828
rect 35300 58774 35302 58826
rect 35302 58774 35354 58826
rect 35354 58774 35356 58826
rect 35300 58772 35356 58774
rect 35404 58826 35460 58828
rect 35404 58774 35406 58826
rect 35406 58774 35458 58826
rect 35458 58774 35460 58826
rect 35404 58772 35460 58774
rect 35196 57258 35252 57260
rect 35196 57206 35198 57258
rect 35198 57206 35250 57258
rect 35250 57206 35252 57258
rect 35196 57204 35252 57206
rect 35300 57258 35356 57260
rect 35300 57206 35302 57258
rect 35302 57206 35354 57258
rect 35354 57206 35356 57258
rect 35300 57204 35356 57206
rect 35404 57258 35460 57260
rect 35404 57206 35406 57258
rect 35406 57206 35458 57258
rect 35458 57206 35460 57258
rect 35404 57204 35460 57206
rect 35196 55690 35252 55692
rect 35196 55638 35198 55690
rect 35198 55638 35250 55690
rect 35250 55638 35252 55690
rect 35196 55636 35252 55638
rect 35300 55690 35356 55692
rect 35300 55638 35302 55690
rect 35302 55638 35354 55690
rect 35354 55638 35356 55690
rect 35300 55636 35356 55638
rect 35404 55690 35460 55692
rect 35404 55638 35406 55690
rect 35406 55638 35458 55690
rect 35458 55638 35460 55690
rect 35404 55636 35460 55638
rect 36876 75068 36932 75124
rect 37660 75122 37716 75124
rect 37660 75070 37662 75122
rect 37662 75070 37714 75122
rect 37714 75070 37716 75122
rect 37660 75068 37716 75070
rect 37996 75852 38052 75908
rect 41020 76690 41076 76692
rect 41020 76638 41022 76690
rect 41022 76638 41074 76690
rect 41074 76638 41076 76690
rect 41020 76636 41076 76638
rect 42028 76690 42084 76692
rect 42028 76638 42030 76690
rect 42030 76638 42082 76690
rect 42082 76638 42084 76690
rect 42028 76636 42084 76638
rect 35196 54122 35252 54124
rect 35196 54070 35198 54122
rect 35198 54070 35250 54122
rect 35250 54070 35252 54122
rect 35196 54068 35252 54070
rect 35300 54122 35356 54124
rect 35300 54070 35302 54122
rect 35302 54070 35354 54122
rect 35354 54070 35356 54122
rect 35300 54068 35356 54070
rect 35404 54122 35460 54124
rect 35404 54070 35406 54122
rect 35406 54070 35458 54122
rect 35458 54070 35460 54122
rect 35404 54068 35460 54070
rect 35196 52554 35252 52556
rect 35196 52502 35198 52554
rect 35198 52502 35250 52554
rect 35250 52502 35252 52554
rect 35196 52500 35252 52502
rect 35300 52554 35356 52556
rect 35300 52502 35302 52554
rect 35302 52502 35354 52554
rect 35354 52502 35356 52554
rect 35300 52500 35356 52502
rect 35404 52554 35460 52556
rect 35404 52502 35406 52554
rect 35406 52502 35458 52554
rect 35458 52502 35460 52554
rect 35404 52500 35460 52502
rect 35196 50986 35252 50988
rect 35196 50934 35198 50986
rect 35198 50934 35250 50986
rect 35250 50934 35252 50986
rect 35196 50932 35252 50934
rect 35300 50986 35356 50988
rect 35300 50934 35302 50986
rect 35302 50934 35354 50986
rect 35354 50934 35356 50986
rect 35300 50932 35356 50934
rect 35404 50986 35460 50988
rect 35404 50934 35406 50986
rect 35406 50934 35458 50986
rect 35458 50934 35460 50986
rect 35404 50932 35460 50934
rect 35196 49418 35252 49420
rect 35196 49366 35198 49418
rect 35198 49366 35250 49418
rect 35250 49366 35252 49418
rect 35196 49364 35252 49366
rect 35300 49418 35356 49420
rect 35300 49366 35302 49418
rect 35302 49366 35354 49418
rect 35354 49366 35356 49418
rect 35300 49364 35356 49366
rect 35404 49418 35460 49420
rect 35404 49366 35406 49418
rect 35406 49366 35458 49418
rect 35458 49366 35460 49418
rect 35404 49364 35460 49366
rect 35196 47850 35252 47852
rect 35196 47798 35198 47850
rect 35198 47798 35250 47850
rect 35250 47798 35252 47850
rect 35196 47796 35252 47798
rect 35300 47850 35356 47852
rect 35300 47798 35302 47850
rect 35302 47798 35354 47850
rect 35354 47798 35356 47850
rect 35300 47796 35356 47798
rect 35404 47850 35460 47852
rect 35404 47798 35406 47850
rect 35406 47798 35458 47850
rect 35458 47798 35460 47850
rect 35404 47796 35460 47798
rect 35196 46282 35252 46284
rect 35196 46230 35198 46282
rect 35198 46230 35250 46282
rect 35250 46230 35252 46282
rect 35196 46228 35252 46230
rect 35300 46282 35356 46284
rect 35300 46230 35302 46282
rect 35302 46230 35354 46282
rect 35354 46230 35356 46282
rect 35300 46228 35356 46230
rect 35404 46282 35460 46284
rect 35404 46230 35406 46282
rect 35406 46230 35458 46282
rect 35458 46230 35460 46282
rect 35404 46228 35460 46230
rect 35196 44714 35252 44716
rect 35196 44662 35198 44714
rect 35198 44662 35250 44714
rect 35250 44662 35252 44714
rect 35196 44660 35252 44662
rect 35300 44714 35356 44716
rect 35300 44662 35302 44714
rect 35302 44662 35354 44714
rect 35354 44662 35356 44714
rect 35300 44660 35356 44662
rect 35404 44714 35460 44716
rect 35404 44662 35406 44714
rect 35406 44662 35458 44714
rect 35458 44662 35460 44714
rect 35404 44660 35460 44662
rect 35196 43146 35252 43148
rect 35196 43094 35198 43146
rect 35198 43094 35250 43146
rect 35250 43094 35252 43146
rect 35196 43092 35252 43094
rect 35300 43146 35356 43148
rect 35300 43094 35302 43146
rect 35302 43094 35354 43146
rect 35354 43094 35356 43146
rect 35300 43092 35356 43094
rect 35404 43146 35460 43148
rect 35404 43094 35406 43146
rect 35406 43094 35458 43146
rect 35458 43094 35460 43146
rect 35404 43092 35460 43094
rect 35196 41578 35252 41580
rect 35196 41526 35198 41578
rect 35198 41526 35250 41578
rect 35250 41526 35252 41578
rect 35196 41524 35252 41526
rect 35300 41578 35356 41580
rect 35300 41526 35302 41578
rect 35302 41526 35354 41578
rect 35354 41526 35356 41578
rect 35300 41524 35356 41526
rect 35404 41578 35460 41580
rect 35404 41526 35406 41578
rect 35406 41526 35458 41578
rect 35458 41526 35460 41578
rect 35404 41524 35460 41526
rect 35196 40010 35252 40012
rect 35196 39958 35198 40010
rect 35198 39958 35250 40010
rect 35250 39958 35252 40010
rect 35196 39956 35252 39958
rect 35300 40010 35356 40012
rect 35300 39958 35302 40010
rect 35302 39958 35354 40010
rect 35354 39958 35356 40010
rect 35300 39956 35356 39958
rect 35404 40010 35460 40012
rect 35404 39958 35406 40010
rect 35406 39958 35458 40010
rect 35458 39958 35460 40010
rect 35404 39956 35460 39958
rect 35196 38442 35252 38444
rect 35196 38390 35198 38442
rect 35198 38390 35250 38442
rect 35250 38390 35252 38442
rect 35196 38388 35252 38390
rect 35300 38442 35356 38444
rect 35300 38390 35302 38442
rect 35302 38390 35354 38442
rect 35354 38390 35356 38442
rect 35300 38388 35356 38390
rect 35404 38442 35460 38444
rect 35404 38390 35406 38442
rect 35406 38390 35458 38442
rect 35458 38390 35460 38442
rect 35404 38388 35460 38390
rect 35196 36874 35252 36876
rect 35196 36822 35198 36874
rect 35198 36822 35250 36874
rect 35250 36822 35252 36874
rect 35196 36820 35252 36822
rect 35300 36874 35356 36876
rect 35300 36822 35302 36874
rect 35302 36822 35354 36874
rect 35354 36822 35356 36874
rect 35300 36820 35356 36822
rect 35404 36874 35460 36876
rect 35404 36822 35406 36874
rect 35406 36822 35458 36874
rect 35458 36822 35460 36874
rect 35404 36820 35460 36822
rect 35196 35306 35252 35308
rect 35196 35254 35198 35306
rect 35198 35254 35250 35306
rect 35250 35254 35252 35306
rect 35196 35252 35252 35254
rect 35300 35306 35356 35308
rect 35300 35254 35302 35306
rect 35302 35254 35354 35306
rect 35354 35254 35356 35306
rect 35300 35252 35356 35254
rect 35404 35306 35460 35308
rect 35404 35254 35406 35306
rect 35406 35254 35458 35306
rect 35458 35254 35460 35306
rect 35404 35252 35460 35254
rect 35196 33738 35252 33740
rect 35196 33686 35198 33738
rect 35198 33686 35250 33738
rect 35250 33686 35252 33738
rect 35196 33684 35252 33686
rect 35300 33738 35356 33740
rect 35300 33686 35302 33738
rect 35302 33686 35354 33738
rect 35354 33686 35356 33738
rect 35300 33684 35356 33686
rect 35404 33738 35460 33740
rect 35404 33686 35406 33738
rect 35406 33686 35458 33738
rect 35458 33686 35460 33738
rect 35404 33684 35460 33686
rect 35196 32170 35252 32172
rect 35196 32118 35198 32170
rect 35198 32118 35250 32170
rect 35250 32118 35252 32170
rect 35196 32116 35252 32118
rect 35300 32170 35356 32172
rect 35300 32118 35302 32170
rect 35302 32118 35354 32170
rect 35354 32118 35356 32170
rect 35300 32116 35356 32118
rect 35404 32170 35460 32172
rect 35404 32118 35406 32170
rect 35406 32118 35458 32170
rect 35458 32118 35460 32170
rect 35404 32116 35460 32118
rect 35196 30602 35252 30604
rect 35196 30550 35198 30602
rect 35198 30550 35250 30602
rect 35250 30550 35252 30602
rect 35196 30548 35252 30550
rect 35300 30602 35356 30604
rect 35300 30550 35302 30602
rect 35302 30550 35354 30602
rect 35354 30550 35356 30602
rect 35300 30548 35356 30550
rect 35404 30602 35460 30604
rect 35404 30550 35406 30602
rect 35406 30550 35458 30602
rect 35458 30550 35460 30602
rect 35404 30548 35460 30550
rect 34972 29148 35028 29204
rect 35196 29034 35252 29036
rect 35196 28982 35198 29034
rect 35198 28982 35250 29034
rect 35250 28982 35252 29034
rect 35196 28980 35252 28982
rect 35300 29034 35356 29036
rect 35300 28982 35302 29034
rect 35302 28982 35354 29034
rect 35354 28982 35356 29034
rect 35300 28980 35356 28982
rect 35404 29034 35460 29036
rect 35404 28982 35406 29034
rect 35406 28982 35458 29034
rect 35458 28982 35460 29034
rect 35404 28980 35460 28982
rect 33516 27804 33572 27860
rect 34524 27916 34580 27972
rect 33404 27692 33460 27748
rect 31836 24780 31892 24836
rect 31836 22764 31892 22820
rect 33180 24556 33236 24612
rect 32956 21868 33012 21924
rect 31388 20860 31444 20916
rect 31612 20018 31668 20020
rect 31612 19966 31614 20018
rect 31614 19966 31666 20018
rect 31666 19966 31668 20018
rect 31612 19964 31668 19966
rect 31164 18060 31220 18116
rect 32172 19740 32228 19796
rect 32620 19906 32676 19908
rect 32620 19854 32622 19906
rect 32622 19854 32674 19906
rect 32674 19854 32676 19906
rect 32620 19852 32676 19854
rect 31836 19292 31892 19348
rect 31276 17554 31332 17556
rect 31276 17502 31278 17554
rect 31278 17502 31330 17554
rect 31330 17502 31332 17554
rect 31276 17500 31332 17502
rect 29708 17052 29764 17108
rect 29484 16882 29540 16884
rect 29484 16830 29486 16882
rect 29486 16830 29538 16882
rect 29538 16830 29540 16882
rect 29484 16828 29540 16830
rect 29260 16492 29316 16548
rect 28588 14700 28644 14756
rect 29708 15596 29764 15652
rect 29484 14530 29540 14532
rect 29484 14478 29486 14530
rect 29486 14478 29538 14530
rect 29538 14478 29540 14530
rect 29484 14476 29540 14478
rect 30828 14476 30884 14532
rect 32284 17276 32340 17332
rect 32508 18338 32564 18340
rect 32508 18286 32510 18338
rect 32510 18286 32562 18338
rect 32562 18286 32564 18338
rect 32508 18284 32564 18286
rect 32732 17052 32788 17108
rect 31836 16044 31892 16100
rect 29708 13916 29764 13972
rect 28476 13858 28532 13860
rect 28476 13806 28478 13858
rect 28478 13806 28530 13858
rect 28530 13806 28532 13858
rect 28476 13804 28532 13806
rect 29036 13858 29092 13860
rect 29036 13806 29038 13858
rect 29038 13806 29090 13858
rect 29090 13806 29092 13858
rect 29036 13804 29092 13806
rect 28588 13468 28644 13524
rect 28364 12796 28420 12852
rect 28588 12572 28644 12628
rect 29372 12572 29428 12628
rect 29484 12850 29540 12852
rect 29484 12798 29486 12850
rect 29486 12798 29538 12850
rect 29538 12798 29540 12850
rect 29484 12796 29540 12798
rect 30268 13916 30324 13972
rect 30940 14252 30996 14308
rect 29932 13858 29988 13860
rect 29932 13806 29934 13858
rect 29934 13806 29986 13858
rect 29986 13806 29988 13858
rect 29932 13804 29988 13806
rect 28588 11676 28644 11732
rect 27916 10780 27972 10836
rect 28476 10610 28532 10612
rect 28476 10558 28478 10610
rect 28478 10558 28530 10610
rect 28530 10558 28532 10610
rect 28476 10556 28532 10558
rect 27804 9938 27860 9940
rect 27804 9886 27806 9938
rect 27806 9886 27858 9938
rect 27858 9886 27860 9938
rect 27804 9884 27860 9886
rect 28028 10108 28084 10164
rect 27804 9436 27860 9492
rect 27468 8876 27524 8932
rect 27356 8370 27412 8372
rect 27356 8318 27358 8370
rect 27358 8318 27410 8370
rect 27410 8318 27412 8370
rect 27356 8316 27412 8318
rect 27580 8034 27636 8036
rect 27580 7982 27582 8034
rect 27582 7982 27634 8034
rect 27634 7982 27636 8034
rect 27580 7980 27636 7982
rect 27244 6690 27300 6692
rect 27244 6638 27246 6690
rect 27246 6638 27298 6690
rect 27298 6638 27300 6690
rect 27244 6636 27300 6638
rect 27692 7586 27748 7588
rect 27692 7534 27694 7586
rect 27694 7534 27746 7586
rect 27746 7534 27748 7586
rect 27692 7532 27748 7534
rect 27692 7250 27748 7252
rect 27692 7198 27694 7250
rect 27694 7198 27746 7250
rect 27746 7198 27748 7250
rect 27692 7196 27748 7198
rect 28588 9100 28644 9156
rect 28140 8482 28196 8484
rect 28140 8430 28142 8482
rect 28142 8430 28194 8482
rect 28194 8430 28196 8482
rect 28140 8428 28196 8430
rect 28140 8146 28196 8148
rect 28140 8094 28142 8146
rect 28142 8094 28194 8146
rect 28194 8094 28196 8146
rect 28140 8092 28196 8094
rect 27804 6860 27860 6916
rect 27916 6636 27972 6692
rect 27804 6300 27860 6356
rect 28028 6578 28084 6580
rect 28028 6526 28030 6578
rect 28030 6526 28082 6578
rect 28082 6526 28084 6578
rect 28028 6524 28084 6526
rect 28812 8930 28868 8932
rect 28812 8878 28814 8930
rect 28814 8878 28866 8930
rect 28866 8878 28868 8930
rect 28812 8876 28868 8878
rect 28588 8092 28644 8148
rect 28364 7532 28420 7588
rect 28476 7362 28532 7364
rect 28476 7310 28478 7362
rect 28478 7310 28530 7362
rect 28530 7310 28532 7362
rect 28476 7308 28532 7310
rect 28252 6860 28308 6916
rect 28364 6412 28420 6468
rect 28140 6076 28196 6132
rect 27244 5628 27300 5684
rect 27244 5180 27300 5236
rect 26460 5068 26516 5124
rect 26460 4284 26516 4340
rect 26908 3388 26964 3444
rect 26684 3164 26740 3220
rect 26684 2604 26740 2660
rect 25900 1596 25956 1652
rect 27132 4508 27188 4564
rect 27916 5852 27972 5908
rect 27692 5682 27748 5684
rect 27692 5630 27694 5682
rect 27694 5630 27746 5682
rect 27746 5630 27748 5682
rect 27692 5628 27748 5630
rect 27804 5516 27860 5572
rect 28252 6188 28308 6244
rect 29932 11676 29988 11732
rect 30380 11282 30436 11284
rect 30380 11230 30382 11282
rect 30382 11230 30434 11282
rect 30434 11230 30436 11282
rect 30380 11228 30436 11230
rect 30156 11170 30212 11172
rect 30156 11118 30158 11170
rect 30158 11118 30210 11170
rect 30210 11118 30212 11170
rect 30156 11116 30212 11118
rect 32508 16098 32564 16100
rect 32508 16046 32510 16098
rect 32510 16046 32562 16098
rect 32562 16046 32564 16098
rect 32508 16044 32564 16046
rect 34076 27074 34132 27076
rect 34076 27022 34078 27074
rect 34078 27022 34130 27074
rect 34130 27022 34132 27074
rect 34076 27020 34132 27022
rect 33404 22988 33460 23044
rect 34300 23548 34356 23604
rect 35756 28028 35812 28084
rect 34972 27244 35028 27300
rect 34748 23938 34804 23940
rect 34748 23886 34750 23938
rect 34750 23886 34802 23938
rect 34802 23886 34804 23938
rect 34748 23884 34804 23886
rect 35308 27858 35364 27860
rect 35308 27806 35310 27858
rect 35310 27806 35362 27858
rect 35362 27806 35364 27858
rect 35308 27804 35364 27806
rect 35196 27466 35252 27468
rect 35196 27414 35198 27466
rect 35198 27414 35250 27466
rect 35250 27414 35252 27466
rect 35196 27412 35252 27414
rect 35300 27466 35356 27468
rect 35300 27414 35302 27466
rect 35302 27414 35354 27466
rect 35354 27414 35356 27466
rect 35300 27412 35356 27414
rect 35404 27466 35460 27468
rect 35404 27414 35406 27466
rect 35406 27414 35458 27466
rect 35458 27414 35460 27466
rect 35404 27412 35460 27414
rect 34972 26962 35028 26964
rect 34972 26910 34974 26962
rect 34974 26910 35026 26962
rect 35026 26910 35028 26962
rect 34972 26908 35028 26910
rect 35420 26796 35476 26852
rect 35196 26514 35252 26516
rect 35196 26462 35198 26514
rect 35198 26462 35250 26514
rect 35250 26462 35252 26514
rect 35196 26460 35252 26462
rect 35644 26962 35700 26964
rect 35644 26910 35646 26962
rect 35646 26910 35698 26962
rect 35698 26910 35700 26962
rect 35644 26908 35700 26910
rect 35196 25898 35252 25900
rect 35196 25846 35198 25898
rect 35198 25846 35250 25898
rect 35250 25846 35252 25898
rect 35196 25844 35252 25846
rect 35300 25898 35356 25900
rect 35300 25846 35302 25898
rect 35302 25846 35354 25898
rect 35354 25846 35356 25898
rect 35300 25844 35356 25846
rect 35404 25898 35460 25900
rect 35404 25846 35406 25898
rect 35406 25846 35458 25898
rect 35458 25846 35460 25898
rect 35404 25844 35460 25846
rect 35532 25452 35588 25508
rect 35420 24892 35476 24948
rect 35196 24330 35252 24332
rect 35196 24278 35198 24330
rect 35198 24278 35250 24330
rect 35250 24278 35252 24330
rect 35196 24276 35252 24278
rect 35300 24330 35356 24332
rect 35300 24278 35302 24330
rect 35302 24278 35354 24330
rect 35354 24278 35356 24330
rect 35300 24276 35356 24278
rect 35404 24330 35460 24332
rect 35404 24278 35406 24330
rect 35406 24278 35458 24330
rect 35458 24278 35460 24330
rect 35404 24276 35460 24278
rect 35084 23714 35140 23716
rect 35084 23662 35086 23714
rect 35086 23662 35138 23714
rect 35138 23662 35140 23714
rect 35084 23660 35140 23662
rect 34188 23154 34244 23156
rect 34188 23102 34190 23154
rect 34190 23102 34242 23154
rect 34242 23102 34244 23154
rect 34188 23100 34244 23102
rect 33292 20860 33348 20916
rect 33516 20636 33572 20692
rect 34860 23100 34916 23156
rect 34748 21532 34804 21588
rect 34524 21474 34580 21476
rect 34524 21422 34526 21474
rect 34526 21422 34578 21474
rect 34578 21422 34580 21474
rect 34524 21420 34580 21422
rect 34636 20412 34692 20468
rect 34412 20242 34468 20244
rect 34412 20190 34414 20242
rect 34414 20190 34466 20242
rect 34466 20190 34468 20242
rect 34412 20188 34468 20190
rect 34860 21308 34916 21364
rect 35308 23100 35364 23156
rect 37660 28476 37716 28532
rect 36652 28364 36708 28420
rect 36204 27074 36260 27076
rect 36204 27022 36206 27074
rect 36206 27022 36258 27074
rect 36258 27022 36260 27074
rect 36204 27020 36260 27022
rect 35980 26460 36036 26516
rect 35644 23826 35700 23828
rect 35644 23774 35646 23826
rect 35646 23774 35698 23826
rect 35698 23774 35700 23826
rect 35644 23772 35700 23774
rect 35980 23548 36036 23604
rect 35756 23154 35812 23156
rect 35756 23102 35758 23154
rect 35758 23102 35810 23154
rect 35810 23102 35812 23154
rect 35756 23100 35812 23102
rect 36428 25394 36484 25396
rect 36428 25342 36430 25394
rect 36430 25342 36482 25394
rect 36482 25342 36484 25394
rect 36428 25340 36484 25342
rect 37100 28082 37156 28084
rect 37100 28030 37102 28082
rect 37102 28030 37154 28082
rect 37154 28030 37156 28082
rect 37100 28028 37156 28030
rect 36652 27858 36708 27860
rect 36652 27806 36654 27858
rect 36654 27806 36706 27858
rect 36706 27806 36708 27858
rect 36652 27804 36708 27806
rect 36988 27074 37044 27076
rect 36988 27022 36990 27074
rect 36990 27022 37042 27074
rect 37042 27022 37044 27074
rect 36988 27020 37044 27022
rect 37324 25676 37380 25732
rect 37772 25618 37828 25620
rect 37772 25566 37774 25618
rect 37774 25566 37826 25618
rect 37826 25566 37828 25618
rect 37772 25564 37828 25566
rect 40124 75628 40180 75684
rect 38892 29148 38948 29204
rect 38556 28476 38612 28532
rect 40908 75682 40964 75684
rect 40908 75630 40910 75682
rect 40910 75630 40962 75682
rect 40962 75630 40964 75682
rect 40908 75628 40964 75630
rect 44156 76636 44212 76692
rect 45836 76636 45892 76692
rect 46172 76636 46228 76692
rect 41132 39058 41188 39060
rect 41132 39006 41134 39058
rect 41134 39006 41186 39058
rect 41186 39006 41188 39058
rect 41132 39004 41188 39006
rect 40796 38892 40852 38948
rect 41692 38834 41748 38836
rect 41692 38782 41694 38834
rect 41694 38782 41746 38834
rect 41746 38782 41748 38834
rect 41692 38780 41748 38782
rect 41580 38722 41636 38724
rect 41580 38670 41582 38722
rect 41582 38670 41634 38722
rect 41634 38670 41636 38722
rect 41580 38668 41636 38670
rect 39116 28028 39172 28084
rect 38332 26124 38388 26180
rect 38444 25900 38500 25956
rect 38332 25788 38388 25844
rect 37324 25340 37380 25396
rect 37436 24556 37492 24612
rect 37212 24332 37268 24388
rect 37884 24722 37940 24724
rect 37884 24670 37886 24722
rect 37886 24670 37938 24722
rect 37938 24670 37940 24722
rect 37884 24668 37940 24670
rect 37884 24220 37940 24276
rect 37212 23884 37268 23940
rect 36540 23548 36596 23604
rect 36764 23548 36820 23604
rect 35532 22876 35588 22932
rect 35196 22762 35252 22764
rect 35196 22710 35198 22762
rect 35198 22710 35250 22762
rect 35250 22710 35252 22762
rect 35196 22708 35252 22710
rect 35300 22762 35356 22764
rect 35300 22710 35302 22762
rect 35302 22710 35354 22762
rect 35354 22710 35356 22762
rect 35300 22708 35356 22710
rect 35404 22762 35460 22764
rect 35404 22710 35406 22762
rect 35406 22710 35458 22762
rect 35458 22710 35460 22762
rect 35404 22708 35460 22710
rect 36204 22876 36260 22932
rect 35084 21586 35140 21588
rect 35084 21534 35086 21586
rect 35086 21534 35138 21586
rect 35138 21534 35140 21586
rect 35084 21532 35140 21534
rect 35308 22370 35364 22372
rect 35308 22318 35310 22370
rect 35310 22318 35362 22370
rect 35362 22318 35364 22370
rect 35308 22316 35364 22318
rect 35756 22316 35812 22372
rect 35308 21308 35364 21364
rect 35196 21194 35252 21196
rect 35196 21142 35198 21194
rect 35198 21142 35250 21194
rect 35250 21142 35252 21194
rect 35196 21140 35252 21142
rect 35300 21194 35356 21196
rect 35300 21142 35302 21194
rect 35302 21142 35354 21194
rect 35354 21142 35356 21194
rect 35300 21140 35356 21142
rect 35404 21194 35460 21196
rect 35404 21142 35406 21194
rect 35406 21142 35458 21194
rect 35458 21142 35460 21194
rect 35404 21140 35460 21142
rect 35420 20972 35476 21028
rect 34860 20802 34916 20804
rect 34860 20750 34862 20802
rect 34862 20750 34914 20802
rect 34914 20750 34916 20802
rect 34860 20748 34916 20750
rect 35196 20690 35252 20692
rect 35196 20638 35198 20690
rect 35198 20638 35250 20690
rect 35250 20638 35252 20690
rect 35196 20636 35252 20638
rect 35756 21586 35812 21588
rect 35756 21534 35758 21586
rect 35758 21534 35810 21586
rect 35810 21534 35812 21586
rect 35756 21532 35812 21534
rect 35980 20972 36036 21028
rect 36204 21308 36260 21364
rect 35756 20802 35812 20804
rect 35756 20750 35758 20802
rect 35758 20750 35810 20802
rect 35810 20750 35812 20802
rect 35756 20748 35812 20750
rect 35532 20690 35588 20692
rect 35532 20638 35534 20690
rect 35534 20638 35586 20690
rect 35586 20638 35588 20690
rect 35532 20636 35588 20638
rect 34748 20188 34804 20244
rect 35644 20412 35700 20468
rect 33852 19740 33908 19796
rect 33740 19628 33796 19684
rect 33516 18338 33572 18340
rect 33516 18286 33518 18338
rect 33518 18286 33570 18338
rect 33570 18286 33572 18338
rect 33516 18284 33572 18286
rect 34076 19068 34132 19124
rect 33628 18060 33684 18116
rect 33180 17836 33236 17892
rect 33740 17948 33796 18004
rect 35308 20076 35364 20132
rect 34748 19964 34804 20020
rect 35532 20130 35588 20132
rect 35532 20078 35534 20130
rect 35534 20078 35586 20130
rect 35586 20078 35588 20130
rect 35532 20076 35588 20078
rect 35420 20018 35476 20020
rect 35420 19966 35422 20018
rect 35422 19966 35474 20018
rect 35474 19966 35476 20018
rect 35420 19964 35476 19966
rect 34300 19906 34356 19908
rect 34300 19854 34302 19906
rect 34302 19854 34354 19906
rect 34354 19854 34356 19906
rect 34300 19852 34356 19854
rect 33404 17778 33460 17780
rect 33404 17726 33406 17778
rect 33406 17726 33458 17778
rect 33458 17726 33460 17778
rect 33404 17724 33460 17726
rect 36652 21868 36708 21924
rect 36540 21586 36596 21588
rect 36540 21534 36542 21586
rect 36542 21534 36594 21586
rect 36594 21534 36596 21586
rect 36540 21532 36596 21534
rect 36428 20802 36484 20804
rect 36428 20750 36430 20802
rect 36430 20750 36482 20802
rect 36482 20750 36484 20802
rect 36428 20748 36484 20750
rect 36540 20636 36596 20692
rect 36428 19964 36484 20020
rect 35196 19626 35252 19628
rect 35196 19574 35198 19626
rect 35198 19574 35250 19626
rect 35250 19574 35252 19626
rect 35196 19572 35252 19574
rect 35300 19626 35356 19628
rect 35300 19574 35302 19626
rect 35302 19574 35354 19626
rect 35354 19574 35356 19626
rect 35300 19572 35356 19574
rect 35404 19626 35460 19628
rect 35404 19574 35406 19626
rect 35406 19574 35458 19626
rect 35458 19574 35460 19626
rect 35404 19572 35460 19574
rect 35756 19628 35812 19684
rect 35756 19292 35812 19348
rect 36428 19516 36484 19572
rect 35420 19122 35476 19124
rect 35420 19070 35422 19122
rect 35422 19070 35474 19122
rect 35474 19070 35476 19122
rect 35420 19068 35476 19070
rect 34748 18396 34804 18452
rect 35532 18956 35588 19012
rect 35196 18058 35252 18060
rect 35196 18006 35198 18058
rect 35198 18006 35250 18058
rect 35250 18006 35252 18058
rect 35196 18004 35252 18006
rect 35300 18058 35356 18060
rect 35300 18006 35302 18058
rect 35302 18006 35354 18058
rect 35354 18006 35356 18058
rect 35300 18004 35356 18006
rect 35404 18058 35460 18060
rect 35404 18006 35406 18058
rect 35406 18006 35458 18058
rect 35458 18006 35460 18058
rect 35404 18004 35460 18006
rect 34412 17724 34468 17780
rect 34748 17778 34804 17780
rect 34748 17726 34750 17778
rect 34750 17726 34802 17778
rect 34802 17726 34804 17778
rect 34748 17724 34804 17726
rect 35084 17724 35140 17780
rect 32284 14588 32340 14644
rect 32508 14418 32564 14420
rect 32508 14366 32510 14418
rect 32510 14366 32562 14418
rect 32562 14366 32564 14418
rect 32508 14364 32564 14366
rect 31276 13746 31332 13748
rect 31276 13694 31278 13746
rect 31278 13694 31330 13746
rect 31330 13694 31332 13746
rect 31276 13692 31332 13694
rect 31164 13580 31220 13636
rect 31612 13746 31668 13748
rect 31612 13694 31614 13746
rect 31614 13694 31666 13746
rect 31666 13694 31668 13746
rect 31612 13692 31668 13694
rect 31500 12684 31556 12740
rect 31612 12572 31668 12628
rect 31948 13746 32004 13748
rect 31948 13694 31950 13746
rect 31950 13694 32002 13746
rect 32002 13694 32004 13746
rect 31948 13692 32004 13694
rect 32172 13580 32228 13636
rect 32620 13580 32676 13636
rect 32508 13468 32564 13524
rect 31052 11004 31108 11060
rect 31948 11900 32004 11956
rect 32508 12348 32564 12404
rect 32508 12066 32564 12068
rect 32508 12014 32510 12066
rect 32510 12014 32562 12066
rect 32562 12014 32564 12066
rect 32508 12012 32564 12014
rect 29708 10556 29764 10612
rect 29484 9714 29540 9716
rect 29484 9662 29486 9714
rect 29486 9662 29538 9714
rect 29538 9662 29540 9714
rect 29484 9660 29540 9662
rect 29260 9602 29316 9604
rect 29260 9550 29262 9602
rect 29262 9550 29314 9602
rect 29314 9550 29316 9602
rect 29260 9548 29316 9550
rect 31276 10498 31332 10500
rect 31276 10446 31278 10498
rect 31278 10446 31330 10498
rect 31330 10446 31332 10498
rect 31276 10444 31332 10446
rect 32508 11788 32564 11844
rect 31836 11282 31892 11284
rect 31836 11230 31838 11282
rect 31838 11230 31890 11282
rect 31890 11230 31892 11282
rect 31836 11228 31892 11230
rect 31612 10220 31668 10276
rect 32060 10332 32116 10388
rect 31724 10108 31780 10164
rect 32172 10108 32228 10164
rect 29708 9324 29764 9380
rect 29932 8428 29988 8484
rect 29596 8316 29652 8372
rect 30044 8316 30100 8372
rect 30268 8428 30324 8484
rect 29596 7868 29652 7924
rect 29484 7420 29540 7476
rect 29372 7362 29428 7364
rect 29372 7310 29374 7362
rect 29374 7310 29426 7362
rect 29426 7310 29428 7362
rect 29372 7308 29428 7310
rect 28700 6524 28756 6580
rect 29148 6860 29204 6916
rect 28700 6300 28756 6356
rect 28588 6188 28644 6244
rect 28588 5404 28644 5460
rect 27468 2940 27524 2996
rect 27916 3948 27972 4004
rect 27804 2828 27860 2884
rect 27580 1820 27636 1876
rect 28700 4338 28756 4340
rect 28700 4286 28702 4338
rect 28702 4286 28754 4338
rect 28754 4286 28756 4338
rect 28700 4284 28756 4286
rect 28364 3948 28420 4004
rect 28476 3612 28532 3668
rect 27244 1260 27300 1316
rect 28588 3442 28644 3444
rect 28588 3390 28590 3442
rect 28590 3390 28642 3442
rect 28642 3390 28644 3442
rect 28588 3388 28644 3390
rect 28588 2492 28644 2548
rect 29260 6578 29316 6580
rect 29260 6526 29262 6578
rect 29262 6526 29314 6578
rect 29314 6526 29316 6578
rect 29260 6524 29316 6526
rect 29372 6412 29428 6468
rect 32508 10834 32564 10836
rect 32508 10782 32510 10834
rect 32510 10782 32562 10834
rect 32562 10782 32564 10834
rect 32508 10780 32564 10782
rect 30492 9324 30548 9380
rect 29820 7196 29876 7252
rect 29708 6860 29764 6916
rect 29148 5964 29204 6020
rect 29260 5852 29316 5908
rect 29372 5964 29428 6020
rect 29260 5628 29316 5684
rect 28924 2940 28980 2996
rect 28812 2380 28868 2436
rect 29260 5122 29316 5124
rect 29260 5070 29262 5122
rect 29262 5070 29314 5122
rect 29314 5070 29316 5122
rect 29260 5068 29316 5070
rect 29708 6300 29764 6356
rect 29708 6076 29764 6132
rect 29708 5516 29764 5572
rect 29596 5346 29652 5348
rect 29596 5294 29598 5346
rect 29598 5294 29650 5346
rect 29650 5294 29652 5346
rect 29596 5292 29652 5294
rect 30156 6524 30212 6580
rect 30044 6466 30100 6468
rect 30044 6414 30046 6466
rect 30046 6414 30098 6466
rect 30098 6414 30100 6466
rect 30044 6412 30100 6414
rect 30044 5852 30100 5908
rect 30268 5794 30324 5796
rect 30268 5742 30270 5794
rect 30270 5742 30322 5794
rect 30322 5742 30324 5794
rect 30268 5740 30324 5742
rect 30156 5628 30212 5684
rect 30268 5346 30324 5348
rect 30268 5294 30270 5346
rect 30270 5294 30322 5346
rect 30322 5294 30324 5346
rect 30268 5292 30324 5294
rect 30156 5122 30212 5124
rect 30156 5070 30158 5122
rect 30158 5070 30210 5122
rect 30210 5070 30212 5122
rect 30156 5068 30212 5070
rect 29260 3836 29316 3892
rect 29260 3276 29316 3332
rect 29260 2268 29316 2324
rect 29148 1596 29204 1652
rect 30044 4898 30100 4900
rect 30044 4846 30046 4898
rect 30046 4846 30098 4898
rect 30098 4846 30100 4898
rect 30044 4844 30100 4846
rect 31164 9212 31220 9268
rect 31836 9212 31892 9268
rect 32620 9772 32676 9828
rect 32508 9548 32564 9604
rect 32284 8428 32340 8484
rect 32396 8652 32452 8708
rect 30828 7756 30884 7812
rect 30492 6076 30548 6132
rect 30492 5292 30548 5348
rect 31276 7586 31332 7588
rect 31276 7534 31278 7586
rect 31278 7534 31330 7586
rect 31330 7534 31332 7586
rect 31276 7532 31332 7534
rect 30940 7474 30996 7476
rect 30940 7422 30942 7474
rect 30942 7422 30994 7474
rect 30994 7422 30996 7474
rect 30940 7420 30996 7422
rect 30828 6300 30884 6356
rect 30940 6412 30996 6468
rect 32060 7586 32116 7588
rect 32060 7534 32062 7586
rect 32062 7534 32114 7586
rect 32114 7534 32116 7586
rect 32060 7532 32116 7534
rect 31724 7420 31780 7476
rect 31052 6076 31108 6132
rect 31052 5906 31108 5908
rect 31052 5854 31054 5906
rect 31054 5854 31106 5906
rect 31106 5854 31108 5906
rect 31052 5852 31108 5854
rect 31388 6300 31444 6356
rect 32956 13746 33012 13748
rect 32956 13694 32958 13746
rect 32958 13694 33010 13746
rect 33010 13694 33012 13746
rect 32956 13692 33012 13694
rect 32844 13468 32900 13524
rect 33404 15596 33460 15652
rect 33404 14364 33460 14420
rect 33404 14028 33460 14084
rect 33628 13970 33684 13972
rect 33628 13918 33630 13970
rect 33630 13918 33682 13970
rect 33682 13918 33684 13970
rect 33628 13916 33684 13918
rect 33292 13132 33348 13188
rect 32956 11394 33012 11396
rect 32956 11342 32958 11394
rect 32958 11342 33010 11394
rect 33010 11342 33012 11394
rect 32956 11340 33012 11342
rect 32956 10108 33012 10164
rect 33180 10108 33236 10164
rect 33292 11116 33348 11172
rect 34300 17554 34356 17556
rect 34300 17502 34302 17554
rect 34302 17502 34354 17554
rect 34354 17502 34356 17554
rect 34300 17500 34356 17502
rect 36092 17442 36148 17444
rect 36092 17390 36094 17442
rect 36094 17390 36146 17442
rect 36146 17390 36148 17442
rect 36092 17388 36148 17390
rect 35980 17164 36036 17220
rect 35420 17106 35476 17108
rect 35420 17054 35422 17106
rect 35422 17054 35474 17106
rect 35474 17054 35476 17106
rect 35420 17052 35476 17054
rect 33852 14812 33908 14868
rect 34076 14028 34132 14084
rect 37772 24108 37828 24164
rect 37324 22316 37380 22372
rect 36988 20690 37044 20692
rect 36988 20638 36990 20690
rect 36990 20638 37042 20690
rect 37042 20638 37044 20690
rect 36988 20636 37044 20638
rect 36764 18956 36820 19012
rect 36428 18844 36484 18900
rect 37100 17724 37156 17780
rect 36988 17554 37044 17556
rect 36988 17502 36990 17554
rect 36990 17502 37042 17554
rect 37042 17502 37044 17554
rect 36988 17500 37044 17502
rect 36316 17164 36372 17220
rect 36988 17164 37044 17220
rect 36204 16940 36260 16996
rect 35196 16490 35252 16492
rect 35196 16438 35198 16490
rect 35198 16438 35250 16490
rect 35250 16438 35252 16490
rect 35196 16436 35252 16438
rect 35300 16490 35356 16492
rect 35300 16438 35302 16490
rect 35302 16438 35354 16490
rect 35354 16438 35356 16490
rect 35300 16436 35356 16438
rect 35404 16490 35460 16492
rect 35404 16438 35406 16490
rect 35406 16438 35458 16490
rect 35458 16438 35460 16490
rect 35404 16436 35460 16438
rect 36988 16994 37044 16996
rect 36988 16942 36990 16994
rect 36990 16942 37042 16994
rect 37042 16942 37044 16994
rect 36988 16940 37044 16942
rect 36540 16828 36596 16884
rect 37436 22876 37492 22932
rect 37772 23826 37828 23828
rect 37772 23774 37774 23826
rect 37774 23774 37826 23826
rect 37826 23774 37828 23826
rect 37772 23772 37828 23774
rect 37660 23548 37716 23604
rect 37660 23324 37716 23380
rect 37772 22370 37828 22372
rect 37772 22318 37774 22370
rect 37774 22318 37826 22370
rect 37826 22318 37828 22370
rect 37772 22316 37828 22318
rect 37324 20578 37380 20580
rect 37324 20526 37326 20578
rect 37326 20526 37378 20578
rect 37378 20526 37380 20578
rect 37324 20524 37380 20526
rect 38108 23324 38164 23380
rect 38668 25788 38724 25844
rect 40348 28082 40404 28084
rect 40348 28030 40350 28082
rect 40350 28030 40402 28082
rect 40402 28030 40404 28082
rect 40348 28028 40404 28030
rect 40012 27356 40068 27412
rect 38780 25564 38836 25620
rect 38892 26124 38948 26180
rect 39452 25228 39508 25284
rect 38892 24332 38948 24388
rect 38556 22876 38612 22932
rect 38332 22204 38388 22260
rect 38556 22652 38612 22708
rect 37884 20076 37940 20132
rect 37996 19740 38052 19796
rect 37660 19180 37716 19236
rect 37324 18844 37380 18900
rect 37772 18284 37828 18340
rect 37436 18172 37492 18228
rect 37324 17388 37380 17444
rect 37548 17164 37604 17220
rect 38332 19234 38388 19236
rect 38332 19182 38334 19234
rect 38334 19182 38386 19234
rect 38386 19182 38388 19234
rect 38332 19180 38388 19182
rect 37884 17666 37940 17668
rect 37884 17614 37886 17666
rect 37886 17614 37938 17666
rect 37938 17614 37940 17666
rect 37884 17612 37940 17614
rect 36764 16268 36820 16324
rect 35980 15596 36036 15652
rect 35196 14922 35252 14924
rect 35196 14870 35198 14922
rect 35198 14870 35250 14922
rect 35250 14870 35252 14922
rect 35196 14868 35252 14870
rect 35300 14922 35356 14924
rect 35300 14870 35302 14922
rect 35302 14870 35354 14922
rect 35354 14870 35356 14922
rect 35300 14868 35356 14870
rect 35404 14922 35460 14924
rect 35404 14870 35406 14922
rect 35406 14870 35458 14922
rect 35458 14870 35460 14922
rect 35404 14868 35460 14870
rect 35532 14306 35588 14308
rect 35532 14254 35534 14306
rect 35534 14254 35586 14306
rect 35586 14254 35588 14306
rect 35532 14252 35588 14254
rect 34972 14028 35028 14084
rect 35756 15260 35812 15316
rect 37548 16716 37604 16772
rect 37324 16210 37380 16212
rect 37324 16158 37326 16210
rect 37326 16158 37378 16210
rect 37378 16158 37380 16210
rect 37324 16156 37380 16158
rect 37996 16940 38052 16996
rect 37996 16322 38052 16324
rect 37996 16270 37998 16322
rect 37998 16270 38050 16322
rect 38050 16270 38052 16322
rect 37996 16268 38052 16270
rect 37996 15202 38052 15204
rect 37996 15150 37998 15202
rect 37998 15150 38050 15202
rect 38050 15150 38052 15202
rect 37996 15148 38052 15150
rect 37996 14700 38052 14756
rect 36764 14252 36820 14308
rect 35308 13970 35364 13972
rect 35308 13918 35310 13970
rect 35310 13918 35362 13970
rect 35362 13918 35364 13970
rect 35308 13916 35364 13918
rect 35196 13354 35252 13356
rect 35196 13302 35198 13354
rect 35198 13302 35250 13354
rect 35250 13302 35252 13354
rect 35196 13300 35252 13302
rect 35300 13354 35356 13356
rect 35300 13302 35302 13354
rect 35302 13302 35354 13354
rect 35354 13302 35356 13354
rect 35300 13300 35356 13302
rect 35404 13354 35460 13356
rect 35404 13302 35406 13354
rect 35406 13302 35458 13354
rect 35458 13302 35460 13354
rect 35404 13300 35460 13302
rect 35644 13746 35700 13748
rect 35644 13694 35646 13746
rect 35646 13694 35698 13746
rect 35698 13694 35700 13746
rect 35644 13692 35700 13694
rect 34300 13020 34356 13076
rect 34636 12348 34692 12404
rect 35084 12402 35140 12404
rect 35084 12350 35086 12402
rect 35086 12350 35138 12402
rect 35138 12350 35140 12402
rect 35084 12348 35140 12350
rect 35980 13916 36036 13972
rect 37660 13804 37716 13860
rect 36988 13244 37044 13300
rect 36428 13074 36484 13076
rect 36428 13022 36430 13074
rect 36430 13022 36482 13074
rect 36482 13022 36484 13074
rect 36428 13020 36484 13022
rect 35644 12290 35700 12292
rect 35644 12238 35646 12290
rect 35646 12238 35698 12290
rect 35698 12238 35700 12290
rect 35644 12236 35700 12238
rect 36204 12290 36260 12292
rect 36204 12238 36206 12290
rect 36206 12238 36258 12290
rect 36258 12238 36260 12290
rect 36204 12236 36260 12238
rect 37772 13244 37828 13300
rect 37772 13074 37828 13076
rect 37772 13022 37774 13074
rect 37774 13022 37826 13074
rect 37826 13022 37828 13074
rect 37772 13020 37828 13022
rect 37996 13746 38052 13748
rect 37996 13694 37998 13746
rect 37998 13694 38050 13746
rect 38050 13694 38052 13746
rect 37996 13692 38052 13694
rect 37884 12796 37940 12852
rect 36988 11900 37044 11956
rect 37100 12572 37156 12628
rect 35196 11786 35252 11788
rect 35196 11734 35198 11786
rect 35198 11734 35250 11786
rect 35250 11734 35252 11786
rect 35196 11732 35252 11734
rect 35300 11786 35356 11788
rect 35300 11734 35302 11786
rect 35302 11734 35354 11786
rect 35354 11734 35356 11786
rect 35300 11732 35356 11734
rect 35404 11786 35460 11788
rect 35404 11734 35406 11786
rect 35406 11734 35458 11786
rect 35458 11734 35460 11786
rect 35404 11732 35460 11734
rect 33740 11452 33796 11508
rect 36428 11564 36484 11620
rect 33516 10668 33572 10724
rect 33292 10444 33348 10500
rect 36428 11340 36484 11396
rect 37884 12348 37940 12404
rect 37548 12178 37604 12180
rect 37548 12126 37550 12178
rect 37550 12126 37602 12178
rect 37602 12126 37604 12178
rect 37548 12124 37604 12126
rect 33068 9996 33124 10052
rect 33964 10050 34020 10052
rect 33964 9998 33966 10050
rect 33966 9998 34018 10050
rect 34018 9998 34020 10050
rect 33964 9996 34020 9998
rect 33516 9772 33572 9828
rect 33180 9714 33236 9716
rect 33180 9662 33182 9714
rect 33182 9662 33234 9714
rect 33234 9662 33236 9714
rect 33180 9660 33236 9662
rect 33292 9324 33348 9380
rect 32732 8876 32788 8932
rect 32956 9212 33012 9268
rect 37212 10892 37268 10948
rect 36988 10780 37044 10836
rect 35196 10218 35252 10220
rect 35196 10166 35198 10218
rect 35198 10166 35250 10218
rect 35250 10166 35252 10218
rect 35196 10164 35252 10166
rect 35300 10218 35356 10220
rect 35300 10166 35302 10218
rect 35302 10166 35354 10218
rect 35354 10166 35356 10218
rect 35300 10164 35356 10166
rect 35404 10218 35460 10220
rect 35404 10166 35406 10218
rect 35406 10166 35458 10218
rect 35458 10166 35460 10218
rect 35404 10164 35460 10166
rect 35756 10050 35812 10052
rect 35756 9998 35758 10050
rect 35758 9998 35810 10050
rect 35810 9998 35812 10050
rect 35756 9996 35812 9998
rect 34188 9436 34244 9492
rect 33852 8258 33908 8260
rect 33852 8206 33854 8258
rect 33854 8206 33906 8258
rect 33906 8206 33908 8258
rect 33852 8204 33908 8206
rect 32956 7420 33012 7476
rect 32172 6300 32228 6356
rect 31836 5740 31892 5796
rect 31276 5292 31332 5348
rect 31052 5180 31108 5236
rect 30604 4956 30660 5012
rect 30716 5068 30772 5124
rect 31836 5292 31892 5348
rect 31276 5122 31332 5124
rect 31276 5070 31278 5122
rect 31278 5070 31330 5122
rect 31330 5070 31332 5122
rect 31276 5068 31332 5070
rect 32172 6076 32228 6132
rect 32620 5906 32676 5908
rect 32620 5854 32622 5906
rect 32622 5854 32674 5906
rect 32674 5854 32676 5906
rect 32620 5852 32676 5854
rect 32172 5740 32228 5796
rect 30940 4732 30996 4788
rect 30044 4060 30100 4116
rect 29932 3500 29988 3556
rect 29932 3052 29988 3108
rect 30268 3724 30324 3780
rect 31836 4732 31892 4788
rect 31276 4450 31332 4452
rect 31276 4398 31278 4450
rect 31278 4398 31330 4450
rect 31330 4398 31332 4450
rect 31276 4396 31332 4398
rect 31388 4284 31444 4340
rect 30940 4060 30996 4116
rect 31164 3612 31220 3668
rect 30492 2716 30548 2772
rect 31836 4226 31892 4228
rect 31836 4174 31838 4226
rect 31838 4174 31890 4226
rect 31890 4174 31892 4226
rect 31836 4172 31892 4174
rect 31836 3948 31892 4004
rect 31612 3330 31668 3332
rect 31612 3278 31614 3330
rect 31614 3278 31666 3330
rect 31666 3278 31668 3330
rect 31612 3276 31668 3278
rect 32620 5404 32676 5460
rect 32396 4284 32452 4340
rect 32508 4620 32564 4676
rect 32732 4508 32788 4564
rect 33292 7868 33348 7924
rect 33404 7980 33460 8036
rect 34860 9602 34916 9604
rect 34860 9550 34862 9602
rect 34862 9550 34914 9602
rect 34914 9550 34916 9602
rect 34860 9548 34916 9550
rect 36204 9826 36260 9828
rect 36204 9774 36206 9826
rect 36206 9774 36258 9826
rect 36258 9774 36260 9826
rect 36204 9772 36260 9774
rect 37436 10556 37492 10612
rect 37324 9826 37380 9828
rect 37324 9774 37326 9826
rect 37326 9774 37378 9826
rect 37378 9774 37380 9826
rect 37324 9772 37380 9774
rect 36540 9714 36596 9716
rect 36540 9662 36542 9714
rect 36542 9662 36594 9714
rect 36594 9662 36596 9714
rect 36540 9660 36596 9662
rect 34748 8764 34804 8820
rect 35196 8650 35252 8652
rect 35196 8598 35198 8650
rect 35198 8598 35250 8650
rect 35250 8598 35252 8650
rect 35196 8596 35252 8598
rect 35300 8650 35356 8652
rect 35300 8598 35302 8650
rect 35302 8598 35354 8650
rect 35354 8598 35356 8650
rect 35300 8596 35356 8598
rect 35404 8650 35460 8652
rect 35404 8598 35406 8650
rect 35406 8598 35458 8650
rect 35458 8598 35460 8650
rect 35404 8596 35460 8598
rect 35420 8204 35476 8260
rect 34300 8146 34356 8148
rect 34300 8094 34302 8146
rect 34302 8094 34354 8146
rect 34354 8094 34356 8146
rect 34300 8092 34356 8094
rect 34524 8034 34580 8036
rect 34524 7982 34526 8034
rect 34526 7982 34578 8034
rect 34578 7982 34580 8034
rect 34524 7980 34580 7982
rect 33068 6300 33124 6356
rect 33180 6130 33236 6132
rect 33180 6078 33182 6130
rect 33182 6078 33234 6130
rect 33234 6078 33236 6130
rect 33180 6076 33236 6078
rect 33740 7474 33796 7476
rect 33740 7422 33742 7474
rect 33742 7422 33794 7474
rect 33794 7422 33796 7474
rect 33740 7420 33796 7422
rect 33404 6524 33460 6580
rect 33740 6578 33796 6580
rect 33740 6526 33742 6578
rect 33742 6526 33794 6578
rect 33794 6526 33796 6578
rect 33740 6524 33796 6526
rect 33964 6578 34020 6580
rect 33964 6526 33966 6578
rect 33966 6526 34018 6578
rect 34018 6526 34020 6578
rect 33964 6524 34020 6526
rect 33852 6466 33908 6468
rect 33852 6414 33854 6466
rect 33854 6414 33906 6466
rect 33906 6414 33908 6466
rect 33852 6412 33908 6414
rect 34412 7308 34468 7364
rect 34076 6412 34132 6468
rect 34412 6524 34468 6580
rect 33740 6076 33796 6132
rect 34412 6076 34468 6132
rect 33516 4956 33572 5012
rect 33740 5628 33796 5684
rect 34300 5628 34356 5684
rect 33628 4172 33684 4228
rect 32172 1596 32228 1652
rect 32508 2604 32564 2660
rect 34972 7868 35028 7924
rect 34860 7196 34916 7252
rect 35196 7308 35252 7364
rect 35420 7308 35476 7364
rect 35868 8876 35924 8932
rect 35532 7196 35588 7252
rect 35196 7082 35252 7084
rect 35196 7030 35198 7082
rect 35198 7030 35250 7082
rect 35250 7030 35252 7082
rect 35196 7028 35252 7030
rect 35300 7082 35356 7084
rect 35300 7030 35302 7082
rect 35302 7030 35354 7082
rect 35354 7030 35356 7082
rect 35300 7028 35356 7030
rect 35404 7082 35460 7084
rect 35404 7030 35406 7082
rect 35406 7030 35458 7082
rect 35458 7030 35460 7082
rect 35404 7028 35460 7030
rect 34972 6524 35028 6580
rect 35084 5964 35140 6020
rect 36092 7644 36148 7700
rect 35868 7532 35924 7588
rect 35756 7308 35812 7364
rect 34412 5516 34468 5572
rect 34076 5180 34132 5236
rect 33740 1372 33796 1428
rect 33852 5068 33908 5124
rect 35196 5514 35252 5516
rect 35196 5462 35198 5514
rect 35198 5462 35250 5514
rect 35250 5462 35252 5514
rect 35196 5460 35252 5462
rect 35300 5514 35356 5516
rect 35300 5462 35302 5514
rect 35302 5462 35354 5514
rect 35354 5462 35356 5514
rect 35300 5460 35356 5462
rect 35404 5514 35460 5516
rect 35404 5462 35406 5514
rect 35406 5462 35458 5514
rect 35458 5462 35460 5514
rect 35404 5460 35460 5462
rect 35084 4172 35140 4228
rect 35196 3946 35252 3948
rect 35196 3894 35198 3946
rect 35198 3894 35250 3946
rect 35250 3894 35252 3946
rect 35196 3892 35252 3894
rect 35300 3946 35356 3948
rect 35300 3894 35302 3946
rect 35302 3894 35354 3946
rect 35354 3894 35356 3946
rect 35300 3892 35356 3894
rect 35404 3946 35460 3948
rect 35404 3894 35406 3946
rect 35406 3894 35458 3946
rect 35458 3894 35460 3946
rect 35404 3892 35460 3894
rect 34972 3388 35028 3444
rect 35308 3442 35364 3444
rect 35308 3390 35310 3442
rect 35310 3390 35362 3442
rect 35362 3390 35364 3442
rect 35308 3388 35364 3390
rect 38556 19234 38612 19236
rect 38556 19182 38558 19234
rect 38558 19182 38610 19234
rect 38610 19182 38612 19234
rect 38556 19180 38612 19182
rect 38332 17052 38388 17108
rect 38556 17442 38612 17444
rect 38556 17390 38558 17442
rect 38558 17390 38610 17442
rect 38610 17390 38612 17442
rect 38556 17388 38612 17390
rect 39452 23548 39508 23604
rect 39340 23212 39396 23268
rect 39004 21980 39060 22036
rect 39228 21420 39284 21476
rect 39004 20748 39060 20804
rect 39900 26236 39956 26292
rect 41468 28028 41524 28084
rect 40572 26962 40628 26964
rect 40572 26910 40574 26962
rect 40574 26910 40626 26962
rect 40626 26910 40628 26962
rect 40572 26908 40628 26910
rect 41020 26290 41076 26292
rect 41020 26238 41022 26290
rect 41022 26238 41074 26290
rect 41074 26238 41076 26290
rect 41020 26236 41076 26238
rect 40348 25676 40404 25732
rect 40348 25506 40404 25508
rect 40348 25454 40350 25506
rect 40350 25454 40402 25506
rect 40402 25454 40404 25506
rect 40348 25452 40404 25454
rect 40236 25340 40292 25396
rect 39788 23996 39844 24052
rect 40348 23660 40404 23716
rect 40460 23548 40516 23604
rect 40124 23212 40180 23268
rect 41020 23996 41076 24052
rect 40908 23154 40964 23156
rect 40908 23102 40910 23154
rect 40910 23102 40962 23154
rect 40962 23102 40964 23154
rect 40908 23100 40964 23102
rect 40348 22652 40404 22708
rect 40908 22652 40964 22708
rect 39788 22316 39844 22372
rect 40572 22428 40628 22484
rect 39788 21868 39844 21924
rect 40348 21868 40404 21924
rect 40124 20748 40180 20804
rect 40012 20690 40068 20692
rect 40012 20638 40014 20690
rect 40014 20638 40066 20690
rect 40066 20638 40068 20690
rect 40012 20636 40068 20638
rect 39676 20578 39732 20580
rect 39676 20526 39678 20578
rect 39678 20526 39730 20578
rect 39730 20526 39732 20578
rect 39676 20524 39732 20526
rect 39564 20412 39620 20468
rect 38780 20188 38836 20244
rect 39228 19292 39284 19348
rect 39340 19234 39396 19236
rect 39340 19182 39342 19234
rect 39342 19182 39394 19234
rect 39394 19182 39396 19234
rect 39340 19180 39396 19182
rect 39564 19068 39620 19124
rect 39116 19010 39172 19012
rect 39116 18958 39118 19010
rect 39118 18958 39170 19010
rect 39170 18958 39172 19010
rect 39116 18956 39172 18958
rect 39004 18284 39060 18340
rect 38780 17724 38836 17780
rect 39900 19180 39956 19236
rect 39676 18060 39732 18116
rect 39004 17666 39060 17668
rect 39004 17614 39006 17666
rect 39006 17614 39058 17666
rect 39058 17614 39060 17666
rect 39004 17612 39060 17614
rect 40460 20636 40516 20692
rect 40908 20636 40964 20692
rect 40572 20524 40628 20580
rect 40684 20412 40740 20468
rect 40572 19180 40628 19236
rect 40684 19964 40740 20020
rect 40460 19122 40516 19124
rect 40460 19070 40462 19122
rect 40462 19070 40514 19122
rect 40514 19070 40516 19122
rect 40460 19068 40516 19070
rect 40572 18844 40628 18900
rect 40236 18172 40292 18228
rect 39788 17666 39844 17668
rect 39788 17614 39790 17666
rect 39790 17614 39842 17666
rect 39842 17614 39844 17666
rect 39788 17612 39844 17614
rect 38780 17554 38836 17556
rect 38780 17502 38782 17554
rect 38782 17502 38834 17554
rect 38834 17502 38836 17554
rect 38780 17500 38836 17502
rect 38780 16994 38836 16996
rect 38780 16942 38782 16994
rect 38782 16942 38834 16994
rect 38834 16942 38836 16994
rect 38780 16940 38836 16942
rect 38332 16658 38388 16660
rect 38332 16606 38334 16658
rect 38334 16606 38386 16658
rect 38386 16606 38388 16658
rect 38332 16604 38388 16606
rect 38220 15932 38276 15988
rect 38556 16828 38612 16884
rect 38780 16210 38836 16212
rect 38780 16158 38782 16210
rect 38782 16158 38834 16210
rect 38834 16158 38836 16210
rect 38780 16156 38836 16158
rect 38444 15372 38500 15428
rect 38892 15202 38948 15204
rect 38892 15150 38894 15202
rect 38894 15150 38946 15202
rect 38946 15150 38948 15202
rect 38892 15148 38948 15150
rect 39004 15036 39060 15092
rect 39676 17554 39732 17556
rect 39676 17502 39678 17554
rect 39678 17502 39730 17554
rect 39730 17502 39732 17554
rect 39676 17500 39732 17502
rect 39564 17164 39620 17220
rect 39228 16882 39284 16884
rect 39228 16830 39230 16882
rect 39230 16830 39282 16882
rect 39282 16830 39284 16882
rect 39228 16828 39284 16830
rect 39564 16828 39620 16884
rect 39228 16604 39284 16660
rect 39452 15932 39508 15988
rect 39900 17164 39956 17220
rect 40348 17164 40404 17220
rect 40796 19628 40852 19684
rect 41692 26962 41748 26964
rect 41692 26910 41694 26962
rect 41694 26910 41746 26962
rect 41746 26910 41748 26962
rect 41692 26908 41748 26910
rect 41356 23996 41412 24052
rect 41244 23266 41300 23268
rect 41244 23214 41246 23266
rect 41246 23214 41298 23266
rect 41298 23214 41300 23266
rect 41244 23212 41300 23214
rect 41244 22764 41300 22820
rect 41356 22876 41412 22932
rect 41244 22258 41300 22260
rect 41244 22206 41246 22258
rect 41246 22206 41298 22258
rect 41298 22206 41300 22258
rect 41244 22204 41300 22206
rect 41244 21868 41300 21924
rect 41244 21644 41300 21700
rect 41132 20018 41188 20020
rect 41132 19966 41134 20018
rect 41134 19966 41186 20018
rect 41186 19966 41188 20018
rect 41132 19964 41188 19966
rect 41356 20130 41412 20132
rect 41356 20078 41358 20130
rect 41358 20078 41410 20130
rect 41410 20078 41412 20130
rect 41356 20076 41412 20078
rect 41244 19628 41300 19684
rect 41132 19180 41188 19236
rect 40796 18620 40852 18676
rect 40908 17500 40964 17556
rect 41020 18508 41076 18564
rect 41244 18844 41300 18900
rect 42252 40348 42308 40404
rect 42924 39340 42980 39396
rect 42700 38946 42756 38948
rect 42700 38894 42702 38946
rect 42702 38894 42754 38946
rect 42754 38894 42756 38946
rect 42700 38892 42756 38894
rect 42588 38834 42644 38836
rect 42588 38782 42590 38834
rect 42590 38782 42642 38834
rect 42642 38782 42644 38834
rect 42588 38780 42644 38782
rect 43260 41804 43316 41860
rect 43260 40348 43316 40404
rect 43708 38834 43764 38836
rect 43708 38782 43710 38834
rect 43710 38782 43762 38834
rect 43762 38782 43764 38834
rect 43708 38780 43764 38782
rect 42924 27132 42980 27188
rect 41916 26908 41972 26964
rect 43036 27074 43092 27076
rect 43036 27022 43038 27074
rect 43038 27022 43090 27074
rect 43090 27022 43092 27074
rect 43036 27020 43092 27022
rect 41804 26460 41860 26516
rect 41916 25676 41972 25732
rect 41804 25452 41860 25508
rect 41692 25340 41748 25396
rect 42588 26514 42644 26516
rect 42588 26462 42590 26514
rect 42590 26462 42642 26514
rect 42642 26462 42644 26514
rect 42588 26460 42644 26462
rect 43820 27186 43876 27188
rect 43820 27134 43822 27186
rect 43822 27134 43874 27186
rect 43874 27134 43876 27186
rect 43820 27132 43876 27134
rect 45052 36370 45108 36372
rect 45052 36318 45054 36370
rect 45054 36318 45106 36370
rect 45106 36318 45108 36370
rect 45052 36316 45108 36318
rect 44716 36204 44772 36260
rect 45164 35644 45220 35700
rect 45164 35084 45220 35140
rect 44380 34690 44436 34692
rect 44380 34638 44382 34690
rect 44382 34638 44434 34690
rect 44434 34638 44436 34690
rect 44380 34636 44436 34638
rect 45276 34802 45332 34804
rect 45276 34750 45278 34802
rect 45278 34750 45330 34802
rect 45330 34750 45332 34802
rect 45276 34748 45332 34750
rect 45164 34636 45220 34692
rect 45276 34076 45332 34132
rect 45164 33234 45220 33236
rect 45164 33182 45166 33234
rect 45166 33182 45218 33234
rect 45218 33182 45220 33234
rect 45164 33180 45220 33182
rect 47852 76636 47908 76692
rect 48188 76636 48244 76692
rect 47404 76354 47460 76356
rect 47404 76302 47406 76354
rect 47406 76302 47458 76354
rect 47458 76302 47460 76354
rect 47404 76300 47460 76302
rect 49196 76690 49252 76692
rect 49196 76638 49198 76690
rect 49198 76638 49250 76690
rect 49250 76638 49252 76690
rect 49196 76636 49252 76638
rect 48636 76300 48692 76356
rect 47628 75682 47684 75684
rect 47628 75630 47630 75682
rect 47630 75630 47682 75682
rect 47682 75630 47684 75682
rect 47628 75628 47684 75630
rect 45612 36370 45668 36372
rect 45612 36318 45614 36370
rect 45614 36318 45666 36370
rect 45666 36318 45668 36370
rect 45612 36316 45668 36318
rect 45724 35698 45780 35700
rect 45724 35646 45726 35698
rect 45726 35646 45778 35698
rect 45778 35646 45780 35698
rect 45724 35644 45780 35646
rect 46620 36204 46676 36260
rect 45948 35698 46004 35700
rect 45948 35646 45950 35698
rect 45950 35646 46002 35698
rect 46002 35646 46004 35698
rect 45948 35644 46004 35646
rect 45724 35084 45780 35140
rect 46060 35196 46116 35252
rect 46284 34972 46340 35028
rect 44828 31612 44884 31668
rect 45052 31666 45108 31668
rect 45052 31614 45054 31666
rect 45054 31614 45106 31666
rect 45106 31614 45108 31666
rect 45052 31612 45108 31614
rect 44268 31500 44324 31556
rect 44716 30994 44772 30996
rect 44716 30942 44718 30994
rect 44718 30942 44770 30994
rect 44770 30942 44772 30994
rect 44716 30940 44772 30942
rect 44940 30492 44996 30548
rect 45724 34300 45780 34356
rect 45836 34130 45892 34132
rect 45836 34078 45838 34130
rect 45838 34078 45890 34130
rect 45890 34078 45892 34130
rect 45836 34076 45892 34078
rect 45724 33234 45780 33236
rect 45724 33182 45726 33234
rect 45726 33182 45778 33234
rect 45778 33182 45780 33234
rect 45724 33180 45780 33182
rect 46060 33292 46116 33348
rect 46620 34748 46676 34804
rect 46508 34300 46564 34356
rect 46508 34130 46564 34132
rect 46508 34078 46510 34130
rect 46510 34078 46562 34130
rect 46562 34078 46564 34130
rect 46508 34076 46564 34078
rect 45500 31554 45556 31556
rect 45500 31502 45502 31554
rect 45502 31502 45554 31554
rect 45554 31502 45556 31554
rect 45500 31500 45556 31502
rect 44828 30098 44884 30100
rect 44828 30046 44830 30098
rect 44830 30046 44882 30098
rect 44882 30046 44884 30098
rect 44828 30044 44884 30046
rect 45164 30044 45220 30100
rect 45388 29986 45444 29988
rect 45388 29934 45390 29986
rect 45390 29934 45442 29986
rect 45442 29934 45444 29986
rect 45388 29932 45444 29934
rect 44828 29538 44884 29540
rect 44828 29486 44830 29538
rect 44830 29486 44882 29538
rect 44882 29486 44884 29538
rect 44828 29484 44884 29486
rect 44604 28588 44660 28644
rect 44828 27580 44884 27636
rect 45052 27634 45108 27636
rect 45052 27582 45054 27634
rect 45054 27582 45106 27634
rect 45106 27582 45108 27634
rect 45052 27580 45108 27582
rect 44940 26962 44996 26964
rect 44940 26910 44942 26962
rect 44942 26910 44994 26962
rect 44994 26910 44996 26962
rect 44940 26908 44996 26910
rect 44156 26684 44212 26740
rect 43708 26460 43764 26516
rect 42364 25452 42420 25508
rect 41692 23996 41748 24052
rect 42028 23884 42084 23940
rect 43708 25564 43764 25620
rect 43036 25340 43092 25396
rect 43372 25506 43428 25508
rect 43372 25454 43374 25506
rect 43374 25454 43426 25506
rect 43426 25454 43428 25506
rect 43372 25452 43428 25454
rect 43372 25116 43428 25172
rect 42700 23938 42756 23940
rect 42700 23886 42702 23938
rect 42702 23886 42754 23938
rect 42754 23886 42756 23938
rect 42700 23884 42756 23886
rect 41580 23324 41636 23380
rect 41692 23266 41748 23268
rect 41692 23214 41694 23266
rect 41694 23214 41746 23266
rect 41746 23214 41748 23266
rect 41692 23212 41748 23214
rect 41804 23100 41860 23156
rect 41692 22930 41748 22932
rect 41692 22878 41694 22930
rect 41694 22878 41746 22930
rect 41746 22878 41748 22930
rect 41692 22876 41748 22878
rect 41804 22204 41860 22260
rect 42028 23324 42084 23380
rect 42252 23042 42308 23044
rect 42252 22990 42254 23042
rect 42254 22990 42306 23042
rect 42306 22990 42308 23042
rect 42252 22988 42308 22990
rect 43372 23378 43428 23380
rect 43372 23326 43374 23378
rect 43374 23326 43426 23378
rect 43426 23326 43428 23378
rect 43372 23324 43428 23326
rect 42476 23100 42532 23156
rect 42812 23266 42868 23268
rect 42812 23214 42814 23266
rect 42814 23214 42866 23266
rect 42866 23214 42868 23266
rect 42812 23212 42868 23214
rect 42028 20748 42084 20804
rect 41916 20076 41972 20132
rect 42140 20412 42196 20468
rect 41580 19516 41636 19572
rect 41804 19404 41860 19460
rect 41692 19292 41748 19348
rect 41580 18956 41636 19012
rect 41580 17948 41636 18004
rect 41356 17388 41412 17444
rect 41468 16994 41524 16996
rect 41468 16942 41470 16994
rect 41470 16942 41522 16994
rect 41522 16942 41524 16994
rect 41468 16940 41524 16942
rect 40236 15820 40292 15876
rect 39228 15260 39284 15316
rect 39116 14700 39172 14756
rect 38556 14252 38612 14308
rect 38444 13916 38500 13972
rect 38220 13858 38276 13860
rect 38220 13806 38222 13858
rect 38222 13806 38274 13858
rect 38274 13806 38276 13858
rect 38220 13804 38276 13806
rect 38332 13580 38388 13636
rect 38220 13468 38276 13524
rect 38780 13858 38836 13860
rect 38780 13806 38782 13858
rect 38782 13806 38834 13858
rect 38834 13806 38836 13858
rect 38780 13804 38836 13806
rect 39116 14140 39172 14196
rect 39900 15314 39956 15316
rect 39900 15262 39902 15314
rect 39902 15262 39954 15314
rect 39954 15262 39956 15314
rect 39900 15260 39956 15262
rect 40124 14140 40180 14196
rect 41916 18450 41972 18452
rect 41916 18398 41918 18450
rect 41918 18398 41970 18450
rect 41970 18398 41972 18450
rect 41916 18396 41972 18398
rect 42028 17724 42084 17780
rect 41916 16882 41972 16884
rect 41916 16830 41918 16882
rect 41918 16830 41970 16882
rect 41970 16830 41972 16882
rect 41916 16828 41972 16830
rect 42140 16044 42196 16100
rect 42252 16828 42308 16884
rect 41804 15260 41860 15316
rect 41580 14812 41636 14868
rect 41244 14588 41300 14644
rect 41468 14140 41524 14196
rect 39676 13468 39732 13524
rect 39116 12908 39172 12964
rect 39564 12962 39620 12964
rect 39564 12910 39566 12962
rect 39566 12910 39618 12962
rect 39618 12910 39620 12962
rect 39564 12908 39620 12910
rect 38108 11340 38164 11396
rect 38220 11228 38276 11284
rect 37660 10892 37716 10948
rect 38332 10780 38388 10836
rect 39564 12124 39620 12180
rect 39452 11228 39508 11284
rect 39340 10834 39396 10836
rect 39340 10782 39342 10834
rect 39342 10782 39394 10834
rect 39394 10782 39396 10834
rect 39340 10780 39396 10782
rect 39676 11116 39732 11172
rect 38892 10610 38948 10612
rect 38892 10558 38894 10610
rect 38894 10558 38946 10610
rect 38946 10558 38948 10610
rect 38892 10556 38948 10558
rect 38780 9884 38836 9940
rect 37100 8764 37156 8820
rect 36204 6636 36260 6692
rect 36092 6578 36148 6580
rect 36092 6526 36094 6578
rect 36094 6526 36146 6578
rect 36146 6526 36148 6578
rect 36092 6524 36148 6526
rect 35868 6412 35924 6468
rect 36092 5852 36148 5908
rect 36316 5404 36372 5460
rect 36428 5292 36484 5348
rect 36540 4396 36596 4452
rect 36092 3612 36148 3668
rect 34524 1820 34580 1876
rect 37100 8146 37156 8148
rect 37100 8094 37102 8146
rect 37102 8094 37154 8146
rect 37154 8094 37156 8146
rect 37100 8092 37156 8094
rect 36988 7644 37044 7700
rect 36876 5404 36932 5460
rect 37436 7196 37492 7252
rect 37772 6972 37828 7028
rect 36876 3612 36932 3668
rect 35980 2044 36036 2100
rect 36540 2268 36596 2324
rect 37100 4060 37156 4116
rect 36988 2828 37044 2884
rect 37212 3500 37268 3556
rect 36876 2156 36932 2212
rect 37548 5404 37604 5460
rect 37660 5180 37716 5236
rect 39788 9826 39844 9828
rect 39788 9774 39790 9826
rect 39790 9774 39842 9826
rect 39842 9774 39844 9826
rect 39788 9772 39844 9774
rect 38668 9212 38724 9268
rect 38220 9154 38276 9156
rect 38220 9102 38222 9154
rect 38222 9102 38274 9154
rect 38274 9102 38276 9154
rect 38220 9100 38276 9102
rect 39676 9602 39732 9604
rect 39676 9550 39678 9602
rect 39678 9550 39730 9602
rect 39730 9550 39732 9602
rect 39676 9548 39732 9550
rect 38892 9212 38948 9268
rect 38780 9100 38836 9156
rect 38668 8988 38724 9044
rect 40796 13746 40852 13748
rect 40796 13694 40798 13746
rect 40798 13694 40850 13746
rect 40850 13694 40852 13746
rect 40796 13692 40852 13694
rect 40236 13580 40292 13636
rect 41356 13634 41412 13636
rect 41356 13582 41358 13634
rect 41358 13582 41410 13634
rect 41410 13582 41412 13634
rect 41356 13580 41412 13582
rect 40908 13356 40964 13412
rect 41804 13692 41860 13748
rect 41916 12908 41972 12964
rect 41244 12402 41300 12404
rect 41244 12350 41246 12402
rect 41246 12350 41298 12402
rect 41298 12350 41300 12402
rect 41244 12348 41300 12350
rect 40236 11676 40292 11732
rect 40236 10834 40292 10836
rect 40236 10782 40238 10834
rect 40238 10782 40290 10834
rect 40290 10782 40292 10834
rect 40236 10780 40292 10782
rect 41020 11564 41076 11620
rect 38556 6860 38612 6916
rect 38108 5068 38164 5124
rect 38220 6524 38276 6580
rect 38780 7586 38836 7588
rect 38780 7534 38782 7586
rect 38782 7534 38834 7586
rect 38834 7534 38836 7586
rect 38780 7532 38836 7534
rect 39564 8092 39620 8148
rect 39228 6860 39284 6916
rect 39340 6748 39396 6804
rect 38780 6076 38836 6132
rect 38668 5292 38724 5348
rect 39004 5628 39060 5684
rect 39004 5010 39060 5012
rect 39004 4958 39006 5010
rect 39006 4958 39058 5010
rect 39058 4958 39060 5010
rect 39004 4956 39060 4958
rect 37324 2940 37380 2996
rect 38556 4732 38612 4788
rect 39228 4508 39284 4564
rect 39116 4450 39172 4452
rect 39116 4398 39118 4450
rect 39118 4398 39170 4450
rect 39170 4398 39172 4450
rect 39116 4396 39172 4398
rect 39116 3778 39172 3780
rect 39116 3726 39118 3778
rect 39118 3726 39170 3778
rect 39170 3726 39172 3778
rect 39116 3724 39172 3726
rect 38668 3612 38724 3668
rect 39900 7644 39956 7700
rect 39900 6972 39956 7028
rect 40124 6802 40180 6804
rect 40124 6750 40126 6802
rect 40126 6750 40178 6802
rect 40178 6750 40180 6802
rect 40124 6748 40180 6750
rect 40124 6076 40180 6132
rect 40124 5180 40180 5236
rect 40012 4844 40068 4900
rect 40460 5794 40516 5796
rect 40460 5742 40462 5794
rect 40462 5742 40514 5794
rect 40514 5742 40516 5794
rect 40460 5740 40516 5742
rect 40348 4620 40404 4676
rect 40348 3612 40404 3668
rect 40236 3500 40292 3556
rect 41356 11282 41412 11284
rect 41356 11230 41358 11282
rect 41358 11230 41410 11282
rect 41410 11230 41412 11282
rect 41356 11228 41412 11230
rect 42140 11228 42196 11284
rect 42588 22204 42644 22260
rect 42476 21698 42532 21700
rect 42476 21646 42478 21698
rect 42478 21646 42530 21698
rect 42530 21646 42532 21698
rect 42476 21644 42532 21646
rect 42476 16828 42532 16884
rect 42700 22092 42756 22148
rect 43372 22652 43428 22708
rect 42812 21868 42868 21924
rect 43260 21474 43316 21476
rect 43260 21422 43262 21474
rect 43262 21422 43314 21474
rect 43314 21422 43316 21474
rect 43260 21420 43316 21422
rect 42924 21084 42980 21140
rect 42924 20802 42980 20804
rect 42924 20750 42926 20802
rect 42926 20750 42978 20802
rect 42978 20750 42980 20802
rect 42924 20748 42980 20750
rect 42812 19292 42868 19348
rect 42588 16156 42644 16212
rect 43036 18620 43092 18676
rect 44044 25618 44100 25620
rect 44044 25566 44046 25618
rect 44046 25566 44098 25618
rect 44098 25566 44100 25618
rect 44044 25564 44100 25566
rect 43596 25228 43652 25284
rect 44156 25452 44212 25508
rect 44044 24892 44100 24948
rect 43596 24220 43652 24276
rect 43708 23996 43764 24052
rect 43596 23324 43652 23380
rect 43596 23100 43652 23156
rect 44828 26684 44884 26740
rect 44604 26514 44660 26516
rect 44604 26462 44606 26514
rect 44606 26462 44658 26514
rect 44658 26462 44660 26514
rect 44604 26460 44660 26462
rect 44380 26348 44436 26404
rect 44940 26402 44996 26404
rect 44940 26350 44942 26402
rect 44942 26350 44994 26402
rect 44994 26350 44996 26402
rect 44940 26348 44996 26350
rect 45052 26290 45108 26292
rect 45052 26238 45054 26290
rect 45054 26238 45106 26290
rect 45106 26238 45108 26290
rect 45052 26236 45108 26238
rect 44828 25788 44884 25844
rect 45388 25676 45444 25732
rect 44940 25394 44996 25396
rect 44940 25342 44942 25394
rect 44942 25342 44994 25394
rect 44994 25342 44996 25394
rect 44940 25340 44996 25342
rect 44156 24220 44212 24276
rect 44044 23100 44100 23156
rect 44268 22876 44324 22932
rect 44156 22540 44212 22596
rect 43820 22092 43876 22148
rect 44268 22146 44324 22148
rect 44268 22094 44270 22146
rect 44270 22094 44322 22146
rect 44322 22094 44324 22146
rect 44268 22092 44324 22094
rect 44156 21868 44212 21924
rect 43596 20412 43652 20468
rect 43708 20860 43764 20916
rect 44492 21420 44548 21476
rect 45276 24892 45332 24948
rect 45724 31106 45780 31108
rect 45724 31054 45726 31106
rect 45726 31054 45778 31106
rect 45778 31054 45780 31106
rect 45724 31052 45780 31054
rect 45948 31612 46004 31668
rect 45948 30994 46004 30996
rect 45948 30942 45950 30994
rect 45950 30942 46002 30994
rect 46002 30942 46004 30994
rect 45948 30940 46004 30942
rect 46172 31778 46228 31780
rect 46172 31726 46174 31778
rect 46174 31726 46226 31778
rect 46226 31726 46228 31778
rect 46172 31724 46228 31726
rect 46396 31106 46452 31108
rect 46396 31054 46398 31106
rect 46398 31054 46450 31106
rect 46450 31054 46452 31106
rect 46396 31052 46452 31054
rect 46172 30994 46228 30996
rect 46172 30942 46174 30994
rect 46174 30942 46226 30994
rect 46226 30942 46228 30994
rect 46172 30940 46228 30942
rect 46172 30210 46228 30212
rect 46172 30158 46174 30210
rect 46174 30158 46226 30210
rect 46226 30158 46228 30210
rect 46172 30156 46228 30158
rect 46620 30268 46676 30324
rect 46060 30098 46116 30100
rect 46060 30046 46062 30098
rect 46062 30046 46114 30098
rect 46114 30046 46116 30098
rect 46060 30044 46116 30046
rect 46060 29820 46116 29876
rect 46956 34972 47012 35028
rect 46844 34914 46900 34916
rect 46844 34862 46846 34914
rect 46846 34862 46898 34914
rect 46898 34862 46900 34914
rect 46844 34860 46900 34862
rect 47068 34076 47124 34132
rect 47292 31106 47348 31108
rect 47292 31054 47294 31106
rect 47294 31054 47346 31106
rect 47346 31054 47348 31106
rect 47292 31052 47348 31054
rect 47068 30882 47124 30884
rect 47068 30830 47070 30882
rect 47070 30830 47122 30882
rect 47122 30830 47124 30882
rect 47068 30828 47124 30830
rect 46956 30492 47012 30548
rect 47292 30268 47348 30324
rect 46172 27580 46228 27636
rect 46396 27186 46452 27188
rect 46396 27134 46398 27186
rect 46398 27134 46450 27186
rect 46450 27134 46452 27186
rect 46396 27132 46452 27134
rect 46060 26684 46116 26740
rect 46060 26402 46116 26404
rect 46060 26350 46062 26402
rect 46062 26350 46114 26402
rect 46114 26350 46116 26402
rect 46060 26348 46116 26350
rect 46284 26290 46340 26292
rect 46284 26238 46286 26290
rect 46286 26238 46338 26290
rect 46338 26238 46340 26290
rect 46284 26236 46340 26238
rect 46508 26290 46564 26292
rect 46508 26238 46510 26290
rect 46510 26238 46562 26290
rect 46562 26238 46564 26290
rect 46508 26236 46564 26238
rect 45724 25676 45780 25732
rect 45724 25506 45780 25508
rect 45724 25454 45726 25506
rect 45726 25454 45778 25506
rect 45778 25454 45780 25506
rect 45724 25452 45780 25454
rect 45948 25004 46004 25060
rect 45612 24444 45668 24500
rect 44828 23826 44884 23828
rect 44828 23774 44830 23826
rect 44830 23774 44882 23826
rect 44882 23774 44884 23826
rect 44828 23772 44884 23774
rect 44940 23548 44996 23604
rect 44828 23436 44884 23492
rect 44828 22652 44884 22708
rect 44940 22258 44996 22260
rect 44940 22206 44942 22258
rect 44942 22206 44994 22258
rect 44994 22206 44996 22258
rect 44940 22204 44996 22206
rect 45388 23826 45444 23828
rect 45388 23774 45390 23826
rect 45390 23774 45442 23826
rect 45442 23774 45444 23826
rect 45388 23772 45444 23774
rect 45500 23714 45556 23716
rect 45500 23662 45502 23714
rect 45502 23662 45554 23714
rect 45554 23662 45556 23714
rect 45500 23660 45556 23662
rect 45276 22540 45332 22596
rect 45388 22764 45444 22820
rect 45276 21196 45332 21252
rect 44828 20802 44884 20804
rect 44828 20750 44830 20802
rect 44830 20750 44882 20802
rect 44882 20750 44884 20802
rect 44828 20748 44884 20750
rect 43484 20076 43540 20132
rect 43932 19740 43988 19796
rect 43372 19404 43428 19460
rect 43372 18508 43428 18564
rect 43148 17948 43204 18004
rect 43036 17442 43092 17444
rect 43036 17390 43038 17442
rect 43038 17390 43090 17442
rect 43090 17390 43092 17442
rect 43036 17388 43092 17390
rect 43036 17052 43092 17108
rect 43036 16828 43092 16884
rect 42924 16716 42980 16772
rect 42812 15874 42868 15876
rect 42812 15822 42814 15874
rect 42814 15822 42866 15874
rect 42866 15822 42868 15874
rect 42812 15820 42868 15822
rect 43372 18060 43428 18116
rect 43596 17612 43652 17668
rect 43484 16268 43540 16324
rect 42364 14364 42420 14420
rect 42476 14306 42532 14308
rect 42476 14254 42478 14306
rect 42478 14254 42530 14306
rect 42530 14254 42532 14306
rect 42476 14252 42532 14254
rect 43372 14642 43428 14644
rect 43372 14590 43374 14642
rect 43374 14590 43426 14642
rect 43426 14590 43428 14642
rect 43372 14588 43428 14590
rect 42700 14530 42756 14532
rect 42700 14478 42702 14530
rect 42702 14478 42754 14530
rect 42754 14478 42756 14530
rect 42700 14476 42756 14478
rect 43260 14418 43316 14420
rect 43260 14366 43262 14418
rect 43262 14366 43314 14418
rect 43314 14366 43316 14418
rect 43260 14364 43316 14366
rect 42924 14140 42980 14196
rect 43260 14140 43316 14196
rect 42588 12348 42644 12404
rect 42588 11004 42644 11060
rect 42140 10498 42196 10500
rect 42140 10446 42142 10498
rect 42142 10446 42194 10498
rect 42194 10446 42196 10498
rect 42140 10444 42196 10446
rect 42140 9714 42196 9716
rect 42140 9662 42142 9714
rect 42142 9662 42194 9714
rect 42194 9662 42196 9714
rect 42140 9660 42196 9662
rect 41132 9212 41188 9268
rect 41020 9100 41076 9156
rect 41356 9100 41412 9156
rect 41132 8428 41188 8484
rect 40908 6972 40964 7028
rect 41244 7980 41300 8036
rect 41244 7644 41300 7700
rect 41468 7644 41524 7700
rect 41580 7980 41636 8036
rect 41468 7362 41524 7364
rect 41468 7310 41470 7362
rect 41470 7310 41522 7362
rect 41522 7310 41524 7362
rect 41468 7308 41524 7310
rect 41580 7084 41636 7140
rect 41692 7532 41748 7588
rect 41132 5964 41188 6020
rect 40908 5852 40964 5908
rect 41020 5628 41076 5684
rect 40684 4844 40740 4900
rect 41020 4956 41076 5012
rect 40908 4562 40964 4564
rect 40908 4510 40910 4562
rect 40910 4510 40962 4562
rect 40962 4510 40964 4562
rect 40908 4508 40964 4510
rect 41132 4284 41188 4340
rect 41356 3612 41412 3668
rect 40460 3276 40516 3332
rect 40572 2492 40628 2548
rect 43036 13356 43092 13412
rect 43932 16716 43988 16772
rect 44156 17724 44212 17780
rect 43932 16492 43988 16548
rect 44044 15874 44100 15876
rect 44044 15822 44046 15874
rect 44046 15822 44098 15874
rect 44098 15822 44100 15874
rect 44044 15820 44100 15822
rect 43484 12908 43540 12964
rect 44268 16492 44324 16548
rect 44268 15148 44324 15204
rect 43372 10444 43428 10500
rect 43372 10108 43428 10164
rect 42924 9548 42980 9604
rect 43596 9884 43652 9940
rect 43596 9266 43652 9268
rect 43596 9214 43598 9266
rect 43598 9214 43650 9266
rect 43650 9214 43652 9266
rect 43596 9212 43652 9214
rect 43596 8764 43652 8820
rect 42924 8428 42980 8484
rect 42924 7980 42980 8036
rect 43036 7644 43092 7700
rect 41916 7308 41972 7364
rect 42252 7420 42308 7476
rect 43708 7420 43764 7476
rect 43820 13580 43876 13636
rect 43148 7084 43204 7140
rect 43036 6972 43092 7028
rect 42476 5906 42532 5908
rect 42476 5854 42478 5906
rect 42478 5854 42530 5906
rect 42530 5854 42532 5906
rect 42476 5852 42532 5854
rect 41916 5292 41972 5348
rect 41916 4338 41972 4340
rect 41916 4286 41918 4338
rect 41918 4286 41970 4338
rect 41970 4286 41972 4338
rect 41916 4284 41972 4286
rect 42476 5404 42532 5460
rect 42476 5122 42532 5124
rect 42476 5070 42478 5122
rect 42478 5070 42530 5122
rect 42530 5070 42532 5122
rect 42476 5068 42532 5070
rect 41804 3612 41860 3668
rect 41916 3836 41972 3892
rect 42700 5740 42756 5796
rect 42588 3724 42644 3780
rect 42700 4060 42756 4116
rect 42252 3388 42308 3444
rect 42476 3500 42532 3556
rect 42812 3724 42868 3780
rect 43260 4284 43316 4340
rect 43036 3388 43092 3444
rect 44492 20130 44548 20132
rect 44492 20078 44494 20130
rect 44494 20078 44546 20130
rect 44546 20078 44548 20130
rect 44492 20076 44548 20078
rect 44716 18396 44772 18452
rect 45276 18450 45332 18452
rect 45276 18398 45278 18450
rect 45278 18398 45330 18450
rect 45330 18398 45332 18450
rect 45276 18396 45332 18398
rect 45052 17836 45108 17892
rect 44940 17724 44996 17780
rect 44940 17500 44996 17556
rect 45276 17724 45332 17780
rect 45388 17612 45444 17668
rect 45052 16940 45108 16996
rect 45276 16994 45332 16996
rect 45276 16942 45278 16994
rect 45278 16942 45330 16994
rect 45330 16942 45332 16994
rect 45276 16940 45332 16942
rect 45612 23154 45668 23156
rect 45612 23102 45614 23154
rect 45614 23102 45666 23154
rect 45666 23102 45668 23154
rect 45612 23100 45668 23102
rect 45836 22988 45892 23044
rect 45836 21868 45892 21924
rect 45836 21586 45892 21588
rect 45836 21534 45838 21586
rect 45838 21534 45890 21586
rect 45890 21534 45892 21586
rect 45836 21532 45892 21534
rect 45724 20188 45780 20244
rect 44828 15820 44884 15876
rect 45500 16210 45556 16212
rect 45500 16158 45502 16210
rect 45502 16158 45554 16210
rect 45554 16158 45556 16210
rect 45500 16156 45556 16158
rect 45500 15708 45556 15764
rect 44828 15148 44884 15204
rect 45500 15314 45556 15316
rect 45500 15262 45502 15314
rect 45502 15262 45554 15314
rect 45554 15262 45556 15314
rect 45500 15260 45556 15262
rect 45388 14924 45444 14980
rect 45500 14476 45556 14532
rect 45388 13468 45444 13524
rect 44044 9660 44100 9716
rect 43932 9266 43988 9268
rect 43932 9214 43934 9266
rect 43934 9214 43986 9266
rect 43986 9214 43988 9266
rect 43932 9212 43988 9214
rect 45052 11004 45108 11060
rect 44380 9548 44436 9604
rect 44156 9266 44212 9268
rect 44156 9214 44158 9266
rect 44158 9214 44210 9266
rect 44210 9214 44212 9266
rect 44156 9212 44212 9214
rect 44380 8204 44436 8260
rect 44156 8034 44212 8036
rect 44156 7982 44158 8034
rect 44158 7982 44210 8034
rect 44210 7982 44212 8034
rect 44156 7980 44212 7982
rect 43932 7474 43988 7476
rect 43932 7422 43934 7474
rect 43934 7422 43986 7474
rect 43986 7422 43988 7474
rect 43932 7420 43988 7422
rect 44268 7532 44324 7588
rect 44940 9154 44996 9156
rect 44940 9102 44942 9154
rect 44942 9102 44994 9154
rect 44994 9102 44996 9154
rect 44940 9100 44996 9102
rect 44940 8818 44996 8820
rect 44940 8766 44942 8818
rect 44942 8766 44994 8818
rect 44994 8766 44996 8818
rect 44940 8764 44996 8766
rect 44828 7868 44884 7924
rect 44268 6748 44324 6804
rect 44380 6860 44436 6916
rect 44268 5852 44324 5908
rect 44268 5068 44324 5124
rect 43596 4284 43652 4340
rect 43708 4172 43764 4228
rect 44268 3724 44324 3780
rect 43932 3612 43988 3668
rect 45612 11004 45668 11060
rect 45612 10108 45668 10164
rect 45276 9212 45332 9268
rect 46060 23660 46116 23716
rect 46284 25116 46340 25172
rect 46732 26402 46788 26404
rect 46732 26350 46734 26402
rect 46734 26350 46786 26402
rect 46786 26350 46788 26402
rect 46732 26348 46788 26350
rect 47068 26908 47124 26964
rect 46844 26684 46900 26740
rect 46956 26572 47012 26628
rect 47292 27074 47348 27076
rect 47292 27022 47294 27074
rect 47294 27022 47346 27074
rect 47346 27022 47348 27074
rect 47292 27020 47348 27022
rect 46956 25676 47012 25732
rect 46508 24892 46564 24948
rect 46956 25116 47012 25172
rect 47516 26514 47572 26516
rect 47516 26462 47518 26514
rect 47518 26462 47570 26514
rect 47570 26462 47572 26514
rect 47516 26460 47572 26462
rect 47628 26402 47684 26404
rect 47628 26350 47630 26402
rect 47630 26350 47682 26402
rect 47682 26350 47684 26402
rect 47628 26348 47684 26350
rect 47740 26684 47796 26740
rect 47516 25788 47572 25844
rect 47964 25676 48020 25732
rect 47292 25116 47348 25172
rect 48188 24946 48244 24948
rect 48188 24894 48190 24946
rect 48190 24894 48242 24946
rect 48242 24894 48244 24946
rect 48188 24892 48244 24894
rect 49980 76188 50036 76244
rect 50556 76858 50612 76860
rect 50556 76806 50558 76858
rect 50558 76806 50610 76858
rect 50610 76806 50612 76858
rect 50556 76804 50612 76806
rect 50660 76858 50716 76860
rect 50660 76806 50662 76858
rect 50662 76806 50714 76858
rect 50714 76806 50716 76858
rect 50660 76804 50716 76806
rect 50764 76858 50820 76860
rect 50764 76806 50766 76858
rect 50766 76806 50818 76858
rect 50818 76806 50820 76858
rect 50764 76804 50820 76806
rect 50204 76636 50260 76692
rect 51212 76690 51268 76692
rect 51212 76638 51214 76690
rect 51214 76638 51266 76690
rect 51266 76638 51268 76690
rect 51212 76636 51268 76638
rect 50540 76354 50596 76356
rect 50540 76302 50542 76354
rect 50542 76302 50594 76354
rect 50594 76302 50596 76354
rect 50540 76300 50596 76302
rect 50092 75740 50148 75796
rect 50764 75794 50820 75796
rect 50764 75742 50766 75794
rect 50766 75742 50818 75794
rect 50818 75742 50820 75794
rect 50764 75740 50820 75742
rect 50316 75682 50372 75684
rect 50316 75630 50318 75682
rect 50318 75630 50370 75682
rect 50370 75630 50372 75682
rect 50316 75628 50372 75630
rect 50556 75290 50612 75292
rect 50556 75238 50558 75290
rect 50558 75238 50610 75290
rect 50610 75238 50612 75290
rect 50556 75236 50612 75238
rect 50660 75290 50716 75292
rect 50660 75238 50662 75290
rect 50662 75238 50714 75290
rect 50714 75238 50716 75290
rect 50660 75236 50716 75238
rect 50764 75290 50820 75292
rect 50764 75238 50766 75290
rect 50766 75238 50818 75290
rect 50818 75238 50820 75290
rect 50764 75236 50820 75238
rect 50556 73722 50612 73724
rect 50556 73670 50558 73722
rect 50558 73670 50610 73722
rect 50610 73670 50612 73722
rect 50556 73668 50612 73670
rect 50660 73722 50716 73724
rect 50660 73670 50662 73722
rect 50662 73670 50714 73722
rect 50714 73670 50716 73722
rect 50660 73668 50716 73670
rect 50764 73722 50820 73724
rect 50764 73670 50766 73722
rect 50766 73670 50818 73722
rect 50818 73670 50820 73722
rect 50764 73668 50820 73670
rect 50556 72154 50612 72156
rect 50556 72102 50558 72154
rect 50558 72102 50610 72154
rect 50610 72102 50612 72154
rect 50556 72100 50612 72102
rect 50660 72154 50716 72156
rect 50660 72102 50662 72154
rect 50662 72102 50714 72154
rect 50714 72102 50716 72154
rect 50660 72100 50716 72102
rect 50764 72154 50820 72156
rect 50764 72102 50766 72154
rect 50766 72102 50818 72154
rect 50818 72102 50820 72154
rect 50764 72100 50820 72102
rect 50556 70586 50612 70588
rect 50556 70534 50558 70586
rect 50558 70534 50610 70586
rect 50610 70534 50612 70586
rect 50556 70532 50612 70534
rect 50660 70586 50716 70588
rect 50660 70534 50662 70586
rect 50662 70534 50714 70586
rect 50714 70534 50716 70586
rect 50660 70532 50716 70534
rect 50764 70586 50820 70588
rect 50764 70534 50766 70586
rect 50766 70534 50818 70586
rect 50818 70534 50820 70586
rect 50764 70532 50820 70534
rect 50556 69018 50612 69020
rect 50556 68966 50558 69018
rect 50558 68966 50610 69018
rect 50610 68966 50612 69018
rect 50556 68964 50612 68966
rect 50660 69018 50716 69020
rect 50660 68966 50662 69018
rect 50662 68966 50714 69018
rect 50714 68966 50716 69018
rect 50660 68964 50716 68966
rect 50764 69018 50820 69020
rect 50764 68966 50766 69018
rect 50766 68966 50818 69018
rect 50818 68966 50820 69018
rect 50764 68964 50820 68966
rect 50556 67450 50612 67452
rect 50556 67398 50558 67450
rect 50558 67398 50610 67450
rect 50610 67398 50612 67450
rect 50556 67396 50612 67398
rect 50660 67450 50716 67452
rect 50660 67398 50662 67450
rect 50662 67398 50714 67450
rect 50714 67398 50716 67450
rect 50660 67396 50716 67398
rect 50764 67450 50820 67452
rect 50764 67398 50766 67450
rect 50766 67398 50818 67450
rect 50818 67398 50820 67450
rect 50764 67396 50820 67398
rect 50556 65882 50612 65884
rect 50556 65830 50558 65882
rect 50558 65830 50610 65882
rect 50610 65830 50612 65882
rect 50556 65828 50612 65830
rect 50660 65882 50716 65884
rect 50660 65830 50662 65882
rect 50662 65830 50714 65882
rect 50714 65830 50716 65882
rect 50660 65828 50716 65830
rect 50764 65882 50820 65884
rect 50764 65830 50766 65882
rect 50766 65830 50818 65882
rect 50818 65830 50820 65882
rect 50764 65828 50820 65830
rect 50556 64314 50612 64316
rect 50556 64262 50558 64314
rect 50558 64262 50610 64314
rect 50610 64262 50612 64314
rect 50556 64260 50612 64262
rect 50660 64314 50716 64316
rect 50660 64262 50662 64314
rect 50662 64262 50714 64314
rect 50714 64262 50716 64314
rect 50660 64260 50716 64262
rect 50764 64314 50820 64316
rect 50764 64262 50766 64314
rect 50766 64262 50818 64314
rect 50818 64262 50820 64314
rect 50764 64260 50820 64262
rect 50556 62746 50612 62748
rect 50556 62694 50558 62746
rect 50558 62694 50610 62746
rect 50610 62694 50612 62746
rect 50556 62692 50612 62694
rect 50660 62746 50716 62748
rect 50660 62694 50662 62746
rect 50662 62694 50714 62746
rect 50714 62694 50716 62746
rect 50660 62692 50716 62694
rect 50764 62746 50820 62748
rect 50764 62694 50766 62746
rect 50766 62694 50818 62746
rect 50818 62694 50820 62746
rect 50764 62692 50820 62694
rect 50556 61178 50612 61180
rect 50556 61126 50558 61178
rect 50558 61126 50610 61178
rect 50610 61126 50612 61178
rect 50556 61124 50612 61126
rect 50660 61178 50716 61180
rect 50660 61126 50662 61178
rect 50662 61126 50714 61178
rect 50714 61126 50716 61178
rect 50660 61124 50716 61126
rect 50764 61178 50820 61180
rect 50764 61126 50766 61178
rect 50766 61126 50818 61178
rect 50818 61126 50820 61178
rect 50764 61124 50820 61126
rect 50556 59610 50612 59612
rect 50556 59558 50558 59610
rect 50558 59558 50610 59610
rect 50610 59558 50612 59610
rect 50556 59556 50612 59558
rect 50660 59610 50716 59612
rect 50660 59558 50662 59610
rect 50662 59558 50714 59610
rect 50714 59558 50716 59610
rect 50660 59556 50716 59558
rect 50764 59610 50820 59612
rect 50764 59558 50766 59610
rect 50766 59558 50818 59610
rect 50818 59558 50820 59610
rect 50764 59556 50820 59558
rect 50556 58042 50612 58044
rect 50556 57990 50558 58042
rect 50558 57990 50610 58042
rect 50610 57990 50612 58042
rect 50556 57988 50612 57990
rect 50660 58042 50716 58044
rect 50660 57990 50662 58042
rect 50662 57990 50714 58042
rect 50714 57990 50716 58042
rect 50660 57988 50716 57990
rect 50764 58042 50820 58044
rect 50764 57990 50766 58042
rect 50766 57990 50818 58042
rect 50818 57990 50820 58042
rect 50764 57988 50820 57990
rect 50556 56474 50612 56476
rect 50556 56422 50558 56474
rect 50558 56422 50610 56474
rect 50610 56422 50612 56474
rect 50556 56420 50612 56422
rect 50660 56474 50716 56476
rect 50660 56422 50662 56474
rect 50662 56422 50714 56474
rect 50714 56422 50716 56474
rect 50660 56420 50716 56422
rect 50764 56474 50820 56476
rect 50764 56422 50766 56474
rect 50766 56422 50818 56474
rect 50818 56422 50820 56474
rect 50764 56420 50820 56422
rect 50556 54906 50612 54908
rect 50556 54854 50558 54906
rect 50558 54854 50610 54906
rect 50610 54854 50612 54906
rect 50556 54852 50612 54854
rect 50660 54906 50716 54908
rect 50660 54854 50662 54906
rect 50662 54854 50714 54906
rect 50714 54854 50716 54906
rect 50660 54852 50716 54854
rect 50764 54906 50820 54908
rect 50764 54854 50766 54906
rect 50766 54854 50818 54906
rect 50818 54854 50820 54906
rect 50764 54852 50820 54854
rect 50556 53338 50612 53340
rect 50556 53286 50558 53338
rect 50558 53286 50610 53338
rect 50610 53286 50612 53338
rect 50556 53284 50612 53286
rect 50660 53338 50716 53340
rect 50660 53286 50662 53338
rect 50662 53286 50714 53338
rect 50714 53286 50716 53338
rect 50660 53284 50716 53286
rect 50764 53338 50820 53340
rect 50764 53286 50766 53338
rect 50766 53286 50818 53338
rect 50818 53286 50820 53338
rect 50764 53284 50820 53286
rect 50556 51770 50612 51772
rect 50556 51718 50558 51770
rect 50558 51718 50610 51770
rect 50610 51718 50612 51770
rect 50556 51716 50612 51718
rect 50660 51770 50716 51772
rect 50660 51718 50662 51770
rect 50662 51718 50714 51770
rect 50714 51718 50716 51770
rect 50660 51716 50716 51718
rect 50764 51770 50820 51772
rect 50764 51718 50766 51770
rect 50766 51718 50818 51770
rect 50818 51718 50820 51770
rect 50764 51716 50820 51718
rect 50556 50202 50612 50204
rect 50556 50150 50558 50202
rect 50558 50150 50610 50202
rect 50610 50150 50612 50202
rect 50556 50148 50612 50150
rect 50660 50202 50716 50204
rect 50660 50150 50662 50202
rect 50662 50150 50714 50202
rect 50714 50150 50716 50202
rect 50660 50148 50716 50150
rect 50764 50202 50820 50204
rect 50764 50150 50766 50202
rect 50766 50150 50818 50202
rect 50818 50150 50820 50202
rect 50764 50148 50820 50150
rect 50556 48634 50612 48636
rect 50556 48582 50558 48634
rect 50558 48582 50610 48634
rect 50610 48582 50612 48634
rect 50556 48580 50612 48582
rect 50660 48634 50716 48636
rect 50660 48582 50662 48634
rect 50662 48582 50714 48634
rect 50714 48582 50716 48634
rect 50660 48580 50716 48582
rect 50764 48634 50820 48636
rect 50764 48582 50766 48634
rect 50766 48582 50818 48634
rect 50818 48582 50820 48634
rect 50764 48580 50820 48582
rect 50556 47066 50612 47068
rect 50556 47014 50558 47066
rect 50558 47014 50610 47066
rect 50610 47014 50612 47066
rect 50556 47012 50612 47014
rect 50660 47066 50716 47068
rect 50660 47014 50662 47066
rect 50662 47014 50714 47066
rect 50714 47014 50716 47066
rect 50660 47012 50716 47014
rect 50764 47066 50820 47068
rect 50764 47014 50766 47066
rect 50766 47014 50818 47066
rect 50818 47014 50820 47066
rect 50764 47012 50820 47014
rect 50556 45498 50612 45500
rect 50556 45446 50558 45498
rect 50558 45446 50610 45498
rect 50610 45446 50612 45498
rect 50556 45444 50612 45446
rect 50660 45498 50716 45500
rect 50660 45446 50662 45498
rect 50662 45446 50714 45498
rect 50714 45446 50716 45498
rect 50660 45444 50716 45446
rect 50764 45498 50820 45500
rect 50764 45446 50766 45498
rect 50766 45446 50818 45498
rect 50818 45446 50820 45498
rect 50764 45444 50820 45446
rect 50556 43930 50612 43932
rect 50556 43878 50558 43930
rect 50558 43878 50610 43930
rect 50610 43878 50612 43930
rect 50556 43876 50612 43878
rect 50660 43930 50716 43932
rect 50660 43878 50662 43930
rect 50662 43878 50714 43930
rect 50714 43878 50716 43930
rect 50660 43876 50716 43878
rect 50764 43930 50820 43932
rect 50764 43878 50766 43930
rect 50766 43878 50818 43930
rect 50818 43878 50820 43930
rect 50764 43876 50820 43878
rect 50556 42362 50612 42364
rect 50556 42310 50558 42362
rect 50558 42310 50610 42362
rect 50610 42310 50612 42362
rect 50556 42308 50612 42310
rect 50660 42362 50716 42364
rect 50660 42310 50662 42362
rect 50662 42310 50714 42362
rect 50714 42310 50716 42362
rect 50660 42308 50716 42310
rect 50764 42362 50820 42364
rect 50764 42310 50766 42362
rect 50766 42310 50818 42362
rect 50818 42310 50820 42362
rect 50764 42308 50820 42310
rect 50556 40794 50612 40796
rect 50556 40742 50558 40794
rect 50558 40742 50610 40794
rect 50610 40742 50612 40794
rect 50556 40740 50612 40742
rect 50660 40794 50716 40796
rect 50660 40742 50662 40794
rect 50662 40742 50714 40794
rect 50714 40742 50716 40794
rect 50660 40740 50716 40742
rect 50764 40794 50820 40796
rect 50764 40742 50766 40794
rect 50766 40742 50818 40794
rect 50818 40742 50820 40794
rect 50764 40740 50820 40742
rect 50556 39226 50612 39228
rect 50556 39174 50558 39226
rect 50558 39174 50610 39226
rect 50610 39174 50612 39226
rect 50556 39172 50612 39174
rect 50660 39226 50716 39228
rect 50660 39174 50662 39226
rect 50662 39174 50714 39226
rect 50714 39174 50716 39226
rect 50660 39172 50716 39174
rect 50764 39226 50820 39228
rect 50764 39174 50766 39226
rect 50766 39174 50818 39226
rect 50818 39174 50820 39226
rect 50764 39172 50820 39174
rect 50316 38668 50372 38724
rect 52892 76636 52948 76692
rect 51996 40236 52052 40292
rect 51660 38668 51716 38724
rect 51884 40012 51940 40068
rect 51884 39004 51940 39060
rect 49532 29820 49588 29876
rect 49868 30268 49924 30324
rect 49308 28588 49364 28644
rect 49084 27074 49140 27076
rect 49084 27022 49086 27074
rect 49086 27022 49138 27074
rect 49138 27022 49140 27074
rect 49084 27020 49140 27022
rect 49644 27132 49700 27188
rect 49756 26962 49812 26964
rect 49756 26910 49758 26962
rect 49758 26910 49810 26962
rect 49810 26910 49812 26962
rect 49756 26908 49812 26910
rect 48860 26684 48916 26740
rect 48860 26402 48916 26404
rect 48860 26350 48862 26402
rect 48862 26350 48914 26402
rect 48914 26350 48916 26402
rect 48860 26348 48916 26350
rect 48748 26290 48804 26292
rect 48748 26238 48750 26290
rect 48750 26238 48802 26290
rect 48802 26238 48804 26290
rect 48748 26236 48804 26238
rect 48636 24892 48692 24948
rect 46396 23714 46452 23716
rect 46396 23662 46398 23714
rect 46398 23662 46450 23714
rect 46450 23662 46452 23714
rect 46396 23660 46452 23662
rect 46060 23100 46116 23156
rect 46060 22876 46116 22932
rect 46396 23100 46452 23156
rect 46284 22988 46340 23044
rect 46172 21532 46228 21588
rect 46060 18396 46116 18452
rect 45836 16268 45892 16324
rect 45724 9884 45780 9940
rect 45836 15708 45892 15764
rect 46620 22316 46676 22372
rect 47740 24668 47796 24724
rect 47068 23660 47124 23716
rect 47180 23378 47236 23380
rect 47180 23326 47182 23378
rect 47182 23326 47234 23378
rect 47234 23326 47236 23378
rect 47180 23324 47236 23326
rect 47068 22652 47124 22708
rect 46732 21980 46788 22036
rect 47516 23660 47572 23716
rect 47516 22652 47572 22708
rect 48860 24722 48916 24724
rect 48860 24670 48862 24722
rect 48862 24670 48914 24722
rect 48914 24670 48916 24722
rect 48860 24668 48916 24670
rect 48300 24220 48356 24276
rect 47852 23884 47908 23940
rect 48748 23826 48804 23828
rect 48748 23774 48750 23826
rect 48750 23774 48802 23826
rect 48802 23774 48804 23826
rect 48748 23772 48804 23774
rect 47852 23154 47908 23156
rect 47852 23102 47854 23154
rect 47854 23102 47906 23154
rect 47906 23102 47908 23154
rect 47852 23100 47908 23102
rect 48076 22988 48132 23044
rect 47404 22370 47460 22372
rect 47404 22318 47406 22370
rect 47406 22318 47458 22370
rect 47458 22318 47460 22370
rect 47404 22316 47460 22318
rect 47068 22258 47124 22260
rect 47068 22206 47070 22258
rect 47070 22206 47122 22258
rect 47122 22206 47124 22258
rect 47068 22204 47124 22206
rect 46956 21532 47012 21588
rect 46620 21474 46676 21476
rect 46620 21422 46622 21474
rect 46622 21422 46674 21474
rect 46674 21422 46676 21474
rect 46620 21420 46676 21422
rect 46508 21308 46564 21364
rect 46620 20802 46676 20804
rect 46620 20750 46622 20802
rect 46622 20750 46674 20802
rect 46674 20750 46676 20802
rect 46620 20748 46676 20750
rect 46172 17554 46228 17556
rect 46172 17502 46174 17554
rect 46174 17502 46226 17554
rect 46226 17502 46228 17554
rect 46172 17500 46228 17502
rect 46284 18396 46340 18452
rect 46620 20018 46676 20020
rect 46620 19966 46622 20018
rect 46622 19966 46674 20018
rect 46674 19966 46676 20018
rect 46620 19964 46676 19966
rect 46620 18844 46676 18900
rect 46620 18396 46676 18452
rect 46172 16098 46228 16100
rect 46172 16046 46174 16098
rect 46174 16046 46226 16098
rect 46226 16046 46228 16098
rect 46172 16044 46228 16046
rect 46396 16940 46452 16996
rect 46508 15484 46564 15540
rect 47068 21196 47124 21252
rect 47292 22146 47348 22148
rect 47292 22094 47294 22146
rect 47294 22094 47346 22146
rect 47346 22094 47348 22146
rect 47292 22092 47348 22094
rect 47404 21980 47460 22036
rect 47628 21980 47684 22036
rect 48076 22652 48132 22708
rect 47964 22092 48020 22148
rect 47180 20972 47236 21028
rect 47180 20802 47236 20804
rect 47180 20750 47182 20802
rect 47182 20750 47234 20802
rect 47234 20750 47236 20802
rect 47180 20748 47236 20750
rect 47740 20972 47796 21028
rect 47068 19852 47124 19908
rect 46844 18620 46900 18676
rect 46732 17724 46788 17780
rect 47404 18450 47460 18452
rect 47404 18398 47406 18450
rect 47406 18398 47458 18450
rect 47458 18398 47460 18450
rect 47404 18396 47460 18398
rect 47404 17948 47460 18004
rect 47292 16882 47348 16884
rect 47292 16830 47294 16882
rect 47294 16830 47346 16882
rect 47346 16830 47348 16882
rect 47292 16828 47348 16830
rect 47180 15708 47236 15764
rect 47180 15538 47236 15540
rect 47180 15486 47182 15538
rect 47182 15486 47234 15538
rect 47234 15486 47236 15538
rect 47180 15484 47236 15486
rect 47516 17500 47572 17556
rect 47404 15372 47460 15428
rect 48076 21532 48132 21588
rect 48300 21756 48356 21812
rect 48188 19906 48244 19908
rect 48188 19854 48190 19906
rect 48190 19854 48242 19906
rect 48242 19854 48244 19906
rect 48188 19852 48244 19854
rect 47740 15372 47796 15428
rect 47740 15148 47796 15204
rect 47964 15538 48020 15540
rect 47964 15486 47966 15538
rect 47966 15486 48018 15538
rect 48018 15486 48020 15538
rect 47964 15484 48020 15486
rect 48860 23154 48916 23156
rect 48860 23102 48862 23154
rect 48862 23102 48914 23154
rect 48914 23102 48916 23154
rect 48860 23100 48916 23102
rect 48748 21756 48804 21812
rect 48636 21644 48692 21700
rect 48412 20300 48468 20356
rect 48524 20748 48580 20804
rect 48748 20748 48804 20804
rect 48860 20018 48916 20020
rect 48860 19966 48862 20018
rect 48862 19966 48914 20018
rect 48914 19966 48916 20018
rect 48860 19964 48916 19966
rect 49196 26572 49252 26628
rect 49308 26460 49364 26516
rect 49532 26460 49588 26516
rect 49420 23548 49476 23604
rect 49420 22876 49476 22932
rect 49308 22764 49364 22820
rect 49084 22316 49140 22372
rect 49084 21868 49140 21924
rect 49084 21532 49140 21588
rect 49420 22092 49476 22148
rect 49644 23714 49700 23716
rect 49644 23662 49646 23714
rect 49646 23662 49698 23714
rect 49698 23662 49700 23714
rect 49644 23660 49700 23662
rect 50092 29148 50148 29204
rect 49868 23660 49924 23716
rect 50092 26348 50148 26404
rect 50556 37658 50612 37660
rect 50556 37606 50558 37658
rect 50558 37606 50610 37658
rect 50610 37606 50612 37658
rect 50556 37604 50612 37606
rect 50660 37658 50716 37660
rect 50660 37606 50662 37658
rect 50662 37606 50714 37658
rect 50714 37606 50716 37658
rect 50660 37604 50716 37606
rect 50764 37658 50820 37660
rect 50764 37606 50766 37658
rect 50766 37606 50818 37658
rect 50818 37606 50820 37658
rect 50764 37604 50820 37606
rect 50556 36090 50612 36092
rect 50556 36038 50558 36090
rect 50558 36038 50610 36090
rect 50610 36038 50612 36090
rect 50556 36036 50612 36038
rect 50660 36090 50716 36092
rect 50660 36038 50662 36090
rect 50662 36038 50714 36090
rect 50714 36038 50716 36090
rect 50660 36036 50716 36038
rect 50764 36090 50820 36092
rect 50764 36038 50766 36090
rect 50766 36038 50818 36090
rect 50818 36038 50820 36090
rect 50764 36036 50820 36038
rect 50556 34522 50612 34524
rect 50556 34470 50558 34522
rect 50558 34470 50610 34522
rect 50610 34470 50612 34522
rect 50556 34468 50612 34470
rect 50660 34522 50716 34524
rect 50660 34470 50662 34522
rect 50662 34470 50714 34522
rect 50714 34470 50716 34522
rect 50660 34468 50716 34470
rect 50764 34522 50820 34524
rect 50764 34470 50766 34522
rect 50766 34470 50818 34522
rect 50818 34470 50820 34522
rect 50764 34468 50820 34470
rect 50556 32954 50612 32956
rect 50556 32902 50558 32954
rect 50558 32902 50610 32954
rect 50610 32902 50612 32954
rect 50556 32900 50612 32902
rect 50660 32954 50716 32956
rect 50660 32902 50662 32954
rect 50662 32902 50714 32954
rect 50714 32902 50716 32954
rect 50660 32900 50716 32902
rect 50764 32954 50820 32956
rect 50764 32902 50766 32954
rect 50766 32902 50818 32954
rect 50818 32902 50820 32954
rect 50764 32900 50820 32902
rect 51324 31948 51380 32004
rect 51100 31778 51156 31780
rect 51100 31726 51102 31778
rect 51102 31726 51154 31778
rect 51154 31726 51156 31778
rect 51100 31724 51156 31726
rect 50556 31386 50612 31388
rect 50556 31334 50558 31386
rect 50558 31334 50610 31386
rect 50610 31334 50612 31386
rect 50556 31332 50612 31334
rect 50660 31386 50716 31388
rect 50660 31334 50662 31386
rect 50662 31334 50714 31386
rect 50714 31334 50716 31386
rect 50660 31332 50716 31334
rect 50764 31386 50820 31388
rect 50764 31334 50766 31386
rect 50766 31334 50818 31386
rect 50818 31334 50820 31386
rect 50764 31332 50820 31334
rect 50316 31106 50372 31108
rect 50316 31054 50318 31106
rect 50318 31054 50370 31106
rect 50370 31054 50372 31106
rect 50316 31052 50372 31054
rect 51100 30994 51156 30996
rect 51100 30942 51102 30994
rect 51102 30942 51154 30994
rect 51154 30942 51156 30994
rect 51100 30940 51156 30942
rect 50540 30828 50596 30884
rect 50652 30210 50708 30212
rect 50652 30158 50654 30210
rect 50654 30158 50706 30210
rect 50706 30158 50708 30210
rect 50652 30156 50708 30158
rect 50764 30098 50820 30100
rect 50764 30046 50766 30098
rect 50766 30046 50818 30098
rect 50818 30046 50820 30098
rect 50764 30044 50820 30046
rect 50556 29818 50612 29820
rect 50556 29766 50558 29818
rect 50558 29766 50610 29818
rect 50610 29766 50612 29818
rect 50556 29764 50612 29766
rect 50660 29818 50716 29820
rect 50660 29766 50662 29818
rect 50662 29766 50714 29818
rect 50714 29766 50716 29818
rect 50660 29764 50716 29766
rect 50764 29818 50820 29820
rect 50764 29766 50766 29818
rect 50766 29766 50818 29818
rect 50818 29766 50820 29818
rect 50764 29764 50820 29766
rect 50316 29372 50372 29428
rect 50316 28588 50372 28644
rect 50428 29260 50484 29316
rect 50556 28250 50612 28252
rect 50556 28198 50558 28250
rect 50558 28198 50610 28250
rect 50610 28198 50612 28250
rect 50556 28196 50612 28198
rect 50660 28250 50716 28252
rect 50660 28198 50662 28250
rect 50662 28198 50714 28250
rect 50714 28198 50716 28250
rect 50660 28196 50716 28198
rect 50764 28250 50820 28252
rect 50764 28198 50766 28250
rect 50766 28198 50818 28250
rect 50818 28198 50820 28250
rect 50764 28196 50820 28198
rect 51212 30770 51268 30772
rect 51212 30718 51214 30770
rect 51214 30718 51266 30770
rect 51266 30718 51268 30770
rect 51212 30716 51268 30718
rect 51436 31836 51492 31892
rect 51436 31164 51492 31220
rect 50876 27468 50932 27524
rect 50764 27186 50820 27188
rect 50764 27134 50766 27186
rect 50766 27134 50818 27186
rect 50818 27134 50820 27186
rect 50764 27132 50820 27134
rect 51212 27132 51268 27188
rect 51324 27468 51380 27524
rect 50556 26682 50612 26684
rect 50556 26630 50558 26682
rect 50558 26630 50610 26682
rect 50610 26630 50612 26682
rect 50556 26628 50612 26630
rect 50660 26682 50716 26684
rect 50660 26630 50662 26682
rect 50662 26630 50714 26682
rect 50714 26630 50716 26682
rect 50660 26628 50716 26630
rect 50764 26682 50820 26684
rect 50764 26630 50766 26682
rect 50766 26630 50818 26682
rect 50818 26630 50820 26682
rect 50764 26628 50820 26630
rect 51212 26684 51268 26740
rect 50428 26460 50484 26516
rect 50092 23436 50148 23492
rect 49868 23042 49924 23044
rect 49868 22990 49870 23042
rect 49870 22990 49922 23042
rect 49922 22990 49924 23042
rect 49868 22988 49924 22990
rect 49868 22540 49924 22596
rect 49868 21698 49924 21700
rect 49868 21646 49870 21698
rect 49870 21646 49922 21698
rect 49922 21646 49924 21698
rect 49868 21644 49924 21646
rect 49196 20748 49252 20804
rect 48300 15148 48356 15204
rect 46620 13634 46676 13636
rect 46620 13582 46622 13634
rect 46622 13582 46674 13634
rect 46674 13582 46676 13634
rect 46620 13580 46676 13582
rect 45836 9548 45892 9604
rect 46956 9772 47012 9828
rect 46060 9266 46116 9268
rect 46060 9214 46062 9266
rect 46062 9214 46114 9266
rect 46114 9214 46116 9266
rect 46060 9212 46116 9214
rect 45276 8204 45332 8260
rect 45948 7868 46004 7924
rect 45724 6972 45780 7028
rect 45276 6300 45332 6356
rect 44492 5906 44548 5908
rect 44492 5854 44494 5906
rect 44494 5854 44546 5906
rect 44546 5854 44548 5906
rect 44492 5852 44548 5854
rect 44828 5404 44884 5460
rect 44604 3724 44660 3780
rect 45612 6018 45668 6020
rect 45612 5966 45614 6018
rect 45614 5966 45666 6018
rect 45666 5966 45668 6018
rect 45612 5964 45668 5966
rect 45388 4844 45444 4900
rect 45500 4508 45556 4564
rect 45276 3554 45332 3556
rect 45276 3502 45278 3554
rect 45278 3502 45330 3554
rect 45330 3502 45332 3554
rect 45276 3500 45332 3502
rect 45164 3442 45220 3444
rect 45164 3390 45166 3442
rect 45166 3390 45218 3442
rect 45218 3390 45220 3442
rect 45164 3388 45220 3390
rect 46844 7474 46900 7476
rect 46844 7422 46846 7474
rect 46846 7422 46898 7474
rect 46898 7422 46900 7474
rect 46844 7420 46900 7422
rect 47404 7084 47460 7140
rect 46284 6300 46340 6356
rect 45948 5516 46004 5572
rect 46508 4956 46564 5012
rect 46396 4508 46452 4564
rect 46732 5964 46788 6020
rect 46956 5906 47012 5908
rect 46956 5854 46958 5906
rect 46958 5854 47010 5906
rect 47010 5854 47012 5906
rect 46956 5852 47012 5854
rect 46620 4450 46676 4452
rect 46620 4398 46622 4450
rect 46622 4398 46674 4450
rect 46674 4398 46676 4450
rect 46620 4396 46676 4398
rect 46732 5404 46788 5460
rect 46844 5122 46900 5124
rect 46844 5070 46846 5122
rect 46846 5070 46898 5122
rect 46898 5070 46900 5122
rect 46844 5068 46900 5070
rect 47740 6018 47796 6020
rect 47740 5966 47742 6018
rect 47742 5966 47794 6018
rect 47794 5966 47796 6018
rect 47740 5964 47796 5966
rect 47516 5180 47572 5236
rect 47404 4508 47460 4564
rect 47180 3388 47236 3444
rect 47628 4396 47684 4452
rect 47964 5516 48020 5572
rect 48412 9660 48468 9716
rect 48524 17388 48580 17444
rect 48748 15932 48804 15988
rect 48748 15426 48804 15428
rect 48748 15374 48750 15426
rect 48750 15374 48802 15426
rect 48802 15374 48804 15426
rect 48748 15372 48804 15374
rect 49420 20802 49476 20804
rect 49420 20750 49422 20802
rect 49422 20750 49474 20802
rect 49474 20750 49476 20802
rect 49420 20748 49476 20750
rect 49756 20802 49812 20804
rect 49756 20750 49758 20802
rect 49758 20750 49810 20802
rect 49810 20750 49812 20802
rect 49756 20748 49812 20750
rect 49420 20130 49476 20132
rect 49420 20078 49422 20130
rect 49422 20078 49474 20130
rect 49474 20078 49476 20130
rect 49420 20076 49476 20078
rect 49756 20300 49812 20356
rect 48972 15596 49028 15652
rect 48972 15372 49028 15428
rect 49420 15372 49476 15428
rect 50092 20748 50148 20804
rect 50092 20018 50148 20020
rect 50092 19966 50094 20018
rect 50094 19966 50146 20018
rect 50146 19966 50148 20018
rect 50092 19964 50148 19966
rect 50204 19852 50260 19908
rect 49084 15036 49140 15092
rect 48860 14028 48916 14084
rect 48748 12796 48804 12852
rect 48524 8204 48580 8260
rect 48412 7196 48468 7252
rect 49980 17724 50036 17780
rect 50556 25114 50612 25116
rect 50556 25062 50558 25114
rect 50558 25062 50610 25114
rect 50610 25062 50612 25114
rect 50556 25060 50612 25062
rect 50660 25114 50716 25116
rect 50660 25062 50662 25114
rect 50662 25062 50714 25114
rect 50714 25062 50716 25114
rect 50660 25060 50716 25062
rect 50764 25114 50820 25116
rect 50764 25062 50766 25114
rect 50766 25062 50818 25114
rect 50818 25062 50820 25114
rect 50764 25060 50820 25062
rect 50556 23546 50612 23548
rect 50556 23494 50558 23546
rect 50558 23494 50610 23546
rect 50610 23494 50612 23546
rect 50556 23492 50612 23494
rect 50660 23546 50716 23548
rect 50660 23494 50662 23546
rect 50662 23494 50714 23546
rect 50714 23494 50716 23546
rect 50660 23492 50716 23494
rect 50764 23546 50820 23548
rect 50764 23494 50766 23546
rect 50766 23494 50818 23546
rect 50818 23494 50820 23546
rect 50764 23492 50820 23494
rect 50428 22652 50484 22708
rect 50876 22146 50932 22148
rect 50876 22094 50878 22146
rect 50878 22094 50930 22146
rect 50930 22094 50932 22146
rect 50876 22092 50932 22094
rect 50556 21978 50612 21980
rect 50556 21926 50558 21978
rect 50558 21926 50610 21978
rect 50610 21926 50612 21978
rect 50556 21924 50612 21926
rect 50660 21978 50716 21980
rect 50660 21926 50662 21978
rect 50662 21926 50714 21978
rect 50714 21926 50716 21978
rect 50660 21924 50716 21926
rect 50764 21978 50820 21980
rect 50764 21926 50766 21978
rect 50766 21926 50818 21978
rect 50818 21926 50820 21978
rect 50764 21924 50820 21926
rect 50652 21644 50708 21700
rect 50556 20410 50612 20412
rect 50556 20358 50558 20410
rect 50558 20358 50610 20410
rect 50610 20358 50612 20410
rect 50556 20356 50612 20358
rect 50660 20410 50716 20412
rect 50660 20358 50662 20410
rect 50662 20358 50714 20410
rect 50714 20358 50716 20410
rect 50660 20356 50716 20358
rect 50764 20410 50820 20412
rect 50764 20358 50766 20410
rect 50766 20358 50818 20410
rect 50818 20358 50820 20410
rect 50764 20356 50820 20358
rect 51100 24892 51156 24948
rect 51212 20748 51268 20804
rect 51324 20914 51380 20916
rect 51324 20862 51326 20914
rect 51326 20862 51378 20914
rect 51378 20862 51380 20914
rect 51324 20860 51380 20862
rect 50876 20076 50932 20132
rect 50876 19852 50932 19908
rect 50556 18842 50612 18844
rect 50556 18790 50558 18842
rect 50558 18790 50610 18842
rect 50610 18790 50612 18842
rect 50556 18788 50612 18790
rect 50660 18842 50716 18844
rect 50660 18790 50662 18842
rect 50662 18790 50714 18842
rect 50714 18790 50716 18842
rect 50660 18788 50716 18790
rect 50764 18842 50820 18844
rect 50764 18790 50766 18842
rect 50766 18790 50818 18842
rect 50818 18790 50820 18842
rect 50764 18788 50820 18790
rect 50540 17500 50596 17556
rect 50988 17948 51044 18004
rect 50988 17500 51044 17556
rect 50764 17388 50820 17444
rect 49980 17276 50036 17332
rect 50556 17274 50612 17276
rect 50556 17222 50558 17274
rect 50558 17222 50610 17274
rect 50610 17222 50612 17274
rect 50556 17220 50612 17222
rect 50660 17274 50716 17276
rect 50660 17222 50662 17274
rect 50662 17222 50714 17274
rect 50714 17222 50716 17274
rect 50660 17220 50716 17222
rect 50764 17274 50820 17276
rect 50764 17222 50766 17274
rect 50766 17222 50818 17274
rect 50818 17222 50820 17274
rect 50764 17220 50820 17222
rect 50988 16940 51044 16996
rect 51324 19852 51380 19908
rect 51436 19628 51492 19684
rect 51772 30210 51828 30212
rect 51772 30158 51774 30210
rect 51774 30158 51826 30210
rect 51826 30158 51828 30210
rect 51772 30156 51828 30158
rect 51772 23436 51828 23492
rect 51660 21868 51716 21924
rect 51660 21532 51716 21588
rect 51772 20860 51828 20916
rect 51212 18508 51268 18564
rect 51660 20524 51716 20580
rect 51436 18060 51492 18116
rect 51772 19852 51828 19908
rect 51324 17724 51380 17780
rect 51660 19068 51716 19124
rect 50428 15874 50484 15876
rect 50428 15822 50430 15874
rect 50430 15822 50482 15874
rect 50482 15822 50484 15874
rect 50428 15820 50484 15822
rect 50556 15706 50612 15708
rect 50556 15654 50558 15706
rect 50558 15654 50610 15706
rect 50610 15654 50612 15706
rect 50556 15652 50612 15654
rect 50660 15706 50716 15708
rect 50660 15654 50662 15706
rect 50662 15654 50714 15706
rect 50714 15654 50716 15706
rect 50660 15652 50716 15654
rect 50764 15706 50820 15708
rect 50764 15654 50766 15706
rect 50766 15654 50818 15706
rect 50818 15654 50820 15706
rect 50764 15652 50820 15654
rect 50652 15426 50708 15428
rect 50652 15374 50654 15426
rect 50654 15374 50706 15426
rect 50706 15374 50708 15426
rect 50652 15372 50708 15374
rect 51436 16380 51492 16436
rect 51212 15372 51268 15428
rect 50428 14364 50484 14420
rect 51324 15820 51380 15876
rect 51660 15202 51716 15204
rect 51660 15150 51662 15202
rect 51662 15150 51714 15202
rect 51714 15150 51716 15202
rect 51660 15148 51716 15150
rect 51324 14530 51380 14532
rect 51324 14478 51326 14530
rect 51326 14478 51378 14530
rect 51378 14478 51380 14530
rect 51324 14476 51380 14478
rect 50876 14252 50932 14308
rect 50556 14138 50612 14140
rect 50556 14086 50558 14138
rect 50558 14086 50610 14138
rect 50610 14086 50612 14138
rect 50556 14084 50612 14086
rect 50660 14138 50716 14140
rect 50660 14086 50662 14138
rect 50662 14086 50714 14138
rect 50714 14086 50716 14138
rect 50660 14084 50716 14086
rect 50764 14138 50820 14140
rect 50764 14086 50766 14138
rect 50766 14086 50818 14138
rect 50818 14086 50820 14138
rect 50764 14084 50820 14086
rect 50556 12570 50612 12572
rect 50556 12518 50558 12570
rect 50558 12518 50610 12570
rect 50610 12518 50612 12570
rect 50556 12516 50612 12518
rect 50660 12570 50716 12572
rect 50660 12518 50662 12570
rect 50662 12518 50714 12570
rect 50714 12518 50716 12570
rect 50660 12516 50716 12518
rect 50764 12570 50820 12572
rect 50764 12518 50766 12570
rect 50766 12518 50818 12570
rect 50818 12518 50820 12570
rect 50764 12516 50820 12518
rect 50556 11002 50612 11004
rect 50556 10950 50558 11002
rect 50558 10950 50610 11002
rect 50610 10950 50612 11002
rect 50556 10948 50612 10950
rect 50660 11002 50716 11004
rect 50660 10950 50662 11002
rect 50662 10950 50714 11002
rect 50714 10950 50716 11002
rect 50660 10948 50716 10950
rect 50764 11002 50820 11004
rect 50764 10950 50766 11002
rect 50766 10950 50818 11002
rect 50818 10950 50820 11002
rect 50764 10948 50820 10950
rect 50556 9434 50612 9436
rect 50556 9382 50558 9434
rect 50558 9382 50610 9434
rect 50610 9382 50612 9434
rect 50556 9380 50612 9382
rect 50660 9434 50716 9436
rect 50660 9382 50662 9434
rect 50662 9382 50714 9434
rect 50714 9382 50716 9434
rect 50660 9380 50716 9382
rect 50764 9434 50820 9436
rect 50764 9382 50766 9434
rect 50766 9382 50818 9434
rect 50818 9382 50820 9434
rect 50764 9380 50820 9382
rect 49868 7644 49924 7700
rect 50204 8988 50260 9044
rect 49084 6636 49140 6692
rect 49532 7420 49588 7476
rect 48636 6578 48692 6580
rect 48636 6526 48638 6578
rect 48638 6526 48690 6578
rect 48690 6526 48692 6578
rect 48636 6524 48692 6526
rect 48188 5964 48244 6020
rect 48748 6076 48804 6132
rect 48972 5852 49028 5908
rect 48748 5628 48804 5684
rect 48300 5292 48356 5348
rect 47964 3836 48020 3892
rect 48076 5068 48132 5124
rect 48972 4284 49028 4340
rect 48524 3836 48580 3892
rect 49196 5740 49252 5796
rect 49196 5068 49252 5124
rect 49308 5404 49364 5460
rect 50556 7866 50612 7868
rect 50556 7814 50558 7866
rect 50558 7814 50610 7866
rect 50610 7814 50612 7866
rect 50556 7812 50612 7814
rect 50660 7866 50716 7868
rect 50660 7814 50662 7866
rect 50662 7814 50714 7866
rect 50714 7814 50716 7866
rect 50660 7812 50716 7814
rect 50764 7866 50820 7868
rect 50764 7814 50766 7866
rect 50766 7814 50818 7866
rect 50818 7814 50820 7866
rect 50764 7812 50820 7814
rect 49532 5068 49588 5124
rect 49644 6524 49700 6580
rect 49756 5794 49812 5796
rect 49756 5742 49758 5794
rect 49758 5742 49810 5794
rect 49810 5742 49812 5794
rect 49756 5740 49812 5742
rect 49868 5180 49924 5236
rect 49084 4060 49140 4116
rect 49308 4060 49364 4116
rect 49196 3276 49252 3332
rect 49196 2492 49252 2548
rect 49868 3836 49924 3892
rect 49868 3612 49924 3668
rect 50092 3500 50148 3556
rect 49644 3442 49700 3444
rect 49644 3390 49646 3442
rect 49646 3390 49698 3442
rect 49698 3390 49700 3442
rect 49644 3388 49700 3390
rect 51212 6524 51268 6580
rect 50764 6412 50820 6468
rect 50556 6298 50612 6300
rect 50556 6246 50558 6298
rect 50558 6246 50610 6298
rect 50610 6246 50612 6298
rect 50556 6244 50612 6246
rect 50660 6298 50716 6300
rect 50660 6246 50662 6298
rect 50662 6246 50714 6298
rect 50714 6246 50716 6298
rect 50660 6244 50716 6246
rect 50764 6298 50820 6300
rect 50764 6246 50766 6298
rect 50766 6246 50818 6298
rect 50818 6246 50820 6298
rect 50764 6244 50820 6246
rect 51212 6300 51268 6356
rect 50876 5516 50932 5572
rect 50428 5122 50484 5124
rect 50428 5070 50430 5122
rect 50430 5070 50482 5122
rect 50482 5070 50484 5122
rect 50428 5068 50484 5070
rect 50316 4956 50372 5012
rect 50556 4730 50612 4732
rect 50556 4678 50558 4730
rect 50558 4678 50610 4730
rect 50610 4678 50612 4730
rect 50556 4676 50612 4678
rect 50660 4730 50716 4732
rect 50660 4678 50662 4730
rect 50662 4678 50714 4730
rect 50714 4678 50716 4730
rect 50660 4676 50716 4678
rect 50764 4730 50820 4732
rect 50764 4678 50766 4730
rect 50766 4678 50818 4730
rect 50818 4678 50820 4730
rect 50764 4676 50820 4678
rect 50540 4114 50596 4116
rect 50540 4062 50542 4114
rect 50542 4062 50594 4114
rect 50594 4062 50596 4114
rect 50540 4060 50596 4062
rect 50540 3724 50596 3780
rect 50876 3388 50932 3444
rect 50204 3276 50260 3332
rect 50556 3162 50612 3164
rect 50556 3110 50558 3162
rect 50558 3110 50610 3162
rect 50610 3110 50612 3162
rect 50556 3108 50612 3110
rect 50660 3162 50716 3164
rect 50660 3110 50662 3162
rect 50662 3110 50714 3162
rect 50714 3110 50716 3162
rect 50660 3108 50716 3110
rect 50764 3162 50820 3164
rect 50764 3110 50766 3162
rect 50766 3110 50818 3162
rect 50818 3110 50820 3162
rect 50764 3108 50820 3110
rect 51996 38780 52052 38836
rect 52332 33404 52388 33460
rect 52332 32284 52388 32340
rect 52332 31052 52388 31108
rect 52220 22316 52276 22372
rect 52108 21308 52164 21364
rect 52108 17778 52164 17780
rect 52108 17726 52110 17778
rect 52110 17726 52162 17778
rect 52162 17726 52164 17778
rect 52108 17724 52164 17726
rect 52108 16940 52164 16996
rect 52780 36652 52836 36708
rect 52780 31890 52836 31892
rect 52780 31838 52782 31890
rect 52782 31838 52834 31890
rect 52834 31838 52836 31890
rect 52780 31836 52836 31838
rect 52892 34300 52948 34356
rect 53116 33458 53172 33460
rect 53116 33406 53118 33458
rect 53118 33406 53170 33458
rect 53170 33406 53172 33458
rect 53116 33404 53172 33406
rect 53004 33346 53060 33348
rect 53004 33294 53006 33346
rect 53006 33294 53058 33346
rect 53058 33294 53060 33346
rect 53004 33292 53060 33294
rect 52780 31218 52836 31220
rect 52780 31166 52782 31218
rect 52782 31166 52834 31218
rect 52834 31166 52836 31218
rect 52780 31164 52836 31166
rect 52780 22540 52836 22596
rect 52556 19964 52612 20020
rect 53900 76690 53956 76692
rect 53900 76638 53902 76690
rect 53902 76638 53954 76690
rect 53954 76638 53956 76690
rect 53900 76636 53956 76638
rect 55132 76690 55188 76692
rect 55132 76638 55134 76690
rect 55134 76638 55186 76690
rect 55186 76638 55188 76690
rect 55132 76636 55188 76638
rect 54908 76524 54964 76580
rect 55580 76524 55636 76580
rect 54460 71484 54516 71540
rect 53340 33404 53396 33460
rect 53228 22428 53284 22484
rect 53116 21586 53172 21588
rect 53116 21534 53118 21586
rect 53118 21534 53170 21586
rect 53170 21534 53172 21586
rect 53116 21532 53172 21534
rect 54236 40124 54292 40180
rect 54124 36092 54180 36148
rect 54012 35698 54068 35700
rect 54012 35646 54014 35698
rect 54014 35646 54066 35698
rect 54066 35646 54068 35698
rect 54012 35644 54068 35646
rect 53788 34972 53844 35028
rect 53900 34914 53956 34916
rect 53900 34862 53902 34914
rect 53902 34862 53954 34914
rect 53954 34862 53956 34914
rect 53900 34860 53956 34862
rect 54236 35810 54292 35812
rect 54236 35758 54238 35810
rect 54238 35758 54290 35810
rect 54290 35758 54292 35810
rect 54236 35756 54292 35758
rect 54124 33458 54180 33460
rect 54124 33406 54126 33458
rect 54126 33406 54178 33458
rect 54178 33406 54180 33458
rect 54124 33404 54180 33406
rect 53676 22316 53732 22372
rect 53788 21868 53844 21924
rect 53676 21474 53732 21476
rect 53676 21422 53678 21474
rect 53678 21422 53730 21474
rect 53730 21422 53732 21474
rect 53676 21420 53732 21422
rect 53340 20860 53396 20916
rect 53452 20748 53508 20804
rect 52780 19068 52836 19124
rect 52780 18732 52836 18788
rect 52556 18508 52612 18564
rect 52444 17948 52500 18004
rect 53004 18284 53060 18340
rect 52668 17388 52724 17444
rect 52556 15372 52612 15428
rect 52108 14754 52164 14756
rect 52108 14702 52110 14754
rect 52110 14702 52162 14754
rect 52162 14702 52164 14754
rect 52108 14700 52164 14702
rect 52892 14700 52948 14756
rect 52668 14530 52724 14532
rect 52668 14478 52670 14530
rect 52670 14478 52722 14530
rect 52722 14478 52724 14530
rect 52668 14476 52724 14478
rect 52220 13746 52276 13748
rect 52220 13694 52222 13746
rect 52222 13694 52274 13746
rect 52274 13694 52276 13746
rect 52220 13692 52276 13694
rect 51996 6524 52052 6580
rect 51884 6412 51940 6468
rect 51548 6076 51604 6132
rect 52108 6076 52164 6132
rect 51324 5234 51380 5236
rect 51324 5182 51326 5234
rect 51326 5182 51378 5234
rect 51378 5182 51380 5234
rect 51324 5180 51380 5182
rect 52444 5740 52500 5796
rect 52556 11564 52612 11620
rect 53564 20188 53620 20244
rect 53340 20018 53396 20020
rect 53340 19966 53342 20018
rect 53342 19966 53394 20018
rect 53394 19966 53396 20018
rect 53340 19964 53396 19966
rect 53228 19068 53284 19124
rect 53228 18732 53284 18788
rect 53116 17164 53172 17220
rect 54236 22482 54292 22484
rect 54236 22430 54238 22482
rect 54238 22430 54290 22482
rect 54290 22430 54292 22482
rect 54236 22428 54292 22430
rect 56924 76636 56980 76692
rect 57596 76412 57652 76468
rect 55916 75628 55972 75684
rect 55244 71484 55300 71540
rect 55804 45276 55860 45332
rect 55580 41858 55636 41860
rect 55580 41806 55582 41858
rect 55582 41806 55634 41858
rect 55634 41806 55636 41858
rect 55580 41804 55636 41806
rect 55468 41692 55524 41748
rect 55244 40572 55300 40628
rect 54908 40012 54964 40068
rect 55356 35868 55412 35924
rect 54908 35756 54964 35812
rect 55692 35586 55748 35588
rect 55692 35534 55694 35586
rect 55694 35534 55746 35586
rect 55746 35534 55748 35586
rect 55692 35532 55748 35534
rect 55020 35196 55076 35252
rect 55356 35026 55412 35028
rect 55356 34974 55358 35026
rect 55358 34974 55410 35026
rect 55410 34974 55412 35026
rect 55356 34972 55412 34974
rect 54684 31500 54740 31556
rect 54572 21756 54628 21812
rect 54348 21644 54404 21700
rect 54460 21420 54516 21476
rect 54124 20860 54180 20916
rect 55132 31500 55188 31556
rect 54460 20636 54516 20692
rect 54348 20242 54404 20244
rect 54348 20190 54350 20242
rect 54350 20190 54402 20242
rect 54402 20190 54404 20242
rect 54348 20188 54404 20190
rect 54908 20860 54964 20916
rect 54796 20076 54852 20132
rect 55020 19516 55076 19572
rect 54796 19068 54852 19124
rect 53676 18284 53732 18340
rect 53676 18060 53732 18116
rect 53340 17276 53396 17332
rect 53228 13804 53284 13860
rect 52892 9212 52948 9268
rect 53004 10892 53060 10948
rect 53340 10108 53396 10164
rect 53004 6300 53060 6356
rect 53452 7980 53508 8036
rect 53004 6076 53060 6132
rect 51436 3724 51492 3780
rect 51660 4844 51716 4900
rect 51212 3276 51268 3332
rect 51324 3612 51380 3668
rect 51772 3836 51828 3892
rect 51660 3554 51716 3556
rect 51660 3502 51662 3554
rect 51662 3502 51714 3554
rect 51714 3502 51716 3554
rect 51660 3500 51716 3502
rect 51996 3500 52052 3556
rect 52780 4844 52836 4900
rect 52668 4060 52724 4116
rect 52332 3388 52388 3444
rect 53004 3612 53060 3668
rect 53228 3500 53284 3556
rect 53340 3612 53396 3668
rect 53676 4620 53732 4676
rect 53900 13916 53956 13972
rect 57036 75628 57092 75684
rect 56140 41858 56196 41860
rect 56140 41806 56142 41858
rect 56142 41806 56194 41858
rect 56194 41806 56196 41858
rect 56140 41804 56196 41806
rect 57036 46956 57092 47012
rect 56700 43596 56756 43652
rect 58044 76748 58100 76804
rect 58156 75404 58212 75460
rect 55916 23436 55972 23492
rect 56028 21810 56084 21812
rect 56028 21758 56030 21810
rect 56030 21758 56082 21810
rect 56082 21758 56084 21810
rect 56028 21756 56084 21758
rect 55580 21698 55636 21700
rect 55580 21646 55582 21698
rect 55582 21646 55634 21698
rect 55634 21646 55636 21698
rect 55580 21644 55636 21646
rect 55580 20860 55636 20916
rect 56252 40796 56308 40852
rect 56812 41746 56868 41748
rect 56812 41694 56814 41746
rect 56814 41694 56866 41746
rect 56866 41694 56868 41746
rect 56812 41692 56868 41694
rect 57708 41746 57764 41748
rect 57708 41694 57710 41746
rect 57710 41694 57762 41746
rect 57762 41694 57764 41746
rect 57708 41692 57764 41694
rect 57484 41468 57540 41524
rect 56588 40796 56644 40852
rect 56252 40236 56308 40292
rect 56812 39228 56868 39284
rect 56812 35922 56868 35924
rect 56812 35870 56814 35922
rect 56814 35870 56866 35922
rect 56866 35870 56868 35922
rect 56812 35868 56868 35870
rect 56700 35532 56756 35588
rect 56140 20860 56196 20916
rect 55244 20690 55300 20692
rect 55244 20638 55246 20690
rect 55246 20638 55298 20690
rect 55298 20638 55300 20690
rect 55244 20636 55300 20638
rect 56252 20690 56308 20692
rect 56252 20638 56254 20690
rect 56254 20638 56306 20690
rect 56306 20638 56308 20690
rect 56252 20636 56308 20638
rect 55468 19068 55524 19124
rect 55132 18450 55188 18452
rect 55132 18398 55134 18450
rect 55134 18398 55186 18450
rect 55186 18398 55188 18450
rect 55132 18396 55188 18398
rect 54796 17276 54852 17332
rect 54460 14924 54516 14980
rect 54684 15260 54740 15316
rect 54572 14700 54628 14756
rect 54796 14588 54852 14644
rect 54236 13858 54292 13860
rect 54236 13806 54238 13858
rect 54238 13806 54290 13858
rect 54290 13806 54292 13858
rect 54236 13804 54292 13806
rect 54236 13132 54292 13188
rect 53900 7420 53956 7476
rect 53900 5180 53956 5236
rect 55132 13970 55188 13972
rect 55132 13918 55134 13970
rect 55134 13918 55186 13970
rect 55186 13918 55188 13970
rect 55132 13916 55188 13918
rect 56700 20130 56756 20132
rect 56700 20078 56702 20130
rect 56702 20078 56754 20130
rect 56754 20078 56756 20130
rect 56700 20076 56756 20078
rect 55804 20018 55860 20020
rect 55804 19966 55806 20018
rect 55806 19966 55858 20018
rect 55858 19966 55860 20018
rect 55804 19964 55860 19966
rect 56588 19516 56644 19572
rect 56140 19068 56196 19124
rect 55020 9324 55076 9380
rect 56028 11676 56084 11732
rect 55244 7532 55300 7588
rect 55356 11340 55412 11396
rect 55244 5234 55300 5236
rect 55244 5182 55246 5234
rect 55246 5182 55298 5234
rect 55298 5182 55300 5234
rect 55244 5180 55300 5182
rect 56028 11228 56084 11284
rect 56700 18338 56756 18340
rect 56700 18286 56702 18338
rect 56702 18286 56754 18338
rect 56754 18286 56756 18338
rect 56700 18284 56756 18286
rect 58828 76466 58884 76468
rect 58828 76414 58830 76466
rect 58830 76414 58882 76466
rect 58882 76414 58884 76466
rect 58828 76412 58884 76414
rect 59836 76690 59892 76692
rect 59836 76638 59838 76690
rect 59838 76638 59890 76690
rect 59890 76638 59892 76690
rect 59836 76636 59892 76638
rect 59612 76412 59668 76468
rect 58940 75292 58996 75348
rect 59388 75458 59444 75460
rect 59388 75406 59390 75458
rect 59390 75406 59442 75458
rect 59442 75406 59444 75458
rect 59388 75404 59444 75406
rect 60284 75516 60340 75572
rect 61628 76972 61684 77028
rect 62860 76972 62916 77028
rect 61964 76860 62020 76916
rect 58492 45276 58548 45332
rect 58604 53788 58660 53844
rect 58492 42866 58548 42868
rect 58492 42814 58494 42866
rect 58494 42814 58546 42866
rect 58546 42814 58548 42866
rect 58492 42812 58548 42814
rect 58380 41692 58436 41748
rect 58156 38892 58212 38948
rect 57484 23100 57540 23156
rect 57932 37100 57988 37156
rect 57148 20914 57204 20916
rect 57148 20862 57150 20914
rect 57150 20862 57202 20914
rect 57202 20862 57204 20914
rect 57148 20860 57204 20862
rect 57372 19122 57428 19124
rect 57372 19070 57374 19122
rect 57374 19070 57426 19122
rect 57426 19070 57428 19122
rect 57372 19068 57428 19070
rect 57148 18450 57204 18452
rect 57148 18398 57150 18450
rect 57150 18398 57202 18450
rect 57202 18398 57204 18450
rect 57148 18396 57204 18398
rect 57148 17612 57204 17668
rect 59500 43708 59556 43764
rect 61180 75570 61236 75572
rect 61180 75518 61182 75570
rect 61182 75518 61234 75570
rect 61234 75518 61236 75570
rect 61180 75516 61236 75518
rect 60508 75292 60564 75348
rect 61068 75404 61124 75460
rect 61292 75292 61348 75348
rect 61740 75682 61796 75684
rect 61740 75630 61742 75682
rect 61742 75630 61794 75682
rect 61794 75630 61796 75682
rect 61740 75628 61796 75630
rect 61516 75516 61572 75572
rect 60956 67228 61012 67284
rect 59948 42812 60004 42868
rect 59724 41244 59780 41300
rect 59836 40514 59892 40516
rect 59836 40462 59838 40514
rect 59838 40462 59890 40514
rect 59890 40462 59892 40514
rect 59836 40460 59892 40462
rect 58716 40348 58772 40404
rect 60060 40402 60116 40404
rect 60060 40350 60062 40402
rect 60062 40350 60114 40402
rect 60114 40350 60116 40402
rect 60060 40348 60116 40350
rect 61068 41074 61124 41076
rect 61068 41022 61070 41074
rect 61070 41022 61122 41074
rect 61122 41022 61124 41074
rect 61068 41020 61124 41022
rect 60956 40460 61012 40516
rect 60508 40348 60564 40404
rect 58604 31724 58660 31780
rect 58828 33180 58884 33236
rect 58828 30156 58884 30212
rect 58940 31612 58996 31668
rect 58940 29372 58996 29428
rect 59612 30940 59668 30996
rect 58716 17666 58772 17668
rect 58716 17614 58718 17666
rect 58718 17614 58770 17666
rect 58770 17614 58772 17666
rect 58716 17612 58772 17614
rect 58380 17442 58436 17444
rect 58380 17390 58382 17442
rect 58382 17390 58434 17442
rect 58434 17390 58436 17442
rect 58380 17388 58436 17390
rect 58828 17276 58884 17332
rect 57932 16940 57988 16996
rect 57148 14812 57204 14868
rect 57932 15148 57988 15204
rect 56140 11116 56196 11172
rect 57148 10108 57204 10164
rect 56028 5852 56084 5908
rect 56588 9884 56644 9940
rect 56140 5180 56196 5236
rect 53788 4172 53844 4228
rect 53900 4114 53956 4116
rect 53900 4062 53902 4114
rect 53902 4062 53954 4114
rect 53954 4062 53956 4114
rect 53900 4060 53956 4062
rect 53676 3554 53732 3556
rect 53676 3502 53678 3554
rect 53678 3502 53730 3554
rect 53730 3502 53732 3554
rect 53676 3500 53732 3502
rect 54684 4060 54740 4116
rect 54236 3724 54292 3780
rect 55356 3500 55412 3556
rect 56028 3666 56084 3668
rect 56028 3614 56030 3666
rect 56030 3614 56082 3666
rect 56082 3614 56084 3666
rect 56028 3612 56084 3614
rect 56812 6636 56868 6692
rect 56588 3612 56644 3668
rect 56700 5628 56756 5684
rect 56924 5906 56980 5908
rect 56924 5854 56926 5906
rect 56926 5854 56978 5906
rect 56978 5854 56980 5906
rect 56924 5852 56980 5854
rect 59612 9772 59668 9828
rect 59948 27356 60004 27412
rect 60732 40236 60788 40292
rect 60508 37660 60564 37716
rect 60508 34972 60564 35028
rect 60172 25676 60228 25732
rect 61068 40402 61124 40404
rect 61068 40350 61070 40402
rect 61070 40350 61122 40402
rect 61122 40350 61124 40402
rect 61068 40348 61124 40350
rect 61292 67228 61348 67284
rect 62076 76466 62132 76468
rect 62076 76414 62078 76466
rect 62078 76414 62130 76466
rect 62130 76414 62132 76466
rect 62076 76412 62132 76414
rect 62076 75404 62132 75460
rect 61852 58156 61908 58212
rect 61292 40460 61348 40516
rect 61516 41298 61572 41300
rect 61516 41246 61518 41298
rect 61518 41246 61570 41298
rect 61570 41246 61572 41298
rect 61516 41244 61572 41246
rect 61628 41020 61684 41076
rect 61180 39676 61236 39732
rect 62076 42700 62132 42756
rect 62188 46956 62244 47012
rect 62748 76412 62804 76468
rect 62972 76636 63028 76692
rect 63980 76690 64036 76692
rect 63980 76638 63982 76690
rect 63982 76638 64034 76690
rect 64034 76638 64036 76690
rect 63980 76636 64036 76638
rect 63756 75516 63812 75572
rect 62188 41580 62244 41636
rect 62188 41356 62244 41412
rect 62412 41186 62468 41188
rect 62412 41134 62414 41186
rect 62414 41134 62466 41186
rect 62466 41134 62468 41186
rect 62412 41132 62468 41134
rect 61740 29596 61796 29652
rect 62636 41804 62692 41860
rect 62636 41356 62692 41412
rect 62748 41132 62804 41188
rect 62188 40236 62244 40292
rect 62636 39730 62692 39732
rect 62636 39678 62638 39730
rect 62638 39678 62690 39730
rect 62690 39678 62692 39730
rect 62636 39676 62692 39678
rect 63308 41580 63364 41636
rect 62972 41186 63028 41188
rect 62972 41134 62974 41186
rect 62974 41134 63026 41186
rect 63026 41134 63028 41186
rect 62972 41132 63028 41134
rect 67004 76972 67060 77028
rect 67788 76972 67844 77028
rect 65324 75740 65380 75796
rect 65548 75458 65604 75460
rect 65548 75406 65550 75458
rect 65550 75406 65602 75458
rect 65602 75406 65604 75458
rect 65548 75404 65604 75406
rect 65324 73388 65380 73444
rect 63756 43260 63812 43316
rect 64876 67228 64932 67284
rect 63420 41916 63476 41972
rect 64540 41970 64596 41972
rect 64540 41918 64542 41970
rect 64542 41918 64594 41970
rect 64594 41918 64596 41970
rect 64540 41916 64596 41918
rect 64876 41916 64932 41972
rect 63644 41858 63700 41860
rect 63644 41806 63646 41858
rect 63646 41806 63698 41858
rect 63698 41806 63700 41858
rect 63644 41804 63700 41806
rect 64204 41132 64260 41188
rect 63196 40236 63252 40292
rect 63644 39394 63700 39396
rect 63644 39342 63646 39394
rect 63646 39342 63698 39394
rect 63698 39342 63700 39394
rect 63644 39340 63700 39342
rect 62972 38722 63028 38724
rect 62972 38670 62974 38722
rect 62974 38670 63026 38722
rect 63026 38670 63028 38722
rect 62972 38668 63028 38670
rect 63532 38668 63588 38724
rect 62860 36540 62916 36596
rect 62076 28476 62132 28532
rect 61404 28252 61460 28308
rect 61292 27244 61348 27300
rect 62860 28476 62916 28532
rect 63084 26236 63140 26292
rect 63196 34076 63252 34132
rect 63308 25618 63364 25620
rect 63308 25566 63310 25618
rect 63310 25566 63362 25618
rect 63362 25566 63364 25618
rect 63308 25564 63364 25566
rect 63196 25116 63252 25172
rect 61292 24444 61348 24500
rect 63308 24108 63364 24164
rect 60620 23660 60676 23716
rect 63420 23548 63476 23604
rect 64876 41186 64932 41188
rect 64876 41134 64878 41186
rect 64878 41134 64930 41186
rect 64930 41134 64932 41186
rect 64876 41132 64932 41134
rect 64428 40908 64484 40964
rect 65212 67228 65268 67284
rect 65916 76074 65972 76076
rect 65916 76022 65918 76074
rect 65918 76022 65970 76074
rect 65970 76022 65972 76074
rect 65916 76020 65972 76022
rect 66020 76074 66076 76076
rect 66020 76022 66022 76074
rect 66022 76022 66074 76074
rect 66074 76022 66076 76074
rect 66020 76020 66076 76022
rect 66124 76074 66180 76076
rect 66124 76022 66126 76074
rect 66126 76022 66178 76074
rect 66178 76022 66180 76074
rect 66124 76020 66180 76022
rect 65996 75794 66052 75796
rect 65996 75742 65998 75794
rect 65998 75742 66050 75794
rect 66050 75742 66052 75794
rect 65996 75740 66052 75742
rect 65916 74506 65972 74508
rect 65916 74454 65918 74506
rect 65918 74454 65970 74506
rect 65970 74454 65972 74506
rect 65916 74452 65972 74454
rect 66020 74506 66076 74508
rect 66020 74454 66022 74506
rect 66022 74454 66074 74506
rect 66074 74454 66076 74506
rect 66020 74452 66076 74454
rect 66124 74506 66180 74508
rect 66124 74454 66126 74506
rect 66126 74454 66178 74506
rect 66178 74454 66180 74506
rect 66124 74452 66180 74454
rect 65916 72938 65972 72940
rect 65916 72886 65918 72938
rect 65918 72886 65970 72938
rect 65970 72886 65972 72938
rect 65916 72884 65972 72886
rect 66020 72938 66076 72940
rect 66020 72886 66022 72938
rect 66022 72886 66074 72938
rect 66074 72886 66076 72938
rect 66020 72884 66076 72886
rect 66124 72938 66180 72940
rect 66124 72886 66126 72938
rect 66126 72886 66178 72938
rect 66178 72886 66180 72938
rect 66124 72884 66180 72886
rect 65916 71370 65972 71372
rect 65916 71318 65918 71370
rect 65918 71318 65970 71370
rect 65970 71318 65972 71370
rect 65916 71316 65972 71318
rect 66020 71370 66076 71372
rect 66020 71318 66022 71370
rect 66022 71318 66074 71370
rect 66074 71318 66076 71370
rect 66020 71316 66076 71318
rect 66124 71370 66180 71372
rect 66124 71318 66126 71370
rect 66126 71318 66178 71370
rect 66178 71318 66180 71370
rect 66124 71316 66180 71318
rect 65916 69802 65972 69804
rect 65916 69750 65918 69802
rect 65918 69750 65970 69802
rect 65970 69750 65972 69802
rect 65916 69748 65972 69750
rect 66020 69802 66076 69804
rect 66020 69750 66022 69802
rect 66022 69750 66074 69802
rect 66074 69750 66076 69802
rect 66020 69748 66076 69750
rect 66124 69802 66180 69804
rect 66124 69750 66126 69802
rect 66126 69750 66178 69802
rect 66178 69750 66180 69802
rect 66124 69748 66180 69750
rect 65916 68234 65972 68236
rect 65916 68182 65918 68234
rect 65918 68182 65970 68234
rect 65970 68182 65972 68234
rect 65916 68180 65972 68182
rect 66020 68234 66076 68236
rect 66020 68182 66022 68234
rect 66022 68182 66074 68234
rect 66074 68182 66076 68234
rect 66020 68180 66076 68182
rect 66124 68234 66180 68236
rect 66124 68182 66126 68234
rect 66126 68182 66178 68234
rect 66178 68182 66180 68234
rect 66124 68180 66180 68182
rect 65212 56140 65268 56196
rect 65324 41916 65380 41972
rect 65324 41020 65380 41076
rect 65100 40514 65156 40516
rect 65100 40462 65102 40514
rect 65102 40462 65154 40514
rect 65154 40462 65156 40514
rect 65100 40460 65156 40462
rect 64316 39394 64372 39396
rect 64316 39342 64318 39394
rect 64318 39342 64370 39394
rect 64370 39342 64372 39394
rect 64316 39340 64372 39342
rect 64316 38780 64372 38836
rect 63868 27916 63924 27972
rect 65212 38834 65268 38836
rect 65212 38782 65214 38834
rect 65214 38782 65266 38834
rect 65266 38782 65268 38834
rect 65212 38780 65268 38782
rect 64876 27804 64932 27860
rect 65916 66666 65972 66668
rect 65916 66614 65918 66666
rect 65918 66614 65970 66666
rect 65970 66614 65972 66666
rect 65916 66612 65972 66614
rect 66020 66666 66076 66668
rect 66020 66614 66022 66666
rect 66022 66614 66074 66666
rect 66074 66614 66076 66666
rect 66020 66612 66076 66614
rect 66124 66666 66180 66668
rect 66124 66614 66126 66666
rect 66126 66614 66178 66666
rect 66178 66614 66180 66666
rect 66124 66612 66180 66614
rect 65916 65098 65972 65100
rect 65916 65046 65918 65098
rect 65918 65046 65970 65098
rect 65970 65046 65972 65098
rect 65916 65044 65972 65046
rect 66020 65098 66076 65100
rect 66020 65046 66022 65098
rect 66022 65046 66074 65098
rect 66074 65046 66076 65098
rect 66020 65044 66076 65046
rect 66124 65098 66180 65100
rect 66124 65046 66126 65098
rect 66126 65046 66178 65098
rect 66178 65046 66180 65098
rect 66124 65044 66180 65046
rect 65916 63530 65972 63532
rect 65916 63478 65918 63530
rect 65918 63478 65970 63530
rect 65970 63478 65972 63530
rect 65916 63476 65972 63478
rect 66020 63530 66076 63532
rect 66020 63478 66022 63530
rect 66022 63478 66074 63530
rect 66074 63478 66076 63530
rect 66020 63476 66076 63478
rect 66124 63530 66180 63532
rect 66124 63478 66126 63530
rect 66126 63478 66178 63530
rect 66178 63478 66180 63530
rect 66124 63476 66180 63478
rect 66892 75404 66948 75460
rect 68348 76636 68404 76692
rect 65916 61962 65972 61964
rect 65916 61910 65918 61962
rect 65918 61910 65970 61962
rect 65970 61910 65972 61962
rect 65916 61908 65972 61910
rect 66020 61962 66076 61964
rect 66020 61910 66022 61962
rect 66022 61910 66074 61962
rect 66074 61910 66076 61962
rect 66020 61908 66076 61910
rect 66124 61962 66180 61964
rect 66124 61910 66126 61962
rect 66126 61910 66178 61962
rect 66178 61910 66180 61962
rect 66124 61908 66180 61910
rect 65916 60394 65972 60396
rect 65916 60342 65918 60394
rect 65918 60342 65970 60394
rect 65970 60342 65972 60394
rect 65916 60340 65972 60342
rect 66020 60394 66076 60396
rect 66020 60342 66022 60394
rect 66022 60342 66074 60394
rect 66074 60342 66076 60394
rect 66020 60340 66076 60342
rect 66124 60394 66180 60396
rect 66124 60342 66126 60394
rect 66126 60342 66178 60394
rect 66178 60342 66180 60394
rect 66124 60340 66180 60342
rect 65916 58826 65972 58828
rect 65916 58774 65918 58826
rect 65918 58774 65970 58826
rect 65970 58774 65972 58826
rect 65916 58772 65972 58774
rect 66020 58826 66076 58828
rect 66020 58774 66022 58826
rect 66022 58774 66074 58826
rect 66074 58774 66076 58826
rect 66020 58772 66076 58774
rect 66124 58826 66180 58828
rect 66124 58774 66126 58826
rect 66126 58774 66178 58826
rect 66178 58774 66180 58826
rect 66124 58772 66180 58774
rect 65916 57258 65972 57260
rect 65916 57206 65918 57258
rect 65918 57206 65970 57258
rect 65970 57206 65972 57258
rect 65916 57204 65972 57206
rect 66020 57258 66076 57260
rect 66020 57206 66022 57258
rect 66022 57206 66074 57258
rect 66074 57206 66076 57258
rect 66020 57204 66076 57206
rect 66124 57258 66180 57260
rect 66124 57206 66126 57258
rect 66126 57206 66178 57258
rect 66178 57206 66180 57258
rect 66124 57204 66180 57206
rect 65916 55690 65972 55692
rect 65916 55638 65918 55690
rect 65918 55638 65970 55690
rect 65970 55638 65972 55690
rect 65916 55636 65972 55638
rect 66020 55690 66076 55692
rect 66020 55638 66022 55690
rect 66022 55638 66074 55690
rect 66074 55638 66076 55690
rect 66020 55636 66076 55638
rect 66124 55690 66180 55692
rect 66124 55638 66126 55690
rect 66126 55638 66178 55690
rect 66178 55638 66180 55690
rect 66124 55636 66180 55638
rect 65916 54122 65972 54124
rect 65916 54070 65918 54122
rect 65918 54070 65970 54122
rect 65970 54070 65972 54122
rect 65916 54068 65972 54070
rect 66020 54122 66076 54124
rect 66020 54070 66022 54122
rect 66022 54070 66074 54122
rect 66074 54070 66076 54122
rect 66020 54068 66076 54070
rect 66124 54122 66180 54124
rect 66124 54070 66126 54122
rect 66126 54070 66178 54122
rect 66178 54070 66180 54122
rect 66124 54068 66180 54070
rect 65916 52554 65972 52556
rect 65916 52502 65918 52554
rect 65918 52502 65970 52554
rect 65970 52502 65972 52554
rect 65916 52500 65972 52502
rect 66020 52554 66076 52556
rect 66020 52502 66022 52554
rect 66022 52502 66074 52554
rect 66074 52502 66076 52554
rect 66020 52500 66076 52502
rect 66124 52554 66180 52556
rect 66124 52502 66126 52554
rect 66126 52502 66178 52554
rect 66178 52502 66180 52554
rect 66124 52500 66180 52502
rect 65916 50986 65972 50988
rect 65916 50934 65918 50986
rect 65918 50934 65970 50986
rect 65970 50934 65972 50986
rect 65916 50932 65972 50934
rect 66020 50986 66076 50988
rect 66020 50934 66022 50986
rect 66022 50934 66074 50986
rect 66074 50934 66076 50986
rect 66020 50932 66076 50934
rect 66124 50986 66180 50988
rect 66124 50934 66126 50986
rect 66126 50934 66178 50986
rect 66178 50934 66180 50986
rect 66124 50932 66180 50934
rect 65916 49418 65972 49420
rect 65916 49366 65918 49418
rect 65918 49366 65970 49418
rect 65970 49366 65972 49418
rect 65916 49364 65972 49366
rect 66020 49418 66076 49420
rect 66020 49366 66022 49418
rect 66022 49366 66074 49418
rect 66074 49366 66076 49418
rect 66020 49364 66076 49366
rect 66124 49418 66180 49420
rect 66124 49366 66126 49418
rect 66126 49366 66178 49418
rect 66178 49366 66180 49418
rect 66124 49364 66180 49366
rect 65916 47850 65972 47852
rect 65916 47798 65918 47850
rect 65918 47798 65970 47850
rect 65970 47798 65972 47850
rect 65916 47796 65972 47798
rect 66020 47850 66076 47852
rect 66020 47798 66022 47850
rect 66022 47798 66074 47850
rect 66074 47798 66076 47850
rect 66020 47796 66076 47798
rect 66124 47850 66180 47852
rect 66124 47798 66126 47850
rect 66126 47798 66178 47850
rect 66178 47798 66180 47850
rect 66124 47796 66180 47798
rect 65916 46282 65972 46284
rect 65916 46230 65918 46282
rect 65918 46230 65970 46282
rect 65970 46230 65972 46282
rect 65916 46228 65972 46230
rect 66020 46282 66076 46284
rect 66020 46230 66022 46282
rect 66022 46230 66074 46282
rect 66074 46230 66076 46282
rect 66020 46228 66076 46230
rect 66124 46282 66180 46284
rect 66124 46230 66126 46282
rect 66126 46230 66178 46282
rect 66178 46230 66180 46282
rect 66124 46228 66180 46230
rect 65916 44714 65972 44716
rect 65916 44662 65918 44714
rect 65918 44662 65970 44714
rect 65970 44662 65972 44714
rect 65916 44660 65972 44662
rect 66020 44714 66076 44716
rect 66020 44662 66022 44714
rect 66022 44662 66074 44714
rect 66074 44662 66076 44714
rect 66020 44660 66076 44662
rect 66124 44714 66180 44716
rect 66124 44662 66126 44714
rect 66126 44662 66178 44714
rect 66178 44662 66180 44714
rect 66124 44660 66180 44662
rect 65916 43146 65972 43148
rect 65916 43094 65918 43146
rect 65918 43094 65970 43146
rect 65970 43094 65972 43146
rect 65916 43092 65972 43094
rect 66020 43146 66076 43148
rect 66020 43094 66022 43146
rect 66022 43094 66074 43146
rect 66074 43094 66076 43146
rect 66020 43092 66076 43094
rect 66124 43146 66180 43148
rect 66124 43094 66126 43146
rect 66126 43094 66178 43146
rect 66178 43094 66180 43146
rect 66124 43092 66180 43094
rect 65916 41578 65972 41580
rect 65916 41526 65918 41578
rect 65918 41526 65970 41578
rect 65970 41526 65972 41578
rect 65916 41524 65972 41526
rect 66020 41578 66076 41580
rect 66020 41526 66022 41578
rect 66022 41526 66074 41578
rect 66074 41526 66076 41578
rect 66020 41524 66076 41526
rect 66124 41578 66180 41580
rect 66124 41526 66126 41578
rect 66126 41526 66178 41578
rect 66178 41526 66180 41578
rect 66124 41524 66180 41526
rect 65660 41186 65716 41188
rect 65660 41134 65662 41186
rect 65662 41134 65714 41186
rect 65714 41134 65716 41186
rect 65660 41132 65716 41134
rect 65772 41074 65828 41076
rect 65772 41022 65774 41074
rect 65774 41022 65826 41074
rect 65826 41022 65828 41074
rect 65772 41020 65828 41022
rect 66332 40572 66388 40628
rect 65660 39618 65716 39620
rect 65660 39566 65662 39618
rect 65662 39566 65714 39618
rect 65714 39566 65716 39618
rect 65660 39564 65716 39566
rect 65916 40010 65972 40012
rect 65916 39958 65918 40010
rect 65918 39958 65970 40010
rect 65970 39958 65972 40010
rect 65916 39956 65972 39958
rect 66020 40010 66076 40012
rect 66020 39958 66022 40010
rect 66022 39958 66074 40010
rect 66074 39958 66076 40010
rect 66020 39956 66076 39958
rect 66124 40010 66180 40012
rect 66124 39958 66126 40010
rect 66126 39958 66178 40010
rect 66178 39958 66180 40010
rect 66124 39956 66180 39958
rect 65436 35756 65492 35812
rect 66332 38780 66388 38836
rect 65324 27244 65380 27300
rect 63868 26124 63924 26180
rect 63756 24892 63812 24948
rect 63980 25116 64036 25172
rect 63532 23212 63588 23268
rect 61628 22092 61684 22148
rect 61292 21420 61348 21476
rect 57932 7756 57988 7812
rect 60172 19740 60228 19796
rect 57148 5852 57204 5908
rect 59500 8204 59556 8260
rect 60284 12908 60340 12964
rect 57932 5682 57988 5684
rect 57932 5630 57934 5682
rect 57934 5630 57986 5682
rect 57986 5630 57988 5682
rect 57932 5628 57988 5630
rect 59388 5628 59444 5684
rect 58156 5234 58212 5236
rect 58156 5182 58158 5234
rect 58158 5182 58210 5234
rect 58210 5182 58212 5234
rect 58156 5180 58212 5182
rect 58716 4844 58772 4900
rect 57596 4114 57652 4116
rect 57596 4062 57598 4114
rect 57598 4062 57650 4114
rect 57650 4062 57652 4114
rect 57596 4060 57652 4062
rect 58156 3724 58212 3780
rect 58044 3666 58100 3668
rect 58044 3614 58046 3666
rect 58046 3614 58098 3666
rect 58098 3614 58100 3666
rect 58044 3612 58100 3614
rect 57372 3388 57428 3444
rect 59052 3666 59108 3668
rect 59052 3614 59054 3666
rect 59054 3614 59106 3666
rect 59106 3614 59108 3666
rect 59052 3612 59108 3614
rect 61292 6636 61348 6692
rect 59948 5068 60004 5124
rect 60060 6412 60116 6468
rect 59500 3500 59556 3556
rect 59724 3388 59780 3444
rect 61516 6466 61572 6468
rect 61516 6414 61518 6466
rect 61518 6414 61570 6466
rect 61570 6414 61572 6466
rect 61516 6412 61572 6414
rect 60844 5682 60900 5684
rect 60844 5630 60846 5682
rect 60846 5630 60898 5682
rect 60898 5630 60900 5682
rect 60844 5628 60900 5630
rect 60732 5180 60788 5236
rect 60508 5122 60564 5124
rect 60508 5070 60510 5122
rect 60510 5070 60562 5122
rect 60562 5070 60564 5122
rect 60508 5068 60564 5070
rect 61516 4898 61572 4900
rect 61516 4846 61518 4898
rect 61518 4846 61570 4898
rect 61570 4846 61572 4898
rect 61516 4844 61572 4846
rect 65916 38442 65972 38444
rect 65916 38390 65918 38442
rect 65918 38390 65970 38442
rect 65970 38390 65972 38442
rect 65916 38388 65972 38390
rect 66020 38442 66076 38444
rect 66020 38390 66022 38442
rect 66022 38390 66074 38442
rect 66074 38390 66076 38442
rect 66020 38388 66076 38390
rect 66124 38442 66180 38444
rect 66124 38390 66126 38442
rect 66126 38390 66178 38442
rect 66178 38390 66180 38442
rect 66124 38388 66180 38390
rect 65916 36874 65972 36876
rect 65916 36822 65918 36874
rect 65918 36822 65970 36874
rect 65970 36822 65972 36874
rect 65916 36820 65972 36822
rect 66020 36874 66076 36876
rect 66020 36822 66022 36874
rect 66022 36822 66074 36874
rect 66074 36822 66076 36874
rect 66020 36820 66076 36822
rect 66124 36874 66180 36876
rect 66124 36822 66126 36874
rect 66126 36822 66178 36874
rect 66178 36822 66180 36874
rect 66124 36820 66180 36822
rect 65916 35306 65972 35308
rect 65916 35254 65918 35306
rect 65918 35254 65970 35306
rect 65970 35254 65972 35306
rect 65916 35252 65972 35254
rect 66020 35306 66076 35308
rect 66020 35254 66022 35306
rect 66022 35254 66074 35306
rect 66074 35254 66076 35306
rect 66020 35252 66076 35254
rect 66124 35306 66180 35308
rect 66124 35254 66126 35306
rect 66126 35254 66178 35306
rect 66178 35254 66180 35306
rect 66124 35252 66180 35254
rect 65916 33738 65972 33740
rect 65916 33686 65918 33738
rect 65918 33686 65970 33738
rect 65970 33686 65972 33738
rect 65916 33684 65972 33686
rect 66020 33738 66076 33740
rect 66020 33686 66022 33738
rect 66022 33686 66074 33738
rect 66074 33686 66076 33738
rect 66020 33684 66076 33686
rect 66124 33738 66180 33740
rect 66124 33686 66126 33738
rect 66126 33686 66178 33738
rect 66178 33686 66180 33738
rect 66124 33684 66180 33686
rect 65916 32170 65972 32172
rect 65916 32118 65918 32170
rect 65918 32118 65970 32170
rect 65970 32118 65972 32170
rect 65916 32116 65972 32118
rect 66020 32170 66076 32172
rect 66020 32118 66022 32170
rect 66022 32118 66074 32170
rect 66074 32118 66076 32170
rect 66020 32116 66076 32118
rect 66124 32170 66180 32172
rect 66124 32118 66126 32170
rect 66126 32118 66178 32170
rect 66178 32118 66180 32170
rect 66124 32116 66180 32118
rect 65916 30602 65972 30604
rect 65916 30550 65918 30602
rect 65918 30550 65970 30602
rect 65970 30550 65972 30602
rect 65916 30548 65972 30550
rect 66020 30602 66076 30604
rect 66020 30550 66022 30602
rect 66022 30550 66074 30602
rect 66074 30550 66076 30602
rect 66020 30548 66076 30550
rect 66124 30602 66180 30604
rect 66124 30550 66126 30602
rect 66126 30550 66178 30602
rect 66178 30550 66180 30602
rect 66124 30548 66180 30550
rect 65916 29034 65972 29036
rect 65916 28982 65918 29034
rect 65918 28982 65970 29034
rect 65970 28982 65972 29034
rect 65916 28980 65972 28982
rect 66020 29034 66076 29036
rect 66020 28982 66022 29034
rect 66022 28982 66074 29034
rect 66074 28982 66076 29034
rect 66020 28980 66076 28982
rect 66124 29034 66180 29036
rect 66124 28982 66126 29034
rect 66126 28982 66178 29034
rect 66178 28982 66180 29034
rect 66124 28980 66180 28982
rect 65916 27466 65972 27468
rect 65916 27414 65918 27466
rect 65918 27414 65970 27466
rect 65970 27414 65972 27466
rect 65916 27412 65972 27414
rect 66020 27466 66076 27468
rect 66020 27414 66022 27466
rect 66022 27414 66074 27466
rect 66074 27414 66076 27466
rect 66020 27412 66076 27414
rect 66124 27466 66180 27468
rect 66124 27414 66126 27466
rect 66126 27414 66178 27466
rect 66178 27414 66180 27466
rect 66124 27412 66180 27414
rect 65916 25898 65972 25900
rect 65916 25846 65918 25898
rect 65918 25846 65970 25898
rect 65970 25846 65972 25898
rect 65916 25844 65972 25846
rect 66020 25898 66076 25900
rect 66020 25846 66022 25898
rect 66022 25846 66074 25898
rect 66074 25846 66076 25898
rect 66020 25844 66076 25846
rect 66124 25898 66180 25900
rect 66124 25846 66126 25898
rect 66126 25846 66178 25898
rect 66178 25846 66180 25898
rect 66124 25844 66180 25846
rect 65916 24330 65972 24332
rect 65916 24278 65918 24330
rect 65918 24278 65970 24330
rect 65970 24278 65972 24330
rect 65916 24276 65972 24278
rect 66020 24330 66076 24332
rect 66020 24278 66022 24330
rect 66022 24278 66074 24330
rect 66074 24278 66076 24330
rect 66020 24276 66076 24278
rect 66124 24330 66180 24332
rect 66124 24278 66126 24330
rect 66126 24278 66178 24330
rect 66178 24278 66180 24330
rect 66124 24276 66180 24278
rect 65916 22762 65972 22764
rect 65916 22710 65918 22762
rect 65918 22710 65970 22762
rect 65970 22710 65972 22762
rect 65916 22708 65972 22710
rect 66020 22762 66076 22764
rect 66020 22710 66022 22762
rect 66022 22710 66074 22762
rect 66074 22710 66076 22762
rect 66020 22708 66076 22710
rect 66124 22762 66180 22764
rect 66124 22710 66126 22762
rect 66126 22710 66178 22762
rect 66178 22710 66180 22762
rect 66124 22708 66180 22710
rect 65660 21756 65716 21812
rect 66556 39676 66612 39732
rect 66780 39564 66836 39620
rect 67452 40626 67508 40628
rect 67452 40574 67454 40626
rect 67454 40574 67506 40626
rect 67506 40574 67508 40626
rect 67452 40572 67508 40574
rect 69692 76972 69748 77028
rect 69356 76690 69412 76692
rect 69356 76638 69358 76690
rect 69358 76638 69410 76690
rect 69410 76638 69412 76690
rect 69356 76636 69412 76638
rect 68684 75628 68740 75684
rect 68124 58828 68180 58884
rect 68572 71820 68628 71876
rect 67676 40572 67732 40628
rect 67116 39730 67172 39732
rect 67116 39678 67118 39730
rect 67118 39678 67170 39730
rect 67170 39678 67172 39730
rect 67116 39676 67172 39678
rect 66556 38050 66612 38052
rect 66556 37998 66558 38050
rect 66558 37998 66610 38050
rect 66610 37998 66612 38050
rect 66556 37996 66612 37998
rect 66444 21532 66500 21588
rect 63420 21196 63476 21252
rect 65916 21194 65972 21196
rect 63644 21084 63700 21140
rect 65916 21142 65918 21194
rect 65918 21142 65970 21194
rect 65970 21142 65972 21194
rect 65916 21140 65972 21142
rect 66020 21194 66076 21196
rect 66020 21142 66022 21194
rect 66022 21142 66074 21194
rect 66074 21142 66076 21194
rect 66020 21140 66076 21142
rect 66124 21194 66180 21196
rect 66124 21142 66126 21194
rect 66126 21142 66178 21194
rect 66178 21142 66180 21194
rect 66124 21140 66180 21142
rect 63420 6690 63476 6692
rect 63420 6638 63422 6690
rect 63422 6638 63474 6690
rect 63474 6638 63476 6690
rect 63420 6636 63476 6638
rect 62748 6412 62804 6468
rect 61628 4508 61684 4564
rect 62524 4562 62580 4564
rect 62524 4510 62526 4562
rect 62526 4510 62578 4562
rect 62578 4510 62580 4562
rect 62524 4508 62580 4510
rect 62076 3836 62132 3892
rect 61404 3724 61460 3780
rect 60956 3554 61012 3556
rect 60956 3502 60958 3554
rect 60958 3502 61010 3554
rect 61010 3502 61012 3554
rect 60956 3500 61012 3502
rect 61852 3554 61908 3556
rect 61852 3502 61854 3554
rect 61854 3502 61906 3554
rect 61906 3502 61908 3554
rect 61852 3500 61908 3502
rect 67004 39340 67060 39396
rect 67564 39394 67620 39396
rect 67564 39342 67566 39394
rect 67566 39342 67618 39394
rect 67618 39342 67620 39394
rect 67564 39340 67620 39342
rect 67900 40514 67956 40516
rect 67900 40462 67902 40514
rect 67902 40462 67954 40514
rect 67954 40462 67956 40514
rect 67900 40460 67956 40462
rect 67340 38668 67396 38724
rect 66892 22652 66948 22708
rect 67788 37436 67844 37492
rect 68684 42812 68740 42868
rect 68348 41020 68404 41076
rect 68124 38668 68180 38724
rect 68572 38834 68628 38836
rect 68572 38782 68574 38834
rect 68574 38782 68626 38834
rect 68626 38782 68628 38834
rect 68572 38780 68628 38782
rect 68348 38050 68404 38052
rect 68348 37998 68350 38050
rect 68350 37998 68402 38050
rect 68402 37998 68404 38050
rect 68348 37996 68404 37998
rect 68460 37490 68516 37492
rect 68460 37438 68462 37490
rect 68462 37438 68514 37490
rect 68514 37438 68516 37490
rect 68460 37436 68516 37438
rect 68124 37154 68180 37156
rect 68124 37102 68126 37154
rect 68126 37102 68178 37154
rect 68178 37102 68180 37154
rect 68124 37100 68180 37102
rect 68012 34972 68068 35028
rect 68684 37100 68740 37156
rect 68796 36594 68852 36596
rect 68796 36542 68798 36594
rect 68798 36542 68850 36594
rect 68850 36542 68852 36594
rect 68796 36540 68852 36542
rect 69916 58828 69972 58884
rect 69580 41356 69636 41412
rect 69580 40626 69636 40628
rect 69580 40574 69582 40626
rect 69582 40574 69634 40626
rect 69634 40574 69636 40626
rect 69580 40572 69636 40574
rect 69804 40572 69860 40628
rect 69468 39676 69524 39732
rect 69580 39618 69636 39620
rect 69580 39566 69582 39618
rect 69582 39566 69634 39618
rect 69634 39566 69636 39618
rect 69580 39564 69636 39566
rect 69020 38834 69076 38836
rect 69020 38782 69022 38834
rect 69022 38782 69074 38834
rect 69074 38782 69076 38834
rect 69020 38780 69076 38782
rect 69356 38668 69412 38724
rect 68908 32172 68964 32228
rect 69020 38556 69076 38612
rect 69244 38444 69300 38500
rect 69468 38332 69524 38388
rect 69132 36540 69188 36596
rect 69244 36428 69300 36484
rect 69132 30716 69188 30772
rect 70028 40572 70084 40628
rect 71708 77084 71764 77140
rect 70924 76972 70980 77028
rect 70364 76524 70420 76580
rect 70476 74060 70532 74116
rect 71596 76578 71652 76580
rect 71596 76526 71598 76578
rect 71598 76526 71650 76578
rect 71650 76526 71652 76578
rect 71596 76524 71652 76526
rect 70588 67228 70644 67284
rect 71148 67228 71204 67284
rect 70476 43484 70532 43540
rect 70588 41692 70644 41748
rect 70364 41132 70420 41188
rect 70252 40626 70308 40628
rect 70252 40574 70254 40626
rect 70254 40574 70306 40626
rect 70306 40574 70308 40626
rect 70252 40572 70308 40574
rect 71148 45276 71204 45332
rect 70812 41804 70868 41860
rect 70924 41244 70980 41300
rect 70812 40796 70868 40852
rect 70140 38444 70196 38500
rect 70252 39618 70308 39620
rect 70252 39566 70254 39618
rect 70254 39566 70306 39618
rect 70306 39566 70308 39618
rect 70252 39564 70308 39566
rect 70812 40348 70868 40404
rect 70700 39618 70756 39620
rect 70700 39566 70702 39618
rect 70702 39566 70754 39618
rect 70754 39566 70756 39618
rect 70700 39564 70756 39566
rect 70476 38780 70532 38836
rect 70700 38834 70756 38836
rect 70700 38782 70702 38834
rect 70702 38782 70754 38834
rect 70754 38782 70756 38834
rect 70700 38780 70756 38782
rect 70924 39506 70980 39508
rect 70924 39454 70926 39506
rect 70926 39454 70978 39506
rect 70978 39454 70980 39506
rect 70924 39452 70980 39454
rect 70924 38668 70980 38724
rect 70140 37548 70196 37604
rect 70028 37436 70084 37492
rect 69692 36482 69748 36484
rect 69692 36430 69694 36482
rect 69694 36430 69746 36482
rect 69746 36430 69748 36482
rect 69692 36428 69748 36430
rect 69580 29372 69636 29428
rect 68796 28252 68852 28308
rect 70588 38444 70644 38500
rect 70476 37548 70532 37604
rect 70588 37436 70644 37492
rect 73052 76972 73108 77028
rect 73164 77084 73220 77140
rect 72156 68684 72212 68740
rect 72044 51436 72100 51492
rect 71372 41692 71428 41748
rect 71484 41132 71540 41188
rect 71372 39730 71428 39732
rect 71372 39678 71374 39730
rect 71374 39678 71426 39730
rect 71426 39678 71428 39730
rect 71372 39676 71428 39678
rect 71932 46172 71988 46228
rect 73724 77084 73780 77140
rect 74284 76972 74340 77028
rect 74060 76578 74116 76580
rect 74060 76526 74062 76578
rect 74062 76526 74114 76578
rect 74114 76526 74116 76578
rect 74060 76524 74116 76526
rect 74508 77084 74564 77140
rect 75068 77084 75124 77140
rect 74620 76636 74676 76692
rect 72716 62076 72772 62132
rect 74060 75404 74116 75460
rect 74956 75122 75012 75124
rect 74956 75070 74958 75122
rect 74958 75070 75010 75122
rect 75010 75070 75012 75122
rect 74956 75068 75012 75070
rect 73948 68796 74004 68852
rect 73052 62076 73108 62132
rect 72156 42924 72212 42980
rect 72268 44604 72324 44660
rect 72044 41468 72100 41524
rect 71932 41298 71988 41300
rect 71932 41246 71934 41298
rect 71934 41246 71986 41298
rect 71986 41246 71988 41298
rect 71932 41244 71988 41246
rect 72156 41132 72212 41188
rect 71708 40348 71764 40404
rect 71596 39564 71652 39620
rect 71372 39452 71428 39508
rect 71372 38668 71428 38724
rect 72044 40908 72100 40964
rect 71260 38444 71316 38500
rect 71372 38050 71428 38052
rect 71372 37998 71374 38050
rect 71374 37998 71426 38050
rect 71426 37998 71428 38050
rect 71372 37996 71428 37998
rect 71596 39004 71652 39060
rect 72156 38780 72212 38836
rect 70812 37548 70868 37604
rect 71148 37490 71204 37492
rect 71148 37438 71150 37490
rect 71150 37438 71202 37490
rect 71202 37438 71204 37490
rect 71148 37436 71204 37438
rect 71260 36594 71316 36596
rect 71260 36542 71262 36594
rect 71262 36542 71314 36594
rect 71314 36542 71316 36594
rect 71260 36540 71316 36542
rect 71484 37490 71540 37492
rect 71484 37438 71486 37490
rect 71486 37438 71538 37490
rect 71538 37438 71540 37490
rect 71484 37436 71540 37438
rect 71372 35922 71428 35924
rect 71372 35870 71374 35922
rect 71374 35870 71426 35922
rect 71426 35870 71428 35922
rect 71372 35868 71428 35870
rect 71372 34860 71428 34916
rect 71148 34242 71204 34244
rect 71148 34190 71150 34242
rect 71150 34190 71202 34242
rect 71202 34190 71204 34242
rect 71148 34188 71204 34190
rect 71260 34076 71316 34132
rect 70924 34018 70980 34020
rect 70924 33966 70926 34018
rect 70926 33966 70978 34018
rect 70978 33966 70980 34018
rect 70924 33964 70980 33966
rect 71708 37548 71764 37604
rect 71708 37212 71764 37268
rect 71708 35586 71764 35588
rect 71708 35534 71710 35586
rect 71710 35534 71762 35586
rect 71762 35534 71764 35586
rect 71708 35532 71764 35534
rect 71820 34690 71876 34692
rect 71820 34638 71822 34690
rect 71822 34638 71874 34690
rect 71874 34638 71876 34690
rect 71820 34636 71876 34638
rect 71708 34130 71764 34132
rect 71708 34078 71710 34130
rect 71710 34078 71762 34130
rect 71762 34078 71764 34130
rect 71708 34076 71764 34078
rect 71596 33122 71652 33124
rect 71596 33070 71598 33122
rect 71598 33070 71650 33122
rect 71650 33070 71652 33122
rect 71596 33068 71652 33070
rect 71708 32956 71764 33012
rect 71820 32844 71876 32900
rect 71148 32396 71204 32452
rect 70924 31836 70980 31892
rect 70924 31106 70980 31108
rect 70924 31054 70926 31106
rect 70926 31054 70978 31106
rect 70978 31054 70980 31106
rect 70924 31052 70980 31054
rect 71708 31836 71764 31892
rect 71484 31500 71540 31556
rect 71372 30882 71428 30884
rect 71372 30830 71374 30882
rect 71374 30830 71426 30882
rect 71426 30830 71428 30882
rect 71372 30828 71428 30830
rect 72940 40178 72996 40180
rect 72940 40126 72942 40178
rect 72942 40126 72994 40178
rect 72994 40126 72996 40178
rect 72940 40124 72996 40126
rect 72940 39676 72996 39732
rect 72380 37772 72436 37828
rect 72268 37548 72324 37604
rect 72604 38444 72660 38500
rect 72156 36482 72212 36484
rect 72156 36430 72158 36482
rect 72158 36430 72210 36482
rect 72210 36430 72212 36482
rect 72156 36428 72212 36430
rect 72156 35644 72212 35700
rect 72268 35532 72324 35588
rect 72156 34188 72212 34244
rect 72492 36876 72548 36932
rect 73164 41074 73220 41076
rect 73164 41022 73166 41074
rect 73166 41022 73218 41074
rect 73218 41022 73220 41074
rect 73164 41020 73220 41022
rect 74844 72268 74900 72324
rect 74060 45164 74116 45220
rect 73724 40572 73780 40628
rect 73388 40290 73444 40292
rect 73388 40238 73390 40290
rect 73390 40238 73442 40290
rect 73442 40238 73444 40290
rect 73388 40236 73444 40238
rect 73276 39506 73332 39508
rect 73276 39454 73278 39506
rect 73278 39454 73330 39506
rect 73330 39454 73332 39506
rect 73276 39452 73332 39454
rect 73052 38050 73108 38052
rect 73052 37998 73054 38050
rect 73054 37998 73106 38050
rect 73106 37998 73108 38050
rect 73052 37996 73108 37998
rect 72828 37548 72884 37604
rect 72828 37378 72884 37380
rect 72828 37326 72830 37378
rect 72830 37326 72882 37378
rect 72882 37326 72884 37378
rect 72828 37324 72884 37326
rect 73276 37324 73332 37380
rect 73500 39564 73556 39620
rect 73836 39506 73892 39508
rect 73836 39454 73838 39506
rect 73838 39454 73890 39506
rect 73890 39454 73892 39506
rect 73836 39452 73892 39454
rect 73500 39004 73556 39060
rect 73500 38668 73556 38724
rect 73500 37826 73556 37828
rect 73500 37774 73502 37826
rect 73502 37774 73554 37826
rect 73554 37774 73556 37826
rect 73500 37772 73556 37774
rect 74172 41244 74228 41300
rect 74284 41186 74340 41188
rect 74284 41134 74286 41186
rect 74286 41134 74338 41186
rect 74338 41134 74340 41186
rect 74284 41132 74340 41134
rect 74284 39564 74340 39620
rect 74060 39340 74116 39396
rect 76076 76748 76132 76804
rect 75404 75516 75460 75572
rect 75628 75628 75684 75684
rect 75404 75010 75460 75012
rect 75404 74958 75406 75010
rect 75406 74958 75458 75010
rect 75458 74958 75460 75010
rect 75404 74956 75460 74958
rect 75292 74114 75348 74116
rect 75292 74062 75294 74114
rect 75294 74062 75346 74114
rect 75346 74062 75348 74114
rect 75292 74060 75348 74062
rect 76076 75516 76132 75572
rect 75964 75010 76020 75012
rect 75964 74958 75966 75010
rect 75966 74958 76018 75010
rect 76018 74958 76020 75010
rect 75964 74956 76020 74958
rect 76188 75068 76244 75124
rect 76300 76412 76356 76468
rect 76748 76354 76804 76356
rect 76748 76302 76750 76354
rect 76750 76302 76802 76354
rect 76802 76302 76804 76354
rect 76748 76300 76804 76302
rect 76524 75628 76580 75684
rect 76972 76748 77028 76804
rect 77308 79100 77364 79156
rect 77084 76412 77140 76468
rect 77196 76860 77252 76916
rect 77308 76690 77364 76692
rect 77308 76638 77310 76690
rect 77310 76638 77362 76690
rect 77362 76638 77364 76690
rect 77308 76636 77364 76638
rect 78764 77980 78820 78036
rect 77868 76466 77924 76468
rect 77868 76414 77870 76466
rect 77870 76414 77922 76466
rect 77922 76414 77924 76466
rect 77868 76412 77924 76414
rect 78204 76076 78260 76132
rect 75628 68796 75684 68852
rect 76748 72380 76804 72436
rect 75180 68684 75236 68740
rect 77532 75068 77588 75124
rect 77644 73554 77700 73556
rect 77644 73502 77646 73554
rect 77646 73502 77698 73554
rect 77698 73502 77700 73554
rect 77644 73500 77700 73502
rect 77644 72434 77700 72436
rect 77644 72382 77646 72434
rect 77646 72382 77698 72434
rect 77698 72382 77700 72434
rect 77644 72380 77700 72382
rect 76972 72268 77028 72324
rect 77644 71260 77700 71316
rect 77644 70978 77700 70980
rect 77644 70926 77646 70978
rect 77646 70926 77698 70978
rect 77698 70926 77700 70978
rect 77644 70924 77700 70926
rect 77420 70754 77476 70756
rect 77420 70702 77422 70754
rect 77422 70702 77474 70754
rect 77474 70702 77476 70754
rect 77420 70700 77476 70702
rect 77644 69020 77700 69076
rect 77420 68626 77476 68628
rect 77420 68574 77422 68626
rect 77422 68574 77474 68626
rect 77474 68574 77476 68626
rect 77420 68572 77476 68574
rect 77644 68514 77700 68516
rect 77644 68462 77646 68514
rect 77646 68462 77698 68514
rect 77698 68462 77700 68514
rect 77644 68460 77700 68462
rect 75404 43596 75460 43652
rect 75292 42924 75348 42980
rect 74732 41858 74788 41860
rect 74732 41806 74734 41858
rect 74734 41806 74786 41858
rect 74786 41806 74788 41858
rect 74732 41804 74788 41806
rect 76300 43484 76356 43540
rect 75740 42028 75796 42084
rect 74620 40626 74676 40628
rect 74620 40574 74622 40626
rect 74622 40574 74674 40626
rect 74674 40574 74676 40626
rect 74620 40572 74676 40574
rect 74508 39676 74564 39732
rect 74396 39340 74452 39396
rect 74172 39004 74228 39060
rect 74172 38668 74228 38724
rect 74508 38556 74564 38612
rect 74284 37996 74340 38052
rect 74172 37938 74228 37940
rect 74172 37886 74174 37938
rect 74174 37886 74226 37938
rect 74226 37886 74228 37938
rect 74172 37884 74228 37886
rect 74060 37772 74116 37828
rect 73948 37324 74004 37380
rect 73164 36876 73220 36932
rect 73164 36482 73220 36484
rect 73164 36430 73166 36482
rect 73166 36430 73218 36482
rect 73218 36430 73220 36482
rect 73164 36428 73220 36430
rect 73052 36258 73108 36260
rect 73052 36206 73054 36258
rect 73054 36206 73106 36258
rect 73106 36206 73108 36258
rect 73052 36204 73108 36206
rect 72156 32396 72212 32452
rect 72268 32060 72324 32116
rect 71260 29036 71316 29092
rect 70700 28082 70756 28084
rect 70700 28030 70702 28082
rect 70702 28030 70754 28082
rect 70754 28030 70756 28082
rect 70700 28028 70756 28030
rect 70700 27804 70756 27860
rect 68796 26012 68852 26068
rect 68684 23100 68740 23156
rect 67676 22428 67732 22484
rect 66668 20748 66724 20804
rect 67228 21644 67284 21700
rect 63756 20636 63812 20692
rect 65916 19626 65972 19628
rect 65916 19574 65918 19626
rect 65918 19574 65970 19626
rect 65970 19574 65972 19626
rect 65916 19572 65972 19574
rect 66020 19626 66076 19628
rect 66020 19574 66022 19626
rect 66022 19574 66074 19626
rect 66074 19574 66076 19626
rect 66020 19572 66076 19574
rect 66124 19626 66180 19628
rect 66124 19574 66126 19626
rect 66126 19574 66178 19626
rect 66178 19574 66180 19626
rect 66124 19572 66180 19574
rect 63756 17052 63812 17108
rect 64540 18620 64596 18676
rect 63868 9660 63924 9716
rect 64428 6466 64484 6468
rect 64428 6414 64430 6466
rect 64430 6414 64482 6466
rect 64482 6414 64484 6466
rect 64428 6412 64484 6414
rect 64428 5234 64484 5236
rect 64428 5182 64430 5234
rect 64430 5182 64482 5234
rect 64482 5182 64484 5234
rect 64428 5180 64484 5182
rect 63756 5068 63812 5124
rect 67788 20860 67844 20916
rect 68908 20188 68964 20244
rect 67788 18956 67844 19012
rect 67900 19852 67956 19908
rect 67228 18396 67284 18452
rect 65916 18058 65972 18060
rect 65916 18006 65918 18058
rect 65918 18006 65970 18058
rect 65970 18006 65972 18058
rect 65916 18004 65972 18006
rect 66020 18058 66076 18060
rect 66020 18006 66022 18058
rect 66022 18006 66074 18058
rect 66074 18006 66076 18058
rect 66020 18004 66076 18006
rect 66124 18058 66180 18060
rect 66124 18006 66126 18058
rect 66126 18006 66178 18058
rect 66178 18006 66180 18058
rect 66124 18004 66180 18006
rect 65916 16490 65972 16492
rect 65916 16438 65918 16490
rect 65918 16438 65970 16490
rect 65970 16438 65972 16490
rect 65916 16436 65972 16438
rect 66020 16490 66076 16492
rect 66020 16438 66022 16490
rect 66022 16438 66074 16490
rect 66074 16438 66076 16490
rect 66020 16436 66076 16438
rect 66124 16490 66180 16492
rect 66124 16438 66126 16490
rect 66126 16438 66178 16490
rect 66178 16438 66180 16490
rect 66124 16436 66180 16438
rect 65916 14922 65972 14924
rect 65916 14870 65918 14922
rect 65918 14870 65970 14922
rect 65970 14870 65972 14922
rect 65916 14868 65972 14870
rect 66020 14922 66076 14924
rect 66020 14870 66022 14922
rect 66022 14870 66074 14922
rect 66074 14870 66076 14922
rect 66020 14868 66076 14870
rect 66124 14922 66180 14924
rect 66124 14870 66126 14922
rect 66126 14870 66178 14922
rect 66178 14870 66180 14922
rect 66124 14868 66180 14870
rect 65916 13354 65972 13356
rect 65916 13302 65918 13354
rect 65918 13302 65970 13354
rect 65970 13302 65972 13354
rect 65916 13300 65972 13302
rect 66020 13354 66076 13356
rect 66020 13302 66022 13354
rect 66022 13302 66074 13354
rect 66074 13302 66076 13354
rect 66020 13300 66076 13302
rect 66124 13354 66180 13356
rect 66124 13302 66126 13354
rect 66126 13302 66178 13354
rect 66178 13302 66180 13354
rect 66124 13300 66180 13302
rect 65916 11786 65972 11788
rect 65916 11734 65918 11786
rect 65918 11734 65970 11786
rect 65970 11734 65972 11786
rect 65916 11732 65972 11734
rect 66020 11786 66076 11788
rect 66020 11734 66022 11786
rect 66022 11734 66074 11786
rect 66074 11734 66076 11786
rect 66020 11732 66076 11734
rect 66124 11786 66180 11788
rect 66124 11734 66126 11786
rect 66126 11734 66178 11786
rect 66178 11734 66180 11786
rect 66124 11732 66180 11734
rect 65916 10218 65972 10220
rect 65916 10166 65918 10218
rect 65918 10166 65970 10218
rect 65970 10166 65972 10218
rect 65916 10164 65972 10166
rect 66020 10218 66076 10220
rect 66020 10166 66022 10218
rect 66022 10166 66074 10218
rect 66074 10166 66076 10218
rect 66020 10164 66076 10166
rect 66124 10218 66180 10220
rect 66124 10166 66126 10218
rect 66126 10166 66178 10218
rect 66178 10166 66180 10218
rect 66124 10164 66180 10166
rect 66556 9212 66612 9268
rect 65916 8650 65972 8652
rect 65916 8598 65918 8650
rect 65918 8598 65970 8650
rect 65970 8598 65972 8650
rect 65916 8596 65972 8598
rect 66020 8650 66076 8652
rect 66020 8598 66022 8650
rect 66022 8598 66074 8650
rect 66074 8598 66076 8650
rect 66020 8596 66076 8598
rect 66124 8650 66180 8652
rect 66124 8598 66126 8650
rect 66126 8598 66178 8650
rect 66178 8598 66180 8650
rect 66124 8596 66180 8598
rect 65916 7082 65972 7084
rect 65916 7030 65918 7082
rect 65918 7030 65970 7082
rect 65970 7030 65972 7082
rect 65916 7028 65972 7030
rect 66020 7082 66076 7084
rect 66020 7030 66022 7082
rect 66022 7030 66074 7082
rect 66074 7030 66076 7082
rect 66020 7028 66076 7030
rect 66124 7082 66180 7084
rect 66124 7030 66126 7082
rect 66126 7030 66178 7082
rect 66178 7030 66180 7082
rect 66124 7028 66180 7030
rect 65916 5514 65972 5516
rect 65916 5462 65918 5514
rect 65918 5462 65970 5514
rect 65970 5462 65972 5514
rect 65916 5460 65972 5462
rect 66020 5514 66076 5516
rect 66020 5462 66022 5514
rect 66022 5462 66074 5514
rect 66074 5462 66076 5514
rect 66020 5460 66076 5462
rect 66124 5514 66180 5516
rect 66124 5462 66126 5514
rect 66126 5462 66178 5514
rect 66178 5462 66180 5514
rect 66124 5460 66180 5462
rect 65548 5068 65604 5124
rect 66332 5180 66388 5236
rect 64092 4060 64148 4116
rect 63868 3666 63924 3668
rect 63868 3614 63870 3666
rect 63870 3614 63922 3666
rect 63922 3614 63924 3666
rect 63868 3612 63924 3614
rect 65916 3946 65972 3948
rect 65916 3894 65918 3946
rect 65918 3894 65970 3946
rect 65970 3894 65972 3946
rect 65916 3892 65972 3894
rect 66020 3946 66076 3948
rect 66020 3894 66022 3946
rect 66022 3894 66074 3946
rect 66074 3894 66076 3946
rect 66020 3892 66076 3894
rect 66124 3946 66180 3948
rect 66124 3894 66126 3946
rect 66126 3894 66178 3946
rect 66178 3894 66180 3946
rect 66124 3892 66180 3894
rect 65548 3724 65604 3780
rect 64540 3612 64596 3668
rect 65660 3666 65716 3668
rect 65660 3614 65662 3666
rect 65662 3614 65714 3666
rect 65714 3614 65716 3666
rect 65660 3612 65716 3614
rect 65436 3500 65492 3556
rect 64764 3388 64820 3444
rect 66668 7698 66724 7700
rect 66668 7646 66670 7698
rect 66670 7646 66722 7698
rect 66722 7646 66724 7698
rect 66668 7644 66724 7646
rect 67116 7196 67172 7252
rect 68796 17388 68852 17444
rect 68908 16268 68964 16324
rect 68796 15036 68852 15092
rect 68460 14364 68516 14420
rect 67340 5516 67396 5572
rect 66780 5068 66836 5124
rect 67564 6076 67620 6132
rect 69580 26348 69636 26404
rect 70924 27858 70980 27860
rect 70924 27806 70926 27858
rect 70926 27806 70978 27858
rect 70978 27806 70980 27858
rect 70924 27804 70980 27806
rect 71708 28754 71764 28756
rect 71708 28702 71710 28754
rect 71710 28702 71762 28754
rect 71762 28702 71764 28754
rect 71708 28700 71764 28702
rect 71932 28588 71988 28644
rect 71820 28140 71876 28196
rect 71372 27580 71428 27636
rect 70924 26514 70980 26516
rect 70924 26462 70926 26514
rect 70926 26462 70978 26514
rect 70978 26462 70980 26514
rect 70924 26460 70980 26462
rect 71260 26348 71316 26404
rect 69468 23324 69524 23380
rect 71148 25900 71204 25956
rect 71036 25228 71092 25284
rect 70812 24668 70868 24724
rect 71372 25340 71428 25396
rect 71372 24610 71428 24612
rect 71372 24558 71374 24610
rect 71374 24558 71426 24610
rect 71426 24558 71428 24610
rect 71372 24556 71428 24558
rect 70700 22988 70756 23044
rect 71372 24332 71428 24388
rect 70588 22540 70644 22596
rect 70924 22652 70980 22708
rect 70364 22204 70420 22260
rect 70028 21810 70084 21812
rect 70028 21758 70030 21810
rect 70030 21758 70082 21810
rect 70082 21758 70084 21810
rect 70028 21756 70084 21758
rect 70364 19292 70420 19348
rect 71932 27916 71988 27972
rect 71932 27356 71988 27412
rect 71708 24946 71764 24948
rect 71708 24894 71710 24946
rect 71710 24894 71762 24946
rect 71762 24894 71764 24946
rect 71708 24892 71764 24894
rect 71260 20636 71316 20692
rect 71708 23378 71764 23380
rect 71708 23326 71710 23378
rect 71710 23326 71762 23378
rect 71762 23326 71764 23378
rect 71708 23324 71764 23326
rect 71708 23100 71764 23156
rect 71708 22316 71764 22372
rect 71596 21420 71652 21476
rect 72268 31500 72324 31556
rect 72156 31388 72212 31444
rect 73388 36988 73444 37044
rect 73500 36876 73556 36932
rect 73276 35644 73332 35700
rect 72828 34412 72884 34468
rect 72940 35196 72996 35252
rect 73052 34690 73108 34692
rect 73052 34638 73054 34690
rect 73054 34638 73106 34690
rect 73106 34638 73108 34690
rect 73052 34636 73108 34638
rect 73164 34412 73220 34468
rect 73164 34242 73220 34244
rect 73164 34190 73166 34242
rect 73166 34190 73218 34242
rect 73218 34190 73220 34242
rect 73164 34188 73220 34190
rect 72716 34130 72772 34132
rect 72716 34078 72718 34130
rect 72718 34078 72770 34130
rect 72770 34078 72772 34130
rect 72716 34076 72772 34078
rect 72940 32956 72996 33012
rect 72604 31836 72660 31892
rect 73052 31778 73108 31780
rect 73052 31726 73054 31778
rect 73054 31726 73106 31778
rect 73106 31726 73108 31778
rect 73052 31724 73108 31726
rect 72716 31388 72772 31444
rect 72156 29708 72212 29764
rect 72828 30156 72884 30212
rect 72716 30098 72772 30100
rect 72716 30046 72718 30098
rect 72718 30046 72770 30098
rect 72770 30046 72772 30098
rect 72716 30044 72772 30046
rect 72604 29932 72660 29988
rect 72716 29820 72772 29876
rect 72716 29314 72772 29316
rect 72716 29262 72718 29314
rect 72718 29262 72770 29314
rect 72770 29262 72772 29314
rect 72716 29260 72772 29262
rect 72604 28924 72660 28980
rect 72380 28642 72436 28644
rect 72380 28590 72382 28642
rect 72382 28590 72434 28642
rect 72434 28590 72436 28642
rect 72380 28588 72436 28590
rect 72268 27916 72324 27972
rect 72380 27074 72436 27076
rect 72380 27022 72382 27074
rect 72382 27022 72434 27074
rect 72434 27022 72436 27074
rect 72380 27020 72436 27022
rect 72380 26796 72436 26852
rect 72716 28530 72772 28532
rect 72716 28478 72718 28530
rect 72718 28478 72770 28530
rect 72770 28478 72772 28530
rect 72716 28476 72772 28478
rect 73052 29932 73108 29988
rect 72940 28924 72996 28980
rect 72828 28140 72884 28196
rect 72940 28476 72996 28532
rect 72716 27970 72772 27972
rect 72716 27918 72718 27970
rect 72718 27918 72770 27970
rect 72770 27918 72772 27970
rect 72716 27916 72772 27918
rect 72604 27244 72660 27300
rect 73276 31500 73332 31556
rect 73948 36988 74004 37044
rect 74060 37100 74116 37156
rect 73612 36204 73668 36260
rect 73612 35308 73668 35364
rect 73500 35196 73556 35252
rect 73612 35084 73668 35140
rect 73500 34802 73556 34804
rect 73500 34750 73502 34802
rect 73502 34750 73554 34802
rect 73554 34750 73556 34802
rect 73500 34748 73556 34750
rect 74508 38050 74564 38052
rect 74508 37998 74510 38050
rect 74510 37998 74562 38050
rect 74562 37998 74564 38050
rect 74508 37996 74564 37998
rect 75180 41298 75236 41300
rect 75180 41246 75182 41298
rect 75182 41246 75234 41298
rect 75234 41246 75236 41298
rect 75180 41244 75236 41246
rect 74956 40348 75012 40404
rect 75068 39788 75124 39844
rect 74956 39452 75012 39508
rect 75292 39900 75348 39956
rect 75404 40124 75460 40180
rect 75292 39564 75348 39620
rect 75628 39676 75684 39732
rect 75068 38892 75124 38948
rect 74956 38220 75012 38276
rect 75068 38556 75124 38612
rect 74284 37436 74340 37492
rect 74284 37266 74340 37268
rect 74284 37214 74286 37266
rect 74286 37214 74338 37266
rect 74338 37214 74340 37266
rect 74284 37212 74340 37214
rect 74620 37266 74676 37268
rect 74620 37214 74622 37266
rect 74622 37214 74674 37266
rect 74674 37214 74676 37266
rect 74620 37212 74676 37214
rect 74508 37154 74564 37156
rect 74508 37102 74510 37154
rect 74510 37102 74562 37154
rect 74562 37102 74564 37154
rect 74508 37100 74564 37102
rect 74284 36988 74340 37044
rect 75068 37266 75124 37268
rect 75068 37214 75070 37266
rect 75070 37214 75122 37266
rect 75122 37214 75124 37266
rect 75068 37212 75124 37214
rect 75180 36988 75236 37044
rect 75852 40124 75908 40180
rect 75404 38556 75460 38612
rect 75964 39788 76020 39844
rect 76076 39676 76132 39732
rect 76188 39506 76244 39508
rect 76188 39454 76190 39506
rect 76190 39454 76242 39506
rect 76242 39454 76244 39506
rect 76188 39452 76244 39454
rect 76524 42866 76580 42868
rect 76524 42814 76526 42866
rect 76526 42814 76578 42866
rect 76578 42814 76580 42866
rect 76524 42812 76580 42814
rect 76412 42700 76468 42756
rect 76412 41244 76468 41300
rect 76748 41356 76804 41412
rect 76524 41020 76580 41076
rect 76524 39618 76580 39620
rect 76524 39566 76526 39618
rect 76526 39566 76578 39618
rect 76578 39566 76580 39618
rect 76524 39564 76580 39566
rect 76412 38892 76468 38948
rect 76076 37884 76132 37940
rect 75404 37266 75460 37268
rect 75404 37214 75406 37266
rect 75406 37214 75458 37266
rect 75458 37214 75460 37266
rect 75404 37212 75460 37214
rect 76188 37378 76244 37380
rect 76188 37326 76190 37378
rect 76190 37326 76242 37378
rect 76242 37326 76244 37378
rect 76188 37324 76244 37326
rect 75516 37100 75572 37156
rect 74732 36540 74788 36596
rect 75628 36370 75684 36372
rect 75628 36318 75630 36370
rect 75630 36318 75682 36370
rect 75682 36318 75684 36370
rect 75628 36316 75684 36318
rect 75068 35980 75124 36036
rect 74060 35308 74116 35364
rect 73836 35196 73892 35252
rect 73724 34130 73780 34132
rect 73724 34078 73726 34130
rect 73726 34078 73778 34130
rect 73778 34078 73780 34130
rect 73724 34076 73780 34078
rect 73948 34412 74004 34468
rect 73948 33570 74004 33572
rect 73948 33518 73950 33570
rect 73950 33518 74002 33570
rect 74002 33518 74004 33570
rect 73948 33516 74004 33518
rect 73836 33458 73892 33460
rect 73836 33406 73838 33458
rect 73838 33406 73890 33458
rect 73890 33406 73892 33458
rect 73836 33404 73892 33406
rect 73724 32732 73780 32788
rect 73948 32844 74004 32900
rect 73500 32450 73556 32452
rect 73500 32398 73502 32450
rect 73502 32398 73554 32450
rect 73554 32398 73556 32450
rect 73500 32396 73556 32398
rect 73724 31778 73780 31780
rect 73724 31726 73726 31778
rect 73726 31726 73778 31778
rect 73778 31726 73780 31778
rect 73724 31724 73780 31726
rect 73500 31276 73556 31332
rect 73836 30994 73892 30996
rect 73836 30942 73838 30994
rect 73838 30942 73890 30994
rect 73890 30942 73892 30994
rect 73836 30940 73892 30942
rect 74284 35532 74340 35588
rect 74172 34690 74228 34692
rect 74172 34638 74174 34690
rect 74174 34638 74226 34690
rect 74226 34638 74228 34690
rect 74172 34636 74228 34638
rect 74284 33292 74340 33348
rect 74620 35420 74676 35476
rect 76412 37826 76468 37828
rect 76412 37774 76414 37826
rect 76414 37774 76466 37826
rect 76466 37774 76468 37826
rect 76412 37772 76468 37774
rect 76748 40908 76804 40964
rect 76748 38892 76804 38948
rect 77644 66780 77700 66836
rect 77644 65660 77700 65716
rect 77644 64706 77700 64708
rect 77644 64654 77646 64706
rect 77646 64654 77698 64706
rect 77698 64654 77700 64706
rect 77644 64652 77700 64654
rect 77420 64594 77476 64596
rect 77420 64542 77422 64594
rect 77422 64542 77474 64594
rect 77474 64542 77476 64594
rect 77420 64540 77476 64542
rect 77644 63980 77700 64036
rect 77420 63922 77476 63924
rect 77420 63870 77422 63922
rect 77422 63870 77474 63922
rect 77474 63870 77476 63922
rect 77420 63868 77476 63870
rect 77644 62914 77700 62916
rect 77644 62862 77646 62914
rect 77646 62862 77698 62914
rect 77698 62862 77700 62914
rect 77644 62860 77700 62862
rect 77644 61570 77700 61572
rect 77644 61518 77646 61570
rect 77646 61518 77698 61570
rect 77698 61518 77700 61570
rect 77644 61516 77700 61518
rect 77868 74002 77924 74004
rect 77868 73950 77870 74002
rect 77870 73950 77922 74002
rect 77922 73950 77924 74002
rect 77868 73948 77924 73950
rect 77868 73442 77924 73444
rect 77868 73390 77870 73442
rect 77870 73390 77922 73442
rect 77922 73390 77924 73442
rect 77868 73388 77924 73390
rect 78652 75516 78708 75572
rect 78092 75404 78148 75460
rect 78204 75122 78260 75124
rect 78204 75070 78206 75122
rect 78206 75070 78258 75122
rect 78258 75070 78260 75122
rect 78204 75068 78260 75070
rect 78764 75068 78820 75124
rect 79100 74956 79156 75012
rect 78316 74620 78372 74676
rect 78092 74114 78148 74116
rect 78092 74062 78094 74114
rect 78094 74062 78146 74114
rect 78146 74062 78148 74114
rect 78092 74060 78148 74062
rect 78204 73554 78260 73556
rect 78204 73502 78206 73554
rect 78206 73502 78258 73554
rect 78258 73502 78260 73554
rect 78204 73500 78260 73502
rect 78204 72434 78260 72436
rect 78204 72382 78206 72434
rect 78206 72382 78258 72434
rect 78258 72382 78260 72434
rect 78204 72380 78260 72382
rect 77868 72322 77924 72324
rect 77868 72270 77870 72322
rect 77870 72270 77922 72322
rect 77922 72270 77924 72322
rect 77868 72268 77924 72270
rect 77868 71874 77924 71876
rect 77868 71822 77870 71874
rect 77870 71822 77922 71874
rect 77922 71822 77924 71874
rect 77868 71820 77924 71822
rect 78204 71260 78260 71316
rect 78204 70754 78260 70756
rect 78204 70702 78206 70754
rect 78206 70702 78258 70754
rect 78258 70702 78260 70754
rect 78204 70700 78260 70702
rect 78204 70140 78260 70196
rect 77868 69186 77924 69188
rect 77868 69134 77870 69186
rect 77870 69134 77922 69186
rect 77922 69134 77924 69186
rect 77868 69132 77924 69134
rect 78204 69020 78260 69076
rect 78204 68626 78260 68628
rect 78204 68574 78206 68626
rect 78206 68574 78258 68626
rect 78258 68574 78260 68626
rect 78204 68572 78260 68574
rect 78204 67900 78260 67956
rect 78764 70924 78820 70980
rect 77868 66050 77924 66052
rect 77868 65998 77870 66050
rect 77870 65998 77922 66050
rect 77922 65998 77924 66050
rect 77868 65996 77924 65998
rect 77868 62188 77924 62244
rect 78204 66780 78260 66836
rect 78204 65660 78260 65716
rect 78204 64594 78260 64596
rect 78204 64542 78206 64594
rect 78206 64542 78258 64594
rect 78258 64542 78260 64594
rect 78204 64540 78260 64542
rect 78204 63922 78260 63924
rect 78204 63870 78206 63922
rect 78206 63870 78258 63922
rect 78258 63870 78260 63922
rect 78204 63868 78260 63870
rect 78204 63420 78260 63476
rect 78204 62860 78260 62916
rect 78204 62300 78260 62356
rect 77420 61180 77476 61236
rect 77868 60898 77924 60900
rect 77868 60846 77870 60898
rect 77870 60846 77922 60898
rect 77922 60846 77924 60898
rect 77868 60844 77924 60846
rect 77644 60786 77700 60788
rect 77644 60734 77646 60786
rect 77646 60734 77698 60786
rect 77698 60734 77700 60786
rect 77644 60732 77700 60734
rect 77644 59106 77700 59108
rect 77644 59054 77646 59106
rect 77646 59054 77698 59106
rect 77698 59054 77700 59106
rect 77644 59052 77700 59054
rect 77420 58940 77476 58996
rect 77868 58210 77924 58212
rect 77868 58158 77870 58210
rect 77870 58158 77922 58210
rect 77922 58158 77924 58210
rect 77868 58156 77924 58158
rect 77644 57820 77700 57876
rect 77644 56754 77700 56756
rect 77644 56702 77646 56754
rect 77646 56702 77698 56754
rect 77698 56702 77700 56754
rect 77644 56700 77700 56702
rect 77868 56194 77924 56196
rect 77868 56142 77870 56194
rect 77870 56142 77922 56194
rect 77922 56142 77924 56194
rect 77868 56140 77924 56142
rect 77308 50316 77364 50372
rect 77644 55580 77700 55636
rect 77644 55074 77700 55076
rect 77644 55022 77646 55074
rect 77646 55022 77698 55074
rect 77698 55022 77700 55074
rect 77644 55020 77700 55022
rect 77868 54012 77924 54068
rect 77868 53788 77924 53844
rect 77644 53340 77700 53396
rect 78204 61180 78260 61236
rect 78204 60786 78260 60788
rect 78204 60734 78206 60786
rect 78206 60734 78258 60786
rect 78258 60734 78260 60786
rect 78204 60732 78260 60734
rect 78204 60060 78260 60116
rect 78204 58940 78260 58996
rect 78204 57820 78260 57876
rect 78204 56754 78260 56756
rect 78204 56702 78206 56754
rect 78206 56702 78258 56754
rect 78258 56702 78260 56754
rect 78204 56700 78260 56702
rect 78204 55580 78260 55636
rect 78204 55020 78260 55076
rect 78204 54460 78260 54516
rect 78204 53340 78260 53396
rect 77644 52834 77700 52836
rect 77644 52782 77646 52834
rect 77646 52782 77698 52834
rect 77698 52782 77700 52834
rect 77644 52780 77700 52782
rect 77644 51100 77700 51156
rect 77644 50482 77700 50484
rect 77644 50430 77646 50482
rect 77646 50430 77698 50482
rect 77698 50430 77700 50482
rect 77644 50428 77700 50430
rect 77868 51490 77924 51492
rect 77868 51438 77870 51490
rect 77870 51438 77922 51490
rect 77922 51438 77924 51490
rect 77868 51436 77924 51438
rect 77868 50370 77924 50372
rect 77868 50318 77870 50370
rect 77870 50318 77922 50370
rect 77922 50318 77924 50370
rect 77868 50316 77924 50318
rect 77644 48914 77700 48916
rect 77644 48862 77646 48914
rect 77646 48862 77698 48914
rect 77698 48862 77700 48914
rect 77644 48860 77700 48862
rect 77420 46844 77476 46900
rect 77868 48354 77924 48356
rect 77868 48302 77870 48354
rect 77870 48302 77922 48354
rect 77922 48302 77924 48354
rect 77868 48300 77924 48302
rect 77644 47740 77700 47796
rect 77644 47346 77700 47348
rect 77644 47294 77646 47346
rect 77646 47294 77698 47346
rect 77698 47294 77700 47346
rect 77644 47292 77700 47294
rect 77868 47234 77924 47236
rect 77868 47182 77870 47234
rect 77870 47182 77922 47234
rect 77922 47182 77924 47234
rect 77868 47180 77924 47182
rect 77532 46172 77588 46228
rect 77644 45500 77700 45556
rect 77308 45276 77364 45332
rect 77644 44994 77700 44996
rect 77644 44942 77646 44994
rect 77646 44942 77698 44994
rect 77698 44942 77700 44994
rect 77644 44940 77700 44942
rect 77868 45218 77924 45220
rect 77868 45166 77870 45218
rect 77870 45166 77922 45218
rect 77922 45166 77924 45218
rect 77868 45164 77924 45166
rect 77756 44604 77812 44660
rect 78204 52780 78260 52836
rect 78204 52220 78260 52276
rect 78204 51100 78260 51156
rect 78204 50482 78260 50484
rect 78204 50430 78206 50482
rect 78206 50430 78258 50482
rect 78258 50430 78260 50482
rect 78204 50428 78260 50430
rect 78204 49980 78260 50036
rect 78204 48914 78260 48916
rect 78204 48862 78206 48914
rect 78206 48862 78258 48914
rect 78258 48862 78260 48914
rect 78204 48860 78260 48862
rect 78204 47740 78260 47796
rect 78092 46956 78148 47012
rect 78204 47346 78260 47348
rect 78204 47294 78206 47346
rect 78206 47294 78258 47346
rect 78258 47294 78260 47346
rect 78204 47292 78260 47294
rect 78204 46620 78260 46676
rect 78204 45500 78260 45556
rect 78204 44940 78260 44996
rect 78204 44380 78260 44436
rect 77868 43650 77924 43652
rect 77868 43598 77870 43650
rect 77870 43598 77922 43650
rect 77922 43598 77924 43650
rect 77868 43596 77924 43598
rect 77084 43538 77140 43540
rect 77084 43486 77086 43538
rect 77086 43486 77138 43538
rect 77138 43486 77140 43538
rect 77084 43484 77140 43486
rect 77644 43260 77700 43316
rect 78204 43260 78260 43316
rect 77308 43036 77364 43092
rect 77084 42812 77140 42868
rect 77420 42642 77476 42644
rect 77420 42590 77422 42642
rect 77422 42590 77474 42642
rect 77474 42590 77476 42642
rect 77420 42588 77476 42590
rect 76972 40124 77028 40180
rect 77084 40908 77140 40964
rect 76972 38834 77028 38836
rect 76972 38782 76974 38834
rect 76974 38782 77026 38834
rect 77026 38782 77028 38834
rect 76972 38780 77028 38782
rect 77196 39116 77252 39172
rect 77420 39004 77476 39060
rect 77756 42028 77812 42084
rect 77980 42140 78036 42196
rect 78092 41298 78148 41300
rect 78092 41246 78094 41298
rect 78094 41246 78146 41298
rect 78146 41246 78148 41298
rect 78092 41244 78148 41246
rect 77644 40908 77700 40964
rect 77644 40572 77700 40628
rect 77980 40236 78036 40292
rect 78540 48300 78596 48356
rect 78540 40796 78596 40852
rect 78764 47180 78820 47236
rect 78092 39900 78148 39956
rect 76412 37490 76468 37492
rect 76412 37438 76414 37490
rect 76414 37438 76466 37490
rect 76466 37438 76468 37490
rect 76412 37436 76468 37438
rect 76076 35980 76132 36036
rect 76188 36988 76244 37044
rect 75628 35756 75684 35812
rect 74620 34412 74676 34468
rect 74620 34076 74676 34132
rect 74396 33180 74452 33236
rect 74172 33068 74228 33124
rect 74396 32060 74452 32116
rect 74284 31948 74340 32004
rect 74844 33740 74900 33796
rect 74844 33458 74900 33460
rect 74844 33406 74846 33458
rect 74846 33406 74898 33458
rect 74898 33406 74900 33458
rect 74844 33404 74900 33406
rect 75292 34636 75348 34692
rect 75068 34188 75124 34244
rect 75292 33852 75348 33908
rect 75180 33628 75236 33684
rect 75068 33516 75124 33572
rect 75292 33346 75348 33348
rect 75292 33294 75294 33346
rect 75294 33294 75346 33346
rect 75346 33294 75348 33346
rect 75292 33292 75348 33294
rect 75068 32620 75124 32676
rect 75180 33180 75236 33236
rect 74844 32338 74900 32340
rect 74844 32286 74846 32338
rect 74846 32286 74898 32338
rect 74898 32286 74900 32338
rect 74844 32284 74900 32286
rect 75068 32284 75124 32340
rect 74956 32172 75012 32228
rect 74172 30994 74228 30996
rect 74172 30942 74174 30994
rect 74174 30942 74226 30994
rect 74226 30942 74228 30994
rect 74172 30940 74228 30942
rect 74060 30322 74116 30324
rect 74060 30270 74062 30322
rect 74062 30270 74114 30322
rect 74114 30270 74116 30322
rect 74060 30268 74116 30270
rect 73500 29932 73556 29988
rect 74620 31666 74676 31668
rect 74620 31614 74622 31666
rect 74622 31614 74674 31666
rect 74674 31614 74676 31666
rect 74620 31612 74676 31614
rect 74508 31554 74564 31556
rect 74508 31502 74510 31554
rect 74510 31502 74562 31554
rect 74562 31502 74564 31554
rect 74508 31500 74564 31502
rect 74508 31106 74564 31108
rect 74508 31054 74510 31106
rect 74510 31054 74562 31106
rect 74562 31054 74564 31106
rect 74508 31052 74564 31054
rect 74844 30994 74900 30996
rect 74844 30942 74846 30994
rect 74846 30942 74898 30994
rect 74898 30942 74900 30994
rect 74844 30940 74900 30942
rect 74732 30268 74788 30324
rect 74508 30044 74564 30100
rect 73724 29596 73780 29652
rect 73724 29426 73780 29428
rect 73724 29374 73726 29426
rect 73726 29374 73778 29426
rect 73778 29374 73780 29426
rect 73724 29372 73780 29374
rect 73612 29148 73668 29204
rect 73388 28924 73444 28980
rect 73724 28476 73780 28532
rect 73500 27858 73556 27860
rect 73500 27806 73502 27858
rect 73502 27806 73554 27858
rect 73554 27806 73556 27858
rect 73500 27804 73556 27806
rect 73164 27132 73220 27188
rect 73388 27244 73444 27300
rect 72380 26460 72436 26516
rect 72268 25452 72324 25508
rect 72380 26290 72436 26292
rect 72380 26238 72382 26290
rect 72382 26238 72434 26290
rect 72434 26238 72436 26290
rect 72380 26236 72436 26238
rect 72156 25116 72212 25172
rect 72156 24892 72212 24948
rect 72380 24498 72436 24500
rect 72380 24446 72382 24498
rect 72382 24446 72434 24498
rect 72434 24446 72436 24498
rect 72380 24444 72436 24446
rect 72156 23714 72212 23716
rect 72156 23662 72158 23714
rect 72158 23662 72210 23714
rect 72210 23662 72212 23714
rect 72156 23660 72212 23662
rect 72156 23324 72212 23380
rect 72156 22482 72212 22484
rect 72156 22430 72158 22482
rect 72158 22430 72210 22482
rect 72210 22430 72212 22482
rect 72156 22428 72212 22430
rect 70588 17724 70644 17780
rect 72156 19180 72212 19236
rect 71372 18396 71428 18452
rect 70252 16604 70308 16660
rect 69356 10892 69412 10948
rect 69020 9324 69076 9380
rect 68572 5068 68628 5124
rect 68124 4844 68180 4900
rect 67452 3778 67508 3780
rect 67452 3726 67454 3778
rect 67454 3726 67506 3778
rect 67506 3726 67508 3778
rect 67452 3724 67508 3726
rect 68348 4114 68404 4116
rect 68348 4062 68350 4114
rect 68350 4062 68402 4114
rect 68402 4062 68404 4114
rect 68348 4060 68404 4062
rect 68796 4060 68852 4116
rect 69804 7644 69860 7700
rect 69020 5628 69076 5684
rect 69356 5516 69412 5572
rect 69356 5234 69412 5236
rect 69356 5182 69358 5234
rect 69358 5182 69410 5234
rect 69410 5182 69412 5234
rect 69356 5180 69412 5182
rect 68908 3500 68964 3556
rect 69468 3724 69524 3780
rect 70476 6412 70532 6468
rect 71036 5906 71092 5908
rect 71036 5854 71038 5906
rect 71038 5854 71090 5906
rect 71090 5854 71092 5906
rect 71036 5852 71092 5854
rect 70476 5516 70532 5572
rect 70812 5628 70868 5684
rect 70476 4284 70532 4340
rect 70476 3948 70532 4004
rect 72492 22204 72548 22260
rect 72716 26460 72772 26516
rect 73836 28364 73892 28420
rect 73052 26962 73108 26964
rect 73052 26910 73054 26962
rect 73054 26910 73106 26962
rect 73106 26910 73108 26962
rect 73052 26908 73108 26910
rect 73052 26572 73108 26628
rect 72940 26178 72996 26180
rect 72940 26126 72942 26178
rect 72942 26126 72994 26178
rect 72994 26126 72996 26178
rect 72940 26124 72996 26126
rect 72940 20914 72996 20916
rect 72940 20862 72942 20914
rect 72942 20862 72994 20914
rect 72994 20862 72996 20914
rect 72940 20860 72996 20862
rect 72380 20188 72436 20244
rect 72716 20802 72772 20804
rect 72716 20750 72718 20802
rect 72718 20750 72770 20802
rect 72770 20750 72772 20802
rect 72716 20748 72772 20750
rect 73612 26796 73668 26852
rect 73276 26012 73332 26068
rect 73500 26012 73556 26068
rect 73276 25506 73332 25508
rect 73276 25454 73278 25506
rect 73278 25454 73330 25506
rect 73330 25454 73332 25506
rect 73276 25452 73332 25454
rect 73500 24722 73556 24724
rect 73500 24670 73502 24722
rect 73502 24670 73554 24722
rect 73554 24670 73556 24722
rect 73500 24668 73556 24670
rect 73948 26908 74004 26964
rect 73276 23938 73332 23940
rect 73276 23886 73278 23938
rect 73278 23886 73330 23938
rect 73330 23886 73332 23938
rect 73276 23884 73332 23886
rect 73612 23938 73668 23940
rect 73612 23886 73614 23938
rect 73614 23886 73666 23938
rect 73666 23886 73668 23938
rect 73612 23884 73668 23886
rect 74956 30210 75012 30212
rect 74956 30158 74958 30210
rect 74958 30158 75010 30210
rect 75010 30158 75012 30210
rect 74956 30156 75012 30158
rect 74956 29538 75012 29540
rect 74956 29486 74958 29538
rect 74958 29486 75010 29538
rect 75010 29486 75012 29538
rect 74956 29484 75012 29486
rect 74284 28642 74340 28644
rect 74284 28590 74286 28642
rect 74286 28590 74338 28642
rect 74338 28590 74340 28642
rect 74284 28588 74340 28590
rect 74396 28476 74452 28532
rect 74172 27970 74228 27972
rect 74172 27918 74174 27970
rect 74174 27918 74226 27970
rect 74226 27918 74228 27970
rect 74172 27916 74228 27918
rect 74284 27858 74340 27860
rect 74284 27806 74286 27858
rect 74286 27806 74338 27858
rect 74338 27806 74340 27858
rect 74284 27804 74340 27806
rect 74508 28418 74564 28420
rect 74508 28366 74510 28418
rect 74510 28366 74562 28418
rect 74562 28366 74564 28418
rect 74508 28364 74564 28366
rect 75740 35420 75796 35476
rect 75516 33964 75572 34020
rect 75292 32396 75348 32452
rect 75180 30940 75236 30996
rect 76300 36706 76356 36708
rect 76300 36654 76302 36706
rect 76302 36654 76354 36706
rect 76354 36654 76356 36706
rect 76300 36652 76356 36654
rect 76524 36988 76580 37044
rect 76748 36988 76804 37044
rect 76300 36316 76356 36372
rect 76300 35868 76356 35924
rect 77308 37660 77364 37716
rect 77532 37436 77588 37492
rect 77644 37772 77700 37828
rect 76748 35756 76804 35812
rect 76972 35980 77028 36036
rect 76300 34300 76356 34356
rect 76524 34972 76580 35028
rect 75852 33628 75908 33684
rect 75740 31890 75796 31892
rect 75740 31838 75742 31890
rect 75742 31838 75794 31890
rect 75794 31838 75796 31890
rect 75740 31836 75796 31838
rect 75628 31276 75684 31332
rect 77196 35868 77252 35924
rect 77420 37154 77476 37156
rect 77420 37102 77422 37154
rect 77422 37102 77474 37154
rect 77474 37102 77476 37154
rect 77420 37100 77476 37102
rect 77420 36652 77476 36708
rect 77420 36316 77476 36372
rect 77308 35698 77364 35700
rect 77308 35646 77310 35698
rect 77310 35646 77362 35698
rect 77362 35646 77364 35698
rect 77308 35644 77364 35646
rect 77868 39116 77924 39172
rect 77980 39004 78036 39060
rect 78204 38780 78260 38836
rect 77756 36652 77812 36708
rect 77532 36092 77588 36148
rect 78428 37324 78484 37380
rect 77532 35810 77588 35812
rect 77532 35758 77534 35810
rect 77534 35758 77586 35810
rect 77586 35758 77588 35810
rect 77532 35756 77588 35758
rect 76412 34018 76468 34020
rect 76412 33966 76414 34018
rect 76414 33966 76466 34018
rect 76466 33966 76468 34018
rect 76412 33964 76468 33966
rect 76860 33628 76916 33684
rect 76748 33516 76804 33572
rect 76860 33404 76916 33460
rect 75964 32732 76020 32788
rect 76636 33122 76692 33124
rect 76636 33070 76638 33122
rect 76638 33070 76690 33122
rect 76690 33070 76692 33122
rect 76636 33068 76692 33070
rect 76860 33068 76916 33124
rect 77084 33628 77140 33684
rect 77308 33292 77364 33348
rect 77868 35084 77924 35140
rect 77532 34524 77588 34580
rect 78204 34524 78260 34580
rect 77532 34242 77588 34244
rect 77532 34190 77534 34242
rect 77534 34190 77586 34242
rect 77586 34190 77588 34242
rect 77532 34188 77588 34190
rect 77980 34076 78036 34132
rect 77868 33852 77924 33908
rect 77644 33628 77700 33684
rect 77756 33740 77812 33796
rect 77868 33516 77924 33572
rect 77532 32674 77588 32676
rect 77532 32622 77534 32674
rect 77534 32622 77586 32674
rect 77586 32622 77588 32674
rect 77532 32620 77588 32622
rect 76412 32396 76468 32452
rect 77420 32396 77476 32452
rect 77308 32060 77364 32116
rect 76860 31778 76916 31780
rect 76860 31726 76862 31778
rect 76862 31726 76914 31778
rect 76914 31726 76916 31778
rect 76860 31724 76916 31726
rect 76636 31554 76692 31556
rect 76636 31502 76638 31554
rect 76638 31502 76690 31554
rect 76690 31502 76692 31554
rect 76636 31500 76692 31502
rect 75516 31106 75572 31108
rect 75516 31054 75518 31106
rect 75518 31054 75570 31106
rect 75570 31054 75572 31106
rect 75516 31052 75572 31054
rect 75404 30380 75460 30436
rect 74396 27580 74452 27636
rect 74732 28588 74788 28644
rect 74396 26684 74452 26740
rect 73836 26236 73892 26292
rect 73836 26012 73892 26068
rect 74060 26066 74116 26068
rect 74060 26014 74062 26066
rect 74062 26014 74114 26066
rect 74114 26014 74116 26066
rect 74060 26012 74116 26014
rect 74172 25676 74228 25732
rect 74284 25564 74340 25620
rect 73836 23324 73892 23380
rect 74172 23772 74228 23828
rect 73500 22092 73556 22148
rect 73948 22370 74004 22372
rect 73948 22318 73950 22370
rect 73950 22318 74002 22370
rect 74002 22318 74004 22370
rect 73948 22316 74004 22318
rect 73612 21980 73668 22036
rect 73276 21586 73332 21588
rect 73276 21534 73278 21586
rect 73278 21534 73330 21586
rect 73330 21534 73332 21586
rect 73276 21532 73332 21534
rect 74060 21586 74116 21588
rect 74060 21534 74062 21586
rect 74062 21534 74114 21586
rect 74114 21534 74116 21586
rect 74060 21532 74116 21534
rect 74396 24220 74452 24276
rect 74732 27858 74788 27860
rect 74732 27806 74734 27858
rect 74734 27806 74786 27858
rect 74786 27806 74788 27858
rect 74732 27804 74788 27806
rect 75180 28530 75236 28532
rect 75180 28478 75182 28530
rect 75182 28478 75234 28530
rect 75234 28478 75236 28530
rect 75180 28476 75236 28478
rect 75068 28364 75124 28420
rect 74956 27970 75012 27972
rect 74956 27918 74958 27970
rect 74958 27918 75010 27970
rect 75010 27918 75012 27970
rect 74956 27916 75012 27918
rect 76188 30156 76244 30212
rect 76636 30994 76692 30996
rect 76636 30942 76638 30994
rect 76638 30942 76690 30994
rect 76690 30942 76692 30994
rect 76636 30940 76692 30942
rect 76524 30828 76580 30884
rect 75404 29314 75460 29316
rect 75404 29262 75406 29314
rect 75406 29262 75458 29314
rect 75458 29262 75460 29314
rect 75404 29260 75460 29262
rect 75404 28924 75460 28980
rect 75292 28364 75348 28420
rect 75404 27916 75460 27972
rect 74620 26962 74676 26964
rect 74620 26910 74622 26962
rect 74622 26910 74674 26962
rect 74674 26910 74676 26962
rect 74620 26908 74676 26910
rect 75068 27132 75124 27188
rect 75404 27692 75460 27748
rect 76636 30210 76692 30212
rect 76636 30158 76638 30210
rect 76638 30158 76690 30210
rect 76690 30158 76692 30210
rect 76636 30156 76692 30158
rect 76972 30156 77028 30212
rect 76524 30044 76580 30100
rect 76412 29820 76468 29876
rect 76076 29538 76132 29540
rect 76076 29486 76078 29538
rect 76078 29486 76130 29538
rect 76130 29486 76132 29538
rect 76076 29484 76132 29486
rect 76524 29484 76580 29540
rect 76188 29314 76244 29316
rect 76188 29262 76190 29314
rect 76190 29262 76242 29314
rect 76242 29262 76244 29314
rect 76188 29260 76244 29262
rect 75740 29202 75796 29204
rect 75740 29150 75742 29202
rect 75742 29150 75794 29202
rect 75794 29150 75796 29202
rect 75740 29148 75796 29150
rect 76524 28924 76580 28980
rect 75628 28642 75684 28644
rect 75628 28590 75630 28642
rect 75630 28590 75682 28642
rect 75682 28590 75684 28642
rect 75628 28588 75684 28590
rect 76860 29148 76916 29204
rect 76636 28642 76692 28644
rect 76636 28590 76638 28642
rect 76638 28590 76690 28642
rect 76690 28590 76692 28642
rect 76636 28588 76692 28590
rect 75852 28476 75908 28532
rect 75516 27356 75572 27412
rect 75628 28364 75684 28420
rect 76188 28530 76244 28532
rect 76188 28478 76190 28530
rect 76190 28478 76242 28530
rect 76242 28478 76244 28530
rect 76188 28476 76244 28478
rect 75964 28082 76020 28084
rect 75964 28030 75966 28082
rect 75966 28030 76018 28082
rect 76018 28030 76020 28082
rect 75964 28028 76020 28030
rect 75852 27970 75908 27972
rect 75852 27918 75854 27970
rect 75854 27918 75906 27970
rect 75906 27918 75908 27970
rect 75852 27916 75908 27918
rect 76188 27970 76244 27972
rect 76188 27918 76190 27970
rect 76190 27918 76242 27970
rect 76242 27918 76244 27970
rect 76188 27916 76244 27918
rect 75628 27244 75684 27300
rect 75964 27692 76020 27748
rect 75516 27132 75572 27188
rect 74844 25340 74900 25396
rect 74620 24220 74676 24276
rect 74732 24108 74788 24164
rect 75964 26908 76020 26964
rect 76636 27804 76692 27860
rect 75628 26684 75684 26740
rect 75516 25506 75572 25508
rect 75516 25454 75518 25506
rect 75518 25454 75570 25506
rect 75570 25454 75572 25506
rect 75516 25452 75572 25454
rect 75404 25340 75460 25396
rect 75292 24162 75348 24164
rect 75292 24110 75294 24162
rect 75294 24110 75346 24162
rect 75346 24110 75348 24162
rect 75292 24108 75348 24110
rect 74620 23826 74676 23828
rect 74620 23774 74622 23826
rect 74622 23774 74674 23826
rect 74674 23774 74676 23826
rect 74620 23772 74676 23774
rect 74844 23660 74900 23716
rect 75404 23938 75460 23940
rect 75404 23886 75406 23938
rect 75406 23886 75458 23938
rect 75458 23886 75460 23938
rect 75404 23884 75460 23886
rect 75068 22930 75124 22932
rect 75068 22878 75070 22930
rect 75070 22878 75122 22930
rect 75122 22878 75124 22930
rect 75068 22876 75124 22878
rect 74284 21532 74340 21588
rect 74284 20972 74340 21028
rect 74956 21868 75012 21924
rect 74844 20860 74900 20916
rect 73836 20076 73892 20132
rect 73052 19404 73108 19460
rect 72268 17836 72324 17892
rect 75964 25564 76020 25620
rect 76188 27298 76244 27300
rect 76188 27246 76190 27298
rect 76190 27246 76242 27298
rect 76242 27246 76244 27298
rect 76188 27244 76244 27246
rect 76300 26402 76356 26404
rect 76300 26350 76302 26402
rect 76302 26350 76354 26402
rect 76354 26350 76356 26402
rect 76300 26348 76356 26350
rect 76188 25452 76244 25508
rect 76524 26684 76580 26740
rect 76076 24556 76132 24612
rect 76524 24668 76580 24724
rect 76188 24162 76244 24164
rect 76188 24110 76190 24162
rect 76190 24110 76242 24162
rect 76242 24110 76244 24162
rect 76188 24108 76244 24110
rect 76076 23884 76132 23940
rect 76524 23772 76580 23828
rect 75740 22316 75796 22372
rect 75628 22204 75684 22260
rect 75964 22204 76020 22260
rect 75180 21698 75236 21700
rect 75180 21646 75182 21698
rect 75182 21646 75234 21698
rect 75234 21646 75236 21698
rect 75180 21644 75236 21646
rect 75516 21586 75572 21588
rect 75516 21534 75518 21586
rect 75518 21534 75570 21586
rect 75570 21534 75572 21586
rect 75516 21532 75572 21534
rect 75292 21420 75348 21476
rect 75852 21868 75908 21924
rect 75068 20524 75124 20580
rect 75628 19964 75684 20020
rect 75852 19292 75908 19348
rect 76860 27298 76916 27300
rect 76860 27246 76862 27298
rect 76862 27246 76914 27298
rect 76914 27246 76916 27298
rect 76860 27244 76916 27246
rect 76972 28140 77028 28196
rect 77420 31836 77476 31892
rect 77420 31106 77476 31108
rect 77420 31054 77422 31106
rect 77422 31054 77474 31106
rect 77474 31054 77476 31106
rect 77420 31052 77476 31054
rect 77196 29932 77252 29988
rect 77308 30268 77364 30324
rect 77196 29202 77252 29204
rect 77196 29150 77198 29202
rect 77198 29150 77250 29202
rect 77250 29150 77252 29202
rect 77196 29148 77252 29150
rect 77756 32786 77812 32788
rect 77756 32734 77758 32786
rect 77758 32734 77810 32786
rect 77810 32734 77812 32786
rect 77756 32732 77812 32734
rect 77756 32508 77812 32564
rect 77644 30994 77700 30996
rect 77644 30942 77646 30994
rect 77646 30942 77698 30994
rect 77698 30942 77700 30994
rect 77644 30940 77700 30942
rect 77644 30380 77700 30436
rect 78540 37212 78596 37268
rect 78764 37324 78820 37380
rect 78540 34524 78596 34580
rect 78652 35644 78708 35700
rect 78428 32396 78484 32452
rect 78204 32060 78260 32116
rect 77980 31276 78036 31332
rect 77084 27692 77140 27748
rect 78092 31052 78148 31108
rect 78876 35308 78932 35364
rect 78988 34188 79044 34244
rect 78764 33740 78820 33796
rect 78316 30604 78372 30660
rect 78316 29036 78372 29092
rect 78540 29820 78596 29876
rect 78428 28700 78484 28756
rect 78204 27970 78260 27972
rect 78204 27918 78206 27970
rect 78206 27918 78258 27970
rect 78258 27918 78260 27970
rect 78204 27916 78260 27918
rect 77756 27580 77812 27636
rect 77532 27244 77588 27300
rect 76748 26460 76804 26516
rect 77084 26684 77140 26740
rect 77756 27020 77812 27076
rect 77084 25676 77140 25732
rect 77420 26348 77476 26404
rect 78540 27916 78596 27972
rect 78876 31836 78932 31892
rect 77868 26684 77924 26740
rect 78092 26796 78148 26852
rect 78092 26236 78148 26292
rect 77756 25730 77812 25732
rect 77756 25678 77758 25730
rect 77758 25678 77810 25730
rect 77810 25678 77812 25730
rect 77756 25676 77812 25678
rect 77196 25116 77252 25172
rect 78540 26796 78596 26852
rect 78204 26124 78260 26180
rect 78764 26460 78820 26516
rect 78204 25340 78260 25396
rect 77644 25228 77700 25284
rect 76860 23826 76916 23828
rect 76860 23774 76862 23826
rect 76862 23774 76914 23826
rect 76914 23774 76916 23826
rect 76860 23772 76916 23774
rect 76748 22428 76804 22484
rect 77196 23212 77252 23268
rect 77868 23324 77924 23380
rect 78204 23660 78260 23716
rect 78316 23884 78372 23940
rect 77084 22316 77140 22372
rect 78092 23548 78148 23604
rect 78204 23100 78260 23156
rect 76412 21868 76468 21924
rect 76636 21868 76692 21924
rect 75404 15932 75460 15988
rect 74396 15036 74452 15092
rect 73052 12684 73108 12740
rect 71708 7586 71764 7588
rect 71708 7534 71710 7586
rect 71710 7534 71762 7586
rect 71762 7534 71764 7586
rect 71708 7532 71764 7534
rect 72380 7532 72436 7588
rect 72268 6466 72324 6468
rect 72268 6414 72270 6466
rect 72270 6414 72322 6466
rect 72322 6414 72324 6466
rect 72268 6412 72324 6414
rect 71708 5794 71764 5796
rect 71708 5742 71710 5794
rect 71710 5742 71762 5794
rect 71762 5742 71764 5794
rect 71708 5740 71764 5742
rect 72268 5740 72324 5796
rect 72828 5180 72884 5236
rect 72156 5068 72212 5124
rect 71708 4226 71764 4228
rect 71708 4174 71710 4226
rect 71710 4174 71762 4226
rect 71762 4174 71764 4226
rect 71708 4172 71764 4174
rect 71260 3666 71316 3668
rect 71260 3614 71262 3666
rect 71262 3614 71314 3666
rect 71314 3614 71316 3666
rect 71260 3612 71316 3614
rect 71484 3388 71540 3444
rect 72268 4898 72324 4900
rect 72268 4846 72270 4898
rect 72270 4846 72322 4898
rect 72322 4846 72324 4898
rect 72268 4844 72324 4846
rect 72268 4172 72324 4228
rect 73276 5682 73332 5684
rect 73276 5630 73278 5682
rect 73278 5630 73330 5682
rect 73330 5630 73332 5682
rect 73276 5628 73332 5630
rect 73724 8316 73780 8372
rect 73724 6636 73780 6692
rect 73836 8092 73892 8148
rect 73836 5404 73892 5460
rect 73388 4956 73444 5012
rect 73500 5292 73556 5348
rect 73052 4172 73108 4228
rect 73276 4114 73332 4116
rect 73276 4062 73278 4114
rect 73278 4062 73330 4114
rect 73330 4062 73332 4114
rect 73276 4060 73332 4062
rect 73948 5068 74004 5124
rect 74172 4172 74228 4228
rect 74060 3948 74116 4004
rect 74956 13074 75012 13076
rect 74956 13022 74958 13074
rect 74958 13022 75010 13074
rect 75010 13022 75012 13074
rect 74956 13020 75012 13022
rect 75628 13020 75684 13076
rect 75292 12738 75348 12740
rect 75292 12686 75294 12738
rect 75294 12686 75346 12738
rect 75346 12686 75348 12738
rect 75292 12684 75348 12686
rect 75516 9996 75572 10052
rect 74956 7532 75012 7588
rect 74508 6300 74564 6356
rect 74396 5852 74452 5908
rect 74620 5404 74676 5460
rect 75292 7644 75348 7700
rect 75404 8764 75460 8820
rect 75404 7532 75460 7588
rect 75292 7474 75348 7476
rect 75292 7422 75294 7474
rect 75294 7422 75346 7474
rect 75346 7422 75348 7474
rect 75292 7420 75348 7422
rect 75180 6748 75236 6804
rect 75404 7196 75460 7252
rect 74956 5404 75012 5460
rect 74956 5068 75012 5124
rect 74508 4956 74564 5012
rect 74508 2940 74564 2996
rect 74284 924 74340 980
rect 75180 5906 75236 5908
rect 75180 5854 75182 5906
rect 75182 5854 75234 5906
rect 75234 5854 75236 5906
rect 75180 5852 75236 5854
rect 75180 4898 75236 4900
rect 75180 4846 75182 4898
rect 75182 4846 75234 4898
rect 75234 4846 75236 4898
rect 75180 4844 75236 4846
rect 75180 4060 75236 4116
rect 75068 3778 75124 3780
rect 75068 3726 75070 3778
rect 75070 3726 75122 3778
rect 75122 3726 75124 3778
rect 75068 3724 75124 3726
rect 75516 6300 75572 6356
rect 75404 5516 75460 5572
rect 75292 3500 75348 3556
rect 75628 5404 75684 5460
rect 75852 8818 75908 8820
rect 75852 8766 75854 8818
rect 75854 8766 75906 8818
rect 75906 8766 75908 8818
rect 75852 8764 75908 8766
rect 76188 20130 76244 20132
rect 76188 20078 76190 20130
rect 76190 20078 76242 20130
rect 76242 20078 76244 20130
rect 76188 20076 76244 20078
rect 76076 20018 76132 20020
rect 76076 19966 76078 20018
rect 76078 19966 76130 20018
rect 76130 19966 76132 20018
rect 76076 19964 76132 19966
rect 76300 18508 76356 18564
rect 76300 13074 76356 13076
rect 76300 13022 76302 13074
rect 76302 13022 76354 13074
rect 76354 13022 76356 13074
rect 76300 13020 76356 13022
rect 76636 20748 76692 20804
rect 76748 21644 76804 21700
rect 77420 22092 77476 22148
rect 77308 21980 77364 22036
rect 77756 22146 77812 22148
rect 77756 22094 77758 22146
rect 77758 22094 77810 22146
rect 77810 22094 77812 22146
rect 77756 22092 77812 22094
rect 76972 20578 77028 20580
rect 76972 20526 76974 20578
rect 76974 20526 77026 20578
rect 77026 20526 77028 20578
rect 76972 20524 77028 20526
rect 78092 21980 78148 22036
rect 76636 19964 76692 20020
rect 77084 19964 77140 20020
rect 77420 19964 77476 20020
rect 76524 19292 76580 19348
rect 76524 18844 76580 18900
rect 76860 19234 76916 19236
rect 76860 19182 76862 19234
rect 76862 19182 76914 19234
rect 76914 19182 76916 19234
rect 76860 19180 76916 19182
rect 77644 19906 77700 19908
rect 77644 19854 77646 19906
rect 77646 19854 77698 19906
rect 77698 19854 77700 19906
rect 77644 19852 77700 19854
rect 77868 20748 77924 20804
rect 77532 19010 77588 19012
rect 77532 18958 77534 19010
rect 77534 18958 77586 19010
rect 77586 18958 77588 19010
rect 77532 18956 77588 18958
rect 77308 18620 77364 18676
rect 76972 18338 77028 18340
rect 76972 18286 76974 18338
rect 76974 18286 77026 18338
rect 77026 18286 77028 18338
rect 76972 18284 77028 18286
rect 77308 18284 77364 18340
rect 77644 17554 77700 17556
rect 77644 17502 77646 17554
rect 77646 17502 77698 17554
rect 77698 17502 77700 17554
rect 77644 17500 77700 17502
rect 77868 18396 77924 18452
rect 77644 16882 77700 16884
rect 77644 16830 77646 16882
rect 77646 16830 77698 16882
rect 77698 16830 77700 16882
rect 77644 16828 77700 16830
rect 77868 15986 77924 15988
rect 77868 15934 77870 15986
rect 77870 15934 77922 15986
rect 77922 15934 77924 15986
rect 77868 15932 77924 15934
rect 77644 15874 77700 15876
rect 77644 15822 77646 15874
rect 77646 15822 77698 15874
rect 77698 15822 77700 15874
rect 77644 15820 77700 15822
rect 77084 15148 77140 15204
rect 76860 14364 76916 14420
rect 76524 11506 76580 11508
rect 76524 11454 76526 11506
rect 76526 11454 76578 11506
rect 76578 11454 76580 11506
rect 76524 11452 76580 11454
rect 76972 10780 77028 10836
rect 76412 9324 76468 9380
rect 75964 7868 76020 7924
rect 76300 7420 76356 7476
rect 76188 6524 76244 6580
rect 76860 8258 76916 8260
rect 76860 8206 76862 8258
rect 76862 8206 76914 8258
rect 76914 8206 76916 8258
rect 76860 8204 76916 8206
rect 78540 22092 78596 22148
rect 78428 21644 78484 21700
rect 78204 20188 78260 20244
rect 78204 19740 78260 19796
rect 78204 18844 78260 18900
rect 78204 17554 78260 17556
rect 78204 17502 78206 17554
rect 78206 17502 78258 17554
rect 78258 17502 78260 17554
rect 78204 17500 78260 17502
rect 78204 16882 78260 16884
rect 78204 16830 78206 16882
rect 78206 16830 78258 16882
rect 78258 16830 78260 16882
rect 78204 16828 78260 16830
rect 78204 16380 78260 16436
rect 78204 15820 78260 15876
rect 78204 15260 78260 15316
rect 77868 14418 77924 14420
rect 77868 14366 77870 14418
rect 77870 14366 77922 14418
rect 77922 14366 77924 14418
rect 77868 14364 77924 14366
rect 77644 14140 77700 14196
rect 77868 13970 77924 13972
rect 77868 13918 77870 13970
rect 77870 13918 77922 13970
rect 77922 13918 77924 13970
rect 77868 13916 77924 13918
rect 77644 13634 77700 13636
rect 77644 13582 77646 13634
rect 77646 13582 77698 13634
rect 77698 13582 77700 13634
rect 77644 13580 77700 13582
rect 77756 12684 77812 12740
rect 78204 14140 78260 14196
rect 78204 13580 78260 13636
rect 78204 13020 78260 13076
rect 78204 11900 78260 11956
rect 78204 11452 78260 11508
rect 77532 10780 77588 10836
rect 77420 9996 77476 10052
rect 77644 9714 77700 9716
rect 77644 9662 77646 9714
rect 77646 9662 77698 9714
rect 77698 9662 77700 9714
rect 77644 9660 77700 9662
rect 77868 9602 77924 9604
rect 77868 9550 77870 9602
rect 77870 9550 77922 9602
rect 77922 9550 77924 9602
rect 77868 9548 77924 9550
rect 77868 9324 77924 9380
rect 76972 8092 77028 8148
rect 76860 7868 76916 7924
rect 76524 7196 76580 7252
rect 76300 5292 76356 5348
rect 76188 5180 76244 5236
rect 75740 5068 75796 5124
rect 76300 5122 76356 5124
rect 76300 5070 76302 5122
rect 76302 5070 76354 5122
rect 76354 5070 76356 5122
rect 76300 5068 76356 5070
rect 75628 4508 75684 4564
rect 76636 6636 76692 6692
rect 76748 6466 76804 6468
rect 76748 6414 76750 6466
rect 76750 6414 76802 6466
rect 76802 6414 76804 6466
rect 76748 6412 76804 6414
rect 76412 4508 76468 4564
rect 76972 4844 77028 4900
rect 77196 4508 77252 4564
rect 76188 3388 76244 3444
rect 77532 8146 77588 8148
rect 77532 8094 77534 8146
rect 77534 8094 77586 8146
rect 77586 8094 77588 8146
rect 77532 8092 77588 8094
rect 77420 7644 77476 7700
rect 77532 7420 77588 7476
rect 78204 9714 78260 9716
rect 78204 9662 78206 9714
rect 78206 9662 78258 9714
rect 78258 9662 78260 9714
rect 78204 9660 78260 9662
rect 78204 8540 78260 8596
rect 78092 8258 78148 8260
rect 78092 8206 78094 8258
rect 78094 8206 78146 8258
rect 78146 8206 78148 8258
rect 78092 8204 78148 8206
rect 77532 6748 77588 6804
rect 77644 5180 77700 5236
rect 77756 6412 77812 6468
rect 78316 6300 78372 6356
rect 78204 4562 78260 4564
rect 78204 4510 78206 4562
rect 78206 4510 78258 4562
rect 78258 4510 78260 4562
rect 78204 4508 78260 4510
rect 77868 3554 77924 3556
rect 77868 3502 77870 3554
rect 77870 3502 77922 3554
rect 77922 3502 77924 3554
rect 77868 3500 77924 3502
rect 78764 21644 78820 21700
rect 78652 9548 78708 9604
rect 75516 1820 75572 1876
<< metal3 >>
rect 79200 79156 80000 79184
rect 77298 79100 77308 79156
rect 77364 79100 80000 79156
rect 79200 79072 80000 79100
rect 79200 78036 80000 78064
rect 78754 77980 78764 78036
rect 78820 77980 80000 78036
rect 79200 77952 80000 77980
rect 0 77364 800 77392
rect 0 77308 2156 77364
rect 2212 77308 2222 77364
rect 0 77280 800 77308
rect 71698 77084 71708 77140
rect 71764 77084 73164 77140
rect 73220 77084 73230 77140
rect 73714 77084 73724 77140
rect 73780 77084 74508 77140
rect 74564 77084 75068 77140
rect 75124 77084 75134 77140
rect 61618 76972 61628 77028
rect 61684 76972 62860 77028
rect 62916 76972 62926 77028
rect 66994 76972 67004 77028
rect 67060 76972 67788 77028
rect 67844 76972 67854 77028
rect 69682 76972 69692 77028
rect 69748 76972 70924 77028
rect 70980 76972 70990 77028
rect 73042 76972 73052 77028
rect 73108 76972 74284 77028
rect 74340 76972 74350 77028
rect 79200 76916 80000 76944
rect 61954 76860 61964 76916
rect 62020 76860 77196 76916
rect 77252 76860 77262 76916
rect 77420 76860 80000 76916
rect 19826 76804 19836 76860
rect 19892 76804 19940 76860
rect 19996 76804 20044 76860
rect 20100 76804 20110 76860
rect 50546 76804 50556 76860
rect 50612 76804 50660 76860
rect 50716 76804 50764 76860
rect 50820 76804 50830 76860
rect 77420 76804 77476 76860
rect 79200 76832 80000 76860
rect 58034 76748 58044 76804
rect 58100 76748 76076 76804
rect 76132 76748 76142 76804
rect 76962 76748 76972 76804
rect 77028 76748 77476 76804
rect 15362 76636 15372 76692
rect 15428 76636 16604 76692
rect 16660 76636 16670 76692
rect 21074 76636 21084 76692
rect 21140 76636 21980 76692
rect 22036 76636 22046 76692
rect 41010 76636 41020 76692
rect 41076 76636 42028 76692
rect 42084 76636 42094 76692
rect 44146 76636 44156 76692
rect 44212 76636 45836 76692
rect 45892 76636 45902 76692
rect 46162 76636 46172 76692
rect 46228 76636 47852 76692
rect 47908 76636 47918 76692
rect 48178 76636 48188 76692
rect 48244 76636 49196 76692
rect 49252 76636 49262 76692
rect 50194 76636 50204 76692
rect 50260 76636 51212 76692
rect 51268 76636 51278 76692
rect 52882 76636 52892 76692
rect 52948 76636 53900 76692
rect 53956 76636 55132 76692
rect 55188 76636 55198 76692
rect 56914 76636 56924 76692
rect 56980 76636 59836 76692
rect 59892 76636 59902 76692
rect 62962 76636 62972 76692
rect 63028 76636 63980 76692
rect 64036 76636 64046 76692
rect 68338 76636 68348 76692
rect 68404 76636 69356 76692
rect 69412 76636 69422 76692
rect 74610 76636 74620 76692
rect 74676 76636 77308 76692
rect 77364 76636 77374 76692
rect 54898 76524 54908 76580
rect 54964 76524 55580 76580
rect 55636 76524 55646 76580
rect 70354 76524 70364 76580
rect 70420 76524 71596 76580
rect 71652 76524 71662 76580
rect 73154 76524 73164 76580
rect 73220 76524 74060 76580
rect 74116 76524 74126 76580
rect 18050 76412 18060 76468
rect 18116 76412 19404 76468
rect 19460 76412 19470 76468
rect 57586 76412 57596 76468
rect 57652 76412 58828 76468
rect 58884 76412 58894 76468
rect 59602 76412 59612 76468
rect 59668 76412 62076 76468
rect 62132 76412 62748 76468
rect 62804 76412 62814 76468
rect 76290 76412 76300 76468
rect 76356 76412 77084 76468
rect 77140 76412 77868 76468
rect 77924 76412 77934 76468
rect 12450 76300 12460 76356
rect 12516 76300 13356 76356
rect 13412 76300 14140 76356
rect 14196 76300 14206 76356
rect 16370 76300 16380 76356
rect 16436 76300 17164 76356
rect 17220 76300 20748 76356
rect 20804 76300 20814 76356
rect 47366 76300 47404 76356
rect 47460 76300 47470 76356
rect 48626 76300 48636 76356
rect 48692 76300 50540 76356
rect 50596 76300 50606 76356
rect 62132 76300 76748 76356
rect 76804 76300 76814 76356
rect 0 76244 800 76272
rect 62132 76244 62188 76300
rect 0 76188 1932 76244
rect 1988 76188 1998 76244
rect 49970 76188 49980 76244
rect 50036 76188 62188 76244
rect 0 76160 800 76188
rect 67172 76076 78204 76132
rect 78260 76076 78270 76132
rect 4466 76020 4476 76076
rect 4532 76020 4580 76076
rect 4636 76020 4684 76076
rect 4740 76020 4750 76076
rect 35186 76020 35196 76076
rect 35252 76020 35300 76076
rect 35356 76020 35404 76076
rect 35460 76020 35470 76076
rect 65906 76020 65916 76076
rect 65972 76020 66020 76076
rect 66076 76020 66124 76076
rect 66180 76020 66190 76076
rect 11890 75852 11900 75908
rect 11956 75852 12572 75908
rect 12628 75852 12638 75908
rect 20626 75852 20636 75908
rect 20692 75852 21980 75908
rect 22036 75852 22046 75908
rect 34962 75852 34972 75908
rect 35028 75852 37996 75908
rect 38052 75852 38062 75908
rect 33618 75740 33628 75796
rect 33684 75740 35196 75796
rect 35252 75740 35262 75796
rect 50082 75740 50092 75796
rect 50148 75740 50764 75796
rect 50820 75740 50830 75796
rect 65314 75740 65324 75796
rect 65380 75740 65996 75796
rect 66052 75740 66062 75796
rect 67172 75684 67228 76076
rect 79200 75796 80000 75824
rect 78988 75740 80000 75796
rect 12562 75628 12572 75684
rect 12628 75628 13580 75684
rect 13636 75628 13646 75684
rect 14690 75628 14700 75684
rect 14756 75628 16492 75684
rect 16548 75628 16558 75684
rect 23762 75628 23772 75684
rect 23828 75628 25228 75684
rect 25284 75628 25900 75684
rect 25956 75628 25966 75684
rect 30146 75628 30156 75684
rect 30212 75628 33516 75684
rect 33572 75628 33582 75684
rect 34738 75628 34748 75684
rect 34804 75628 35532 75684
rect 35588 75628 35598 75684
rect 40114 75628 40124 75684
rect 40180 75628 40908 75684
rect 40964 75628 40974 75684
rect 47170 75628 47180 75684
rect 47236 75628 47628 75684
rect 47684 75628 47694 75684
rect 50306 75628 50316 75684
rect 50372 75628 55916 75684
rect 55972 75628 55982 75684
rect 57026 75628 57036 75684
rect 57092 75628 61740 75684
rect 61796 75628 61806 75684
rect 63756 75628 67228 75684
rect 68674 75628 68684 75684
rect 68740 75628 75628 75684
rect 75684 75628 75694 75684
rect 76486 75628 76524 75684
rect 76580 75628 76590 75684
rect 63756 75572 63812 75628
rect 11554 75516 11564 75572
rect 11620 75516 13916 75572
rect 13972 75516 13982 75572
rect 17938 75516 17948 75572
rect 18004 75516 19180 75572
rect 19236 75516 19246 75572
rect 60274 75516 60284 75572
rect 60340 75516 61180 75572
rect 61236 75516 61516 75572
rect 61572 75516 61582 75572
rect 63746 75516 63756 75572
rect 63812 75516 63822 75572
rect 75394 75516 75404 75572
rect 75460 75516 76076 75572
rect 76132 75516 78652 75572
rect 78708 75516 78718 75572
rect 78988 75460 79044 75740
rect 79200 75712 80000 75740
rect 58146 75404 58156 75460
rect 58212 75404 59388 75460
rect 59444 75404 59454 75460
rect 61058 75404 61068 75460
rect 61124 75404 62076 75460
rect 62132 75404 62142 75460
rect 65538 75404 65548 75460
rect 65604 75404 66892 75460
rect 66948 75404 66958 75460
rect 74050 75404 74060 75460
rect 74116 75404 78092 75460
rect 78148 75404 79044 75460
rect 1922 75292 1932 75348
rect 1988 75292 1998 75348
rect 58930 75292 58940 75348
rect 58996 75292 60508 75348
rect 60564 75292 61292 75348
rect 61348 75292 61358 75348
rect 0 75124 800 75152
rect 1932 75124 1988 75292
rect 19826 75236 19836 75292
rect 19892 75236 19940 75292
rect 19996 75236 20044 75292
rect 20100 75236 20110 75292
rect 50546 75236 50556 75292
rect 50612 75236 50660 75292
rect 50716 75236 50764 75292
rect 50820 75236 50830 75292
rect 0 75068 1988 75124
rect 36866 75068 36876 75124
rect 36932 75068 37660 75124
rect 37716 75068 37726 75124
rect 74946 75068 74956 75124
rect 75012 75068 76188 75124
rect 76244 75068 76254 75124
rect 77522 75068 77532 75124
rect 77588 75068 78204 75124
rect 78260 75068 78764 75124
rect 78820 75068 78830 75124
rect 0 75040 800 75068
rect 75394 74956 75404 75012
rect 75460 74956 75964 75012
rect 76020 74956 79100 75012
rect 79156 74956 79166 75012
rect 11666 74844 11676 74900
rect 11732 74844 13468 74900
rect 13524 74844 14252 74900
rect 14308 74844 14318 74900
rect 18834 74732 18844 74788
rect 18900 74732 19852 74788
rect 19908 74732 20300 74788
rect 20356 74732 20366 74788
rect 31042 74732 31052 74788
rect 31108 74732 35084 74788
rect 35140 74732 35150 74788
rect 79200 74676 80000 74704
rect 78306 74620 78316 74676
rect 78372 74620 80000 74676
rect 79200 74592 80000 74620
rect 4466 74452 4476 74508
rect 4532 74452 4580 74508
rect 4636 74452 4684 74508
rect 4740 74452 4750 74508
rect 35186 74452 35196 74508
rect 35252 74452 35300 74508
rect 35356 74452 35404 74508
rect 35460 74452 35470 74508
rect 65906 74452 65916 74508
rect 65972 74452 66020 74508
rect 66076 74452 66124 74508
rect 66180 74452 66190 74508
rect 1922 74172 1932 74228
rect 1988 74172 1998 74228
rect 0 74004 800 74032
rect 1932 74004 1988 74172
rect 70466 74060 70476 74116
rect 70532 74060 73948 74116
rect 75282 74060 75292 74116
rect 75348 74060 78092 74116
rect 78148 74060 78484 74116
rect 73892 74004 73948 74060
rect 0 73948 1988 74004
rect 12674 73948 12684 74004
rect 12740 73948 14364 74004
rect 14420 73948 14430 74004
rect 18274 73948 18284 74004
rect 18340 73948 20860 74004
rect 20916 73948 20926 74004
rect 73892 73948 77868 74004
rect 77924 73948 77934 74004
rect 0 73920 800 73948
rect 19826 73668 19836 73724
rect 19892 73668 19940 73724
rect 19996 73668 20044 73724
rect 20100 73668 20110 73724
rect 50546 73668 50556 73724
rect 50612 73668 50660 73724
rect 50716 73668 50764 73724
rect 50820 73668 50830 73724
rect 78428 73556 78484 74060
rect 79200 73556 80000 73584
rect 77634 73500 77644 73556
rect 77700 73500 78204 73556
rect 78260 73500 78270 73556
rect 78428 73500 80000 73556
rect 79200 73472 80000 73500
rect 17826 73388 17836 73444
rect 17892 73388 18172 73444
rect 18228 73388 18238 73444
rect 65314 73388 65324 73444
rect 65380 73388 77868 73444
rect 77924 73388 77934 73444
rect 14018 73276 14028 73332
rect 14084 73276 16268 73332
rect 16324 73276 16334 73332
rect 17602 73164 17612 73220
rect 17668 73164 18060 73220
rect 18116 73164 18126 73220
rect 1922 73052 1932 73108
rect 1988 73052 1998 73108
rect 0 72884 800 72912
rect 1932 72884 1988 73052
rect 4466 72884 4476 72940
rect 4532 72884 4580 72940
rect 4636 72884 4684 72940
rect 4740 72884 4750 72940
rect 35186 72884 35196 72940
rect 35252 72884 35300 72940
rect 35356 72884 35404 72940
rect 35460 72884 35470 72940
rect 65906 72884 65916 72940
rect 65972 72884 66020 72940
rect 66076 72884 66124 72940
rect 66180 72884 66190 72940
rect 0 72828 1988 72884
rect 0 72800 800 72828
rect 79200 72436 80000 72464
rect 76738 72380 76748 72436
rect 76804 72380 77252 72436
rect 77634 72380 77644 72436
rect 77700 72380 78204 72436
rect 78260 72380 80000 72436
rect 77196 72324 77252 72380
rect 79200 72352 80000 72380
rect 74834 72268 74844 72324
rect 74900 72268 76972 72324
rect 77028 72268 77038 72324
rect 77196 72268 77868 72324
rect 77924 72268 77934 72324
rect 19826 72100 19836 72156
rect 19892 72100 19940 72156
rect 19996 72100 20044 72156
rect 20100 72100 20110 72156
rect 50546 72100 50556 72156
rect 50612 72100 50660 72156
rect 50716 72100 50764 72156
rect 50820 72100 50830 72156
rect 1922 71932 1932 71988
rect 1988 71932 1998 71988
rect 3154 71932 3164 71988
rect 3220 71932 3948 71988
rect 4004 71932 4014 71988
rect 0 71764 800 71792
rect 1932 71764 1988 71932
rect 2482 71820 2492 71876
rect 2548 71820 2940 71876
rect 2996 71820 4508 71876
rect 4564 71820 5740 71876
rect 5796 71820 5806 71876
rect 68562 71820 68572 71876
rect 68628 71820 77868 71876
rect 77924 71820 77934 71876
rect 0 71708 1988 71764
rect 0 71680 800 71708
rect 54450 71484 54460 71540
rect 54516 71484 55244 71540
rect 55300 71484 55310 71540
rect 4466 71316 4476 71372
rect 4532 71316 4580 71372
rect 4636 71316 4684 71372
rect 4740 71316 4750 71372
rect 35186 71316 35196 71372
rect 35252 71316 35300 71372
rect 35356 71316 35404 71372
rect 35460 71316 35470 71372
rect 65906 71316 65916 71372
rect 65972 71316 66020 71372
rect 66076 71316 66124 71372
rect 66180 71316 66190 71372
rect 79200 71316 80000 71344
rect 77634 71260 77644 71316
rect 77700 71260 78204 71316
rect 78260 71260 80000 71316
rect 79200 71232 80000 71260
rect 77634 70924 77644 70980
rect 77700 70924 78764 70980
rect 78820 70924 78830 70980
rect 77410 70700 77420 70756
rect 77476 70700 78204 70756
rect 78260 70700 78270 70756
rect 0 70644 800 70672
rect 0 70588 1932 70644
rect 1988 70588 1998 70644
rect 0 70560 800 70588
rect 19826 70532 19836 70588
rect 19892 70532 19940 70588
rect 19996 70532 20044 70588
rect 20100 70532 20110 70588
rect 50546 70532 50556 70588
rect 50612 70532 50660 70588
rect 50716 70532 50764 70588
rect 50820 70532 50830 70588
rect 79200 70196 80000 70224
rect 2706 70140 2716 70196
rect 2772 70140 3836 70196
rect 3892 70140 3902 70196
rect 78194 70140 78204 70196
rect 78260 70140 80000 70196
rect 79200 70112 80000 70140
rect 4466 69748 4476 69804
rect 4532 69748 4580 69804
rect 4636 69748 4684 69804
rect 4740 69748 4750 69804
rect 35186 69748 35196 69804
rect 35252 69748 35300 69804
rect 35356 69748 35404 69804
rect 35460 69748 35470 69804
rect 65906 69748 65916 69804
rect 65972 69748 66020 69804
rect 66076 69748 66124 69804
rect 66180 69748 66190 69804
rect 0 69524 800 69552
rect 0 69468 1932 69524
rect 1988 69468 1998 69524
rect 0 69440 800 69468
rect 76738 69132 76748 69188
rect 76804 69132 77868 69188
rect 77924 69132 77934 69188
rect 79200 69076 80000 69104
rect 77634 69020 77644 69076
rect 77700 69020 78204 69076
rect 78260 69020 80000 69076
rect 19826 68964 19836 69020
rect 19892 68964 19940 69020
rect 19996 68964 20044 69020
rect 20100 68964 20110 69020
rect 50546 68964 50556 69020
rect 50612 68964 50660 69020
rect 50716 68964 50764 69020
rect 50820 68964 50830 69020
rect 79200 68992 80000 69020
rect 73938 68796 73948 68852
rect 74004 68796 75628 68852
rect 75684 68796 75694 68852
rect 72146 68684 72156 68740
rect 72212 68684 75180 68740
rect 75236 68684 75246 68740
rect 77410 68572 77420 68628
rect 77476 68572 78204 68628
rect 78260 68572 78270 68628
rect 76850 68460 76860 68516
rect 76916 68460 77644 68516
rect 77700 68460 77710 68516
rect 0 68404 800 68432
rect 0 68348 2716 68404
rect 2772 68348 2782 68404
rect 0 68320 800 68348
rect 4466 68180 4476 68236
rect 4532 68180 4580 68236
rect 4636 68180 4684 68236
rect 4740 68180 4750 68236
rect 35186 68180 35196 68236
rect 35252 68180 35300 68236
rect 35356 68180 35404 68236
rect 35460 68180 35470 68236
rect 65906 68180 65916 68236
rect 65972 68180 66020 68236
rect 66076 68180 66124 68236
rect 66180 68180 66190 68236
rect 79200 67956 80000 67984
rect 78194 67900 78204 67956
rect 78260 67900 80000 67956
rect 79200 67872 80000 67900
rect 19826 67396 19836 67452
rect 19892 67396 19940 67452
rect 19996 67396 20044 67452
rect 20100 67396 20110 67452
rect 50546 67396 50556 67452
rect 50612 67396 50660 67452
rect 50716 67396 50764 67452
rect 50820 67396 50830 67452
rect 0 67284 800 67312
rect 0 67228 1932 67284
rect 1988 67228 1998 67284
rect 60946 67228 60956 67284
rect 61012 67228 61292 67284
rect 61348 67228 61358 67284
rect 64866 67228 64876 67284
rect 64932 67228 65212 67284
rect 65268 67228 65278 67284
rect 70578 67228 70588 67284
rect 70644 67228 71148 67284
rect 71204 67228 71214 67284
rect 0 67200 800 67228
rect 2370 67116 2380 67172
rect 2436 67116 3052 67172
rect 3108 67116 3118 67172
rect 79200 66836 80000 66864
rect 77634 66780 77644 66836
rect 77700 66780 78204 66836
rect 78260 66780 80000 66836
rect 79200 66752 80000 66780
rect 4466 66612 4476 66668
rect 4532 66612 4580 66668
rect 4636 66612 4684 66668
rect 4740 66612 4750 66668
rect 35186 66612 35196 66668
rect 35252 66612 35300 66668
rect 35356 66612 35404 66668
rect 35460 66612 35470 66668
rect 65906 66612 65916 66668
rect 65972 66612 66020 66668
rect 66076 66612 66124 66668
rect 66180 66612 66190 66668
rect 0 66164 800 66192
rect 0 66108 2772 66164
rect 0 66080 800 66108
rect 2716 66052 2772 66108
rect 2706 65996 2716 66052
rect 2772 65996 2782 66052
rect 76626 65996 76636 66052
rect 76692 65996 77868 66052
rect 77924 65996 77934 66052
rect 19826 65828 19836 65884
rect 19892 65828 19940 65884
rect 19996 65828 20044 65884
rect 20100 65828 20110 65884
rect 50546 65828 50556 65884
rect 50612 65828 50660 65884
rect 50716 65828 50764 65884
rect 50820 65828 50830 65884
rect 79200 65716 80000 65744
rect 77634 65660 77644 65716
rect 77700 65660 78204 65716
rect 78260 65660 80000 65716
rect 79200 65632 80000 65660
rect 1922 65212 1932 65268
rect 1988 65212 1998 65268
rect 0 65044 800 65072
rect 1932 65044 1988 65212
rect 4466 65044 4476 65100
rect 4532 65044 4580 65100
rect 4636 65044 4684 65100
rect 4740 65044 4750 65100
rect 35186 65044 35196 65100
rect 35252 65044 35300 65100
rect 35356 65044 35404 65100
rect 35460 65044 35470 65100
rect 65906 65044 65916 65100
rect 65972 65044 66020 65100
rect 66076 65044 66124 65100
rect 66180 65044 66190 65100
rect 0 64988 1988 65044
rect 0 64960 800 64988
rect 77074 64652 77084 64708
rect 77140 64652 77644 64708
rect 77700 64652 77710 64708
rect 79200 64596 80000 64624
rect 3602 64540 3612 64596
rect 3668 64540 4956 64596
rect 5012 64540 5022 64596
rect 77410 64540 77420 64596
rect 77476 64540 78204 64596
rect 78260 64540 80000 64596
rect 79200 64512 80000 64540
rect 19826 64260 19836 64316
rect 19892 64260 19940 64316
rect 19996 64260 20044 64316
rect 20100 64260 20110 64316
rect 50546 64260 50556 64316
rect 50612 64260 50660 64316
rect 50716 64260 50764 64316
rect 50820 64260 50830 64316
rect 76402 63980 76412 64036
rect 76468 63980 77644 64036
rect 77700 63980 77710 64036
rect 0 63924 800 63952
rect 0 63868 1932 63924
rect 1988 63868 1998 63924
rect 2482 63868 2492 63924
rect 2548 63868 2940 63924
rect 2996 63868 3612 63924
rect 3668 63868 3678 63924
rect 77410 63868 77420 63924
rect 77476 63868 78204 63924
rect 78260 63868 78270 63924
rect 0 63840 800 63868
rect 4466 63476 4476 63532
rect 4532 63476 4580 63532
rect 4636 63476 4684 63532
rect 4740 63476 4750 63532
rect 35186 63476 35196 63532
rect 35252 63476 35300 63532
rect 35356 63476 35404 63532
rect 35460 63476 35470 63532
rect 65906 63476 65916 63532
rect 65972 63476 66020 63532
rect 66076 63476 66124 63532
rect 66180 63476 66190 63532
rect 79200 63476 80000 63504
rect 78194 63420 78204 63476
rect 78260 63420 80000 63476
rect 79200 63392 80000 63420
rect 77634 62860 77644 62916
rect 77700 62860 78204 62916
rect 78260 62860 78270 62916
rect 0 62804 800 62832
rect 0 62748 1932 62804
rect 1988 62748 1998 62804
rect 0 62720 800 62748
rect 19826 62692 19836 62748
rect 19892 62692 19940 62748
rect 19996 62692 20044 62748
rect 20100 62692 20110 62748
rect 50546 62692 50556 62748
rect 50612 62692 50660 62748
rect 50716 62692 50764 62748
rect 50820 62692 50830 62748
rect 79200 62356 80000 62384
rect 78194 62300 78204 62356
rect 78260 62300 80000 62356
rect 79200 62272 80000 62300
rect 76178 62188 76188 62244
rect 76244 62188 77868 62244
rect 77924 62188 77934 62244
rect 72706 62076 72716 62132
rect 72772 62076 73052 62132
rect 73108 62076 73118 62132
rect 4466 61908 4476 61964
rect 4532 61908 4580 61964
rect 4636 61908 4684 61964
rect 4740 61908 4750 61964
rect 35186 61908 35196 61964
rect 35252 61908 35300 61964
rect 35356 61908 35404 61964
rect 35460 61908 35470 61964
rect 65906 61908 65916 61964
rect 65972 61908 66020 61964
rect 66076 61908 66124 61964
rect 66180 61908 66190 61964
rect 0 61684 800 61712
rect 0 61628 1932 61684
rect 1988 61628 1998 61684
rect 0 61600 800 61628
rect 2930 61516 2940 61572
rect 2996 61516 3612 61572
rect 3668 61516 3678 61572
rect 75394 61516 75404 61572
rect 75460 61516 77644 61572
rect 77700 61516 77710 61572
rect 3042 61292 3052 61348
rect 3108 61292 4172 61348
rect 4228 61292 4238 61348
rect 79200 61236 80000 61264
rect 77410 61180 77420 61236
rect 77476 61180 78204 61236
rect 78260 61180 80000 61236
rect 19826 61124 19836 61180
rect 19892 61124 19940 61180
rect 19996 61124 20044 61180
rect 20100 61124 20110 61180
rect 50546 61124 50556 61180
rect 50612 61124 50660 61180
rect 50716 61124 50764 61180
rect 50820 61124 50830 61180
rect 79200 61152 80000 61180
rect 76290 60844 76300 60900
rect 76356 60844 77868 60900
rect 77924 60844 77934 60900
rect 77634 60732 77644 60788
rect 77700 60732 78204 60788
rect 78260 60732 78270 60788
rect 0 60564 800 60592
rect 0 60508 2716 60564
rect 2772 60508 2782 60564
rect 0 60480 800 60508
rect 4466 60340 4476 60396
rect 4532 60340 4580 60396
rect 4636 60340 4684 60396
rect 4740 60340 4750 60396
rect 35186 60340 35196 60396
rect 35252 60340 35300 60396
rect 35356 60340 35404 60396
rect 35460 60340 35470 60396
rect 65906 60340 65916 60396
rect 65972 60340 66020 60396
rect 66076 60340 66124 60396
rect 66180 60340 66190 60396
rect 79200 60116 80000 60144
rect 78194 60060 78204 60116
rect 78260 60060 80000 60116
rect 79200 60032 80000 60060
rect 2706 59948 2716 60004
rect 2772 59948 3836 60004
rect 3892 59948 3902 60004
rect 19826 59556 19836 59612
rect 19892 59556 19940 59612
rect 19996 59556 20044 59612
rect 20100 59556 20110 59612
rect 50546 59556 50556 59612
rect 50612 59556 50660 59612
rect 50716 59556 50764 59612
rect 50820 59556 50830 59612
rect 0 59444 800 59472
rect 0 59388 1932 59444
rect 1988 59388 1998 59444
rect 0 59360 800 59388
rect 2146 59164 2156 59220
rect 2212 59164 2940 59220
rect 2996 59164 3500 59220
rect 3556 59164 3566 59220
rect 74946 59052 74956 59108
rect 75012 59052 77644 59108
rect 77700 59052 77710 59108
rect 79200 58996 80000 59024
rect 77410 58940 77420 58996
rect 77476 58940 78204 58996
rect 78260 58940 80000 58996
rect 79200 58912 80000 58940
rect 68114 58828 68124 58884
rect 68180 58828 69916 58884
rect 69972 58828 69982 58884
rect 4466 58772 4476 58828
rect 4532 58772 4580 58828
rect 4636 58772 4684 58828
rect 4740 58772 4750 58828
rect 35186 58772 35196 58828
rect 35252 58772 35300 58828
rect 35356 58772 35404 58828
rect 35460 58772 35470 58828
rect 65906 58772 65916 58828
rect 65972 58772 66020 58828
rect 66076 58772 66124 58828
rect 66180 58772 66190 58828
rect 0 58324 800 58352
rect 0 58268 2772 58324
rect 0 58240 800 58268
rect 2716 58212 2772 58268
rect 2706 58156 2716 58212
rect 2772 58156 2782 58212
rect 61842 58156 61852 58212
rect 61908 58156 77868 58212
rect 77924 58156 77934 58212
rect 19826 57988 19836 58044
rect 19892 57988 19940 58044
rect 19996 57988 20044 58044
rect 20100 57988 20110 58044
rect 50546 57988 50556 58044
rect 50612 57988 50660 58044
rect 50716 57988 50764 58044
rect 50820 57988 50830 58044
rect 79200 57876 80000 57904
rect 77634 57820 77644 57876
rect 77700 57820 78204 57876
rect 78260 57820 80000 57876
rect 79200 57792 80000 57820
rect 1922 57372 1932 57428
rect 1988 57372 1998 57428
rect 0 57204 800 57232
rect 1932 57204 1988 57372
rect 4466 57204 4476 57260
rect 4532 57204 4580 57260
rect 4636 57204 4684 57260
rect 4740 57204 4750 57260
rect 35186 57204 35196 57260
rect 35252 57204 35300 57260
rect 35356 57204 35404 57260
rect 35460 57204 35470 57260
rect 65906 57204 65916 57260
rect 65972 57204 66020 57260
rect 66076 57204 66124 57260
rect 66180 57204 66190 57260
rect 0 57148 1988 57204
rect 0 57120 800 57148
rect 79200 56756 80000 56784
rect 77634 56700 77644 56756
rect 77700 56700 78204 56756
rect 78260 56700 80000 56756
rect 79200 56672 80000 56700
rect 19826 56420 19836 56476
rect 19892 56420 19940 56476
rect 19996 56420 20044 56476
rect 20100 56420 20110 56476
rect 50546 56420 50556 56476
rect 50612 56420 50660 56476
rect 50716 56420 50764 56476
rect 50820 56420 50830 56476
rect 2706 56140 2716 56196
rect 2772 56140 3388 56196
rect 3444 56140 4844 56196
rect 4900 56140 4910 56196
rect 65202 56140 65212 56196
rect 65268 56140 77868 56196
rect 77924 56140 77934 56196
rect 0 56084 800 56112
rect 0 56028 1932 56084
rect 1988 56028 1998 56084
rect 0 56000 800 56028
rect 4466 55636 4476 55692
rect 4532 55636 4580 55692
rect 4636 55636 4684 55692
rect 4740 55636 4750 55692
rect 35186 55636 35196 55692
rect 35252 55636 35300 55692
rect 35356 55636 35404 55692
rect 35460 55636 35470 55692
rect 65906 55636 65916 55692
rect 65972 55636 66020 55692
rect 66076 55636 66124 55692
rect 66180 55636 66190 55692
rect 79200 55636 80000 55664
rect 77634 55580 77644 55636
rect 77700 55580 78204 55636
rect 78260 55580 80000 55636
rect 79200 55552 80000 55580
rect 2706 55020 2716 55076
rect 2772 55020 2782 55076
rect 77634 55020 77644 55076
rect 77700 55020 78204 55076
rect 78260 55020 78270 55076
rect 0 54964 800 54992
rect 2716 54964 2772 55020
rect 0 54908 2772 54964
rect 0 54880 800 54908
rect 19826 54852 19836 54908
rect 19892 54852 19940 54908
rect 19996 54852 20044 54908
rect 20100 54852 20110 54908
rect 50546 54852 50556 54908
rect 50612 54852 50660 54908
rect 50716 54852 50764 54908
rect 50820 54852 50830 54908
rect 79200 54516 80000 54544
rect 78194 54460 78204 54516
rect 78260 54460 80000 54516
rect 79200 54432 80000 54460
rect 4466 54068 4476 54124
rect 4532 54068 4580 54124
rect 4636 54068 4684 54124
rect 4740 54068 4750 54124
rect 35186 54068 35196 54124
rect 35252 54068 35300 54124
rect 35356 54068 35404 54124
rect 35460 54068 35470 54124
rect 65906 54068 65916 54124
rect 65972 54068 66020 54124
rect 66076 54068 66124 54124
rect 66180 54068 66190 54124
rect 72594 54012 72604 54068
rect 72660 54012 77868 54068
rect 77924 54012 77934 54068
rect 0 53844 800 53872
rect 0 53788 1932 53844
rect 1988 53788 1998 53844
rect 58594 53788 58604 53844
rect 58660 53788 77868 53844
rect 77924 53788 77934 53844
rect 0 53760 800 53788
rect 3154 53564 3164 53620
rect 3220 53564 3948 53620
rect 4004 53564 4014 53620
rect 2482 53452 2492 53508
rect 2548 53452 2940 53508
rect 2996 53452 3836 53508
rect 3892 53452 3902 53508
rect 79200 53396 80000 53424
rect 77634 53340 77644 53396
rect 77700 53340 78204 53396
rect 78260 53340 80000 53396
rect 19826 53284 19836 53340
rect 19892 53284 19940 53340
rect 19996 53284 20044 53340
rect 20100 53284 20110 53340
rect 50546 53284 50556 53340
rect 50612 53284 50660 53340
rect 50716 53284 50764 53340
rect 50820 53284 50830 53340
rect 79200 53312 80000 53340
rect 77634 52780 77644 52836
rect 77700 52780 78204 52836
rect 78260 52780 78270 52836
rect 0 52724 800 52752
rect 0 52668 1932 52724
rect 1988 52668 1998 52724
rect 0 52640 800 52668
rect 4466 52500 4476 52556
rect 4532 52500 4580 52556
rect 4636 52500 4684 52556
rect 4740 52500 4750 52556
rect 35186 52500 35196 52556
rect 35252 52500 35300 52556
rect 35356 52500 35404 52556
rect 35460 52500 35470 52556
rect 65906 52500 65916 52556
rect 65972 52500 66020 52556
rect 66076 52500 66124 52556
rect 66180 52500 66190 52556
rect 79200 52276 80000 52304
rect 78194 52220 78204 52276
rect 78260 52220 80000 52276
rect 79200 52192 80000 52220
rect 19826 51716 19836 51772
rect 19892 51716 19940 51772
rect 19996 51716 20044 51772
rect 20100 51716 20110 51772
rect 50546 51716 50556 51772
rect 50612 51716 50660 51772
rect 50716 51716 50764 51772
rect 50820 51716 50830 51772
rect 0 51604 800 51632
rect 0 51548 1932 51604
rect 1988 51548 1998 51604
rect 0 51520 800 51548
rect 72034 51436 72044 51492
rect 72100 51436 77868 51492
rect 77924 51436 77934 51492
rect 79200 51156 80000 51184
rect 77634 51100 77644 51156
rect 77700 51100 78204 51156
rect 78260 51100 80000 51156
rect 79200 51072 80000 51100
rect 4466 50932 4476 50988
rect 4532 50932 4580 50988
rect 4636 50932 4684 50988
rect 4740 50932 4750 50988
rect 35186 50932 35196 50988
rect 35252 50932 35300 50988
rect 35356 50932 35404 50988
rect 35460 50932 35470 50988
rect 65906 50932 65916 50988
rect 65972 50932 66020 50988
rect 66076 50932 66124 50988
rect 66180 50932 66190 50988
rect 1922 50652 1932 50708
rect 1988 50652 1998 50708
rect 0 50484 800 50512
rect 1932 50484 1988 50652
rect 2818 50540 2828 50596
rect 2884 50540 3836 50596
rect 3892 50540 3902 50596
rect 0 50428 1988 50484
rect 77634 50428 77644 50484
rect 77700 50428 78204 50484
rect 78260 50428 78270 50484
rect 0 50400 800 50428
rect 77298 50316 77308 50372
rect 77364 50316 77868 50372
rect 77924 50316 77934 50372
rect 19826 50148 19836 50204
rect 19892 50148 19940 50204
rect 19996 50148 20044 50204
rect 20100 50148 20110 50204
rect 50546 50148 50556 50204
rect 50612 50148 50660 50204
rect 50716 50148 50764 50204
rect 50820 50148 50830 50204
rect 79200 50036 80000 50064
rect 78194 49980 78204 50036
rect 78260 49980 80000 50036
rect 79200 49952 80000 49980
rect 1922 49532 1932 49588
rect 1988 49532 1998 49588
rect 3154 49532 3164 49588
rect 3220 49532 3612 49588
rect 3668 49532 3678 49588
rect 0 49364 800 49392
rect 1932 49364 1988 49532
rect 4466 49364 4476 49420
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4740 49364 4750 49420
rect 35186 49364 35196 49420
rect 35252 49364 35300 49420
rect 35356 49364 35404 49420
rect 35460 49364 35470 49420
rect 65906 49364 65916 49420
rect 65972 49364 66020 49420
rect 66076 49364 66124 49420
rect 66180 49364 66190 49420
rect 0 49308 1988 49364
rect 0 49280 800 49308
rect 2706 48972 2716 49028
rect 2772 48972 3836 49028
rect 3892 48972 3902 49028
rect 79200 48916 80000 48944
rect 77634 48860 77644 48916
rect 77700 48860 78204 48916
rect 78260 48860 80000 48916
rect 79200 48832 80000 48860
rect 19826 48580 19836 48636
rect 19892 48580 19940 48636
rect 19996 48580 20044 48636
rect 20100 48580 20110 48636
rect 50546 48580 50556 48636
rect 50612 48580 50660 48636
rect 50716 48580 50764 48636
rect 50820 48580 50830 48636
rect 77858 48300 77868 48356
rect 77924 48300 78540 48356
rect 78596 48300 78606 48356
rect 0 48244 800 48272
rect 0 48188 1932 48244
rect 1988 48188 1998 48244
rect 0 48160 800 48188
rect 4466 47796 4476 47852
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4740 47796 4750 47852
rect 35186 47796 35196 47852
rect 35252 47796 35300 47852
rect 35356 47796 35404 47852
rect 35460 47796 35470 47852
rect 65906 47796 65916 47852
rect 65972 47796 66020 47852
rect 66076 47796 66124 47852
rect 66180 47796 66190 47852
rect 79200 47796 80000 47824
rect 77634 47740 77644 47796
rect 77700 47740 78204 47796
rect 78260 47740 80000 47796
rect 79200 47712 80000 47740
rect 77634 47292 77644 47348
rect 77700 47292 78204 47348
rect 78260 47292 78270 47348
rect 2706 47180 2716 47236
rect 2772 47180 2782 47236
rect 77858 47180 77868 47236
rect 77924 47180 78764 47236
rect 78820 47180 78830 47236
rect 0 47124 800 47152
rect 2716 47124 2772 47180
rect 0 47068 2772 47124
rect 0 47040 800 47068
rect 19826 47012 19836 47068
rect 19892 47012 19940 47068
rect 19996 47012 20044 47068
rect 20100 47012 20110 47068
rect 50546 47012 50556 47068
rect 50612 47012 50660 47068
rect 50716 47012 50764 47068
rect 50820 47012 50830 47068
rect 57026 46956 57036 47012
rect 57092 46956 62188 47012
rect 62244 46956 62254 47012
rect 74722 46956 74732 47012
rect 74788 46956 78092 47012
rect 78148 46956 78158 47012
rect 74050 46844 74060 46900
rect 74116 46844 77420 46900
rect 77476 46844 77486 46900
rect 79200 46676 80000 46704
rect 78194 46620 78204 46676
rect 78260 46620 80000 46676
rect 79200 46592 80000 46620
rect 4466 46228 4476 46284
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4740 46228 4750 46284
rect 35186 46228 35196 46284
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35460 46228 35470 46284
rect 65906 46228 65916 46284
rect 65972 46228 66020 46284
rect 66076 46228 66124 46284
rect 66180 46228 66190 46284
rect 71922 46172 71932 46228
rect 71988 46172 77532 46228
rect 77588 46172 77598 46228
rect 0 46004 800 46032
rect 0 45948 1932 46004
rect 1988 45948 1998 46004
rect 0 45920 800 45948
rect 2370 45836 2380 45892
rect 2436 45836 3052 45892
rect 3108 45836 3612 45892
rect 3668 45836 3678 45892
rect 2818 45724 2828 45780
rect 2884 45724 3276 45780
rect 3332 45724 4284 45780
rect 4340 45724 4350 45780
rect 79200 45556 80000 45584
rect 77634 45500 77644 45556
rect 77700 45500 78204 45556
rect 78260 45500 80000 45556
rect 19826 45444 19836 45500
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 20100 45444 20110 45500
rect 50546 45444 50556 45500
rect 50612 45444 50660 45500
rect 50716 45444 50764 45500
rect 50820 45444 50830 45500
rect 79200 45472 80000 45500
rect 55794 45276 55804 45332
rect 55860 45276 58492 45332
rect 58548 45276 58558 45332
rect 71138 45276 71148 45332
rect 71204 45276 77308 45332
rect 77364 45276 77374 45332
rect 74050 45164 74060 45220
rect 74116 45164 77868 45220
rect 77924 45164 77934 45220
rect 77634 44940 77644 44996
rect 77700 44940 78204 44996
rect 78260 44940 78270 44996
rect 0 44884 800 44912
rect 0 44828 2716 44884
rect 2772 44828 2782 44884
rect 0 44800 800 44828
rect 4466 44660 4476 44716
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4740 44660 4750 44716
rect 35186 44660 35196 44716
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35460 44660 35470 44716
rect 65906 44660 65916 44716
rect 65972 44660 66020 44716
rect 66076 44660 66124 44716
rect 66180 44660 66190 44716
rect 72258 44604 72268 44660
rect 72324 44604 77756 44660
rect 77812 44604 77822 44660
rect 79200 44436 80000 44464
rect 78194 44380 78204 44436
rect 78260 44380 80000 44436
rect 79200 44352 80000 44380
rect 2706 44044 2716 44100
rect 2772 44044 2782 44100
rect 2716 43988 2772 44044
rect 924 43932 2772 43988
rect 0 43764 800 43792
rect 924 43764 980 43932
rect 19826 43876 19836 43932
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 20100 43876 20110 43932
rect 50546 43876 50556 43932
rect 50612 43876 50660 43932
rect 50716 43876 50764 43932
rect 50820 43876 50830 43932
rect 0 43708 980 43764
rect 57148 43708 59500 43764
rect 59556 43708 59566 43764
rect 0 43680 800 43708
rect 57148 43652 57204 43708
rect 56690 43596 56700 43652
rect 56756 43596 57204 43652
rect 75394 43596 75404 43652
rect 75460 43596 77868 43652
rect 77924 43596 77934 43652
rect 2258 43484 2268 43540
rect 2324 43484 2828 43540
rect 2884 43484 2894 43540
rect 70466 43484 70476 43540
rect 70532 43484 76300 43540
rect 76356 43484 77084 43540
rect 77140 43484 77150 43540
rect 79200 43316 80000 43344
rect 63746 43260 63756 43316
rect 63812 43260 73948 43316
rect 77634 43260 77644 43316
rect 77700 43260 78204 43316
rect 78260 43260 80000 43316
rect 4466 43092 4476 43148
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4740 43092 4750 43148
rect 35186 43092 35196 43148
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35460 43092 35470 43148
rect 65906 43092 65916 43148
rect 65972 43092 66020 43148
rect 66076 43092 66124 43148
rect 66180 43092 66190 43148
rect 73892 43092 73948 43260
rect 79200 43232 80000 43260
rect 73892 43036 77308 43092
rect 77364 43036 77374 43092
rect 72146 42924 72156 42980
rect 72212 42924 75292 42980
rect 75348 42924 75358 42980
rect 1922 42812 1932 42868
rect 1988 42812 1998 42868
rect 58482 42812 58492 42868
rect 58548 42812 59948 42868
rect 60004 42812 60014 42868
rect 68674 42812 68684 42868
rect 68740 42812 76524 42868
rect 76580 42812 77084 42868
rect 77140 42812 77150 42868
rect 0 42644 800 42672
rect 1932 42644 1988 42812
rect 2706 42700 2716 42756
rect 2772 42700 3836 42756
rect 3892 42700 3902 42756
rect 62066 42700 62076 42756
rect 62132 42700 76412 42756
rect 76468 42700 76478 42756
rect 0 42588 1988 42644
rect 77410 42588 77420 42644
rect 77476 42588 77644 42644
rect 77700 42588 77710 42644
rect 0 42560 800 42588
rect 19826 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20110 42364
rect 50546 42308 50556 42364
rect 50612 42308 50660 42364
rect 50716 42308 50764 42364
rect 50820 42308 50830 42364
rect 79200 42196 80000 42224
rect 77970 42140 77980 42196
rect 78036 42140 80000 42196
rect 79200 42112 80000 42140
rect 75730 42028 75740 42084
rect 75796 42028 77756 42084
rect 77812 42028 77822 42084
rect 1698 41916 1708 41972
rect 1764 41916 3836 41972
rect 3892 41916 4732 41972
rect 4788 41916 4798 41972
rect 63410 41916 63420 41972
rect 63476 41916 64540 41972
rect 64596 41916 64606 41972
rect 64866 41916 64876 41972
rect 64932 41916 65324 41972
rect 65380 41916 65390 41972
rect 43250 41804 43260 41860
rect 43316 41804 55580 41860
rect 55636 41804 56140 41860
rect 56196 41804 62188 41860
rect 62626 41804 62636 41860
rect 62692 41804 63644 41860
rect 63700 41804 63710 41860
rect 65660 41804 70812 41860
rect 70868 41804 74732 41860
rect 74788 41804 74844 41860
rect 74900 41804 74910 41860
rect 62132 41748 62188 41804
rect 65660 41748 65716 41804
rect 1922 41692 1932 41748
rect 1988 41692 1998 41748
rect 55458 41692 55468 41748
rect 55524 41692 56812 41748
rect 56868 41692 57708 41748
rect 57764 41692 58380 41748
rect 58436 41692 58446 41748
rect 62132 41692 65716 41748
rect 65772 41692 70588 41748
rect 70644 41692 71372 41748
rect 71428 41692 71438 41748
rect 0 41524 800 41552
rect 1932 41524 1988 41692
rect 62178 41580 62188 41636
rect 62244 41580 63308 41636
rect 63364 41580 63374 41636
rect 4466 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4750 41580
rect 35186 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35470 41580
rect 65772 41524 65828 41692
rect 65906 41524 65916 41580
rect 65972 41524 66020 41580
rect 66076 41524 66124 41580
rect 66180 41524 66190 41580
rect 0 41468 1988 41524
rect 57474 41468 57484 41524
rect 57540 41468 65828 41524
rect 72006 41468 72044 41524
rect 72100 41468 72110 41524
rect 0 41440 800 41468
rect 62178 41356 62188 41412
rect 62244 41356 62636 41412
rect 62692 41356 62702 41412
rect 69570 41356 69580 41412
rect 69636 41356 76748 41412
rect 76804 41356 76814 41412
rect 59714 41244 59724 41300
rect 59780 41244 61516 41300
rect 61572 41244 61582 41300
rect 70914 41244 70924 41300
rect 70980 41244 71932 41300
rect 71988 41244 71998 41300
rect 74162 41244 74172 41300
rect 74228 41244 75180 41300
rect 75236 41244 75246 41300
rect 76402 41244 76412 41300
rect 76468 41244 78092 41300
rect 78148 41244 78158 41300
rect 62402 41132 62412 41188
rect 62468 41132 62748 41188
rect 62804 41132 62972 41188
rect 63028 41132 64204 41188
rect 64260 41132 64270 41188
rect 64866 41132 64876 41188
rect 64932 41132 65660 41188
rect 65716 41132 65726 41188
rect 70354 41132 70364 41188
rect 70420 41132 71484 41188
rect 71540 41132 71550 41188
rect 72146 41132 72156 41188
rect 72212 41132 74284 41188
rect 74340 41132 74350 41188
rect 79200 41076 80000 41104
rect 61058 41020 61068 41076
rect 61124 41020 61628 41076
rect 61684 41020 64484 41076
rect 65314 41020 65324 41076
rect 65380 41020 65772 41076
rect 65828 41020 65838 41076
rect 68338 41020 68348 41076
rect 68404 41020 73164 41076
rect 73220 41020 73230 41076
rect 76514 41020 76524 41076
rect 76580 41020 80000 41076
rect 64428 40964 64484 41020
rect 68348 40964 68404 41020
rect 79200 40992 80000 41020
rect 64418 40908 64428 40964
rect 64484 40908 68404 40964
rect 72006 40908 72044 40964
rect 72100 40908 72110 40964
rect 76738 40908 76748 40964
rect 76804 40908 77084 40964
rect 77140 40908 77150 40964
rect 77606 40908 77644 40964
rect 77700 40908 77710 40964
rect 56242 40796 56252 40852
rect 56308 40796 56588 40852
rect 56644 40796 70812 40852
rect 70868 40796 70878 40852
rect 72482 40796 72492 40852
rect 72548 40796 78540 40852
rect 78596 40796 78606 40852
rect 19826 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20110 40796
rect 50546 40740 50556 40796
rect 50612 40740 50660 40796
rect 50716 40740 50764 40796
rect 50820 40740 50830 40796
rect 2258 40572 2268 40628
rect 2324 40572 5404 40628
rect 5460 40572 5470 40628
rect 55234 40572 55244 40628
rect 55300 40572 62188 40628
rect 66322 40572 66332 40628
rect 66388 40572 67452 40628
rect 67508 40572 67518 40628
rect 67666 40572 67676 40628
rect 67732 40572 69580 40628
rect 69636 40572 69646 40628
rect 69794 40572 69804 40628
rect 69860 40572 70028 40628
rect 70084 40572 70252 40628
rect 70308 40572 70318 40628
rect 73714 40572 73724 40628
rect 73780 40572 74620 40628
rect 74676 40572 77644 40628
rect 77700 40572 77710 40628
rect 4050 40460 4060 40516
rect 4116 40460 4508 40516
rect 4564 40460 5180 40516
rect 5236 40460 5246 40516
rect 59826 40460 59836 40516
rect 59892 40460 60956 40516
rect 61012 40460 61292 40516
rect 61348 40460 61358 40516
rect 0 40404 800 40432
rect 62132 40404 62188 40572
rect 65090 40460 65100 40516
rect 65156 40460 67900 40516
rect 67956 40460 67966 40516
rect 0 40348 1932 40404
rect 1988 40348 1998 40404
rect 3154 40348 3164 40404
rect 3220 40348 4956 40404
rect 5012 40348 26908 40404
rect 26964 40348 26974 40404
rect 42242 40348 42252 40404
rect 42308 40348 43260 40404
rect 43316 40348 43326 40404
rect 58706 40348 58716 40404
rect 58772 40348 60060 40404
rect 60116 40348 60508 40404
rect 60564 40348 61068 40404
rect 61124 40348 61134 40404
rect 62132 40348 70812 40404
rect 70868 40348 71708 40404
rect 71764 40348 71774 40404
rect 74834 40348 74844 40404
rect 74900 40348 74956 40404
rect 75012 40348 75022 40404
rect 0 40320 800 40348
rect 51986 40236 51996 40292
rect 52052 40236 56252 40292
rect 56308 40236 56318 40292
rect 60722 40236 60732 40292
rect 60788 40236 62188 40292
rect 62244 40236 63196 40292
rect 63252 40236 63262 40292
rect 73378 40236 73388 40292
rect 73444 40236 77980 40292
rect 78036 40236 78046 40292
rect 54226 40124 54236 40180
rect 54292 40124 72940 40180
rect 72996 40124 73006 40180
rect 75394 40124 75404 40180
rect 75460 40124 75852 40180
rect 75908 40124 76972 40180
rect 77028 40124 77038 40180
rect 51874 40012 51884 40068
rect 51940 40012 54908 40068
rect 54964 40012 54974 40068
rect 4466 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4750 40012
rect 35186 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35470 40012
rect 65906 39956 65916 40012
rect 65972 39956 66020 40012
rect 66076 39956 66124 40012
rect 66180 39956 66190 40012
rect 79200 39956 80000 39984
rect 75282 39900 75292 39956
rect 75348 39900 78092 39956
rect 78148 39900 78158 39956
rect 78316 39900 80000 39956
rect 78316 39844 78372 39900
rect 79200 39872 80000 39900
rect 75058 39788 75068 39844
rect 75124 39788 75964 39844
rect 76020 39788 78372 39844
rect 61170 39676 61180 39732
rect 61236 39676 62636 39732
rect 62692 39676 62702 39732
rect 66546 39676 66556 39732
rect 66612 39676 67116 39732
rect 67172 39676 67182 39732
rect 69458 39676 69468 39732
rect 69524 39676 71372 39732
rect 71428 39676 71438 39732
rect 72930 39676 72940 39732
rect 72996 39676 74508 39732
rect 74564 39676 74574 39732
rect 75618 39676 75628 39732
rect 75684 39676 76076 39732
rect 76132 39676 76142 39732
rect 2594 39564 2604 39620
rect 2660 39564 3836 39620
rect 3892 39564 4732 39620
rect 4788 39564 4798 39620
rect 65650 39564 65660 39620
rect 65716 39564 66780 39620
rect 66836 39564 66846 39620
rect 69570 39564 69580 39620
rect 69636 39564 70252 39620
rect 70308 39564 70318 39620
rect 70690 39564 70700 39620
rect 70756 39564 71596 39620
rect 71652 39564 71662 39620
rect 73490 39564 73500 39620
rect 73556 39564 74284 39620
rect 74340 39564 74350 39620
rect 75282 39564 75292 39620
rect 75348 39564 76524 39620
rect 76580 39564 76590 39620
rect 70914 39452 70924 39508
rect 70980 39452 71372 39508
rect 71428 39452 71438 39508
rect 73266 39452 73276 39508
rect 73332 39452 73836 39508
rect 73892 39452 74956 39508
rect 75012 39452 75022 39508
rect 76178 39452 76188 39508
rect 76244 39452 76254 39508
rect 5170 39340 5180 39396
rect 5236 39340 42924 39396
rect 42980 39340 42990 39396
rect 63634 39340 63644 39396
rect 63700 39340 64316 39396
rect 64372 39340 64382 39396
rect 66994 39340 67004 39396
rect 67060 39340 67564 39396
rect 67620 39340 67630 39396
rect 74050 39340 74060 39396
rect 74116 39340 74396 39396
rect 74452 39340 74462 39396
rect 0 39284 800 39312
rect 76188 39284 76244 39452
rect 0 39228 1932 39284
rect 1988 39228 1998 39284
rect 56802 39228 56812 39284
rect 56868 39228 76244 39284
rect 0 39200 800 39228
rect 19826 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20110 39228
rect 50546 39172 50556 39228
rect 50612 39172 50660 39228
rect 50716 39172 50764 39228
rect 50820 39172 50830 39228
rect 77186 39116 77196 39172
rect 77252 39116 77868 39172
rect 77924 39116 77934 39172
rect 41122 39004 41132 39060
rect 41188 39004 51884 39060
rect 51940 39004 51950 39060
rect 69458 39004 69468 39060
rect 69524 39004 71596 39060
rect 71652 39004 73500 39060
rect 73556 39004 73566 39060
rect 74162 39004 74172 39060
rect 74228 39004 74508 39060
rect 74564 39004 74574 39060
rect 77410 39004 77420 39060
rect 77476 39004 77980 39060
rect 78036 39004 78046 39060
rect 26898 38892 26908 38948
rect 26964 38892 40796 38948
rect 40852 38892 40862 38948
rect 42690 38892 42700 38948
rect 42756 38892 43708 38948
rect 58146 38892 58156 38948
rect 58212 38892 74284 38948
rect 74340 38892 75068 38948
rect 75124 38892 75134 38948
rect 76402 38892 76412 38948
rect 76468 38892 76748 38948
rect 76804 38892 76814 38948
rect 41682 38780 41692 38836
rect 41748 38780 42588 38836
rect 42644 38780 42654 38836
rect 43652 38780 43708 38892
rect 79200 38836 80000 38864
rect 43764 38780 51996 38836
rect 52052 38780 52062 38836
rect 64306 38780 64316 38836
rect 64372 38780 65212 38836
rect 65268 38780 66332 38836
rect 66388 38780 66398 38836
rect 68562 38780 68572 38836
rect 68628 38780 69020 38836
rect 69076 38780 69086 38836
rect 70466 38780 70476 38836
rect 70532 38780 70542 38836
rect 70690 38780 70700 38836
rect 70756 38780 72156 38836
rect 72212 38780 72222 38836
rect 76934 38780 76972 38836
rect 77028 38780 77038 38836
rect 78194 38780 78204 38836
rect 78260 38780 80000 38836
rect 2930 38668 2940 38724
rect 2996 38668 3276 38724
rect 3332 38668 41580 38724
rect 41636 38668 41646 38724
rect 50306 38668 50316 38724
rect 50372 38668 51660 38724
rect 51716 38668 51726 38724
rect 62962 38668 62972 38724
rect 63028 38668 63532 38724
rect 63588 38668 63598 38724
rect 67330 38668 67340 38724
rect 67396 38668 68124 38724
rect 68180 38668 69356 38724
rect 69412 38668 69422 38724
rect 70476 38612 70532 38780
rect 79200 38752 80000 38780
rect 70914 38668 70924 38724
rect 70980 38668 71372 38724
rect 71428 38668 71438 38724
rect 73490 38668 73500 38724
rect 73556 38668 74172 38724
rect 74228 38668 74238 38724
rect 69010 38556 69020 38612
rect 69076 38556 70532 38612
rect 74498 38556 74508 38612
rect 74564 38556 75068 38612
rect 75124 38556 75404 38612
rect 75460 38556 75470 38612
rect 69234 38444 69244 38500
rect 69300 38444 70140 38500
rect 70196 38444 70206 38500
rect 70578 38444 70588 38500
rect 70644 38444 71260 38500
rect 71316 38444 72604 38500
rect 72660 38444 72670 38500
rect 4466 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4750 38444
rect 35186 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35470 38444
rect 65906 38388 65916 38444
rect 65972 38388 66020 38444
rect 66076 38388 66124 38444
rect 66180 38388 66190 38444
rect 69430 38332 69468 38388
rect 69524 38332 69534 38388
rect 74946 38220 74956 38276
rect 75012 38220 75068 38276
rect 75124 38220 75134 38276
rect 0 38164 800 38192
rect 0 38108 3388 38164
rect 3444 38108 3454 38164
rect 0 38080 800 38108
rect 66546 37996 66556 38052
rect 66612 37996 68348 38052
rect 68404 37996 68414 38052
rect 71362 37996 71372 38052
rect 71428 37996 73052 38052
rect 73108 37996 73118 38052
rect 74274 37996 74284 38052
rect 74340 37996 74508 38052
rect 74564 37996 74574 38052
rect 74162 37884 74172 37940
rect 74228 37884 76076 37940
rect 76132 37884 76142 37940
rect 72370 37772 72380 37828
rect 72436 37772 73500 37828
rect 73556 37772 73566 37828
rect 74050 37772 74060 37828
rect 74116 37772 74172 37828
rect 74228 37772 74238 37828
rect 76402 37772 76412 37828
rect 76468 37772 77644 37828
rect 77700 37772 77710 37828
rect 79200 37716 80000 37744
rect 60498 37660 60508 37716
rect 60564 37660 77308 37716
rect 77364 37660 77374 37716
rect 77858 37660 77868 37716
rect 77924 37660 80000 37716
rect 19826 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20110 37660
rect 50546 37604 50556 37660
rect 50612 37604 50660 37660
rect 50716 37604 50764 37660
rect 50820 37604 50830 37660
rect 79200 37632 80000 37660
rect 70130 37548 70140 37604
rect 70196 37548 70476 37604
rect 70532 37548 70542 37604
rect 70802 37548 70812 37604
rect 70868 37548 71708 37604
rect 71764 37548 72268 37604
rect 72324 37548 72828 37604
rect 72884 37548 72894 37604
rect 67778 37436 67788 37492
rect 67844 37436 68460 37492
rect 68516 37436 70028 37492
rect 70084 37436 70588 37492
rect 70644 37436 71148 37492
rect 71204 37436 71214 37492
rect 71474 37436 71484 37492
rect 71540 37436 74284 37492
rect 74340 37436 74676 37492
rect 76402 37436 76412 37492
rect 76468 37436 77532 37492
rect 77588 37436 77598 37492
rect 2034 37324 2044 37380
rect 2100 37324 26908 37380
rect 26964 37324 26974 37380
rect 72818 37324 72828 37380
rect 72884 37324 73276 37380
rect 73332 37324 73948 37380
rect 74004 37324 74014 37380
rect 74620 37268 74676 37436
rect 76178 37324 76188 37380
rect 76244 37324 78428 37380
rect 78484 37324 78764 37380
rect 78820 37324 78830 37380
rect 71698 37212 71708 37268
rect 71764 37212 74172 37268
rect 74228 37212 74284 37268
rect 74340 37212 74350 37268
rect 74610 37212 74620 37268
rect 74676 37212 75068 37268
rect 75124 37212 75134 37268
rect 75394 37212 75404 37268
rect 75460 37212 76524 37268
rect 76580 37212 78540 37268
rect 78596 37212 78606 37268
rect 57922 37100 57932 37156
rect 57988 37100 68124 37156
rect 68180 37100 68684 37156
rect 68740 37100 68750 37156
rect 74050 37100 74060 37156
rect 74116 37100 74508 37156
rect 74564 37100 74574 37156
rect 75506 37100 75516 37156
rect 75572 37100 77420 37156
rect 77476 37100 77486 37156
rect 0 37044 800 37072
rect 0 36988 1708 37044
rect 1764 36988 2492 37044
rect 2548 36988 2558 37044
rect 73378 36988 73388 37044
rect 73444 36988 73948 37044
rect 74004 36988 74014 37044
rect 74246 36988 74284 37044
rect 74340 36988 74350 37044
rect 75170 36988 75180 37044
rect 75236 36988 76188 37044
rect 76244 36988 76254 37044
rect 76514 36988 76524 37044
rect 76580 36988 76748 37044
rect 76804 36988 76972 37044
rect 77028 36988 77038 37044
rect 0 36960 800 36988
rect 72454 36876 72492 36932
rect 72548 36876 72558 36932
rect 73154 36876 73164 36932
rect 73220 36876 73500 36932
rect 73556 36876 73566 36932
rect 4466 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4750 36876
rect 35186 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35470 36876
rect 65906 36820 65916 36876
rect 65972 36820 66020 36876
rect 66076 36820 66124 36876
rect 66180 36820 66190 36876
rect 52770 36652 52780 36708
rect 52836 36652 76300 36708
rect 76356 36652 76366 36708
rect 77410 36652 77420 36708
rect 77476 36652 77756 36708
rect 77812 36652 77822 36708
rect 79200 36596 80000 36624
rect 50372 36540 62860 36596
rect 62916 36540 68796 36596
rect 68852 36540 69132 36596
rect 69188 36540 69198 36596
rect 71250 36540 71260 36596
rect 71316 36540 74732 36596
rect 74788 36540 80000 36596
rect 26898 36316 26908 36372
rect 26964 36316 45052 36372
rect 45108 36316 45612 36372
rect 45668 36316 45678 36372
rect 50372 36260 50428 36540
rect 79200 36512 80000 36540
rect 69234 36428 69244 36484
rect 69300 36428 69692 36484
rect 69748 36428 69758 36484
rect 72146 36428 72156 36484
rect 72212 36428 73164 36484
rect 73220 36428 73230 36484
rect 75618 36316 75628 36372
rect 75684 36316 76300 36372
rect 76356 36316 77420 36372
rect 77476 36316 77486 36372
rect 2034 36204 2044 36260
rect 2100 36204 44716 36260
rect 44772 36204 44782 36260
rect 46610 36204 46620 36260
rect 46676 36204 50428 36260
rect 73042 36204 73052 36260
rect 73108 36204 73612 36260
rect 73668 36204 73678 36260
rect 54114 36092 54124 36148
rect 54180 36092 77532 36148
rect 77588 36092 77598 36148
rect 19826 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20110 36092
rect 50546 36036 50556 36092
rect 50612 36036 50660 36092
rect 50716 36036 50764 36092
rect 50820 36036 50830 36092
rect 75030 35980 75068 36036
rect 75124 35980 75134 36036
rect 76066 35980 76076 36036
rect 76132 35980 76972 36036
rect 77028 35980 77038 36036
rect 0 35924 800 35952
rect 0 35868 1708 35924
rect 1764 35868 2492 35924
rect 2548 35868 2558 35924
rect 55346 35868 55356 35924
rect 55412 35868 56812 35924
rect 56868 35868 56878 35924
rect 71362 35868 71372 35924
rect 71428 35868 76300 35924
rect 76356 35868 77196 35924
rect 77252 35868 77262 35924
rect 0 35840 800 35868
rect 54226 35756 54236 35812
rect 54292 35756 54908 35812
rect 54964 35756 54974 35812
rect 65426 35756 65436 35812
rect 65492 35756 73948 35812
rect 75618 35756 75628 35812
rect 75684 35756 76748 35812
rect 76804 35756 77532 35812
rect 77588 35756 77598 35812
rect 73892 35700 73948 35756
rect 45154 35644 45164 35700
rect 45220 35644 45724 35700
rect 45780 35644 45790 35700
rect 45938 35644 45948 35700
rect 46004 35644 54012 35700
rect 54068 35644 54078 35700
rect 72146 35644 72156 35700
rect 72212 35644 73276 35700
rect 73332 35644 73342 35700
rect 73892 35644 77308 35700
rect 77364 35644 78652 35700
rect 78708 35644 78718 35700
rect 55682 35532 55692 35588
rect 55748 35532 56700 35588
rect 56756 35532 56766 35588
rect 71698 35532 71708 35588
rect 71764 35532 72268 35588
rect 72324 35532 72334 35588
rect 74274 35532 74284 35588
rect 74340 35532 74620 35588
rect 74676 35532 74686 35588
rect 79200 35476 80000 35504
rect 74498 35420 74508 35476
rect 74564 35420 74620 35476
rect 74676 35420 74686 35476
rect 75730 35420 75740 35476
rect 75796 35420 80000 35476
rect 79200 35392 80000 35420
rect 73602 35308 73612 35364
rect 73668 35308 74060 35364
rect 74116 35308 74126 35364
rect 74284 35308 78876 35364
rect 78932 35308 78942 35364
rect 4466 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4750 35308
rect 35186 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35470 35308
rect 65906 35252 65916 35308
rect 65972 35252 66020 35308
rect 66076 35252 66124 35308
rect 66180 35252 66190 35308
rect 46050 35196 46060 35252
rect 46116 35196 55020 35252
rect 55076 35196 55086 35252
rect 72930 35196 72940 35252
rect 72996 35196 73500 35252
rect 73556 35196 73836 35252
rect 73892 35196 73902 35252
rect 74284 35140 74340 35308
rect 45154 35084 45164 35140
rect 45220 35084 45724 35140
rect 45780 35084 45790 35140
rect 73602 35084 73612 35140
rect 73668 35084 74340 35140
rect 77830 35084 77868 35140
rect 77924 35084 77934 35140
rect 46274 34972 46284 35028
rect 46340 34972 46956 35028
rect 47012 34972 47022 35028
rect 53778 34972 53788 35028
rect 53844 34972 55356 35028
rect 55412 34972 60508 35028
rect 60564 34972 60574 35028
rect 68002 34972 68012 35028
rect 68068 34972 75740 35028
rect 75796 34972 76524 35028
rect 76580 34972 76590 35028
rect 77868 34916 77924 35084
rect 46834 34860 46844 34916
rect 46900 34860 53900 34916
rect 53956 34860 53966 34916
rect 71362 34860 71372 34916
rect 71428 34860 77924 34916
rect 0 34804 800 34832
rect 0 34748 1708 34804
rect 1764 34748 2492 34804
rect 2548 34748 2558 34804
rect 45266 34748 45276 34804
rect 45332 34748 46620 34804
rect 46676 34748 46686 34804
rect 73490 34748 73500 34804
rect 73556 34748 73566 34804
rect 0 34720 800 34748
rect 73500 34692 73556 34748
rect 2034 34636 2044 34692
rect 2100 34636 44380 34692
rect 44436 34636 45164 34692
rect 45220 34636 45230 34692
rect 71810 34636 71820 34692
rect 71876 34636 71886 34692
rect 73042 34636 73052 34692
rect 73108 34636 73276 34692
rect 73332 34636 73342 34692
rect 73500 34636 74172 34692
rect 74228 34636 75292 34692
rect 75348 34636 75358 34692
rect 71820 34580 71876 34636
rect 71820 34524 77532 34580
rect 77588 34524 77598 34580
rect 78194 34524 78204 34580
rect 78260 34524 78540 34580
rect 78596 34524 78606 34580
rect 19826 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20110 34524
rect 50546 34468 50556 34524
rect 50612 34468 50660 34524
rect 50716 34468 50764 34524
rect 50820 34468 50830 34524
rect 72818 34412 72828 34468
rect 72884 34412 73164 34468
rect 73220 34412 73230 34468
rect 73938 34412 73948 34468
rect 74004 34412 74620 34468
rect 74676 34412 74686 34468
rect 79200 34356 80000 34384
rect 45714 34300 45724 34356
rect 45780 34300 46508 34356
rect 46564 34300 46574 34356
rect 52882 34300 52892 34356
rect 52948 34300 76300 34356
rect 76356 34300 76366 34356
rect 76524 34300 80000 34356
rect 76524 34244 76580 34300
rect 79200 34272 80000 34300
rect 71138 34188 71148 34244
rect 71204 34188 72156 34244
rect 72212 34188 73164 34244
rect 73220 34188 73230 34244
rect 73892 34188 75068 34244
rect 75124 34188 76580 34244
rect 77522 34188 77532 34244
rect 77588 34188 78988 34244
rect 79044 34188 79054 34244
rect 45266 34076 45276 34132
rect 45332 34076 45836 34132
rect 45892 34076 45902 34132
rect 46498 34076 46508 34132
rect 46564 34076 47068 34132
rect 47124 34076 47134 34132
rect 63186 34076 63196 34132
rect 63252 34076 71260 34132
rect 71316 34076 71326 34132
rect 71698 34076 71708 34132
rect 71764 34076 72716 34132
rect 72772 34076 73724 34132
rect 73780 34076 73790 34132
rect 73892 34020 73948 34188
rect 74610 34076 74620 34132
rect 74676 34076 77980 34132
rect 78036 34076 78046 34132
rect 70914 33964 70924 34020
rect 70980 33964 73948 34020
rect 75506 33964 75516 34020
rect 75572 33964 76412 34020
rect 76468 33964 76478 34020
rect 75282 33852 75292 33908
rect 75348 33852 77868 33908
rect 77924 33852 77934 33908
rect 74834 33740 74844 33796
rect 74900 33740 77756 33796
rect 77812 33740 78764 33796
rect 78820 33740 78830 33796
rect 0 33684 800 33712
rect 4466 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4750 33740
rect 35186 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35470 33740
rect 65906 33684 65916 33740
rect 65972 33684 66020 33740
rect 66076 33684 66124 33740
rect 66180 33684 66190 33740
rect 0 33628 1708 33684
rect 1764 33628 2492 33684
rect 2548 33628 2558 33684
rect 75058 33628 75068 33684
rect 75124 33628 75180 33684
rect 75236 33628 75246 33684
rect 75842 33628 75852 33684
rect 75908 33628 76860 33684
rect 76916 33628 77084 33684
rect 77140 33628 77644 33684
rect 77700 33628 77710 33684
rect 0 33600 800 33628
rect 73938 33516 73948 33572
rect 74004 33516 75068 33572
rect 75124 33516 75134 33572
rect 76738 33516 76748 33572
rect 76804 33516 77868 33572
rect 77924 33516 77934 33572
rect 52322 33404 52332 33460
rect 52388 33404 53116 33460
rect 53172 33404 53182 33460
rect 53330 33404 53340 33460
rect 53396 33404 54124 33460
rect 54180 33404 54190 33460
rect 73826 33404 73836 33460
rect 73892 33404 74844 33460
rect 74900 33404 74910 33460
rect 76738 33404 76748 33460
rect 76804 33404 76860 33460
rect 76916 33404 76926 33460
rect 2034 33292 2044 33348
rect 2100 33292 8428 33348
rect 46050 33292 46060 33348
rect 46116 33292 53004 33348
rect 53060 33292 53070 33348
rect 74274 33292 74284 33348
rect 74340 33292 74676 33348
rect 75282 33292 75292 33348
rect 75348 33292 77308 33348
rect 77364 33292 77374 33348
rect 8372 33236 8428 33292
rect 74620 33236 74676 33292
rect 79200 33236 80000 33264
rect 8372 33180 45164 33236
rect 45220 33180 45724 33236
rect 45780 33180 45790 33236
rect 58818 33180 58828 33236
rect 58884 33180 74396 33236
rect 74452 33180 74462 33236
rect 74620 33180 75180 33236
rect 75236 33180 80000 33236
rect 79200 33152 80000 33180
rect 2034 33068 2044 33124
rect 2100 33068 28476 33124
rect 28532 33068 28542 33124
rect 71586 33068 71596 33124
rect 71652 33068 73948 33124
rect 74162 33068 74172 33124
rect 74228 33068 76636 33124
rect 76692 33068 76702 33124
rect 76850 33068 76860 33124
rect 76916 33068 76926 33124
rect 73892 33012 73948 33068
rect 76860 33012 76916 33068
rect 71698 32956 71708 33012
rect 71764 32956 72940 33012
rect 72996 32956 73006 33012
rect 73892 32956 76916 33012
rect 19826 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20110 32956
rect 50546 32900 50556 32956
rect 50612 32900 50660 32956
rect 50716 32900 50764 32956
rect 50820 32900 50830 32956
rect 71810 32844 71820 32900
rect 71876 32844 73948 32900
rect 74004 32844 74014 32900
rect 73714 32732 73724 32788
rect 73780 32732 73948 32788
rect 75954 32732 75964 32788
rect 76020 32732 77756 32788
rect 77812 32732 77822 32788
rect 0 32564 800 32592
rect 73892 32564 73948 32732
rect 75058 32620 75068 32676
rect 75124 32620 77532 32676
rect 77588 32620 77598 32676
rect 0 32508 1708 32564
rect 1764 32508 2492 32564
rect 2548 32508 2558 32564
rect 73892 32508 77756 32564
rect 77812 32508 77822 32564
rect 0 32480 800 32508
rect 71138 32396 71148 32452
rect 71204 32396 72156 32452
rect 72212 32396 73500 32452
rect 73556 32396 75292 32452
rect 75348 32396 76412 32452
rect 76468 32396 76478 32452
rect 77410 32396 77420 32452
rect 77476 32396 78428 32452
rect 78484 32396 78494 32452
rect 52322 32284 52332 32340
rect 52388 32284 74844 32340
rect 74900 32284 74910 32340
rect 75058 32284 75068 32340
rect 75124 32284 75162 32340
rect 68898 32172 68908 32228
rect 68964 32172 74956 32228
rect 75012 32172 75022 32228
rect 4466 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4750 32172
rect 35186 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35470 32172
rect 65906 32116 65916 32172
rect 65972 32116 66020 32172
rect 66076 32116 66124 32172
rect 66180 32116 66190 32172
rect 79200 32116 80000 32144
rect 71138 32060 71148 32116
rect 71204 32060 72268 32116
rect 72324 32060 72334 32116
rect 74386 32060 74396 32116
rect 74452 32060 77308 32116
rect 77364 32060 77374 32116
rect 78194 32060 78204 32116
rect 78260 32060 80000 32116
rect 79200 32032 80000 32060
rect 51314 31948 51324 32004
rect 51380 31948 74284 32004
rect 74340 31948 74350 32004
rect 51426 31836 51436 31892
rect 51492 31836 52780 31892
rect 52836 31836 52846 31892
rect 70914 31836 70924 31892
rect 70980 31836 71708 31892
rect 71764 31836 72604 31892
rect 72660 31836 72670 31892
rect 75702 31836 75740 31892
rect 75796 31836 75806 31892
rect 77410 31836 77420 31892
rect 77476 31836 78876 31892
rect 78932 31836 78942 31892
rect 46162 31724 46172 31780
rect 46228 31724 51100 31780
rect 51156 31724 51166 31780
rect 58594 31724 58604 31780
rect 58660 31724 73052 31780
rect 73108 31724 73724 31780
rect 73780 31724 73790 31780
rect 76822 31724 76860 31780
rect 76916 31724 76926 31780
rect 28466 31612 28476 31668
rect 28532 31612 44828 31668
rect 44884 31612 44894 31668
rect 45042 31612 45052 31668
rect 45108 31612 45948 31668
rect 46004 31612 46014 31668
rect 58930 31612 58940 31668
rect 58996 31612 74620 31668
rect 74676 31612 74686 31668
rect 44828 31556 44884 31612
rect 2034 31500 2044 31556
rect 2100 31500 44268 31556
rect 44324 31500 44334 31556
rect 44828 31500 45500 31556
rect 45556 31500 45566 31556
rect 54674 31500 54684 31556
rect 54740 31500 55132 31556
rect 55188 31500 55198 31556
rect 71474 31500 71484 31556
rect 71540 31500 72268 31556
rect 72324 31500 73276 31556
rect 73332 31500 73342 31556
rect 74498 31500 74508 31556
rect 74564 31500 76636 31556
rect 76692 31500 76702 31556
rect 0 31444 800 31472
rect 76860 31444 76916 31724
rect 0 31388 1708 31444
rect 1764 31388 2492 31444
rect 2548 31388 2558 31444
rect 72146 31388 72156 31444
rect 72212 31388 72716 31444
rect 72772 31388 74732 31444
rect 74788 31388 74798 31444
rect 75404 31388 76916 31444
rect 0 31360 800 31388
rect 19826 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20110 31388
rect 50546 31332 50556 31388
rect 50612 31332 50660 31388
rect 50716 31332 50764 31388
rect 50820 31332 50830 31388
rect 75404 31332 75460 31388
rect 73490 31276 73500 31332
rect 73556 31276 75460 31332
rect 75618 31276 75628 31332
rect 75684 31276 77980 31332
rect 78036 31276 78046 31332
rect 51426 31164 51436 31220
rect 51492 31164 52780 31220
rect 52836 31164 52846 31220
rect 73892 31164 78148 31220
rect 73892 31108 73948 31164
rect 78092 31108 78148 31164
rect 2034 31052 2044 31108
rect 2100 31052 26908 31108
rect 26964 31052 26974 31108
rect 45714 31052 45724 31108
rect 45780 31052 46396 31108
rect 46452 31052 47292 31108
rect 47348 31052 47358 31108
rect 50306 31052 50316 31108
rect 50372 31052 52332 31108
rect 52388 31052 52398 31108
rect 70914 31052 70924 31108
rect 70980 31052 73948 31108
rect 74498 31052 74508 31108
rect 74564 31052 75516 31108
rect 75572 31052 75582 31108
rect 77410 31052 77420 31108
rect 77476 31052 77924 31108
rect 78082 31052 78092 31108
rect 78148 31052 78158 31108
rect 74844 30996 74900 31052
rect 44706 30940 44716 30996
rect 44772 30940 45948 30996
rect 46004 30940 46014 30996
rect 46162 30940 46172 30996
rect 46228 30940 51100 30996
rect 51156 30940 51166 30996
rect 59602 30940 59612 30996
rect 59668 30940 73500 30996
rect 73556 30940 73836 30996
rect 73892 30940 74172 30996
rect 74228 30940 74238 30996
rect 74722 30940 74732 30996
rect 74788 30940 74844 30996
rect 74900 30940 74910 30996
rect 75170 30940 75180 30996
rect 75236 30940 76636 30996
rect 76692 30940 77644 30996
rect 77700 30940 77710 30996
rect 1698 30828 1708 30884
rect 1764 30828 2492 30884
rect 2548 30828 2558 30884
rect 47058 30828 47068 30884
rect 47124 30828 50540 30884
rect 50596 30828 50606 30884
rect 71362 30828 71372 30884
rect 71428 30828 71438 30884
rect 76514 30828 76524 30884
rect 76580 30828 77084 30884
rect 77140 30828 77150 30884
rect 71372 30772 71428 30828
rect 77868 30772 77924 31052
rect 79200 30996 80000 31024
rect 51174 30716 51212 30772
rect 51268 30716 51278 30772
rect 69122 30716 69132 30772
rect 69188 30716 70924 30772
rect 70980 30716 70990 30772
rect 71372 30716 77924 30772
rect 78316 30940 80000 30996
rect 78316 30660 78372 30940
rect 79200 30912 80000 30940
rect 78306 30604 78316 30660
rect 78372 30604 78382 30660
rect 4466 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4750 30604
rect 35186 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35470 30604
rect 65906 30548 65916 30604
rect 65972 30548 66020 30604
rect 66076 30548 66124 30604
rect 66180 30548 66190 30604
rect 44930 30492 44940 30548
rect 44996 30492 46956 30548
rect 47012 30492 47022 30548
rect 75394 30380 75404 30436
rect 75460 30380 77644 30436
rect 77700 30380 77710 30436
rect 0 30324 800 30352
rect 0 30268 1708 30324
rect 1764 30268 1774 30324
rect 46610 30268 46620 30324
rect 46676 30268 47292 30324
rect 47348 30268 47358 30324
rect 49858 30268 49868 30324
rect 49924 30268 74060 30324
rect 74116 30268 74126 30324
rect 74722 30268 74732 30324
rect 74788 30268 77308 30324
rect 77364 30268 77374 30324
rect 0 30240 800 30268
rect 46162 30156 46172 30212
rect 46228 30156 50652 30212
rect 50708 30156 50718 30212
rect 51762 30156 51772 30212
rect 51828 30156 58828 30212
rect 58884 30156 58894 30212
rect 71362 30156 71372 30212
rect 71428 30156 72828 30212
rect 72884 30156 72894 30212
rect 74946 30156 74956 30212
rect 75012 30156 76188 30212
rect 76244 30156 76254 30212
rect 76598 30156 76636 30212
rect 76692 30156 76972 30212
rect 77028 30156 77038 30212
rect 51772 30100 51828 30156
rect 26898 30044 26908 30100
rect 26964 30044 44828 30100
rect 44884 30044 44894 30100
rect 45154 30044 45164 30100
rect 45220 30044 46060 30100
rect 46116 30044 46126 30100
rect 50754 30044 50764 30100
rect 50820 30044 51828 30100
rect 72678 30044 72716 30100
rect 72772 30044 72782 30100
rect 74498 30044 74508 30100
rect 74564 30044 76524 30100
rect 76580 30044 76590 30100
rect 44828 29988 44884 30044
rect 44828 29932 45388 29988
rect 45444 29932 45454 29988
rect 72566 29932 72604 29988
rect 72660 29932 73052 29988
rect 73108 29932 73118 29988
rect 73490 29932 73500 29988
rect 73556 29932 77196 29988
rect 77252 29932 77262 29988
rect 79200 29876 80000 29904
rect 46050 29820 46060 29876
rect 46116 29820 49532 29876
rect 49588 29820 49598 29876
rect 72706 29820 72716 29876
rect 72772 29820 76412 29876
rect 76468 29820 76478 29876
rect 78530 29820 78540 29876
rect 78596 29820 80000 29876
rect 19826 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20110 29820
rect 50546 29764 50556 29820
rect 50612 29764 50660 29820
rect 50716 29764 50764 29820
rect 50820 29764 50830 29820
rect 79200 29792 80000 29820
rect 72146 29708 72156 29764
rect 72212 29708 76412 29764
rect 76468 29708 76478 29764
rect 61730 29596 61740 29652
rect 61796 29596 73724 29652
rect 73780 29596 73790 29652
rect 2034 29484 2044 29540
rect 2100 29484 44828 29540
rect 44884 29484 44894 29540
rect 74946 29484 74956 29540
rect 75012 29484 76076 29540
rect 76132 29484 76142 29540
rect 76402 29484 76412 29540
rect 76468 29484 76524 29540
rect 76580 29484 76590 29540
rect 18022 29372 18060 29428
rect 18116 29372 18126 29428
rect 50306 29372 50316 29428
rect 50372 29372 58940 29428
rect 58996 29372 59006 29428
rect 69542 29372 69580 29428
rect 69636 29372 69646 29428
rect 73714 29372 73724 29428
rect 73780 29372 73790 29428
rect 73724 29316 73780 29372
rect 50418 29260 50428 29316
rect 50484 29260 72716 29316
rect 72772 29260 72782 29316
rect 73724 29260 75404 29316
rect 75460 29260 75470 29316
rect 75618 29260 75628 29316
rect 75684 29260 76188 29316
rect 76244 29260 76254 29316
rect 0 29204 800 29232
rect 0 29148 1708 29204
rect 1764 29148 2492 29204
rect 2548 29148 2558 29204
rect 34962 29148 34972 29204
rect 35028 29148 38892 29204
rect 38948 29148 38958 29204
rect 50082 29148 50092 29204
rect 50148 29148 73612 29204
rect 73668 29148 73678 29204
rect 75730 29148 75740 29204
rect 75796 29148 76860 29204
rect 76916 29148 77196 29204
rect 77252 29148 77262 29204
rect 0 29120 800 29148
rect 71250 29036 71260 29092
rect 71316 29036 78316 29092
rect 78372 29036 78382 29092
rect 4466 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4750 29036
rect 35186 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35470 29036
rect 65906 28980 65916 29036
rect 65972 28980 66020 29036
rect 66076 28980 66124 29036
rect 66180 28980 66190 29036
rect 72594 28924 72604 28980
rect 72660 28924 72940 28980
rect 72996 28924 73006 28980
rect 73378 28924 73388 28980
rect 73444 28924 75404 28980
rect 75460 28924 75470 28980
rect 76290 28924 76300 28980
rect 76356 28924 76524 28980
rect 76580 28924 76590 28980
rect 76300 28868 76356 28924
rect 75292 28812 76356 28868
rect 71698 28700 71708 28756
rect 71764 28700 75012 28756
rect 74956 28644 75012 28700
rect 75292 28644 75348 28812
rect 79200 28756 80000 28784
rect 78418 28700 78428 28756
rect 78484 28700 80000 28756
rect 79200 28672 80000 28700
rect 2034 28588 2044 28644
rect 2100 28588 44604 28644
rect 44660 28588 44670 28644
rect 49298 28588 49308 28644
rect 49364 28588 50316 28644
rect 50372 28588 50382 28644
rect 71922 28588 71932 28644
rect 71988 28588 72380 28644
rect 72436 28588 74284 28644
rect 74340 28588 74350 28644
rect 74610 28588 74620 28644
rect 74676 28588 74732 28644
rect 74788 28588 74798 28644
rect 74956 28588 75348 28644
rect 75618 28588 75628 28644
rect 75684 28588 76636 28644
rect 76692 28588 76702 28644
rect 37650 28476 37660 28532
rect 37716 28476 38556 28532
rect 38612 28476 38622 28532
rect 62066 28476 62076 28532
rect 62132 28476 62860 28532
rect 62916 28476 62926 28532
rect 72678 28476 72716 28532
rect 72772 28476 72940 28532
rect 72996 28476 73724 28532
rect 73780 28476 73790 28532
rect 74386 28476 74396 28532
rect 74452 28476 75180 28532
rect 75236 28476 75246 28532
rect 75842 28476 75852 28532
rect 75908 28476 76188 28532
rect 76244 28476 76254 28532
rect 36642 28364 36652 28420
rect 36708 28364 73836 28420
rect 73892 28364 73902 28420
rect 74498 28364 74508 28420
rect 74564 28364 75068 28420
rect 75124 28364 75134 28420
rect 75282 28364 75292 28420
rect 75348 28364 75628 28420
rect 75684 28364 75694 28420
rect 61394 28252 61404 28308
rect 61460 28252 68796 28308
rect 68852 28252 68862 28308
rect 71820 28252 74956 28308
rect 75012 28252 75022 28308
rect 19826 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20110 28252
rect 50546 28196 50556 28252
rect 50612 28196 50660 28252
rect 50716 28196 50764 28252
rect 50820 28196 50830 28252
rect 71820 28196 71876 28252
rect 71810 28140 71820 28196
rect 71876 28140 71886 28196
rect 72818 28140 72828 28196
rect 72884 28140 76972 28196
rect 77028 28140 77038 28196
rect 0 28084 800 28112
rect 0 28028 1708 28084
rect 1764 28028 2492 28084
rect 2548 28028 2558 28084
rect 35746 28028 35756 28084
rect 35812 28028 37100 28084
rect 37156 28028 37166 28084
rect 39106 28028 39116 28084
rect 39172 28028 40348 28084
rect 40404 28028 41468 28084
rect 41524 28028 41534 28084
rect 70690 28028 70700 28084
rect 70756 28028 75964 28084
rect 76020 28028 76030 28084
rect 0 28000 800 28028
rect 34514 27916 34524 27972
rect 34580 27916 63868 27972
rect 63924 27916 63934 27972
rect 71922 27916 71932 27972
rect 71988 27916 72268 27972
rect 72324 27916 72334 27972
rect 72706 27916 72716 27972
rect 72772 27916 74060 27972
rect 74116 27916 74172 27972
rect 74228 27916 74238 27972
rect 74918 27916 74956 27972
rect 75012 27916 75022 27972
rect 75394 27916 75404 27972
rect 75460 27916 75852 27972
rect 75908 27916 75918 27972
rect 76150 27916 76188 27972
rect 76244 27916 76254 27972
rect 76636 27916 78204 27972
rect 78260 27916 78540 27972
rect 78596 27916 78606 27972
rect 76636 27860 76692 27916
rect 33506 27804 33516 27860
rect 33572 27804 35308 27860
rect 35364 27804 36652 27860
rect 36708 27804 36718 27860
rect 64866 27804 64876 27860
rect 64932 27804 70700 27860
rect 70756 27804 70766 27860
rect 70914 27804 70924 27860
rect 70980 27804 70990 27860
rect 73490 27804 73500 27860
rect 73556 27804 74284 27860
rect 74340 27804 74732 27860
rect 74788 27804 74798 27860
rect 76626 27804 76636 27860
rect 76692 27804 76702 27860
rect 70924 27748 70980 27804
rect 5394 27692 5404 27748
rect 5460 27692 33404 27748
rect 33460 27692 33470 27748
rect 70924 27692 75404 27748
rect 75460 27692 75470 27748
rect 75954 27692 75964 27748
rect 76020 27692 77084 27748
rect 77140 27692 77150 27748
rect 79200 27636 80000 27664
rect 2034 27580 2044 27636
rect 2100 27580 44828 27636
rect 44884 27580 44894 27636
rect 45042 27580 45052 27636
rect 45108 27580 46172 27636
rect 46228 27580 46238 27636
rect 71362 27580 71372 27636
rect 71428 27580 74396 27636
rect 74452 27580 74462 27636
rect 76178 27580 76188 27636
rect 76244 27580 76254 27636
rect 77746 27580 77756 27636
rect 77812 27580 80000 27636
rect 76188 27524 76244 27580
rect 79200 27552 80000 27580
rect 50866 27468 50876 27524
rect 50932 27468 51324 27524
rect 51380 27468 51390 27524
rect 73892 27468 76244 27524
rect 4466 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4750 27468
rect 35186 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35470 27468
rect 65906 27412 65916 27468
rect 65972 27412 66020 27468
rect 66076 27412 66124 27468
rect 66180 27412 66190 27468
rect 73892 27412 73948 27468
rect 40002 27356 40012 27412
rect 40068 27356 59948 27412
rect 60004 27356 60014 27412
rect 71922 27356 71932 27412
rect 71988 27356 73948 27412
rect 75478 27356 75516 27412
rect 75572 27356 75582 27412
rect 34962 27244 34972 27300
rect 35028 27244 61292 27300
rect 61348 27244 61358 27300
rect 65314 27244 65324 27300
rect 65380 27244 72604 27300
rect 72660 27244 73388 27300
rect 73444 27244 73454 27300
rect 75618 27244 75628 27300
rect 75684 27244 76188 27300
rect 76244 27244 76254 27300
rect 76850 27244 76860 27300
rect 76916 27244 77532 27300
rect 77588 27244 77598 27300
rect 42914 27132 42924 27188
rect 42980 27132 43820 27188
rect 43876 27132 43886 27188
rect 46386 27132 46396 27188
rect 46452 27132 49644 27188
rect 49700 27132 49710 27188
rect 50372 27132 50764 27188
rect 50820 27132 51212 27188
rect 51268 27132 51278 27188
rect 73126 27132 73164 27188
rect 73220 27132 73230 27188
rect 75058 27132 75068 27188
rect 75124 27132 75516 27188
rect 75572 27132 75582 27188
rect 34066 27020 34076 27076
rect 34132 27020 36204 27076
rect 36260 27020 36988 27076
rect 37044 27020 37054 27076
rect 41916 27020 43036 27076
rect 43092 27020 43102 27076
rect 47282 27020 47292 27076
rect 47348 27020 49084 27076
rect 49140 27020 49150 27076
rect 0 26964 800 26992
rect 41916 26964 41972 27020
rect 50372 26964 50428 27132
rect 72370 27020 72380 27076
rect 72436 27020 77756 27076
rect 77812 27020 77822 27076
rect 0 26908 1708 26964
rect 1764 26908 2492 26964
rect 2548 26908 2558 26964
rect 34962 26908 34972 26964
rect 35028 26908 35644 26964
rect 35700 26908 35710 26964
rect 40562 26908 40572 26964
rect 40628 26908 41692 26964
rect 41748 26908 41916 26964
rect 41972 26908 41982 26964
rect 44930 26908 44940 26964
rect 44996 26908 47068 26964
rect 47124 26908 47134 26964
rect 49746 26908 49756 26964
rect 49812 26908 50428 26964
rect 72706 26908 72716 26964
rect 72772 26908 73052 26964
rect 73108 26908 73118 26964
rect 73612 26908 73948 26964
rect 74004 26908 74014 26964
rect 74610 26908 74620 26964
rect 74676 26908 74732 26964
rect 74788 26908 75964 26964
rect 76020 26908 76030 26964
rect 0 26880 800 26908
rect 73612 26852 73668 26908
rect 35410 26796 35420 26852
rect 35476 26796 56196 26852
rect 56690 26796 56700 26852
rect 56756 26796 72380 26852
rect 72436 26796 72446 26852
rect 73602 26796 73612 26852
rect 73668 26796 73678 26852
rect 75506 26796 75516 26852
rect 75572 26796 77924 26852
rect 78082 26796 78092 26852
rect 78148 26796 78540 26852
rect 78596 26796 78606 26852
rect 44146 26684 44156 26740
rect 44212 26684 44828 26740
rect 44884 26684 44894 26740
rect 46022 26684 46060 26740
rect 46116 26684 46126 26740
rect 46834 26684 46844 26740
rect 46900 26684 47740 26740
rect 47796 26684 47806 26740
rect 48850 26684 48860 26740
rect 48916 26684 48926 26740
rect 51174 26684 51212 26740
rect 51268 26684 51278 26740
rect 19826 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20110 26684
rect 48860 26628 48916 26684
rect 50546 26628 50556 26684
rect 50612 26628 50660 26684
rect 50716 26628 50764 26684
rect 50820 26628 50830 26684
rect 56140 26628 56196 26796
rect 77868 26740 77924 26796
rect 62132 26684 74396 26740
rect 74452 26684 74462 26740
rect 75618 26684 75628 26740
rect 75684 26684 76524 26740
rect 76580 26684 77084 26740
rect 77140 26684 77150 26740
rect 77858 26684 77868 26740
rect 77924 26684 77934 26740
rect 62132 26628 62188 26684
rect 26852 26572 46956 26628
rect 47012 26572 47022 26628
rect 48860 26572 49196 26628
rect 49252 26572 49262 26628
rect 56140 26572 62188 26628
rect 73014 26572 73052 26628
rect 73108 26572 73118 26628
rect 26852 26516 26908 26572
rect 79200 26516 80000 26544
rect 2146 26460 2156 26516
rect 2212 26460 26908 26516
rect 35186 26460 35196 26516
rect 35252 26460 35980 26516
rect 36036 26460 36046 26516
rect 41794 26460 41804 26516
rect 41860 26460 42588 26516
rect 42644 26460 42654 26516
rect 43698 26460 43708 26516
rect 43764 26460 44604 26516
rect 44660 26460 44670 26516
rect 47506 26460 47516 26516
rect 47572 26460 49308 26516
rect 49364 26460 49374 26516
rect 49522 26460 49532 26516
rect 49588 26460 50428 26516
rect 50484 26460 50494 26516
rect 56690 26460 56700 26516
rect 56756 26460 56766 26516
rect 70886 26460 70924 26516
rect 70980 26460 70990 26516
rect 72370 26460 72380 26516
rect 72436 26460 72716 26516
rect 72772 26460 72782 26516
rect 76738 26460 76748 26516
rect 76804 26460 78764 26516
rect 78820 26460 80000 26516
rect 2034 26348 2044 26404
rect 2100 26348 44380 26404
rect 44436 26348 44940 26404
rect 44996 26348 45006 26404
rect 46050 26348 46060 26404
rect 46116 26348 46732 26404
rect 46788 26348 47628 26404
rect 47684 26348 47694 26404
rect 48850 26348 48860 26404
rect 48916 26348 50092 26404
rect 50148 26348 50158 26404
rect 39890 26236 39900 26292
rect 39956 26236 41020 26292
rect 41076 26236 41086 26292
rect 45042 26236 45052 26292
rect 45108 26236 46284 26292
rect 46340 26236 46350 26292
rect 46498 26236 46508 26292
rect 46564 26236 48748 26292
rect 48804 26236 48814 26292
rect 56700 26180 56756 26460
rect 79200 26432 80000 26460
rect 69542 26348 69580 26404
rect 69636 26348 69646 26404
rect 71250 26348 71260 26404
rect 71316 26348 76132 26404
rect 76290 26348 76300 26404
rect 76356 26348 77420 26404
rect 77476 26348 77486 26404
rect 76076 26292 76132 26348
rect 63074 26236 63084 26292
rect 63140 26236 72380 26292
rect 72436 26236 72446 26292
rect 72604 26236 73836 26292
rect 73892 26236 73902 26292
rect 76076 26236 78092 26292
rect 78148 26236 78158 26292
rect 72604 26180 72660 26236
rect 38322 26124 38332 26180
rect 38388 26124 38398 26180
rect 38882 26124 38892 26180
rect 38948 26124 56756 26180
rect 63858 26124 63868 26180
rect 63924 26124 72660 26180
rect 72930 26124 72940 26180
rect 72996 26124 78204 26180
rect 78260 26124 78270 26180
rect 38332 25956 38388 26124
rect 68786 26012 68796 26068
rect 68852 26012 73276 26068
rect 73332 26012 73500 26068
rect 73556 26012 73566 26068
rect 73826 26012 73836 26068
rect 73892 26012 74060 26068
rect 74116 26012 74126 26068
rect 75618 26012 75628 26068
rect 75684 26012 75694 26068
rect 75628 25956 75684 26012
rect 38332 25900 38444 25956
rect 38500 25900 38510 25956
rect 71138 25900 71148 25956
rect 71204 25900 75684 25956
rect 0 25844 800 25872
rect 4466 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4750 25900
rect 35186 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35470 25900
rect 65906 25844 65916 25900
rect 65972 25844 66020 25900
rect 66076 25844 66124 25900
rect 66180 25844 66190 25900
rect 0 25788 1708 25844
rect 1764 25788 2492 25844
rect 2548 25788 2558 25844
rect 38322 25788 38332 25844
rect 38388 25788 38668 25844
rect 38724 25788 38734 25844
rect 44818 25788 44828 25844
rect 44884 25788 47516 25844
rect 47572 25788 47582 25844
rect 0 25760 800 25788
rect 37314 25676 37324 25732
rect 37380 25676 40348 25732
rect 40404 25676 41916 25732
rect 41972 25676 41982 25732
rect 45378 25676 45388 25732
rect 45444 25676 45724 25732
rect 45780 25676 45790 25732
rect 46946 25676 46956 25732
rect 47012 25676 47964 25732
rect 48020 25676 48030 25732
rect 60162 25676 60172 25732
rect 60228 25676 74172 25732
rect 74228 25676 74238 25732
rect 77074 25676 77084 25732
rect 77140 25676 77756 25732
rect 77812 25676 77822 25732
rect 37762 25564 37772 25620
rect 37828 25564 38780 25620
rect 38836 25564 38846 25620
rect 43698 25564 43708 25620
rect 43764 25564 44044 25620
rect 44100 25564 63308 25620
rect 63364 25564 63374 25620
rect 74274 25564 74284 25620
rect 74340 25564 75964 25620
rect 76020 25564 76030 25620
rect 35522 25452 35532 25508
rect 35588 25452 40348 25508
rect 40404 25452 40414 25508
rect 41794 25452 41804 25508
rect 41860 25452 42364 25508
rect 42420 25452 42430 25508
rect 43362 25452 43372 25508
rect 43428 25452 44156 25508
rect 44212 25452 45724 25508
rect 45780 25452 45790 25508
rect 72258 25452 72268 25508
rect 72324 25452 73276 25508
rect 73332 25452 73342 25508
rect 75506 25452 75516 25508
rect 75572 25452 76188 25508
rect 76244 25452 76254 25508
rect 79200 25396 80000 25424
rect 36418 25340 36428 25396
rect 36484 25340 37324 25396
rect 37380 25340 40236 25396
rect 40292 25340 41692 25396
rect 41748 25340 41758 25396
rect 43026 25340 43036 25396
rect 43092 25340 44940 25396
rect 44996 25340 45006 25396
rect 71362 25340 71372 25396
rect 71428 25340 73948 25396
rect 74834 25340 74844 25396
rect 74900 25340 75404 25396
rect 75460 25340 75470 25396
rect 78194 25340 78204 25396
rect 78260 25340 80000 25396
rect 73892 25284 73948 25340
rect 79200 25312 80000 25340
rect 13458 25228 13468 25284
rect 13524 25228 23660 25284
rect 23716 25228 24108 25284
rect 24164 25228 24174 25284
rect 39442 25228 39452 25284
rect 39508 25228 43596 25284
rect 43652 25228 43662 25284
rect 43820 25228 71036 25284
rect 71092 25228 71102 25284
rect 73892 25228 77644 25284
rect 77700 25228 77710 25284
rect 43820 25172 43876 25228
rect 43362 25116 43372 25172
rect 43428 25116 43876 25172
rect 46274 25116 46284 25172
rect 46340 25116 46956 25172
rect 47012 25116 47292 25172
rect 47348 25116 47358 25172
rect 63186 25116 63196 25172
rect 63252 25116 63980 25172
rect 64036 25116 71148 25172
rect 71204 25116 71214 25172
rect 72146 25116 72156 25172
rect 72212 25116 77196 25172
rect 77252 25116 77262 25172
rect 19826 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20110 25116
rect 46284 25060 46340 25116
rect 50546 25060 50556 25116
rect 50612 25060 50660 25116
rect 50716 25060 50764 25116
rect 50820 25060 50830 25116
rect 24322 25004 24332 25060
rect 24388 25004 25228 25060
rect 25284 25004 25294 25060
rect 45938 25004 45948 25060
rect 46004 25004 46340 25060
rect 30268 24892 35420 24948
rect 35476 24892 35486 24948
rect 38612 24892 44044 24948
rect 44100 24892 44110 24948
rect 45266 24892 45276 24948
rect 45332 24892 46508 24948
rect 46564 24892 48188 24948
rect 48244 24892 48254 24948
rect 48626 24892 48636 24948
rect 48692 24892 51100 24948
rect 51156 24892 51166 24948
rect 63746 24892 63756 24948
rect 63812 24892 71708 24948
rect 71764 24892 72156 24948
rect 72212 24892 72222 24948
rect 14242 24780 14252 24836
rect 14308 24780 14812 24836
rect 14868 24780 17164 24836
rect 17220 24780 17230 24836
rect 0 24724 800 24752
rect 0 24668 1708 24724
rect 1764 24668 2492 24724
rect 2548 24668 2558 24724
rect 16594 24668 16604 24724
rect 16660 24668 17500 24724
rect 17556 24668 20636 24724
rect 20692 24668 20702 24724
rect 25554 24668 25564 24724
rect 25620 24668 27020 24724
rect 27076 24668 28476 24724
rect 28532 24668 28542 24724
rect 0 24640 800 24668
rect 30268 24612 30324 24892
rect 38612 24836 38668 24892
rect 31826 24780 31836 24836
rect 31892 24780 38668 24836
rect 30482 24668 30492 24724
rect 30548 24668 37884 24724
rect 37940 24668 37950 24724
rect 47730 24668 47740 24724
rect 47796 24668 48860 24724
rect 48916 24668 70812 24724
rect 70868 24668 70878 24724
rect 73490 24668 73500 24724
rect 73556 24668 76524 24724
rect 76580 24668 76590 24724
rect 17602 24556 17612 24612
rect 17668 24556 18172 24612
rect 18228 24556 18238 24612
rect 18386 24556 18396 24612
rect 18452 24556 18490 24612
rect 24994 24556 25004 24612
rect 25060 24556 25676 24612
rect 25732 24556 25742 24612
rect 26852 24556 30324 24612
rect 33170 24556 33180 24612
rect 33236 24556 37436 24612
rect 37492 24556 37502 24612
rect 71362 24556 71372 24612
rect 71428 24556 76076 24612
rect 76132 24556 76142 24612
rect 12450 24444 12460 24500
rect 12516 24444 23324 24500
rect 23380 24444 23390 24500
rect 4466 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4750 24332
rect 26852 24276 26908 24556
rect 43586 24444 43596 24500
rect 43652 24444 45612 24500
rect 45668 24444 45678 24500
rect 61282 24444 61292 24500
rect 61348 24444 72380 24500
rect 72436 24444 72446 24500
rect 37202 24332 37212 24388
rect 37268 24332 38892 24388
rect 38948 24332 38958 24388
rect 71334 24332 71372 24388
rect 71428 24332 71438 24388
rect 35186 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35470 24332
rect 65906 24276 65916 24332
rect 65972 24276 66020 24332
rect 66076 24276 66124 24332
rect 66180 24276 66190 24332
rect 79200 24276 80000 24304
rect 17714 24220 17724 24276
rect 17780 24220 18396 24276
rect 18452 24220 19740 24276
rect 19796 24220 26908 24276
rect 37874 24220 37884 24276
rect 37940 24220 43596 24276
rect 43652 24220 43662 24276
rect 44146 24220 44156 24276
rect 44212 24220 48300 24276
rect 48356 24220 48366 24276
rect 74386 24220 74396 24276
rect 74452 24220 74620 24276
rect 74676 24220 80000 24276
rect 79200 24192 80000 24220
rect 37762 24108 37772 24164
rect 37828 24108 63308 24164
rect 63364 24108 63374 24164
rect 74722 24108 74732 24164
rect 74788 24108 75292 24164
rect 75348 24108 76188 24164
rect 76244 24108 76254 24164
rect 2034 23996 2044 24052
rect 2100 23996 38668 24052
rect 39778 23996 39788 24052
rect 39844 23996 41020 24052
rect 41076 23996 41086 24052
rect 41346 23996 41356 24052
rect 41412 23996 41692 24052
rect 41748 23996 41758 24052
rect 43698 23996 43708 24052
rect 43764 23996 47908 24052
rect 38612 23940 38668 23996
rect 47852 23940 47908 23996
rect 18022 23884 18060 23940
rect 18116 23884 18126 23940
rect 20738 23884 20748 23940
rect 20804 23884 21196 23940
rect 21252 23884 21262 23940
rect 23986 23884 23996 23940
rect 24052 23884 27468 23940
rect 27524 23884 27534 23940
rect 34738 23884 34748 23940
rect 34804 23884 37212 23940
rect 37268 23884 37278 23940
rect 38612 23884 41188 23940
rect 42018 23884 42028 23940
rect 42084 23884 42700 23940
rect 42756 23884 42766 23940
rect 43652 23884 45444 23940
rect 47842 23884 47852 23940
rect 47908 23884 50428 23940
rect 73238 23884 73276 23940
rect 73332 23884 73342 23940
rect 73602 23884 73612 23940
rect 73668 23884 75404 23940
rect 75460 23884 75470 23940
rect 76066 23884 76076 23940
rect 76132 23884 78316 23940
rect 78372 23884 78382 23940
rect 41132 23828 41188 23884
rect 43652 23828 43708 23884
rect 45388 23828 45444 23884
rect 50372 23828 50428 23884
rect 17154 23772 17164 23828
rect 17220 23772 18508 23828
rect 18564 23772 18574 23828
rect 18722 23772 18732 23828
rect 18788 23772 19516 23828
rect 19572 23772 20412 23828
rect 20468 23772 20478 23828
rect 27906 23772 27916 23828
rect 27972 23772 30492 23828
rect 30548 23772 30558 23828
rect 35634 23772 35644 23828
rect 35700 23772 37772 23828
rect 37828 23772 37838 23828
rect 41132 23772 43708 23828
rect 44818 23772 44828 23828
rect 44884 23772 44894 23828
rect 45378 23772 45388 23828
rect 45444 23772 48748 23828
rect 48804 23772 48814 23828
rect 50372 23772 74172 23828
rect 74228 23772 74238 23828
rect 74610 23772 74620 23828
rect 74676 23772 76524 23828
rect 76580 23772 76860 23828
rect 76916 23772 76926 23828
rect 44828 23716 44884 23772
rect 17938 23660 17948 23716
rect 18004 23660 18396 23716
rect 18452 23660 18462 23716
rect 19404 23660 20524 23716
rect 20580 23660 20590 23716
rect 21634 23660 21644 23716
rect 21700 23660 22316 23716
rect 22372 23660 24220 23716
rect 24276 23660 35084 23716
rect 35140 23660 40348 23716
rect 40404 23660 40414 23716
rect 43652 23660 44884 23716
rect 45490 23660 45500 23716
rect 45556 23660 46060 23716
rect 46116 23660 46126 23716
rect 46386 23660 46396 23716
rect 46452 23660 47068 23716
rect 47124 23660 47134 23716
rect 47506 23660 47516 23716
rect 47572 23660 49644 23716
rect 49700 23660 49868 23716
rect 49924 23660 49934 23716
rect 60610 23660 60620 23716
rect 60676 23660 72156 23716
rect 72212 23660 72222 23716
rect 74834 23660 74844 23716
rect 74900 23660 78204 23716
rect 78260 23660 78270 23716
rect 0 23604 800 23632
rect 19404 23604 19460 23660
rect 43652 23604 43708 23660
rect 0 23548 1708 23604
rect 1764 23548 2492 23604
rect 2548 23548 2558 23604
rect 11554 23548 11564 23604
rect 11620 23548 13468 23604
rect 13524 23548 13534 23604
rect 13794 23548 13804 23604
rect 13860 23548 16268 23604
rect 16324 23548 19404 23604
rect 19460 23548 19470 23604
rect 34290 23548 34300 23604
rect 34356 23548 35980 23604
rect 36036 23548 36540 23604
rect 36596 23548 36606 23604
rect 36754 23548 36764 23604
rect 36820 23548 37660 23604
rect 37716 23548 37726 23604
rect 39442 23548 39452 23604
rect 39508 23548 40460 23604
rect 40516 23548 40526 23604
rect 40684 23548 43708 23604
rect 44930 23548 44940 23604
rect 44996 23548 49420 23604
rect 49476 23548 49486 23604
rect 63410 23548 63420 23604
rect 63476 23548 78092 23604
rect 78148 23548 78158 23604
rect 0 23520 800 23548
rect 19826 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20110 23548
rect 2146 23436 2156 23492
rect 2212 23436 3388 23492
rect 17602 23436 17612 23492
rect 17668 23436 18620 23492
rect 18676 23436 18686 23492
rect 26852 23436 40460 23492
rect 40516 23436 40526 23492
rect 3332 23380 3388 23436
rect 26852 23380 26908 23436
rect 40684 23380 40740 23548
rect 50546 23492 50556 23548
rect 50612 23492 50660 23548
rect 50716 23492 50764 23548
rect 50820 23492 50830 23548
rect 40898 23436 40908 23492
rect 40964 23436 44828 23492
rect 44884 23436 44894 23492
rect 50054 23436 50092 23492
rect 50148 23436 50158 23492
rect 51762 23436 51772 23492
rect 51828 23436 55916 23492
rect 55972 23436 55982 23492
rect 3332 23324 26908 23380
rect 27570 23324 27580 23380
rect 27636 23324 28140 23380
rect 28196 23324 28206 23380
rect 28466 23324 28476 23380
rect 28532 23324 37660 23380
rect 37716 23324 37726 23380
rect 38098 23324 38108 23380
rect 38164 23324 40740 23380
rect 41570 23324 41580 23380
rect 41636 23324 42028 23380
rect 42084 23324 42094 23380
rect 42588 23324 43372 23380
rect 43428 23324 43438 23380
rect 43586 23324 43596 23380
rect 43652 23324 47180 23380
rect 47236 23324 47246 23380
rect 69458 23324 69468 23380
rect 69524 23324 71708 23380
rect 71764 23324 72156 23380
rect 72212 23324 72222 23380
rect 73826 23324 73836 23380
rect 73892 23324 77868 23380
rect 77924 23324 77934 23380
rect 27580 23268 27636 23324
rect 42588 23268 42644 23324
rect 16818 23212 16828 23268
rect 16884 23212 17500 23268
rect 17556 23212 17566 23268
rect 24098 23212 24108 23268
rect 24164 23212 25844 23268
rect 26002 23212 26012 23268
rect 26068 23212 27636 23268
rect 29922 23212 29932 23268
rect 29988 23212 39172 23268
rect 39330 23212 39340 23268
rect 39396 23212 40124 23268
rect 40180 23212 41244 23268
rect 41300 23212 41310 23268
rect 41682 23212 41692 23268
rect 41748 23212 42644 23268
rect 42802 23212 42812 23268
rect 42868 23212 48916 23268
rect 63522 23212 63532 23268
rect 63588 23212 77196 23268
rect 77252 23212 77262 23268
rect 25788 23156 25844 23212
rect 39116 23156 39172 23212
rect 48860 23156 48916 23212
rect 79200 23156 80000 23184
rect 12786 23100 12796 23156
rect 12852 23100 23996 23156
rect 24052 23100 24062 23156
rect 24210 23100 24220 23156
rect 24276 23100 25116 23156
rect 25172 23100 25182 23156
rect 25554 23100 25564 23156
rect 25620 23100 25630 23156
rect 25788 23100 26908 23156
rect 26964 23100 26974 23156
rect 34178 23100 34188 23156
rect 34244 23100 34860 23156
rect 34916 23100 34926 23156
rect 35298 23100 35308 23156
rect 35364 23100 35756 23156
rect 35812 23100 35822 23156
rect 39116 23100 40908 23156
rect 40964 23100 41804 23156
rect 41860 23100 41870 23156
rect 42466 23100 42476 23156
rect 42532 23100 43596 23156
rect 43652 23100 43662 23156
rect 44034 23100 44044 23156
rect 44100 23100 45612 23156
rect 45668 23100 45678 23156
rect 46022 23100 46060 23156
rect 46116 23100 46126 23156
rect 46386 23100 46396 23156
rect 46452 23100 47852 23156
rect 47908 23100 47918 23156
rect 48850 23100 48860 23156
rect 48916 23100 57484 23156
rect 57540 23100 57550 23156
rect 68674 23100 68684 23156
rect 68740 23100 71708 23156
rect 71764 23100 71774 23156
rect 78194 23100 78204 23156
rect 78260 23100 80000 23156
rect 23996 23044 24052 23100
rect 1698 22988 1708 23044
rect 1764 22988 2492 23044
rect 2548 22988 2558 23044
rect 19170 22988 19180 23044
rect 19236 22988 19628 23044
rect 19684 22988 19694 23044
rect 23996 22988 24556 23044
rect 24612 22988 24622 23044
rect 25564 22932 25620 23100
rect 79200 23072 80000 23100
rect 27458 22988 27468 23044
rect 27524 22988 28700 23044
rect 28756 22988 28766 23044
rect 33394 22988 33404 23044
rect 33460 22988 42252 23044
rect 42308 22988 42318 23044
rect 45826 22988 45836 23044
rect 45892 22988 46284 23044
rect 46340 22988 46350 23044
rect 48066 22988 48076 23044
rect 48132 22988 49868 23044
rect 49924 22988 70700 23044
rect 70756 22988 70766 23044
rect 2034 22876 2044 22932
rect 2100 22876 15148 22932
rect 25564 22876 27132 22932
rect 27188 22876 27198 22932
rect 35522 22876 35532 22932
rect 35588 22876 36204 22932
rect 36260 22876 36270 22932
rect 37426 22876 37436 22932
rect 37492 22876 38556 22932
rect 38612 22876 38622 22932
rect 41346 22876 41356 22932
rect 41412 22876 41692 22932
rect 41748 22876 41758 22932
rect 44258 22876 44268 22932
rect 44324 22876 46060 22932
rect 46116 22876 46126 22932
rect 49410 22876 49420 22932
rect 49476 22876 75068 22932
rect 75124 22876 75134 22932
rect 15092 22820 15148 22876
rect 15092 22764 31836 22820
rect 31892 22764 31902 22820
rect 41234 22764 41244 22820
rect 41300 22764 43596 22820
rect 43652 22764 45388 22820
rect 45444 22764 45454 22820
rect 45948 22764 49308 22820
rect 49364 22764 49374 22820
rect 4466 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4750 22764
rect 35186 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35470 22764
rect 45948 22708 46004 22764
rect 65906 22708 65916 22764
rect 65972 22708 66020 22764
rect 66076 22708 66124 22764
rect 66180 22708 66190 22764
rect 38546 22652 38556 22708
rect 38612 22652 40348 22708
rect 40404 22652 40414 22708
rect 40898 22652 40908 22708
rect 40964 22652 43372 22708
rect 43428 22652 44660 22708
rect 44818 22652 44828 22708
rect 44884 22652 46004 22708
rect 47058 22652 47068 22708
rect 47124 22652 47516 22708
rect 47572 22652 47908 22708
rect 48066 22652 48076 22708
rect 48132 22652 50428 22708
rect 50484 22652 62188 22708
rect 66882 22652 66892 22708
rect 66948 22652 70924 22708
rect 70980 22652 70990 22708
rect 44604 22596 44660 22652
rect 47852 22596 47908 22652
rect 62132 22596 62188 22652
rect 30146 22540 30156 22596
rect 30212 22540 44156 22596
rect 44212 22540 44222 22596
rect 44604 22540 45276 22596
rect 45332 22540 45342 22596
rect 47852 22540 49868 22596
rect 49924 22540 52780 22596
rect 52836 22540 52846 22596
rect 62132 22540 70588 22596
rect 70644 22540 70654 22596
rect 0 22484 800 22512
rect 0 22428 1708 22484
rect 1764 22428 1774 22484
rect 19394 22428 19404 22484
rect 19460 22428 20412 22484
rect 20468 22428 20478 22484
rect 40562 22428 40572 22484
rect 40628 22428 50428 22484
rect 53218 22428 53228 22484
rect 53284 22428 54236 22484
rect 54292 22428 54302 22484
rect 67666 22428 67676 22484
rect 67732 22428 72156 22484
rect 72212 22428 72222 22484
rect 76710 22428 76748 22484
rect 76804 22428 76814 22484
rect 0 22400 800 22428
rect 19842 22316 19852 22372
rect 19908 22316 21196 22372
rect 21252 22316 21262 22372
rect 27682 22316 27692 22372
rect 27748 22316 30940 22372
rect 30996 22316 35308 22372
rect 35364 22316 35374 22372
rect 35746 22316 35756 22372
rect 35812 22316 37324 22372
rect 37380 22316 37390 22372
rect 37762 22316 37772 22372
rect 37828 22316 39788 22372
rect 39844 22316 39854 22372
rect 46610 22316 46620 22372
rect 46676 22316 47404 22372
rect 47460 22316 47628 22372
rect 47684 22316 47694 22372
rect 49074 22316 49084 22372
rect 49140 22316 49150 22372
rect 38322 22204 38332 22260
rect 38388 22204 41244 22260
rect 41300 22204 41310 22260
rect 41794 22204 41804 22260
rect 41860 22204 42588 22260
rect 42644 22204 44324 22260
rect 44930 22204 44940 22260
rect 44996 22204 47068 22260
rect 47124 22204 47134 22260
rect 44268 22148 44324 22204
rect 49084 22148 49140 22316
rect 50372 22260 50428 22428
rect 52210 22316 52220 22372
rect 52276 22316 53676 22372
rect 53732 22316 53742 22372
rect 71698 22316 71708 22372
rect 71764 22316 73948 22372
rect 74004 22316 74014 22372
rect 75702 22316 75740 22372
rect 75796 22316 75806 22372
rect 77046 22316 77084 22372
rect 77140 22316 77150 22372
rect 50372 22204 61684 22260
rect 70354 22204 70364 22260
rect 70420 22204 72492 22260
rect 72548 22204 72558 22260
rect 75618 22204 75628 22260
rect 75684 22204 75964 22260
rect 76020 22204 76030 22260
rect 61628 22148 61684 22204
rect 18722 22092 18732 22148
rect 18788 22092 19852 22148
rect 19908 22092 23548 22148
rect 23604 22092 23614 22148
rect 27122 22092 27132 22148
rect 27188 22092 27692 22148
rect 27748 22092 28252 22148
rect 28308 22092 28318 22148
rect 42690 22092 42700 22148
rect 42756 22092 43820 22148
rect 43876 22092 43886 22148
rect 44258 22092 44268 22148
rect 44324 22092 44334 22148
rect 47282 22092 47292 22148
rect 47348 22092 47964 22148
rect 48020 22092 48030 22148
rect 49084 22092 49420 22148
rect 49476 22092 50876 22148
rect 50932 22092 50942 22148
rect 61618 22092 61628 22148
rect 61684 22092 61694 22148
rect 73490 22092 73500 22148
rect 73556 22092 77420 22148
rect 77476 22092 77486 22148
rect 77746 22092 77756 22148
rect 77812 22092 78540 22148
rect 78596 22092 78606 22148
rect 79200 22036 80000 22064
rect 17266 21980 17276 22036
rect 17332 21980 17948 22036
rect 18004 21980 19180 22036
rect 19236 21980 19246 22036
rect 21634 21980 21644 22036
rect 21700 21980 22988 22036
rect 23044 21980 39004 22036
rect 39060 21980 39070 22036
rect 46722 21980 46732 22036
rect 46788 21980 47404 22036
rect 47460 21980 47470 22036
rect 47618 21980 47628 22036
rect 47684 21980 47722 22036
rect 73602 21980 73612 22036
rect 73668 21980 77308 22036
rect 77364 21980 77374 22036
rect 78082 21980 78092 22036
rect 78148 21980 80000 22036
rect 19826 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20110 21980
rect 50546 21924 50556 21980
rect 50612 21924 50660 21980
rect 50716 21924 50764 21980
rect 50820 21924 50830 21980
rect 79200 21952 80000 21980
rect 22082 21868 22092 21924
rect 22148 21868 24332 21924
rect 24388 21868 24398 21924
rect 32946 21868 32956 21924
rect 33012 21868 36652 21924
rect 36708 21868 36718 21924
rect 39778 21868 39788 21924
rect 39844 21868 40348 21924
rect 40404 21868 41244 21924
rect 41300 21868 41310 21924
rect 42802 21868 42812 21924
rect 42868 21868 44156 21924
rect 44212 21868 44222 21924
rect 45826 21868 45836 21924
rect 45892 21868 49084 21924
rect 49140 21868 49150 21924
rect 51650 21868 51660 21924
rect 51716 21868 53788 21924
rect 53844 21868 53854 21924
rect 74918 21868 74956 21924
rect 75012 21868 75022 21924
rect 75842 21868 75852 21924
rect 75908 21868 76412 21924
rect 76468 21868 76636 21924
rect 76692 21868 76702 21924
rect 2146 21756 2156 21812
rect 2212 21756 46004 21812
rect 48290 21756 48300 21812
rect 48356 21756 48748 21812
rect 48804 21756 48814 21812
rect 54562 21756 54572 21812
rect 54628 21756 56028 21812
rect 56084 21756 56094 21812
rect 65650 21756 65660 21812
rect 65716 21756 70028 21812
rect 70084 21756 70094 21812
rect 45948 21700 46004 21756
rect 11666 21644 11676 21700
rect 11732 21644 15596 21700
rect 15652 21644 15662 21700
rect 21858 21644 21868 21700
rect 21924 21644 22316 21700
rect 22372 21644 22382 21700
rect 24434 21644 24444 21700
rect 24500 21644 25676 21700
rect 25732 21644 25742 21700
rect 41234 21644 41244 21700
rect 41300 21644 42476 21700
rect 42532 21644 42542 21700
rect 45948 21644 48132 21700
rect 48626 21644 48636 21700
rect 48692 21644 49868 21700
rect 49924 21644 50652 21700
rect 50708 21644 50718 21700
rect 54338 21644 54348 21700
rect 54404 21644 55580 21700
rect 55636 21644 55646 21700
rect 62132 21644 67228 21700
rect 67284 21644 67294 21700
rect 75170 21644 75180 21700
rect 75236 21644 76748 21700
rect 76804 21644 76814 21700
rect 78418 21644 78428 21700
rect 78484 21644 78764 21700
rect 78820 21644 78830 21700
rect 21868 21588 21924 21644
rect 48076 21588 48132 21644
rect 17154 21532 17164 21588
rect 17220 21532 17948 21588
rect 18004 21532 21924 21588
rect 34738 21532 34748 21588
rect 34804 21532 35084 21588
rect 35140 21532 35150 21588
rect 35746 21532 35756 21588
rect 35812 21532 36540 21588
rect 36596 21532 36606 21588
rect 39452 21532 45836 21588
rect 45892 21532 45902 21588
rect 46162 21532 46172 21588
rect 46228 21532 46956 21588
rect 47012 21532 47022 21588
rect 48066 21532 48076 21588
rect 48132 21532 48142 21588
rect 49074 21532 49084 21588
rect 49140 21532 51660 21588
rect 51716 21532 53116 21588
rect 53172 21532 53182 21588
rect 53452 21532 61348 21588
rect 15586 21420 15596 21476
rect 15652 21420 23548 21476
rect 23604 21420 23996 21476
rect 24052 21420 24062 21476
rect 34486 21420 34524 21476
rect 34580 21420 34590 21476
rect 34860 21420 39228 21476
rect 39284 21420 39294 21476
rect 0 21364 800 21392
rect 34860 21364 34916 21420
rect 39452 21364 39508 21532
rect 46172 21476 46228 21532
rect 53452 21476 53508 21532
rect 61292 21476 61348 21532
rect 43250 21420 43260 21476
rect 43316 21420 44492 21476
rect 44548 21420 46228 21476
rect 46610 21420 46620 21476
rect 46676 21420 53508 21476
rect 53666 21420 53676 21476
rect 53732 21420 54460 21476
rect 54516 21420 54526 21476
rect 61282 21420 61292 21476
rect 61348 21420 61358 21476
rect 62132 21364 62188 21644
rect 66434 21532 66444 21588
rect 66500 21532 73276 21588
rect 73332 21532 74060 21588
rect 74116 21532 74126 21588
rect 74274 21532 74284 21588
rect 74340 21532 75516 21588
rect 75572 21532 75582 21588
rect 71586 21420 71596 21476
rect 71652 21420 75292 21476
rect 75348 21420 75358 21476
rect 0 21308 1708 21364
rect 1764 21308 2492 21364
rect 2548 21308 2558 21364
rect 17714 21308 17724 21364
rect 17780 21308 18396 21364
rect 18452 21308 20748 21364
rect 20804 21308 34860 21364
rect 34916 21308 34926 21364
rect 35298 21308 35308 21364
rect 35364 21308 36204 21364
rect 36260 21308 36270 21364
rect 38612 21308 39508 21364
rect 46498 21308 46508 21364
rect 46564 21308 50428 21364
rect 52098 21308 52108 21364
rect 52164 21308 62188 21364
rect 0 21280 800 21308
rect 4466 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4750 21196
rect 35186 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35470 21196
rect 35410 20972 35420 21028
rect 35476 20972 35980 21028
rect 36036 20972 36046 21028
rect 38612 20916 38668 21308
rect 50372 21252 50428 21308
rect 45266 21196 45276 21252
rect 45332 21196 47068 21252
rect 47124 21196 47134 21252
rect 50372 21196 63420 21252
rect 63476 21196 63486 21252
rect 65906 21140 65916 21196
rect 65972 21140 66020 21196
rect 66076 21140 66124 21196
rect 66180 21140 66190 21196
rect 42914 21084 42924 21140
rect 42980 21084 63644 21140
rect 63700 21084 63710 21140
rect 47170 20972 47180 21028
rect 47236 20972 47740 21028
rect 47796 20972 47806 21028
rect 50372 20972 74284 21028
rect 74340 20972 74350 21028
rect 50372 20916 50428 20972
rect 79200 20916 80000 20944
rect 31378 20860 31388 20916
rect 31444 20860 33292 20916
rect 33348 20860 38668 20916
rect 43698 20860 43708 20916
rect 43764 20860 50428 20916
rect 51314 20860 51324 20916
rect 51380 20860 51772 20916
rect 51828 20860 51838 20916
rect 53330 20860 53340 20916
rect 53396 20860 54124 20916
rect 54180 20860 54908 20916
rect 54964 20860 55580 20916
rect 55636 20860 55646 20916
rect 56130 20860 56140 20916
rect 56196 20860 57148 20916
rect 57204 20860 57214 20916
rect 67778 20860 67788 20916
rect 67844 20860 72940 20916
rect 72996 20860 73006 20916
rect 74834 20860 74844 20916
rect 74900 20860 80000 20916
rect 51772 20804 51828 20860
rect 79200 20832 80000 20860
rect 18610 20748 18620 20804
rect 18676 20748 19068 20804
rect 19124 20748 20188 20804
rect 20244 20748 20254 20804
rect 23650 20748 23660 20804
rect 23716 20748 24780 20804
rect 24836 20748 25340 20804
rect 25396 20748 25406 20804
rect 26002 20748 26012 20804
rect 26068 20748 27244 20804
rect 27300 20748 27310 20804
rect 34850 20748 34860 20804
rect 34916 20748 35756 20804
rect 35812 20748 35822 20804
rect 36418 20748 36428 20804
rect 36484 20748 39004 20804
rect 39060 20748 40124 20804
rect 40180 20748 40190 20804
rect 42018 20748 42028 20804
rect 42084 20748 42924 20804
rect 42980 20748 42990 20804
rect 44818 20748 44828 20804
rect 44884 20748 46620 20804
rect 46676 20748 46686 20804
rect 47142 20748 47180 20804
rect 47236 20748 48524 20804
rect 48580 20748 48590 20804
rect 48738 20748 48748 20804
rect 48804 20748 49196 20804
rect 49252 20748 49420 20804
rect 49476 20748 49756 20804
rect 49812 20748 50092 20804
rect 50148 20748 50158 20804
rect 51202 20748 51212 20804
rect 51268 20748 51716 20804
rect 51772 20748 53452 20804
rect 53508 20748 53518 20804
rect 66658 20748 66668 20804
rect 66724 20748 72716 20804
rect 72772 20748 72782 20804
rect 76626 20748 76636 20804
rect 76692 20748 77868 20804
rect 77924 20748 77934 20804
rect 26338 20636 26348 20692
rect 26404 20636 29036 20692
rect 29092 20636 29102 20692
rect 33506 20636 33516 20692
rect 33572 20636 35196 20692
rect 35252 20636 35262 20692
rect 35522 20636 35532 20692
rect 35588 20636 36540 20692
rect 36596 20636 36988 20692
rect 37044 20636 37054 20692
rect 40002 20636 40012 20692
rect 40068 20636 40460 20692
rect 40516 20636 40908 20692
rect 40964 20636 40974 20692
rect 35532 20580 35588 20636
rect 51660 20580 51716 20748
rect 54450 20636 54460 20692
rect 54516 20636 55244 20692
rect 55300 20636 56252 20692
rect 56308 20636 56318 20692
rect 63746 20636 63756 20692
rect 63812 20636 71260 20692
rect 71316 20636 71326 20692
rect 24882 20524 24892 20580
rect 24948 20524 25564 20580
rect 25620 20524 26124 20580
rect 26180 20524 26190 20580
rect 26674 20524 26684 20580
rect 26740 20524 27356 20580
rect 27412 20524 27916 20580
rect 27972 20524 27982 20580
rect 28466 20524 28476 20580
rect 28532 20524 29596 20580
rect 29652 20524 29662 20580
rect 34972 20524 35588 20580
rect 37314 20524 37324 20580
rect 37380 20524 39676 20580
rect 39732 20524 40572 20580
rect 40628 20524 40638 20580
rect 51650 20524 51660 20580
rect 51716 20524 51726 20580
rect 75058 20524 75068 20580
rect 75124 20524 76972 20580
rect 77028 20524 77038 20580
rect 26684 20468 26740 20524
rect 34972 20468 35028 20524
rect 19058 20412 19068 20468
rect 19124 20412 19404 20468
rect 19460 20412 19470 20468
rect 25890 20412 25900 20468
rect 25956 20412 26740 20468
rect 34626 20412 34636 20468
rect 34692 20412 35028 20468
rect 35634 20412 35644 20468
rect 35700 20412 39564 20468
rect 39620 20412 39630 20468
rect 40674 20412 40684 20468
rect 40740 20412 42140 20468
rect 42196 20412 43596 20468
rect 43652 20412 43662 20468
rect 19826 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20110 20412
rect 50546 20356 50556 20412
rect 50612 20356 50660 20412
rect 50716 20356 50764 20412
rect 50820 20356 50830 20412
rect 2034 20300 2044 20356
rect 2100 20300 3388 20356
rect 48402 20300 48412 20356
rect 48468 20300 49756 20356
rect 49812 20300 49822 20356
rect 0 20244 800 20272
rect 3332 20244 3388 20300
rect 0 20188 1708 20244
rect 1764 20188 2492 20244
rect 2548 20188 2558 20244
rect 3332 20188 33012 20244
rect 34402 20188 34412 20244
rect 34468 20188 34748 20244
rect 34804 20188 34814 20244
rect 38770 20188 38780 20244
rect 38836 20188 45724 20244
rect 45780 20188 45790 20244
rect 53554 20188 53564 20244
rect 53620 20188 54348 20244
rect 54404 20188 54414 20244
rect 68898 20188 68908 20244
rect 68964 20188 72380 20244
rect 72436 20188 72446 20244
rect 77644 20188 78204 20244
rect 78260 20188 78270 20244
rect 0 20160 800 20188
rect 32956 20132 33012 20188
rect 18386 20076 18396 20132
rect 18452 20076 18956 20132
rect 19012 20076 19022 20132
rect 22642 20076 22652 20132
rect 22708 20076 23212 20132
rect 23268 20076 26348 20132
rect 26404 20076 26908 20132
rect 26964 20076 26974 20132
rect 27570 20076 27580 20132
rect 27636 20076 30940 20132
rect 30996 20076 31006 20132
rect 32956 20076 35308 20132
rect 35364 20076 35374 20132
rect 35522 20076 35532 20132
rect 35588 20076 37884 20132
rect 37940 20076 37950 20132
rect 41346 20076 41356 20132
rect 41412 20076 41916 20132
rect 41972 20076 41982 20132
rect 43474 20076 43484 20132
rect 43540 20076 44492 20132
rect 44548 20076 44558 20132
rect 49410 20076 49420 20132
rect 49476 20076 50876 20132
rect 50932 20076 50942 20132
rect 54786 20076 54796 20132
rect 54852 20076 56700 20132
rect 56756 20076 56766 20132
rect 73826 20076 73836 20132
rect 73892 20076 76188 20132
rect 76244 20076 76254 20132
rect 27122 19964 27132 20020
rect 27188 19964 27692 20020
rect 27748 19964 29708 20020
rect 29764 19964 31612 20020
rect 31668 19964 31678 20020
rect 34514 19964 34524 20020
rect 34580 19964 34748 20020
rect 34804 19964 34814 20020
rect 35410 19964 35420 20020
rect 35476 19964 36428 20020
rect 36484 19964 36494 20020
rect 40674 19964 40684 20020
rect 40740 19964 41132 20020
rect 41188 19964 41198 20020
rect 46610 19964 46620 20020
rect 46676 19964 48860 20020
rect 48916 19964 48926 20020
rect 50054 19964 50092 20020
rect 50148 19964 50158 20020
rect 52546 19964 52556 20020
rect 52612 19964 53340 20020
rect 53396 19964 55804 20020
rect 55860 19964 55870 20020
rect 75618 19964 75628 20020
rect 75684 19964 76076 20020
rect 76132 19964 76636 20020
rect 76692 19964 77084 20020
rect 77140 19964 77420 20020
rect 77476 19964 77486 20020
rect 77644 19908 77700 20188
rect 19170 19852 19180 19908
rect 19236 19852 19628 19908
rect 19684 19852 20300 19908
rect 20356 19852 20366 19908
rect 24658 19852 24668 19908
rect 24724 19852 27468 19908
rect 27524 19852 27534 19908
rect 32610 19852 32620 19908
rect 32676 19852 34300 19908
rect 34356 19852 34366 19908
rect 34636 19852 47068 19908
rect 47124 19852 47134 19908
rect 48178 19852 48188 19908
rect 48244 19852 50204 19908
rect 50260 19852 50270 19908
rect 50866 19852 50876 19908
rect 50932 19852 51324 19908
rect 51380 19852 51390 19908
rect 51762 19852 51772 19908
rect 51828 19852 67900 19908
rect 67956 19852 67966 19908
rect 77634 19852 77644 19908
rect 77700 19852 77710 19908
rect 7522 19740 7532 19796
rect 7588 19740 32172 19796
rect 32228 19740 33852 19796
rect 33908 19740 33918 19796
rect 34636 19684 34692 19852
rect 79200 19796 80000 19824
rect 33730 19628 33740 19684
rect 33796 19628 34692 19684
rect 34748 19740 37996 19796
rect 38052 19740 38062 19796
rect 38612 19740 43708 19796
rect 43922 19740 43932 19796
rect 43988 19740 60172 19796
rect 60228 19740 60238 19796
rect 78194 19740 78204 19796
rect 78260 19740 80000 19796
rect 4466 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4750 19628
rect 34748 19572 34804 19740
rect 38612 19684 38668 19740
rect 43652 19684 43708 19740
rect 79200 19712 80000 19740
rect 35746 19628 35756 19684
rect 35812 19628 38668 19684
rect 40786 19628 40796 19684
rect 40852 19628 41244 19684
rect 41300 19628 41310 19684
rect 43652 19628 51436 19684
rect 51492 19628 51502 19684
rect 35186 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35470 19628
rect 65906 19572 65916 19628
rect 65972 19572 66020 19628
rect 66076 19572 66124 19628
rect 66180 19572 66190 19628
rect 19394 19516 19404 19572
rect 19460 19516 24444 19572
rect 24500 19516 24510 19572
rect 28242 19516 28252 19572
rect 28308 19516 34804 19572
rect 36418 19516 36428 19572
rect 36484 19516 41580 19572
rect 41636 19516 41646 19572
rect 55010 19516 55020 19572
rect 55076 19516 56588 19572
rect 56644 19516 56654 19572
rect 21746 19404 21756 19460
rect 21812 19404 22988 19460
rect 23044 19404 25564 19460
rect 25620 19404 28756 19460
rect 22530 19292 22540 19348
rect 22596 19292 25452 19348
rect 25508 19292 26460 19348
rect 26516 19292 26526 19348
rect 28700 19236 28756 19404
rect 31612 19404 41804 19460
rect 41860 19404 43372 19460
rect 43428 19404 43438 19460
rect 73042 19404 73052 19460
rect 73108 19404 77588 19460
rect 20402 19180 20412 19236
rect 20468 19180 20748 19236
rect 20804 19180 21980 19236
rect 22036 19180 22652 19236
rect 22708 19180 22718 19236
rect 27458 19180 27468 19236
rect 27524 19180 28476 19236
rect 28532 19180 28542 19236
rect 28690 19180 28700 19236
rect 28756 19180 28766 19236
rect 0 19124 800 19152
rect 0 19068 1708 19124
rect 1764 19068 2492 19124
rect 2548 19068 2558 19124
rect 21410 19068 21420 19124
rect 21476 19068 23548 19124
rect 23604 19068 23614 19124
rect 25106 19068 25116 19124
rect 25172 19068 25788 19124
rect 25844 19068 25854 19124
rect 27794 19068 27804 19124
rect 27860 19068 28700 19124
rect 28756 19068 30268 19124
rect 30324 19068 30828 19124
rect 30884 19068 30894 19124
rect 0 19040 800 19068
rect 19506 18956 19516 19012
rect 19572 18956 23100 19012
rect 23156 18956 23166 19012
rect 24434 18956 24444 19012
rect 24500 18956 26460 19012
rect 26516 18956 26526 19012
rect 27458 18956 27468 19012
rect 27524 18956 28140 19012
rect 28196 18956 29484 19012
rect 29540 18956 29550 19012
rect 31612 18900 31668 19404
rect 31826 19292 31836 19348
rect 31892 19292 35756 19348
rect 35812 19292 35822 19348
rect 38332 19292 39228 19348
rect 39284 19292 39294 19348
rect 41682 19292 41692 19348
rect 41748 19292 42812 19348
rect 42868 19292 70364 19348
rect 70420 19292 70430 19348
rect 75842 19292 75852 19348
rect 75908 19292 76524 19348
rect 76580 19292 76590 19348
rect 38332 19236 38388 19292
rect 37650 19180 37660 19236
rect 37716 19180 38332 19236
rect 38388 19180 38398 19236
rect 38546 19180 38556 19236
rect 38612 19180 39340 19236
rect 39396 19180 39900 19236
rect 39956 19180 39966 19236
rect 40562 19180 40572 19236
rect 40628 19180 41132 19236
rect 41188 19180 41198 19236
rect 72146 19180 72156 19236
rect 72212 19180 76860 19236
rect 76916 19180 76926 19236
rect 34066 19068 34076 19124
rect 34132 19068 35420 19124
rect 35476 19068 35486 19124
rect 39554 19068 39564 19124
rect 39620 19068 40460 19124
rect 40516 19068 40526 19124
rect 51650 19068 51660 19124
rect 51716 19068 52780 19124
rect 52836 19068 53228 19124
rect 53284 19068 53294 19124
rect 54786 19068 54796 19124
rect 54852 19068 55468 19124
rect 55524 19068 55534 19124
rect 56130 19068 56140 19124
rect 56196 19068 57372 19124
rect 57428 19068 57438 19124
rect 77532 19012 77588 19404
rect 35522 18956 35532 19012
rect 35588 18956 36764 19012
rect 36820 18956 36830 19012
rect 39106 18956 39116 19012
rect 39172 18956 41580 19012
rect 41636 18956 41646 19012
rect 41804 18956 67788 19012
rect 67844 18956 67854 19012
rect 77522 18956 77532 19012
rect 77588 18956 77598 19012
rect 41804 18900 41860 18956
rect 20514 18844 20524 18900
rect 20580 18844 21532 18900
rect 21588 18844 23884 18900
rect 23940 18844 31668 18900
rect 36418 18844 36428 18900
rect 36484 18844 37324 18900
rect 37380 18844 37390 18900
rect 40562 18844 40572 18900
rect 40628 18844 41244 18900
rect 41300 18844 41860 18900
rect 43652 18844 46620 18900
rect 46676 18844 46686 18900
rect 76514 18844 76524 18900
rect 76580 18844 78204 18900
rect 78260 18844 78270 18900
rect 19826 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20110 18844
rect 43652 18788 43708 18844
rect 50546 18788 50556 18844
rect 50612 18788 50660 18844
rect 50716 18788 50764 18844
rect 50820 18788 50830 18844
rect 26852 18732 28308 18788
rect 29474 18732 29484 18788
rect 29540 18732 43708 18788
rect 52770 18732 52780 18788
rect 52836 18732 53228 18788
rect 53284 18732 53294 18788
rect 26852 18676 26908 18732
rect 28252 18676 28308 18732
rect 79200 18676 80000 18704
rect 18162 18620 18172 18676
rect 18228 18620 19180 18676
rect 19236 18620 19246 18676
rect 20178 18620 20188 18676
rect 20244 18620 20636 18676
rect 20692 18620 21644 18676
rect 21700 18620 26908 18676
rect 27794 18620 27804 18676
rect 27860 18620 27870 18676
rect 28252 18620 40796 18676
rect 40852 18620 43036 18676
rect 43092 18620 43102 18676
rect 46834 18620 46844 18676
rect 46900 18620 64540 18676
rect 64596 18620 64606 18676
rect 77298 18620 77308 18676
rect 77364 18620 80000 18676
rect 14018 18508 14028 18564
rect 14084 18508 16716 18564
rect 16772 18508 16782 18564
rect 18610 18508 18620 18564
rect 18676 18508 19628 18564
rect 19684 18508 19694 18564
rect 27804 18452 27860 18620
rect 79200 18592 80000 18620
rect 28690 18508 28700 18564
rect 28756 18508 41020 18564
rect 41076 18508 43372 18564
rect 43428 18508 43438 18564
rect 51202 18508 51212 18564
rect 51268 18508 52556 18564
rect 52612 18508 52622 18564
rect 76290 18508 76300 18564
rect 76356 18508 77924 18564
rect 77868 18452 77924 18508
rect 26450 18396 26460 18452
rect 26516 18396 27860 18452
rect 32284 18396 34748 18452
rect 34804 18396 34814 18452
rect 41906 18396 41916 18452
rect 41972 18396 44716 18452
rect 44772 18396 44782 18452
rect 45266 18396 45276 18452
rect 45332 18396 46060 18452
rect 46116 18396 46284 18452
rect 46340 18396 46350 18452
rect 46610 18396 46620 18452
rect 46676 18396 47404 18452
rect 47460 18396 47470 18452
rect 55122 18396 55132 18452
rect 55188 18396 57148 18452
rect 57204 18396 57214 18452
rect 67218 18396 67228 18452
rect 67284 18396 71372 18452
rect 71428 18396 71438 18452
rect 77858 18396 77868 18452
rect 77924 18396 77934 18452
rect 32284 18340 32340 18396
rect 19282 18284 19292 18340
rect 19348 18284 20636 18340
rect 20692 18284 20702 18340
rect 24658 18284 24668 18340
rect 24724 18284 25340 18340
rect 25396 18284 25406 18340
rect 27122 18284 27132 18340
rect 27188 18284 32340 18340
rect 32498 18284 32508 18340
rect 32564 18284 33516 18340
rect 33572 18284 33582 18340
rect 37762 18284 37772 18340
rect 37828 18284 39004 18340
rect 39060 18284 39070 18340
rect 52994 18284 53004 18340
rect 53060 18284 53676 18340
rect 53732 18284 56700 18340
rect 56756 18284 56766 18340
rect 76962 18284 76972 18340
rect 77028 18284 77308 18340
rect 77364 18284 77374 18340
rect 18050 18172 18060 18228
rect 18116 18172 21980 18228
rect 22036 18172 22046 18228
rect 22306 18172 22316 18228
rect 22372 18172 25676 18228
rect 25732 18172 35588 18228
rect 37426 18172 37436 18228
rect 37492 18172 40236 18228
rect 40292 18172 40302 18228
rect 26562 18060 26572 18116
rect 26628 18060 30716 18116
rect 30772 18060 30782 18116
rect 31154 18060 31164 18116
rect 31220 18060 33628 18116
rect 33684 18060 33694 18116
rect 0 18004 800 18032
rect 4466 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4750 18060
rect 35186 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35470 18060
rect 35532 18004 35588 18172
rect 39666 18060 39676 18116
rect 39732 18060 43372 18116
rect 43428 18060 43438 18116
rect 51426 18060 51436 18116
rect 51492 18060 53676 18116
rect 53732 18060 53742 18116
rect 65906 18004 65916 18060
rect 65972 18004 66020 18060
rect 66076 18004 66124 18060
rect 66180 18004 66190 18060
rect 0 17948 1708 18004
rect 1764 17948 2492 18004
rect 2548 17948 2558 18004
rect 9986 17948 9996 18004
rect 10052 17948 33740 18004
rect 33796 17948 33806 18004
rect 35532 17948 41580 18004
rect 41636 17948 43148 18004
rect 43204 17948 43214 18004
rect 47394 17948 47404 18004
rect 47460 17948 50988 18004
rect 51044 17948 52444 18004
rect 52500 17948 52510 18004
rect 0 17920 800 17948
rect 2034 17836 2044 17892
rect 2100 17836 26908 17892
rect 28466 17836 28476 17892
rect 28532 17836 33180 17892
rect 33236 17836 33246 17892
rect 45042 17836 45052 17892
rect 45108 17836 72268 17892
rect 72324 17836 72334 17892
rect 26852 17668 26908 17836
rect 28130 17724 28140 17780
rect 28196 17724 28588 17780
rect 28644 17724 33404 17780
rect 33460 17724 34412 17780
rect 34468 17724 34478 17780
rect 34738 17724 34748 17780
rect 34804 17724 35084 17780
rect 35140 17724 35150 17780
rect 37090 17724 37100 17780
rect 37156 17724 38780 17780
rect 38836 17724 38846 17780
rect 42018 17724 42028 17780
rect 42084 17724 44156 17780
rect 44212 17724 44940 17780
rect 44996 17724 45006 17780
rect 45266 17724 45276 17780
rect 45332 17724 46732 17780
rect 46788 17724 46798 17780
rect 49970 17724 49980 17780
rect 50036 17724 51324 17780
rect 51380 17724 52108 17780
rect 52164 17724 52174 17780
rect 56252 17724 70588 17780
rect 70644 17724 70654 17780
rect 56252 17668 56308 17724
rect 19394 17612 19404 17668
rect 19460 17612 20188 17668
rect 20244 17612 20254 17668
rect 26852 17612 37884 17668
rect 37940 17612 37950 17668
rect 38994 17612 39004 17668
rect 39060 17612 39788 17668
rect 39844 17612 39854 17668
rect 43586 17612 43596 17668
rect 43652 17612 45388 17668
rect 45444 17612 45454 17668
rect 45612 17612 56308 17668
rect 57138 17612 57148 17668
rect 57204 17612 58716 17668
rect 58772 17612 58782 17668
rect 45612 17556 45668 17612
rect 79200 17556 80000 17584
rect 18722 17500 18732 17556
rect 18788 17500 19292 17556
rect 19348 17500 20860 17556
rect 20916 17500 20926 17556
rect 21858 17500 21868 17556
rect 21924 17500 25116 17556
rect 25172 17500 25182 17556
rect 30370 17500 30380 17556
rect 30436 17500 31276 17556
rect 31332 17500 31342 17556
rect 34290 17500 34300 17556
rect 34356 17500 36988 17556
rect 37044 17500 37054 17556
rect 38770 17500 38780 17556
rect 38836 17500 39676 17556
rect 39732 17500 40908 17556
rect 40964 17500 40974 17556
rect 44930 17500 44940 17556
rect 44996 17500 45668 17556
rect 46162 17500 46172 17556
rect 46228 17500 47516 17556
rect 47572 17500 47582 17556
rect 50530 17500 50540 17556
rect 50596 17500 50988 17556
rect 51044 17500 51054 17556
rect 77634 17500 77644 17556
rect 77700 17500 78204 17556
rect 78260 17500 80000 17556
rect 79200 17472 80000 17500
rect 1698 17388 1708 17444
rect 1764 17388 2492 17444
rect 2548 17388 2558 17444
rect 36082 17388 36092 17444
rect 36148 17388 37324 17444
rect 37380 17388 37390 17444
rect 38546 17388 38556 17444
rect 38612 17388 41356 17444
rect 41412 17388 41422 17444
rect 43026 17388 43036 17444
rect 43092 17388 48524 17444
rect 48580 17388 48590 17444
rect 50754 17388 50764 17444
rect 50820 17388 52668 17444
rect 52724 17388 52734 17444
rect 58370 17388 58380 17444
rect 58436 17388 68796 17444
rect 68852 17388 68862 17444
rect 29250 17276 29260 17332
rect 29316 17276 32284 17332
rect 32340 17276 38668 17332
rect 19826 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20110 17276
rect 38612 17220 38668 17276
rect 39116 17276 49980 17332
rect 50036 17276 50046 17332
rect 53116 17276 53340 17332
rect 53396 17276 54796 17332
rect 54852 17276 58828 17332
rect 58884 17276 58894 17332
rect 39116 17220 39172 17276
rect 50546 17220 50556 17276
rect 50612 17220 50660 17276
rect 50716 17220 50764 17276
rect 50820 17220 50830 17276
rect 53116 17220 53172 17276
rect 35970 17164 35980 17220
rect 36036 17164 36316 17220
rect 36372 17164 36382 17220
rect 36978 17164 36988 17220
rect 37044 17164 37548 17220
rect 37604 17164 37614 17220
rect 38612 17164 39172 17220
rect 39554 17164 39564 17220
rect 39620 17164 39900 17220
rect 39956 17164 39966 17220
rect 40338 17164 40348 17220
rect 40404 17164 49588 17220
rect 53106 17164 53116 17220
rect 53172 17164 53182 17220
rect 49532 17108 49588 17164
rect 2034 17052 2044 17108
rect 2100 17052 26908 17108
rect 29698 17052 29708 17108
rect 29764 17052 32732 17108
rect 32788 17052 35420 17108
rect 35476 17052 38332 17108
rect 38388 17052 38398 17108
rect 43026 17052 43036 17108
rect 43092 17052 45332 17108
rect 49532 17052 63756 17108
rect 63812 17052 63822 17108
rect 26852 16996 26908 17052
rect 45276 16996 45332 17052
rect 26852 16940 36036 16996
rect 36194 16940 36204 16996
rect 36260 16940 36988 16996
rect 37044 16940 37054 16996
rect 37986 16940 37996 16996
rect 38052 16940 38780 16996
rect 38836 16940 38846 16996
rect 41458 16940 41468 16996
rect 41524 16940 45052 16996
rect 45108 16940 45118 16996
rect 45266 16940 45276 16996
rect 45332 16940 45342 16996
rect 46386 16940 46396 16996
rect 46452 16940 50428 16996
rect 50978 16940 50988 16996
rect 51044 16940 52108 16996
rect 52164 16940 52174 16996
rect 57922 16940 57932 16996
rect 57988 16940 57998 16996
rect 0 16884 800 16912
rect 35980 16884 36036 16940
rect 50372 16884 50428 16940
rect 57932 16884 57988 16940
rect 0 16828 1708 16884
rect 1764 16828 1774 16884
rect 28130 16828 28140 16884
rect 28196 16828 29484 16884
rect 29540 16828 29550 16884
rect 35980 16828 36540 16884
rect 36596 16828 37604 16884
rect 38546 16828 38556 16884
rect 38612 16828 39228 16884
rect 39284 16828 39294 16884
rect 39554 16828 39564 16884
rect 39620 16828 41916 16884
rect 41972 16828 41982 16884
rect 42242 16828 42252 16884
rect 42308 16828 42476 16884
rect 42532 16828 43036 16884
rect 43092 16828 43102 16884
rect 47254 16828 47292 16884
rect 47348 16828 47358 16884
rect 50372 16828 57988 16884
rect 77634 16828 77644 16884
rect 77700 16828 78204 16884
rect 78260 16828 78270 16884
rect 0 16800 800 16828
rect 37548 16772 37604 16828
rect 37538 16716 37548 16772
rect 37604 16716 37614 16772
rect 42914 16716 42924 16772
rect 42980 16716 43932 16772
rect 43988 16716 43998 16772
rect 38322 16604 38332 16660
rect 38388 16604 39228 16660
rect 39284 16604 39294 16660
rect 50372 16604 70252 16660
rect 70308 16604 70318 16660
rect 50372 16548 50428 16604
rect 28242 16492 28252 16548
rect 28308 16492 29260 16548
rect 29316 16492 29326 16548
rect 43922 16492 43932 16548
rect 43988 16492 44268 16548
rect 44324 16492 50428 16548
rect 4466 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4750 16492
rect 35186 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35470 16492
rect 65906 16436 65916 16492
rect 65972 16436 66020 16492
rect 66076 16436 66124 16492
rect 66180 16436 66190 16492
rect 79200 16436 80000 16464
rect 25554 16380 25564 16436
rect 25620 16380 26572 16436
rect 26628 16380 27804 16436
rect 27860 16380 31332 16436
rect 31276 16324 31332 16380
rect 35532 16380 51436 16436
rect 51492 16380 51502 16436
rect 78194 16380 78204 16436
rect 78260 16380 80000 16436
rect 35532 16324 35588 16380
rect 79200 16352 80000 16380
rect 2034 16268 2044 16324
rect 2100 16268 26908 16324
rect 31276 16268 35588 16324
rect 36754 16268 36764 16324
rect 36820 16268 37996 16324
rect 38052 16268 38062 16324
rect 43474 16268 43484 16324
rect 43540 16268 45836 16324
rect 45892 16268 68908 16324
rect 68964 16268 68974 16324
rect 26852 16212 26908 16268
rect 26852 16156 37324 16212
rect 37380 16156 37390 16212
rect 38612 16156 38780 16212
rect 38836 16156 38846 16212
rect 42578 16156 42588 16212
rect 42644 16156 45500 16212
rect 45556 16156 45566 16212
rect 1922 16044 1932 16100
rect 1988 16044 28476 16100
rect 28532 16044 28542 16100
rect 31826 16044 31836 16100
rect 31892 16044 32508 16100
rect 32564 16044 32574 16100
rect 38612 15988 38668 16156
rect 42130 16044 42140 16100
rect 42196 16044 46172 16100
rect 46228 16044 46238 16100
rect 5954 15932 5964 15988
rect 6020 15932 27132 15988
rect 27188 15932 27198 15988
rect 28578 15932 28588 15988
rect 28644 15932 38220 15988
rect 38276 15932 38668 15988
rect 39442 15932 39452 15988
rect 39508 15932 48748 15988
rect 48804 15932 48814 15988
rect 75394 15932 75404 15988
rect 75460 15932 77868 15988
rect 77924 15932 77934 15988
rect 25666 15820 25676 15876
rect 25732 15820 27356 15876
rect 27412 15820 27422 15876
rect 40226 15820 40236 15876
rect 40292 15820 42812 15876
rect 42868 15820 42878 15876
rect 44034 15820 44044 15876
rect 44100 15820 44828 15876
rect 44884 15820 44894 15876
rect 47180 15820 50428 15876
rect 50484 15820 51324 15876
rect 51380 15820 51390 15876
rect 77634 15820 77644 15876
rect 77700 15820 78204 15876
rect 78260 15820 78270 15876
rect 0 15764 800 15792
rect 47180 15764 47236 15820
rect 0 15708 1708 15764
rect 1764 15708 2492 15764
rect 2548 15708 2558 15764
rect 26786 15708 26796 15764
rect 0 15680 800 15708
rect 19826 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20110 15708
rect 26852 15652 26908 15764
rect 45490 15708 45500 15764
rect 45556 15708 45836 15764
rect 45892 15708 45902 15764
rect 47170 15708 47180 15764
rect 47236 15708 47246 15764
rect 50546 15652 50556 15708
rect 50612 15652 50660 15708
rect 50716 15652 50764 15708
rect 50820 15652 50830 15708
rect 26852 15596 27692 15652
rect 27748 15596 28028 15652
rect 28084 15596 29708 15652
rect 29764 15596 29774 15652
rect 33394 15596 33404 15652
rect 33460 15596 35980 15652
rect 36036 15596 48972 15652
rect 49028 15596 49038 15652
rect 26002 15484 26012 15540
rect 26068 15484 27468 15540
rect 27524 15484 28140 15540
rect 28196 15484 43708 15540
rect 46498 15484 46508 15540
rect 46564 15484 47180 15540
rect 47236 15484 47246 15540
rect 47954 15484 47964 15540
rect 48020 15484 49028 15540
rect 43652 15428 43708 15484
rect 48972 15428 49028 15484
rect 2034 15372 2044 15428
rect 2100 15372 38444 15428
rect 38500 15372 38510 15428
rect 43652 15372 47404 15428
rect 47460 15372 47470 15428
rect 47730 15372 47740 15428
rect 47796 15372 48748 15428
rect 48804 15372 48814 15428
rect 48962 15372 48972 15428
rect 49028 15372 49420 15428
rect 49476 15372 50652 15428
rect 50708 15372 50718 15428
rect 51202 15372 51212 15428
rect 51268 15372 52556 15428
rect 52612 15372 52622 15428
rect 79200 15316 80000 15344
rect 27794 15260 27804 15316
rect 27860 15260 28476 15316
rect 28532 15260 28542 15316
rect 35746 15260 35756 15316
rect 35812 15260 39228 15316
rect 39284 15260 39294 15316
rect 39890 15260 39900 15316
rect 39956 15260 41804 15316
rect 41860 15260 41870 15316
rect 45490 15260 45500 15316
rect 45556 15260 54684 15316
rect 54740 15260 54750 15316
rect 78194 15260 78204 15316
rect 78260 15260 80000 15316
rect 79200 15232 80000 15260
rect 37986 15148 37996 15204
rect 38052 15148 38892 15204
rect 38948 15148 38958 15204
rect 44258 15148 44268 15204
rect 44324 15148 44828 15204
rect 44884 15148 44894 15204
rect 47730 15148 47740 15204
rect 47796 15148 48300 15204
rect 48356 15148 48366 15204
rect 51650 15148 51660 15204
rect 51716 15148 57932 15204
rect 57988 15148 57998 15204
rect 77046 15148 77084 15204
rect 77140 15148 77150 15204
rect 38994 15036 39004 15092
rect 39060 15036 49084 15092
rect 49140 15036 49150 15092
rect 68786 15036 68796 15092
rect 68852 15036 74396 15092
rect 74452 15036 74462 15092
rect 45378 14924 45388 14980
rect 45444 14924 54460 14980
rect 54516 14924 54526 14980
rect 4466 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4750 14924
rect 35186 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35470 14924
rect 65906 14868 65916 14924
rect 65972 14868 66020 14924
rect 66076 14868 66124 14924
rect 66180 14868 66190 14924
rect 21858 14812 21868 14868
rect 21924 14812 24892 14868
rect 24948 14812 24958 14868
rect 28812 14812 33852 14868
rect 33908 14812 33918 14868
rect 41570 14812 41580 14868
rect 41636 14812 57148 14868
rect 57204 14812 57214 14868
rect 2146 14700 2156 14756
rect 2212 14700 28588 14756
rect 28644 14700 28654 14756
rect 0 14644 800 14672
rect 28812 14644 28868 14812
rect 37986 14700 37996 14756
rect 38052 14700 39116 14756
rect 39172 14700 39182 14756
rect 52098 14700 52108 14756
rect 52164 14700 52892 14756
rect 52948 14700 54572 14756
rect 54628 14700 54638 14756
rect 0 14588 1708 14644
rect 1764 14588 2492 14644
rect 2548 14588 2558 14644
rect 10098 14588 10108 14644
rect 10164 14588 28868 14644
rect 29260 14588 32284 14644
rect 32340 14588 32350 14644
rect 41234 14588 41244 14644
rect 41300 14588 43372 14644
rect 43428 14588 54796 14644
rect 54852 14588 54862 14644
rect 0 14560 800 14588
rect 29260 14532 29316 14588
rect 6962 14476 6972 14532
rect 7028 14476 29316 14532
rect 29474 14476 29484 14532
rect 29540 14476 30828 14532
rect 30884 14476 30894 14532
rect 42690 14476 42700 14532
rect 42756 14476 45500 14532
rect 45556 14476 45566 14532
rect 51314 14476 51324 14532
rect 51380 14476 52668 14532
rect 52724 14476 52734 14532
rect 32498 14364 32508 14420
rect 32564 14364 33404 14420
rect 33460 14364 33470 14420
rect 42354 14364 42364 14420
rect 42420 14364 43260 14420
rect 43316 14364 43326 14420
rect 50418 14364 50428 14420
rect 50484 14364 68460 14420
rect 68516 14364 68526 14420
rect 76850 14364 76860 14420
rect 76916 14364 77868 14420
rect 77924 14364 77934 14420
rect 18946 14252 18956 14308
rect 19012 14252 19740 14308
rect 19796 14252 19806 14308
rect 20066 14252 20076 14308
rect 20132 14252 21420 14308
rect 21476 14252 22876 14308
rect 22932 14252 22942 14308
rect 30930 14252 30940 14308
rect 30996 14252 35532 14308
rect 35588 14252 35598 14308
rect 36754 14252 36764 14308
rect 36820 14252 36830 14308
rect 38546 14252 38556 14308
rect 38612 14252 42476 14308
rect 42532 14252 42542 14308
rect 50372 14252 50876 14308
rect 50932 14252 50942 14308
rect 36764 14196 36820 14252
rect 26852 14140 36820 14196
rect 39106 14140 39116 14196
rect 39172 14140 40124 14196
rect 40180 14140 41468 14196
rect 41524 14140 42924 14196
rect 42980 14140 43260 14196
rect 43316 14140 43326 14196
rect 19826 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20110 14140
rect 26852 13972 26908 14140
rect 50372 14084 50428 14252
rect 79200 14196 80000 14224
rect 77634 14140 77644 14196
rect 77700 14140 78204 14196
rect 78260 14140 80000 14196
rect 50546 14084 50556 14140
rect 50612 14084 50660 14140
rect 50716 14084 50764 14140
rect 50820 14084 50830 14140
rect 79200 14112 80000 14140
rect 33394 14028 33404 14084
rect 33460 14028 34076 14084
rect 34132 14028 34972 14084
rect 35028 14028 48860 14084
rect 48916 14028 50428 14084
rect 2034 13916 2044 13972
rect 2100 13916 26908 13972
rect 29698 13916 29708 13972
rect 29764 13916 30268 13972
rect 30324 13916 30334 13972
rect 33618 13916 33628 13972
rect 33684 13916 35308 13972
rect 35364 13916 35980 13972
rect 36036 13916 36046 13972
rect 37436 13916 38444 13972
rect 38500 13916 38668 13972
rect 53890 13916 53900 13972
rect 53956 13916 55132 13972
rect 55188 13916 55198 13972
rect 76738 13916 76748 13972
rect 76804 13916 77868 13972
rect 77924 13916 77934 13972
rect 30268 13860 30324 13916
rect 37436 13860 37492 13916
rect 38612 13860 38668 13916
rect 18610 13804 18620 13860
rect 18676 13804 19180 13860
rect 19236 13804 19246 13860
rect 23538 13804 23548 13860
rect 23604 13804 25900 13860
rect 25956 13804 25966 13860
rect 26852 13804 27020 13860
rect 27076 13804 27086 13860
rect 28466 13804 28476 13860
rect 28532 13804 29036 13860
rect 29092 13804 29932 13860
rect 29988 13804 29998 13860
rect 30268 13804 37492 13860
rect 37650 13804 37660 13860
rect 37716 13804 38220 13860
rect 38276 13804 38286 13860
rect 38612 13804 38780 13860
rect 38836 13804 38846 13860
rect 53218 13804 53228 13860
rect 53284 13804 54236 13860
rect 54292 13804 54302 13860
rect 19506 13692 19516 13748
rect 19572 13692 20300 13748
rect 20356 13692 20366 13748
rect 22530 13692 22540 13748
rect 22596 13692 24892 13748
rect 24948 13692 24958 13748
rect 26852 13636 26908 13804
rect 28476 13748 28532 13804
rect 35532 13748 35588 13804
rect 27122 13692 27132 13748
rect 27188 13692 28532 13748
rect 31266 13692 31276 13748
rect 31332 13692 31612 13748
rect 31668 13692 31678 13748
rect 31938 13692 31948 13748
rect 32004 13692 32956 13748
rect 33012 13692 33022 13748
rect 35532 13692 35644 13748
rect 35700 13692 35710 13748
rect 37986 13692 37996 13748
rect 38052 13692 40796 13748
rect 40852 13692 40862 13748
rect 41794 13692 41804 13748
rect 41860 13692 52220 13748
rect 52276 13692 52286 13748
rect 31612 13636 31668 13692
rect 18050 13580 18060 13636
rect 18116 13580 19068 13636
rect 19124 13580 19134 13636
rect 24658 13580 24668 13636
rect 24724 13580 26908 13636
rect 27682 13580 27692 13636
rect 27748 13580 31164 13636
rect 31220 13580 31230 13636
rect 31612 13580 32172 13636
rect 32228 13580 32238 13636
rect 32610 13580 32620 13636
rect 32676 13580 38332 13636
rect 38388 13580 38398 13636
rect 40226 13580 40236 13636
rect 40292 13580 41356 13636
rect 41412 13580 41422 13636
rect 43810 13580 43820 13636
rect 43876 13580 46620 13636
rect 46676 13580 46686 13636
rect 77634 13580 77644 13636
rect 77700 13580 78204 13636
rect 78260 13580 78270 13636
rect 0 13524 800 13552
rect 0 13468 1708 13524
rect 1764 13468 2492 13524
rect 2548 13468 2558 13524
rect 25442 13468 25452 13524
rect 25508 13468 28588 13524
rect 28644 13468 28654 13524
rect 32498 13468 32508 13524
rect 32564 13468 32844 13524
rect 32900 13468 32910 13524
rect 38210 13468 38220 13524
rect 38276 13468 39676 13524
rect 39732 13468 39742 13524
rect 43036 13468 45388 13524
rect 45444 13468 45454 13524
rect 0 13440 800 13468
rect 39676 13412 39732 13468
rect 43036 13412 43092 13468
rect 39676 13356 40908 13412
rect 40964 13356 40974 13412
rect 43026 13356 43036 13412
rect 43092 13356 43102 13412
rect 4466 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4750 13356
rect 35186 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35470 13356
rect 65906 13300 65916 13356
rect 65972 13300 66020 13356
rect 66076 13300 66124 13356
rect 66180 13300 66190 13356
rect 36978 13244 36988 13300
rect 37044 13244 37772 13300
rect 37828 13244 37838 13300
rect 33282 13132 33292 13188
rect 33348 13132 54236 13188
rect 54292 13132 54302 13188
rect 79200 13076 80000 13104
rect 6626 13020 6636 13076
rect 6692 13020 34300 13076
rect 34356 13020 34366 13076
rect 36418 13020 36428 13076
rect 36484 13020 37772 13076
rect 37828 13020 37838 13076
rect 74946 13020 74956 13076
rect 75012 13020 75628 13076
rect 75684 13020 75740 13076
rect 75796 13020 76300 13076
rect 76356 13020 76366 13076
rect 78194 13020 78204 13076
rect 78260 13020 80000 13076
rect 79200 12992 80000 13020
rect 39106 12908 39116 12964
rect 39172 12908 39564 12964
rect 39620 12908 41916 12964
rect 41972 12908 41982 12964
rect 43474 12908 43484 12964
rect 43540 12908 60284 12964
rect 60340 12908 60350 12964
rect 25778 12796 25788 12852
rect 25844 12796 28364 12852
rect 28420 12796 29484 12852
rect 29540 12796 29550 12852
rect 37874 12796 37884 12852
rect 37940 12796 48748 12852
rect 48804 12796 48814 12852
rect 31490 12684 31500 12740
rect 31556 12684 73052 12740
rect 73108 12684 73118 12740
rect 75282 12684 75292 12740
rect 75348 12684 77756 12740
rect 77812 12684 77822 12740
rect 28578 12572 28588 12628
rect 28644 12572 29372 12628
rect 29428 12572 31612 12628
rect 31668 12572 37100 12628
rect 37156 12572 37166 12628
rect 19826 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20110 12572
rect 50546 12516 50556 12572
rect 50612 12516 50660 12572
rect 50716 12516 50764 12572
rect 50820 12516 50830 12572
rect 0 12404 800 12432
rect 0 12348 1708 12404
rect 1764 12348 2492 12404
rect 2548 12348 2558 12404
rect 3332 12348 26908 12404
rect 32498 12348 32508 12404
rect 32564 12348 34636 12404
rect 34692 12348 34702 12404
rect 35074 12348 35084 12404
rect 35140 12348 37884 12404
rect 37940 12348 37950 12404
rect 41234 12348 41244 12404
rect 41300 12348 42588 12404
rect 42644 12348 42654 12404
rect 0 12320 800 12348
rect 3332 12292 3388 12348
rect 2146 12236 2156 12292
rect 2212 12236 3388 12292
rect 26852 12292 26908 12348
rect 26852 12236 35644 12292
rect 35700 12236 36204 12292
rect 36260 12236 36270 12292
rect 37538 12124 37548 12180
rect 37604 12124 39564 12180
rect 39620 12124 39630 12180
rect 9874 12012 9884 12068
rect 9940 12012 11788 12068
rect 11844 12012 11854 12068
rect 23426 12012 23436 12068
rect 23492 12012 25340 12068
rect 25396 12012 25406 12068
rect 31948 12012 32508 12068
rect 32564 12012 32574 12068
rect 31948 11956 32004 12012
rect 79200 11956 80000 11984
rect 31938 11900 31948 11956
rect 32004 11900 32014 11956
rect 32508 11900 36988 11956
rect 37044 11900 37054 11956
rect 78194 11900 78204 11956
rect 78260 11900 80000 11956
rect 32508 11844 32564 11900
rect 79200 11872 80000 11900
rect 12674 11788 12684 11844
rect 12740 11788 15372 11844
rect 15428 11788 16604 11844
rect 16660 11788 16670 11844
rect 32498 11788 32508 11844
rect 32564 11788 32574 11844
rect 4466 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4750 11788
rect 35186 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35470 11788
rect 65906 11732 65916 11788
rect 65972 11732 66020 11788
rect 66076 11732 66124 11788
rect 66180 11732 66190 11788
rect 26852 11676 28588 11732
rect 28644 11676 29932 11732
rect 29988 11676 29998 11732
rect 40226 11676 40236 11732
rect 40292 11676 56028 11732
rect 56084 11676 56094 11732
rect 26852 11620 26908 11676
rect 26226 11564 26236 11620
rect 26292 11564 26908 11620
rect 36418 11564 36428 11620
rect 36484 11564 41020 11620
rect 41076 11564 41086 11620
rect 50372 11564 52556 11620
rect 52612 11564 52622 11620
rect 50372 11508 50428 11564
rect 13682 11452 13692 11508
rect 13748 11452 14476 11508
rect 14532 11452 15596 11508
rect 15652 11452 15662 11508
rect 19954 11452 19964 11508
rect 20020 11452 20748 11508
rect 20804 11452 21756 11508
rect 21812 11452 21822 11508
rect 33730 11452 33740 11508
rect 33796 11452 50428 11508
rect 76514 11452 76524 11508
rect 76580 11452 78204 11508
rect 78260 11452 78270 11508
rect 32946 11340 32956 11396
rect 33012 11340 36428 11396
rect 36484 11340 36494 11396
rect 38098 11340 38108 11396
rect 38164 11340 40068 11396
rect 44482 11340 44492 11396
rect 44548 11340 55356 11396
rect 55412 11340 55422 11396
rect 0 11284 800 11312
rect 0 11228 1708 11284
rect 1764 11228 2492 11284
rect 2548 11228 2558 11284
rect 22642 11228 22652 11284
rect 22708 11228 24892 11284
rect 24948 11228 24958 11284
rect 30370 11228 30380 11284
rect 30436 11228 31836 11284
rect 31892 11228 31902 11284
rect 38210 11228 38220 11284
rect 38276 11228 39452 11284
rect 39508 11228 39518 11284
rect 0 11200 800 11228
rect 40012 11172 40068 11340
rect 41346 11228 41356 11284
rect 41412 11228 42140 11284
rect 42196 11228 42206 11284
rect 47012 11228 56028 11284
rect 56084 11228 56094 11284
rect 47012 11172 47068 11228
rect 2034 11116 2044 11172
rect 2100 11116 2110 11172
rect 11554 11116 11564 11172
rect 11620 11116 12012 11172
rect 12068 11116 12460 11172
rect 12516 11116 12526 11172
rect 13010 11116 13020 11172
rect 13076 11116 13468 11172
rect 13524 11116 13534 11172
rect 18946 11116 18956 11172
rect 19012 11116 19740 11172
rect 19796 11116 19806 11172
rect 27122 11116 27132 11172
rect 27188 11116 30156 11172
rect 30212 11116 30222 11172
rect 33282 11116 33292 11172
rect 33348 11116 39676 11172
rect 39732 11116 39742 11172
rect 40012 11116 47068 11172
rect 50372 11116 56140 11172
rect 56196 11116 56206 11172
rect 2044 10836 2100 11116
rect 50372 11060 50428 11116
rect 31042 11004 31052 11060
rect 31108 11004 42588 11060
rect 42644 11004 42654 11060
rect 45042 11004 45052 11060
rect 45108 11004 45612 11060
rect 45668 11004 50428 11060
rect 19826 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20110 11004
rect 50546 10948 50556 11004
rect 50612 10948 50660 11004
rect 50716 10948 50764 11004
rect 50820 10948 50830 11004
rect 2370 10892 2380 10948
rect 2436 10892 9996 10948
rect 10052 10892 10062 10948
rect 17798 10892 17836 10948
rect 17892 10892 17902 10948
rect 25218 10892 25228 10948
rect 25284 10892 26684 10948
rect 26740 10892 26750 10948
rect 26852 10892 37212 10948
rect 37268 10892 37660 10948
rect 37716 10892 37726 10948
rect 52994 10892 53004 10948
rect 53060 10892 69356 10948
rect 69412 10892 69422 10948
rect 26852 10836 26908 10892
rect 79200 10836 80000 10864
rect 2044 10780 26908 10836
rect 27906 10780 27916 10836
rect 27972 10780 32508 10836
rect 32564 10780 36988 10836
rect 37044 10780 38332 10836
rect 38388 10780 38398 10836
rect 39330 10780 39340 10836
rect 39396 10780 40236 10836
rect 40292 10780 40302 10836
rect 76962 10780 76972 10836
rect 77028 10780 77532 10836
rect 77588 10780 80000 10836
rect 79200 10752 80000 10780
rect 33506 10668 33516 10724
rect 33572 10668 44492 10724
rect 44548 10668 44558 10724
rect 17714 10556 17724 10612
rect 17780 10556 18284 10612
rect 18340 10556 18350 10612
rect 28466 10556 28476 10612
rect 28532 10556 29708 10612
rect 29764 10556 29774 10612
rect 37426 10556 37436 10612
rect 37492 10556 38892 10612
rect 38948 10556 38958 10612
rect 9426 10444 9436 10500
rect 9492 10444 10332 10500
rect 10388 10444 10398 10500
rect 13794 10444 13804 10500
rect 13860 10444 14476 10500
rect 14532 10444 14542 10500
rect 22978 10444 22988 10500
rect 23044 10444 25340 10500
rect 25396 10444 25406 10500
rect 31266 10444 31276 10500
rect 31332 10444 33292 10500
rect 33348 10444 33358 10500
rect 42130 10444 42140 10500
rect 42196 10444 43372 10500
rect 43428 10444 43438 10500
rect 26226 10332 26236 10388
rect 26292 10332 32060 10388
rect 32116 10332 32126 10388
rect 25778 10220 25788 10276
rect 25844 10220 31612 10276
rect 31668 10220 31678 10276
rect 0 10164 800 10192
rect 4466 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4750 10220
rect 35186 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35470 10220
rect 65906 10164 65916 10220
rect 65972 10164 66020 10220
rect 66076 10164 66124 10220
rect 66180 10164 66190 10220
rect 0 10108 1708 10164
rect 1764 10108 2492 10164
rect 2548 10108 2558 10164
rect 11778 10108 11788 10164
rect 11844 10108 13020 10164
rect 13076 10108 13086 10164
rect 13346 10108 13356 10164
rect 13412 10108 14028 10164
rect 14084 10108 28028 10164
rect 28084 10108 28094 10164
rect 31714 10108 31724 10164
rect 31780 10108 32172 10164
rect 32228 10108 32956 10164
rect 33012 10108 33180 10164
rect 33236 10108 33246 10164
rect 43362 10108 43372 10164
rect 43428 10108 45612 10164
rect 45668 10108 45678 10164
rect 53330 10108 53340 10164
rect 53396 10108 57148 10164
rect 57204 10108 57214 10164
rect 0 10080 800 10108
rect 2034 9996 2044 10052
rect 2100 9996 10108 10052
rect 10164 9996 10174 10052
rect 33058 9996 33068 10052
rect 33124 9996 33964 10052
rect 34020 9996 34030 10052
rect 35746 9996 35756 10052
rect 35812 9996 44436 10052
rect 75506 9996 75516 10052
rect 75572 9996 77420 10052
rect 77476 9996 77486 10052
rect 13794 9884 13804 9940
rect 13860 9884 14140 9940
rect 14196 9884 24668 9940
rect 24724 9884 24734 9940
rect 26852 9884 27804 9940
rect 27860 9884 27870 9940
rect 38770 9884 38780 9940
rect 38836 9884 43596 9940
rect 43652 9884 43662 9940
rect 26852 9828 26908 9884
rect 12338 9772 12348 9828
rect 12404 9772 13468 9828
rect 13524 9772 13916 9828
rect 13972 9772 13982 9828
rect 20290 9772 20300 9828
rect 20356 9772 20860 9828
rect 20916 9772 22764 9828
rect 22820 9772 26908 9828
rect 32610 9772 32620 9828
rect 32676 9772 33516 9828
rect 33572 9772 33582 9828
rect 36194 9772 36204 9828
rect 36260 9772 37324 9828
rect 37380 9772 39788 9828
rect 39844 9772 39854 9828
rect 9538 9660 9548 9716
rect 9604 9660 11900 9716
rect 11956 9660 11966 9716
rect 14690 9660 14700 9716
rect 14756 9660 18508 9716
rect 18564 9660 18574 9716
rect 29474 9660 29484 9716
rect 29540 9660 33180 9716
rect 33236 9660 33246 9716
rect 36530 9660 36540 9716
rect 36596 9660 39956 9716
rect 42130 9660 42140 9716
rect 42196 9660 44044 9716
rect 44100 9660 44110 9716
rect 39900 9604 39956 9660
rect 44380 9604 44436 9996
rect 45714 9884 45724 9940
rect 45780 9884 56588 9940
rect 56644 9884 56654 9940
rect 46946 9772 46956 9828
rect 47012 9772 59612 9828
rect 59668 9772 59678 9828
rect 79200 9716 80000 9744
rect 48402 9660 48412 9716
rect 48468 9660 63868 9716
rect 63924 9660 63934 9716
rect 77634 9660 77644 9716
rect 77700 9660 78204 9716
rect 78260 9660 80000 9716
rect 79200 9632 80000 9660
rect 1698 9548 1708 9604
rect 1764 9548 2492 9604
rect 2548 9548 2558 9604
rect 8306 9548 8316 9604
rect 8372 9548 9324 9604
rect 9380 9548 9390 9604
rect 11106 9548 11116 9604
rect 11172 9548 14476 9604
rect 14532 9548 14542 9604
rect 23426 9548 23436 9604
rect 23492 9548 29260 9604
rect 29316 9548 29326 9604
rect 32498 9548 32508 9604
rect 32564 9548 34860 9604
rect 34916 9548 34926 9604
rect 39666 9548 39676 9604
rect 39732 9548 39742 9604
rect 39900 9548 42924 9604
rect 42980 9548 42990 9604
rect 44370 9548 44380 9604
rect 44436 9548 44446 9604
rect 45826 9548 45836 9604
rect 45892 9548 53172 9604
rect 77858 9548 77868 9604
rect 77924 9548 78652 9604
rect 78708 9548 78718 9604
rect 27794 9436 27804 9492
rect 27860 9436 34188 9492
rect 34244 9436 34254 9492
rect 19826 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20110 9436
rect 39676 9380 39732 9548
rect 50546 9380 50556 9436
rect 50612 9380 50660 9436
rect 50716 9380 50764 9436
rect 50820 9380 50830 9436
rect 16706 9324 16716 9380
rect 16772 9324 18620 9380
rect 18676 9324 18686 9380
rect 29698 9324 29708 9380
rect 29764 9324 30492 9380
rect 30548 9324 30558 9380
rect 33282 9324 33292 9380
rect 33348 9324 39732 9380
rect 53116 9268 53172 9548
rect 55010 9324 55020 9380
rect 55076 9324 69020 9380
rect 69076 9324 69086 9380
rect 76402 9324 76412 9380
rect 76468 9324 77868 9380
rect 77924 9324 77934 9380
rect 16146 9212 16156 9268
rect 16212 9212 17612 9268
rect 17668 9212 17678 9268
rect 18386 9212 18396 9268
rect 18452 9212 18844 9268
rect 18900 9212 18910 9268
rect 22306 9212 22316 9268
rect 22372 9212 23548 9268
rect 23604 9212 23614 9268
rect 24658 9212 24668 9268
rect 24724 9212 25228 9268
rect 25284 9212 31164 9268
rect 31220 9212 31836 9268
rect 31892 9212 32956 9268
rect 33012 9212 33022 9268
rect 33180 9212 38668 9268
rect 38724 9212 38734 9268
rect 38882 9212 38892 9268
rect 38948 9212 41132 9268
rect 41188 9212 41198 9268
rect 43586 9212 43596 9268
rect 43652 9212 43932 9268
rect 43988 9212 43998 9268
rect 44146 9212 44156 9268
rect 44212 9212 45276 9268
rect 45332 9212 46060 9268
rect 46116 9212 52892 9268
rect 52948 9212 52958 9268
rect 53116 9212 66556 9268
rect 66612 9212 66622 9268
rect 33180 9156 33236 9212
rect 28578 9100 28588 9156
rect 28644 9100 33236 9156
rect 38210 9100 38220 9156
rect 38276 9100 38780 9156
rect 38836 9100 38846 9156
rect 41010 9100 41020 9156
rect 41076 9100 41356 9156
rect 41412 9100 44940 9156
rect 44996 9100 45006 9156
rect 0 9044 800 9072
rect 0 8988 1708 9044
rect 1764 8988 1774 9044
rect 15586 8988 15596 9044
rect 15652 8988 17388 9044
rect 17444 8988 17454 9044
rect 18722 8988 18732 9044
rect 18788 8988 19404 9044
rect 19460 8988 22092 9044
rect 22148 8988 23212 9044
rect 23268 8988 23660 9044
rect 23716 8988 25340 9044
rect 25396 8988 25900 9044
rect 25956 8988 25966 9044
rect 26786 8988 26796 9044
rect 26852 8988 28868 9044
rect 38658 8988 38668 9044
rect 38724 8988 50204 9044
rect 50260 8988 50270 9044
rect 0 8960 800 8988
rect 28812 8932 28868 8988
rect 9314 8876 9324 8932
rect 9380 8876 10332 8932
rect 10388 8876 10398 8932
rect 13794 8876 13804 8932
rect 13860 8876 14588 8932
rect 14644 8876 14654 8932
rect 19506 8876 19516 8932
rect 19572 8876 20076 8932
rect 20132 8876 20142 8932
rect 21410 8876 21420 8932
rect 21476 8876 26348 8932
rect 26404 8876 26414 8932
rect 26674 8876 26684 8932
rect 26740 8876 27468 8932
rect 27524 8876 27534 8932
rect 28802 8876 28812 8932
rect 28868 8876 32732 8932
rect 32788 8876 32798 8932
rect 34524 8876 35868 8932
rect 35924 8876 35934 8932
rect 34524 8820 34580 8876
rect 18722 8764 18732 8820
rect 18788 8764 20188 8820
rect 20244 8764 20254 8820
rect 26562 8764 26572 8820
rect 26628 8764 34580 8820
rect 34738 8764 34748 8820
rect 34804 8764 37100 8820
rect 37156 8764 37166 8820
rect 43586 8764 43596 8820
rect 43652 8764 44940 8820
rect 44996 8764 45006 8820
rect 75394 8764 75404 8820
rect 75460 8764 75852 8820
rect 75908 8764 75918 8820
rect 20402 8652 20412 8708
rect 20468 8652 32396 8708
rect 32452 8652 32462 8708
rect 4466 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4750 8652
rect 35186 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35470 8652
rect 65906 8596 65916 8652
rect 65972 8596 66020 8652
rect 66076 8596 66124 8652
rect 66180 8596 66190 8652
rect 79200 8596 80000 8624
rect 14914 8540 14924 8596
rect 14980 8540 15372 8596
rect 15428 8540 15438 8596
rect 16370 8540 16380 8596
rect 16436 8540 28196 8596
rect 78194 8540 78204 8596
rect 78260 8540 80000 8596
rect 28140 8484 28196 8540
rect 79200 8512 80000 8540
rect 8866 8428 8876 8484
rect 8932 8428 13132 8484
rect 13188 8428 13198 8484
rect 16706 8428 16716 8484
rect 16772 8428 19180 8484
rect 19236 8428 19246 8484
rect 25890 8428 25900 8484
rect 25956 8428 27972 8484
rect 28130 8428 28140 8484
rect 28196 8428 28206 8484
rect 28364 8428 29932 8484
rect 29988 8428 29998 8484
rect 30258 8428 30268 8484
rect 30324 8428 32284 8484
rect 32340 8428 32350 8484
rect 41122 8428 41132 8484
rect 41188 8428 42924 8484
rect 42980 8428 42990 8484
rect 27916 8372 27972 8428
rect 28364 8372 28420 8428
rect 16482 8316 16492 8372
rect 16548 8316 17836 8372
rect 17892 8316 18620 8372
rect 18676 8316 18686 8372
rect 19590 8316 19628 8372
rect 19684 8316 19694 8372
rect 19954 8316 19964 8372
rect 20020 8316 20188 8372
rect 20244 8316 20254 8372
rect 26898 8316 26908 8372
rect 26964 8316 27356 8372
rect 27412 8316 27422 8372
rect 27916 8316 28420 8372
rect 29586 8316 29596 8372
rect 29652 8316 30044 8372
rect 30100 8316 73724 8372
rect 73780 8316 73790 8372
rect 10994 8204 11004 8260
rect 11060 8204 12012 8260
rect 12068 8204 12572 8260
rect 12628 8204 12638 8260
rect 19394 8204 19404 8260
rect 19460 8204 20076 8260
rect 20132 8204 22316 8260
rect 22372 8204 22382 8260
rect 25554 8204 25564 8260
rect 25620 8204 26012 8260
rect 26068 8204 27020 8260
rect 27076 8204 27086 8260
rect 33842 8204 33852 8260
rect 33908 8204 35420 8260
rect 35476 8204 35486 8260
rect 44370 8204 44380 8260
rect 44436 8204 45276 8260
rect 45332 8204 45342 8260
rect 48514 8204 48524 8260
rect 48580 8204 59500 8260
rect 59556 8204 59566 8260
rect 76850 8204 76860 8260
rect 76916 8204 78092 8260
rect 78148 8204 78158 8260
rect 45276 8148 45332 8204
rect 9426 8092 9436 8148
rect 9492 8092 11900 8148
rect 11956 8092 11966 8148
rect 13010 8092 13020 8148
rect 13076 8092 14252 8148
rect 14308 8092 15036 8148
rect 15092 8092 16044 8148
rect 16100 8092 20188 8148
rect 20244 8092 20254 8148
rect 24658 8092 24668 8148
rect 24724 8092 25788 8148
rect 25844 8092 25854 8148
rect 26226 8092 26236 8148
rect 26292 8092 26572 8148
rect 26628 8092 26638 8148
rect 28130 8092 28140 8148
rect 28196 8092 28588 8148
rect 28644 8092 28654 8148
rect 34290 8092 34300 8148
rect 34356 8092 37100 8148
rect 37156 8092 39564 8148
rect 39620 8092 39630 8148
rect 45276 8092 73836 8148
rect 73892 8092 73902 8148
rect 76962 8092 76972 8148
rect 77028 8092 77532 8148
rect 77588 8092 77598 8148
rect 15810 7980 15820 8036
rect 15876 7980 18508 8036
rect 18564 7980 18574 8036
rect 19618 7980 19628 8036
rect 19684 7980 20692 8036
rect 27570 7980 27580 8036
rect 27636 7980 27646 8036
rect 0 7924 800 7952
rect 19628 7924 19684 7980
rect 0 7868 1708 7924
rect 1764 7868 2492 7924
rect 2548 7868 2558 7924
rect 14326 7868 14364 7924
rect 14420 7868 14430 7924
rect 17938 7868 17948 7924
rect 18004 7868 19684 7924
rect 0 7840 800 7868
rect 19826 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20110 7868
rect 20636 7812 20692 7980
rect 27580 7924 27636 7980
rect 20962 7868 20972 7924
rect 21028 7868 27636 7924
rect 28140 7812 28196 8092
rect 33394 7980 33404 8036
rect 33460 7980 34524 8036
rect 34580 7980 34590 8036
rect 41234 7980 41244 8036
rect 41300 7980 41580 8036
rect 41636 7980 41646 8036
rect 42914 7980 42924 8036
rect 42980 7980 44156 8036
rect 44212 7980 44222 8036
rect 50372 7980 53452 8036
rect 53508 7980 53518 8036
rect 50372 7924 50428 7980
rect 9650 7756 9660 7812
rect 9716 7756 10556 7812
rect 10612 7756 13692 7812
rect 13748 7756 14924 7812
rect 14980 7756 14990 7812
rect 17798 7756 17836 7812
rect 17892 7756 17902 7812
rect 18386 7756 18396 7812
rect 18452 7756 18956 7812
rect 19012 7756 19022 7812
rect 20626 7756 20636 7812
rect 20692 7756 21644 7812
rect 21700 7756 25340 7812
rect 25396 7756 26460 7812
rect 26516 7756 26526 7812
rect 26852 7756 28196 7812
rect 29148 7868 29596 7924
rect 29652 7868 29662 7924
rect 33282 7868 33292 7924
rect 33348 7868 34972 7924
rect 35028 7868 35038 7924
rect 38612 7868 44828 7924
rect 44884 7868 45948 7924
rect 46004 7868 50428 7924
rect 75954 7868 75964 7924
rect 76020 7868 76860 7924
rect 76916 7868 76926 7924
rect 26852 7700 26908 7756
rect 29148 7700 29204 7868
rect 38612 7812 38668 7868
rect 50546 7812 50556 7868
rect 50612 7812 50660 7868
rect 50716 7812 50764 7868
rect 50820 7812 50830 7868
rect 2034 7644 2044 7700
rect 2100 7644 6636 7700
rect 6692 7644 6702 7700
rect 18834 7644 18844 7700
rect 18900 7644 20300 7700
rect 20356 7644 20366 7700
rect 26338 7644 26348 7700
rect 26404 7644 26908 7700
rect 27468 7644 29204 7700
rect 29260 7756 30660 7812
rect 30818 7756 30828 7812
rect 30884 7756 38668 7812
rect 57922 7756 57932 7812
rect 57988 7756 67228 7812
rect 27468 7588 27524 7644
rect 17602 7532 17612 7588
rect 17668 7532 19740 7588
rect 19796 7532 19806 7588
rect 20178 7532 20188 7588
rect 20244 7532 20748 7588
rect 20804 7532 21196 7588
rect 21252 7532 27524 7588
rect 27682 7532 27692 7588
rect 27748 7532 28364 7588
rect 28420 7532 28430 7588
rect 27692 7476 27748 7532
rect 29260 7476 29316 7756
rect 30604 7700 30660 7756
rect 67172 7700 67228 7756
rect 30604 7644 36092 7700
rect 36148 7644 36988 7700
rect 37044 7644 37054 7700
rect 39890 7644 39900 7700
rect 39956 7644 41244 7700
rect 41300 7644 41310 7700
rect 41458 7644 41468 7700
rect 41524 7644 43036 7700
rect 43092 7644 43102 7700
rect 49858 7644 49868 7700
rect 49924 7644 66668 7700
rect 66724 7644 66734 7700
rect 67172 7644 69804 7700
rect 69860 7644 69870 7700
rect 75282 7644 75292 7700
rect 75348 7644 77420 7700
rect 77476 7644 77486 7700
rect 31266 7532 31276 7588
rect 31332 7532 32060 7588
rect 32116 7532 32126 7588
rect 35858 7532 35868 7588
rect 35924 7532 38780 7588
rect 38836 7532 38846 7588
rect 41682 7532 41692 7588
rect 41748 7532 44268 7588
rect 44324 7532 44334 7588
rect 55234 7532 55244 7588
rect 55300 7532 71708 7588
rect 71764 7532 72380 7588
rect 72436 7532 72446 7588
rect 74946 7532 74956 7588
rect 75012 7532 75404 7588
rect 75460 7532 75470 7588
rect 79200 7476 80000 7504
rect 11442 7420 11452 7476
rect 11508 7420 13468 7476
rect 13524 7420 14252 7476
rect 14308 7420 14812 7476
rect 14868 7420 14878 7476
rect 15092 7420 15484 7476
rect 15540 7420 15550 7476
rect 19618 7420 19628 7476
rect 19684 7420 19852 7476
rect 19908 7420 19918 7476
rect 20066 7420 20076 7476
rect 20132 7420 20188 7476
rect 20244 7420 20254 7476
rect 25778 7420 25788 7476
rect 25844 7420 27748 7476
rect 28252 7420 29316 7476
rect 29474 7420 29484 7476
rect 29540 7420 30940 7476
rect 30996 7420 31006 7476
rect 31714 7420 31724 7476
rect 31780 7420 32956 7476
rect 33012 7420 33740 7476
rect 33796 7420 33806 7476
rect 33964 7420 42252 7476
rect 42308 7420 42318 7476
rect 43698 7420 43708 7476
rect 43764 7420 43932 7476
rect 43988 7420 46844 7476
rect 46900 7420 49532 7476
rect 49588 7420 49598 7476
rect 53890 7420 53900 7476
rect 53956 7420 75292 7476
rect 75348 7420 76300 7476
rect 76356 7420 76366 7476
rect 77522 7420 77532 7476
rect 77588 7420 80000 7476
rect 15092 7364 15148 7420
rect 28252 7364 28308 7420
rect 33964 7364 34020 7420
rect 79200 7392 80000 7420
rect 1698 7308 1708 7364
rect 1764 7308 2492 7364
rect 2548 7308 2558 7364
rect 11666 7308 11676 7364
rect 11732 7308 15148 7364
rect 15250 7308 15260 7364
rect 15316 7308 17052 7364
rect 17108 7308 17118 7364
rect 25554 7308 25564 7364
rect 25620 7308 28308 7364
rect 28466 7308 28476 7364
rect 28532 7308 29372 7364
rect 29428 7308 34020 7364
rect 34402 7308 34412 7364
rect 34468 7308 35196 7364
rect 35252 7308 35262 7364
rect 35410 7308 35420 7364
rect 35476 7308 35756 7364
rect 35812 7308 35822 7364
rect 41458 7308 41468 7364
rect 41524 7308 41916 7364
rect 41972 7308 41982 7364
rect 29820 7252 29876 7308
rect 18386 7196 18396 7252
rect 18452 7196 25452 7252
rect 25508 7196 25518 7252
rect 26852 7196 27692 7252
rect 27748 7196 27758 7252
rect 29810 7196 29820 7252
rect 29876 7196 29886 7252
rect 34850 7196 34860 7252
rect 34916 7196 35532 7252
rect 35588 7196 37436 7252
rect 37492 7196 37502 7252
rect 48402 7196 48412 7252
rect 48468 7196 67116 7252
rect 67172 7196 67182 7252
rect 75394 7196 75404 7252
rect 75460 7196 76524 7252
rect 76580 7196 76590 7252
rect 26852 7140 26908 7196
rect 22418 7084 22428 7140
rect 22484 7084 22876 7140
rect 22932 7084 26908 7140
rect 41570 7084 41580 7140
rect 41636 7084 43148 7140
rect 43204 7084 47404 7140
rect 47460 7084 47470 7140
rect 4466 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4750 7084
rect 35186 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35470 7084
rect 65906 7028 65916 7084
rect 65972 7028 66020 7084
rect 66076 7028 66124 7084
rect 66180 7028 66190 7084
rect 23202 6972 23212 7028
rect 23268 6972 23436 7028
rect 23492 6972 23502 7028
rect 24770 6972 24780 7028
rect 24836 6972 25788 7028
rect 25844 6972 25854 7028
rect 37762 6972 37772 7028
rect 37828 6972 39900 7028
rect 39956 6972 40908 7028
rect 40964 6972 40974 7028
rect 43026 6972 43036 7028
rect 43092 6972 45724 7028
rect 45780 6972 45790 7028
rect 7410 6860 7420 6916
rect 7476 6860 10892 6916
rect 10948 6860 10958 6916
rect 11218 6860 11228 6916
rect 11284 6860 14140 6916
rect 14196 6860 14206 6916
rect 24098 6860 24108 6916
rect 24164 6860 26124 6916
rect 26180 6860 26190 6916
rect 27794 6860 27804 6916
rect 27860 6860 28252 6916
rect 28308 6860 29148 6916
rect 29204 6860 29708 6916
rect 29764 6860 38556 6916
rect 38612 6860 38622 6916
rect 39218 6860 39228 6916
rect 39284 6860 44380 6916
rect 44436 6860 44446 6916
rect 0 6804 800 6832
rect 0 6748 1708 6804
rect 1764 6748 1774 6804
rect 2706 6748 2716 6804
rect 2772 6748 7532 6804
rect 7588 6748 7598 6804
rect 8418 6748 8428 6804
rect 8484 6748 9100 6804
rect 9156 6748 9772 6804
rect 9828 6748 9838 6804
rect 9996 6748 18732 6804
rect 18788 6748 18798 6804
rect 22530 6748 22540 6804
rect 22596 6748 23380 6804
rect 0 6720 800 6748
rect 9996 6692 10052 6748
rect 9884 6636 10052 6692
rect 13234 6636 13244 6692
rect 13300 6636 13916 6692
rect 13972 6636 13982 6692
rect 14914 6636 14924 6692
rect 14980 6636 16380 6692
rect 16436 6636 16446 6692
rect 17126 6636 17164 6692
rect 17220 6636 17230 6692
rect 18162 6636 18172 6692
rect 18228 6636 19628 6692
rect 19684 6636 19694 6692
rect 9884 6580 9940 6636
rect 23324 6580 23380 6748
rect 23660 6748 25676 6804
rect 25732 6748 25742 6804
rect 26002 6748 26012 6804
rect 26068 6748 26348 6804
rect 26404 6748 26414 6804
rect 39330 6748 39340 6804
rect 39396 6748 40124 6804
rect 40180 6748 44268 6804
rect 44324 6748 44334 6804
rect 75170 6748 75180 6804
rect 75236 6748 77532 6804
rect 77588 6748 77598 6804
rect 23660 6580 23716 6748
rect 27234 6636 27244 6692
rect 27300 6636 27916 6692
rect 27972 6636 27982 6692
rect 33964 6636 36204 6692
rect 36260 6636 36270 6692
rect 49074 6636 49084 6692
rect 49140 6636 56812 6692
rect 56868 6636 56878 6692
rect 61282 6636 61292 6692
rect 61348 6636 63420 6692
rect 63476 6636 63486 6692
rect 73714 6636 73724 6692
rect 73780 6636 76636 6692
rect 76692 6636 76702 6692
rect 33964 6580 34020 6636
rect 9874 6524 9884 6580
rect 9940 6524 9950 6580
rect 12124 6524 15148 6580
rect 16146 6524 16156 6580
rect 16212 6524 20636 6580
rect 20692 6524 20702 6580
rect 23314 6524 23324 6580
rect 23380 6524 23390 6580
rect 23650 6524 23660 6580
rect 23716 6524 23726 6580
rect 23884 6524 28028 6580
rect 28084 6524 28094 6580
rect 28690 6524 28700 6580
rect 28756 6524 29260 6580
rect 29316 6524 30156 6580
rect 30212 6524 30222 6580
rect 33394 6524 33404 6580
rect 33460 6524 33740 6580
rect 33796 6524 33806 6580
rect 33954 6524 33964 6580
rect 34020 6524 34030 6580
rect 34402 6524 34412 6580
rect 34468 6524 34972 6580
rect 35028 6524 35038 6580
rect 36082 6524 36092 6580
rect 36148 6524 38220 6580
rect 38276 6524 38286 6580
rect 48626 6524 48636 6580
rect 48692 6524 49644 6580
rect 49700 6524 49710 6580
rect 51202 6524 51212 6580
rect 51268 6524 51996 6580
rect 52052 6524 76188 6580
rect 76244 6524 76254 6580
rect 12124 6468 12180 6524
rect 6290 6412 6300 6468
rect 6356 6412 8204 6468
rect 8260 6412 8270 6468
rect 12114 6412 12124 6468
rect 12180 6412 12190 6468
rect 13458 6412 13468 6468
rect 13524 6412 14028 6468
rect 14084 6412 14094 6468
rect 14466 6412 14476 6468
rect 14532 6412 14542 6468
rect 14690 6412 14700 6468
rect 14756 6412 14794 6468
rect 14476 6244 14532 6412
rect 15092 6356 15148 6524
rect 23884 6468 23940 6524
rect 15698 6412 15708 6468
rect 15764 6412 19516 6468
rect 19572 6412 19582 6468
rect 20066 6412 20076 6468
rect 20132 6412 23940 6468
rect 24658 6412 24668 6468
rect 24724 6412 25340 6468
rect 25396 6412 25406 6468
rect 28354 6412 28364 6468
rect 28420 6412 29372 6468
rect 29428 6412 30044 6468
rect 30100 6412 30110 6468
rect 30930 6412 30940 6468
rect 30996 6412 33852 6468
rect 33908 6412 33918 6468
rect 34066 6412 34076 6468
rect 34132 6412 35868 6468
rect 35924 6412 35934 6468
rect 38612 6412 50484 6468
rect 50754 6412 50764 6468
rect 50820 6412 51884 6468
rect 51940 6412 55468 6468
rect 60050 6412 60060 6468
rect 60116 6412 61516 6468
rect 61572 6412 61582 6468
rect 62738 6412 62748 6468
rect 62804 6412 64428 6468
rect 64484 6412 64494 6468
rect 70466 6412 70476 6468
rect 70532 6412 72268 6468
rect 72324 6412 72334 6468
rect 76738 6412 76748 6468
rect 76804 6412 77756 6468
rect 77812 6412 77822 6468
rect 15092 6300 17164 6356
rect 17220 6300 17230 6356
rect 21942 6300 21980 6356
rect 22036 6300 22046 6356
rect 23538 6300 23548 6356
rect 23604 6300 26908 6356
rect 27794 6300 27804 6356
rect 27860 6300 28700 6356
rect 28756 6300 28766 6356
rect 29698 6300 29708 6356
rect 29764 6300 30828 6356
rect 30884 6300 30894 6356
rect 31378 6300 31388 6356
rect 31444 6300 32172 6356
rect 32228 6300 33068 6356
rect 33124 6300 33134 6356
rect 19826 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20110 6300
rect 26852 6244 26908 6300
rect 38612 6244 38668 6412
rect 45266 6300 45276 6356
rect 45332 6300 46284 6356
rect 46340 6300 46350 6356
rect 10434 6188 10444 6244
rect 10500 6188 12236 6244
rect 12292 6188 12302 6244
rect 14476 6188 19068 6244
rect 19124 6188 19134 6244
rect 21522 6188 21532 6244
rect 21588 6188 22820 6244
rect 26852 6188 28252 6244
rect 28308 6188 28318 6244
rect 28578 6188 28588 6244
rect 28644 6188 38668 6244
rect 22764 6132 22820 6188
rect 50428 6132 50484 6412
rect 55412 6356 55468 6412
rect 79200 6356 80000 6384
rect 51202 6300 51212 6356
rect 51268 6300 53004 6356
rect 53060 6300 53070 6356
rect 55412 6300 74508 6356
rect 74564 6300 75516 6356
rect 75572 6300 75582 6356
rect 78306 6300 78316 6356
rect 78372 6300 80000 6356
rect 50546 6244 50556 6300
rect 50612 6244 50660 6300
rect 50716 6244 50764 6300
rect 50820 6244 50830 6300
rect 79200 6272 80000 6300
rect 8306 6076 8316 6132
rect 8372 6076 13244 6132
rect 13300 6076 13310 6132
rect 16146 6076 16156 6132
rect 16212 6076 18788 6132
rect 22764 6076 25788 6132
rect 25844 6076 25854 6132
rect 26852 6076 28140 6132
rect 28196 6076 28206 6132
rect 29148 6076 29708 6132
rect 29764 6076 29774 6132
rect 30482 6076 30492 6132
rect 30548 6076 31052 6132
rect 31108 6076 31118 6132
rect 32162 6076 32172 6132
rect 32228 6076 33180 6132
rect 33236 6076 33246 6132
rect 33730 6076 33740 6132
rect 33796 6076 34412 6132
rect 34468 6076 34478 6132
rect 38612 6076 38780 6132
rect 38836 6076 38846 6132
rect 40114 6076 40124 6132
rect 40180 6076 48748 6132
rect 48804 6076 48814 6132
rect 50428 6076 51548 6132
rect 51604 6076 52108 6132
rect 52164 6076 53004 6132
rect 53060 6076 53070 6132
rect 55412 6076 67564 6132
rect 67620 6076 67630 6132
rect 18732 6020 18788 6076
rect 10658 5964 10668 6020
rect 10724 5964 11228 6020
rect 11284 5964 11294 6020
rect 13010 5964 13020 6020
rect 13076 5964 13580 6020
rect 13636 5964 13646 6020
rect 13906 5964 13916 6020
rect 13972 5964 14812 6020
rect 14868 5964 14878 6020
rect 17154 5964 17164 6020
rect 17220 5964 17388 6020
rect 17444 5964 17454 6020
rect 18732 5964 22764 6020
rect 22820 5964 22830 6020
rect 26852 5908 26908 6076
rect 29148 6020 29204 6076
rect 6738 5852 6748 5908
rect 6804 5852 8652 5908
rect 8708 5852 8718 5908
rect 9874 5852 9884 5908
rect 9940 5852 14476 5908
rect 14532 5852 17276 5908
rect 17332 5852 17342 5908
rect 18946 5852 18956 5908
rect 19012 5852 21196 5908
rect 21252 5852 21262 5908
rect 21522 5852 21532 5908
rect 21588 5852 22204 5908
rect 22260 5852 22270 5908
rect 26562 5852 26572 5908
rect 26628 5852 26908 5908
rect 27692 5964 29148 6020
rect 29204 5964 29214 6020
rect 29362 5964 29372 6020
rect 29428 5964 35084 6020
rect 35140 5964 35150 6020
rect 27692 5796 27748 5964
rect 27906 5852 27916 5908
rect 27972 5852 29260 5908
rect 29316 5852 29326 5908
rect 30034 5852 30044 5908
rect 30100 5852 31052 5908
rect 31108 5852 31118 5908
rect 32610 5852 32620 5908
rect 32676 5852 36092 5908
rect 36148 5852 36158 5908
rect 38612 5796 38668 6076
rect 55412 6020 55468 6076
rect 41122 5964 41132 6020
rect 41188 5964 45612 6020
rect 45668 5964 45678 6020
rect 46722 5964 46732 6020
rect 46788 5964 47740 6020
rect 47796 5964 47806 6020
rect 48178 5964 48188 6020
rect 48244 5964 55468 6020
rect 40898 5852 40908 5908
rect 40964 5852 42476 5908
rect 42532 5852 42542 5908
rect 44258 5852 44268 5908
rect 44324 5852 44492 5908
rect 44548 5852 44558 5908
rect 46946 5852 46956 5908
rect 47012 5852 48972 5908
rect 49028 5852 49038 5908
rect 56018 5852 56028 5908
rect 56084 5852 56924 5908
rect 56980 5852 56990 5908
rect 57138 5852 57148 5908
rect 57204 5852 71036 5908
rect 71092 5852 71102 5908
rect 74386 5852 74396 5908
rect 74452 5852 75180 5908
rect 75236 5852 75246 5908
rect 2034 5740 2044 5796
rect 2100 5740 6972 5796
rect 7028 5740 7038 5796
rect 7186 5740 7196 5796
rect 7252 5740 12460 5796
rect 12516 5740 12526 5796
rect 13122 5740 13132 5796
rect 13188 5740 16828 5796
rect 16884 5740 16894 5796
rect 19506 5740 19516 5796
rect 19572 5740 24220 5796
rect 24276 5740 24286 5796
rect 25442 5740 25452 5796
rect 25508 5740 27748 5796
rect 30258 5740 30268 5796
rect 30324 5740 31836 5796
rect 31892 5740 31902 5796
rect 32162 5740 32172 5796
rect 32228 5740 39284 5796
rect 40450 5740 40460 5796
rect 40516 5740 42700 5796
rect 42756 5740 42766 5796
rect 49186 5740 49196 5796
rect 49252 5740 49756 5796
rect 49812 5740 49822 5796
rect 52434 5740 52444 5796
rect 52500 5740 71708 5796
rect 71764 5740 72268 5796
rect 72324 5740 72334 5796
rect 0 5684 800 5712
rect 39228 5684 39284 5740
rect 0 5628 1708 5684
rect 1764 5628 2492 5684
rect 2548 5628 2558 5684
rect 4274 5628 4284 5684
rect 4340 5628 9548 5684
rect 9604 5628 9614 5684
rect 12562 5628 12572 5684
rect 12628 5628 15372 5684
rect 15428 5628 15438 5684
rect 19394 5628 19404 5684
rect 19460 5628 21868 5684
rect 21924 5628 21934 5684
rect 23426 5628 23436 5684
rect 23492 5628 26012 5684
rect 26068 5628 26078 5684
rect 27234 5628 27244 5684
rect 27300 5628 27692 5684
rect 27748 5628 27758 5684
rect 29250 5628 29260 5684
rect 29316 5628 30156 5684
rect 30212 5628 30222 5684
rect 33730 5628 33740 5684
rect 33796 5628 34300 5684
rect 34356 5628 39004 5684
rect 39060 5628 39070 5684
rect 39228 5628 41020 5684
rect 41076 5628 48748 5684
rect 48804 5628 48814 5684
rect 56690 5628 56700 5684
rect 56756 5628 57932 5684
rect 57988 5628 57998 5684
rect 59378 5628 59388 5684
rect 59444 5628 60844 5684
rect 60900 5628 60910 5684
rect 69010 5628 69020 5684
rect 69076 5628 70532 5684
rect 70802 5628 70812 5684
rect 70868 5628 73276 5684
rect 73332 5628 73342 5684
rect 0 5600 800 5628
rect 70476 5572 70532 5628
rect 7858 5516 7868 5572
rect 7924 5516 9436 5572
rect 9492 5516 9502 5572
rect 13682 5516 13692 5572
rect 13748 5516 14364 5572
rect 14420 5516 14430 5572
rect 14802 5516 14812 5572
rect 14868 5516 17836 5572
rect 17892 5516 17902 5572
rect 21522 5516 21532 5572
rect 21588 5516 27804 5572
rect 27860 5516 27870 5572
rect 29698 5516 29708 5572
rect 29764 5516 34412 5572
rect 34468 5516 34478 5572
rect 45938 5516 45948 5572
rect 46004 5516 47964 5572
rect 48020 5516 48030 5572
rect 50372 5516 50876 5572
rect 50932 5516 50942 5572
rect 67330 5516 67340 5572
rect 67396 5516 69356 5572
rect 69412 5516 69422 5572
rect 70466 5516 70476 5572
rect 70532 5516 75404 5572
rect 75460 5516 75470 5572
rect 4466 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4750 5516
rect 35186 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35470 5516
rect 50372 5460 50428 5516
rect 65906 5460 65916 5516
rect 65972 5460 66020 5516
rect 66076 5460 66124 5516
rect 66180 5460 66190 5516
rect 7410 5404 7420 5460
rect 7476 5404 9156 5460
rect 9314 5404 9324 5460
rect 9380 5404 15260 5460
rect 15316 5404 15326 5460
rect 19954 5404 19964 5460
rect 20020 5404 23660 5460
rect 23716 5404 23726 5460
rect 25442 5404 25452 5460
rect 25508 5404 26348 5460
rect 26404 5404 26414 5460
rect 26674 5404 26684 5460
rect 26740 5404 28420 5460
rect 28578 5404 28588 5460
rect 28644 5404 32620 5460
rect 32676 5404 32686 5460
rect 36306 5404 36316 5460
rect 36372 5404 36876 5460
rect 36932 5404 37548 5460
rect 37604 5404 37614 5460
rect 42466 5404 42476 5460
rect 42532 5404 44828 5460
rect 44884 5404 44894 5460
rect 46722 5404 46732 5460
rect 46788 5404 49308 5460
rect 49364 5404 50428 5460
rect 73826 5404 73836 5460
rect 73892 5404 74620 5460
rect 74676 5404 74686 5460
rect 74946 5404 74956 5460
rect 75012 5404 75628 5460
rect 75684 5404 75694 5460
rect 9100 5348 9156 5404
rect 4946 5292 4956 5348
rect 5012 5292 8876 5348
rect 8932 5292 8942 5348
rect 9100 5292 9548 5348
rect 9604 5292 10108 5348
rect 10164 5292 11340 5348
rect 11396 5292 11406 5348
rect 13234 5292 13244 5348
rect 13300 5292 13692 5348
rect 13748 5292 13758 5348
rect 14018 5292 14028 5348
rect 14084 5292 15148 5348
rect 15204 5292 15214 5348
rect 18386 5292 18396 5348
rect 18452 5292 22204 5348
rect 22260 5292 22270 5348
rect 22418 5292 22428 5348
rect 22484 5292 28196 5348
rect 8194 5180 8204 5236
rect 8260 5180 10668 5236
rect 10724 5180 10734 5236
rect 10882 5180 10892 5236
rect 10948 5180 13580 5236
rect 13636 5180 13646 5236
rect 13906 5180 13916 5236
rect 13972 5180 14364 5236
rect 14420 5180 14430 5236
rect 17378 5180 17388 5236
rect 17444 5180 17780 5236
rect 21634 5180 21644 5236
rect 21700 5180 23884 5236
rect 23940 5180 23950 5236
rect 26002 5180 26012 5236
rect 26068 5180 27244 5236
rect 27300 5180 27310 5236
rect 17724 5124 17780 5180
rect 28140 5124 28196 5292
rect 28364 5236 28420 5404
rect 29586 5292 29596 5348
rect 29652 5292 30268 5348
rect 30324 5292 30492 5348
rect 30548 5292 30558 5348
rect 30716 5292 31276 5348
rect 31332 5292 31342 5348
rect 31826 5292 31836 5348
rect 31892 5292 36428 5348
rect 36484 5292 38668 5348
rect 38724 5292 38734 5348
rect 41906 5292 41916 5348
rect 41972 5292 48300 5348
rect 48356 5292 48366 5348
rect 73490 5292 73500 5348
rect 73556 5292 76300 5348
rect 76356 5292 76366 5348
rect 30716 5236 30772 5292
rect 79200 5236 80000 5264
rect 28364 5180 30772 5236
rect 31042 5180 31052 5236
rect 31108 5180 34076 5236
rect 34132 5180 34142 5236
rect 37650 5180 37660 5236
rect 37716 5180 40124 5236
rect 40180 5180 40190 5236
rect 47506 5180 47516 5236
rect 47572 5180 49868 5236
rect 49924 5180 51324 5236
rect 51380 5180 51390 5236
rect 53890 5180 53900 5236
rect 53956 5180 55244 5236
rect 55300 5180 55310 5236
rect 56130 5180 56140 5236
rect 56196 5180 58156 5236
rect 58212 5180 58222 5236
rect 60722 5180 60732 5236
rect 60788 5180 64428 5236
rect 64484 5180 64494 5236
rect 66322 5180 66332 5236
rect 66388 5180 69356 5236
rect 69412 5180 69422 5236
rect 72818 5180 72828 5236
rect 72884 5180 76188 5236
rect 76244 5180 76254 5236
rect 77634 5180 77644 5236
rect 77700 5180 80000 5236
rect 79200 5152 80000 5180
rect 8754 5068 8764 5124
rect 8820 5068 11564 5124
rect 11620 5068 11630 5124
rect 11890 5068 11900 5124
rect 11956 5068 12460 5124
rect 12516 5068 12526 5124
rect 13010 5068 13020 5124
rect 13076 5068 14140 5124
rect 14196 5068 14700 5124
rect 14756 5068 14766 5124
rect 15372 5068 17500 5124
rect 17556 5068 17566 5124
rect 17724 5068 21924 5124
rect 23314 5068 23324 5124
rect 23380 5068 26460 5124
rect 26516 5068 26526 5124
rect 28140 5068 29260 5124
rect 29316 5068 29326 5124
rect 30146 5068 30156 5124
rect 30212 5068 30716 5124
rect 30772 5068 30782 5124
rect 31266 5068 31276 5124
rect 31332 5068 33852 5124
rect 33908 5068 33918 5124
rect 38098 5068 38108 5124
rect 38164 5068 42476 5124
rect 42532 5068 42542 5124
rect 44258 5068 44268 5124
rect 44324 5068 46844 5124
rect 46900 5068 46910 5124
rect 48066 5068 48076 5124
rect 48132 5068 49196 5124
rect 49252 5068 49262 5124
rect 49522 5068 49532 5124
rect 49588 5068 50428 5124
rect 50484 5068 50494 5124
rect 59938 5068 59948 5124
rect 60004 5068 60508 5124
rect 60564 5068 60574 5124
rect 63746 5068 63756 5124
rect 63812 5068 65548 5124
rect 65604 5068 65614 5124
rect 66770 5068 66780 5124
rect 66836 5068 68572 5124
rect 68628 5068 68638 5124
rect 72146 5068 72156 5124
rect 72212 5068 73948 5124
rect 74004 5068 74014 5124
rect 74946 5068 74956 5124
rect 75012 5068 75740 5124
rect 75796 5068 76300 5124
rect 76356 5068 76366 5124
rect 15372 5012 15428 5068
rect 8418 4956 8428 5012
rect 8484 4956 9044 5012
rect 9202 4956 9212 5012
rect 9268 4956 9884 5012
rect 9940 4956 9950 5012
rect 12562 4956 12572 5012
rect 12628 4956 13916 5012
rect 13972 4956 13982 5012
rect 15362 4956 15372 5012
rect 15428 4956 15438 5012
rect 17938 4956 17948 5012
rect 18004 4956 18172 5012
rect 18228 4956 18284 5012
rect 18340 4956 18350 5012
rect 20374 4956 20412 5012
rect 20468 4956 20478 5012
rect 8988 4900 9044 4956
rect 21868 4900 21924 5068
rect 22082 4956 22092 5012
rect 22148 4956 22540 5012
rect 22596 4956 23548 5012
rect 23604 4956 23614 5012
rect 30594 4956 30604 5012
rect 30660 4956 33516 5012
rect 33572 4956 33582 5012
rect 38994 4956 39004 5012
rect 39060 4956 41020 5012
rect 41076 4956 41086 5012
rect 46498 4956 46508 5012
rect 46564 4956 50316 5012
rect 50372 4956 50382 5012
rect 73378 4956 73388 5012
rect 73444 4956 74508 5012
rect 74564 4956 74574 5012
rect 5170 4844 5180 4900
rect 5236 4844 6412 4900
rect 6468 4844 6478 4900
rect 6850 4844 6860 4900
rect 6916 4844 8652 4900
rect 8708 4844 8718 4900
rect 8988 4844 10332 4900
rect 10388 4844 11676 4900
rect 11732 4844 11742 4900
rect 12338 4844 12348 4900
rect 12404 4844 13468 4900
rect 13524 4844 13534 4900
rect 19292 4844 21700 4900
rect 21858 4844 21868 4900
rect 21924 4844 21934 4900
rect 23174 4844 23212 4900
rect 23268 4844 23278 4900
rect 26852 4844 30044 4900
rect 30100 4844 30110 4900
rect 40002 4844 40012 4900
rect 40068 4844 40684 4900
rect 40740 4844 45388 4900
rect 45444 4844 45454 4900
rect 51650 4844 51660 4900
rect 51716 4844 52780 4900
rect 52836 4844 52846 4900
rect 58706 4844 58716 4900
rect 58772 4844 61516 4900
rect 61572 4844 61582 4900
rect 68114 4844 68124 4900
rect 68180 4844 72268 4900
rect 72324 4844 72334 4900
rect 75170 4844 75180 4900
rect 75236 4844 76972 4900
rect 77028 4844 77038 4900
rect 19292 4788 19348 4844
rect 2034 4732 2044 4788
rect 2100 4732 5964 4788
rect 6020 4732 6030 4788
rect 6178 4732 6188 4788
rect 6244 4732 9772 4788
rect 9828 4732 9838 4788
rect 15138 4732 15148 4788
rect 15204 4732 15484 4788
rect 15540 4732 15550 4788
rect 17042 4732 17052 4788
rect 17108 4732 18284 4788
rect 18340 4732 18350 4788
rect 19058 4732 19068 4788
rect 19124 4732 19292 4788
rect 19348 4732 19358 4788
rect 19826 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20110 4732
rect 21644 4676 21700 4844
rect 26852 4788 26908 4844
rect 22642 4732 22652 4788
rect 22708 4732 26908 4788
rect 30930 4732 30940 4788
rect 30996 4732 31836 4788
rect 31892 4732 38556 4788
rect 38612 4732 38622 4788
rect 50546 4676 50556 4732
rect 50612 4676 50660 4732
rect 50716 4676 50764 4732
rect 50820 4676 50830 4732
rect 7074 4620 7084 4676
rect 7140 4620 7196 4676
rect 7252 4620 7262 4676
rect 21644 4620 22876 4676
rect 22932 4620 22942 4676
rect 32498 4620 32508 4676
rect 32564 4620 40348 4676
rect 40404 4620 40414 4676
rect 53666 4620 53676 4676
rect 53732 4620 55468 4676
rect 0 4564 800 4592
rect 0 4508 1708 4564
rect 1764 4508 2492 4564
rect 2548 4508 2558 4564
rect 7970 4508 7980 4564
rect 8036 4508 8820 4564
rect 9426 4508 9436 4564
rect 9492 4508 14252 4564
rect 14308 4508 14318 4564
rect 16482 4508 16492 4564
rect 16548 4508 19068 4564
rect 19124 4508 20412 4564
rect 20468 4508 20478 4564
rect 22418 4508 22428 4564
rect 22484 4508 22988 4564
rect 23044 4508 24444 4564
rect 24500 4508 24510 4564
rect 27122 4508 27132 4564
rect 27188 4508 32732 4564
rect 32788 4508 32798 4564
rect 39218 4508 39228 4564
rect 39284 4508 40908 4564
rect 40964 4508 40974 4564
rect 45490 4508 45500 4564
rect 45556 4508 46396 4564
rect 46452 4508 47404 4564
rect 47460 4508 47470 4564
rect 0 4480 800 4508
rect 8764 4452 8820 4508
rect 7634 4396 7644 4452
rect 7700 4396 8316 4452
rect 8372 4396 8382 4452
rect 8754 4396 8764 4452
rect 8820 4396 8830 4452
rect 9762 4396 9772 4452
rect 9828 4396 13468 4452
rect 13524 4396 13534 4452
rect 14802 4396 14812 4452
rect 14868 4396 20300 4452
rect 20356 4396 20366 4452
rect 20626 4396 20636 4452
rect 20692 4396 21308 4452
rect 21364 4396 21980 4452
rect 22036 4396 22046 4452
rect 24658 4396 24668 4452
rect 24724 4396 31276 4452
rect 31332 4396 31342 4452
rect 36530 4396 36540 4452
rect 36596 4396 39116 4452
rect 39172 4396 39182 4452
rect 46610 4396 46620 4452
rect 46676 4396 47628 4452
rect 47684 4396 47694 4452
rect 55412 4340 55468 4620
rect 61618 4508 61628 4564
rect 61684 4508 62524 4564
rect 62580 4508 62590 4564
rect 75618 4508 75628 4564
rect 75684 4508 76412 4564
rect 76468 4508 77196 4564
rect 77252 4508 78204 4564
rect 78260 4508 78270 4564
rect 6066 4284 6076 4340
rect 6132 4284 7980 4340
rect 8036 4284 8046 4340
rect 9874 4284 9884 4340
rect 9940 4284 16492 4340
rect 16548 4284 16558 4340
rect 16818 4284 16828 4340
rect 16884 4284 17836 4340
rect 17892 4284 17902 4340
rect 20290 4284 20300 4340
rect 20356 4284 22988 4340
rect 23044 4284 23054 4340
rect 26450 4284 26460 4340
rect 26516 4284 28700 4340
rect 28756 4284 28766 4340
rect 31378 4284 31388 4340
rect 31444 4284 32396 4340
rect 32452 4284 41132 4340
rect 41188 4284 41198 4340
rect 41906 4284 41916 4340
rect 41972 4284 43260 4340
rect 43316 4284 43326 4340
rect 43586 4284 43596 4340
rect 43652 4284 48972 4340
rect 49028 4284 49038 4340
rect 55412 4284 70476 4340
rect 70532 4284 70542 4340
rect 10210 4172 10220 4228
rect 10276 4172 13356 4228
rect 13412 4172 13422 4228
rect 15138 4172 15148 4228
rect 15204 4172 17052 4228
rect 17108 4172 17118 4228
rect 17266 4172 17276 4228
rect 17332 4172 19404 4228
rect 19460 4172 19470 4228
rect 19618 4172 19628 4228
rect 19684 4172 21532 4228
rect 21588 4172 21598 4228
rect 22194 4172 22204 4228
rect 22260 4172 22316 4228
rect 22372 4172 22708 4228
rect 23202 4172 23212 4228
rect 23268 4172 26012 4228
rect 26068 4172 26078 4228
rect 31826 4172 31836 4228
rect 31892 4172 33628 4228
rect 33684 4172 33694 4228
rect 35074 4172 35084 4228
rect 35140 4172 43708 4228
rect 43764 4172 43774 4228
rect 53778 4172 53788 4228
rect 53844 4172 71708 4228
rect 71764 4172 72268 4228
rect 72324 4172 72334 4228
rect 73042 4172 73052 4228
rect 73108 4172 74172 4228
rect 74228 4172 74238 4228
rect 7410 4060 7420 4116
rect 7476 4060 10108 4116
rect 10164 4060 10174 4116
rect 10882 4060 10892 4116
rect 10948 4060 11452 4116
rect 11508 4060 11518 4116
rect 16818 4060 16828 4116
rect 16884 4060 17948 4116
rect 18004 4060 18014 4116
rect 18610 4060 18620 4116
rect 18676 4060 19292 4116
rect 19348 4060 22428 4116
rect 22484 4060 22494 4116
rect 22652 4004 22708 4172
rect 79200 4116 80000 4144
rect 24322 4060 24332 4116
rect 24388 4060 30044 4116
rect 30100 4060 30110 4116
rect 30930 4060 30940 4116
rect 30996 4060 37100 4116
rect 37156 4060 37166 4116
rect 42690 4060 42700 4116
rect 42756 4060 49084 4116
rect 49140 4060 49150 4116
rect 49298 4060 49308 4116
rect 49364 4060 50540 4116
rect 50596 4060 50606 4116
rect 52658 4060 52668 4116
rect 52724 4060 53900 4116
rect 53956 4060 53966 4116
rect 54674 4060 54684 4116
rect 54740 4060 57596 4116
rect 57652 4060 57662 4116
rect 64082 4060 64092 4116
rect 64148 4060 68348 4116
rect 68404 4060 68414 4116
rect 68786 4060 68796 4116
rect 68852 4060 73276 4116
rect 73332 4060 73342 4116
rect 75170 4060 75180 4116
rect 75236 4060 80000 4116
rect 79200 4032 80000 4060
rect 8754 3948 8764 4004
rect 8820 3948 10332 4004
rect 10388 3948 10398 4004
rect 10770 3948 10780 4004
rect 10836 3948 11228 4004
rect 11284 3948 11956 4004
rect 12562 3948 12572 4004
rect 12628 3948 21756 4004
rect 21812 3948 21822 4004
rect 22652 3948 27916 4004
rect 27972 3948 27982 4004
rect 28354 3948 28364 4004
rect 28420 3948 31836 4004
rect 31892 3948 31902 4004
rect 70466 3948 70476 4004
rect 70532 3948 74060 4004
rect 74116 3948 74126 4004
rect 4466 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4750 3948
rect 11900 3892 11956 3948
rect 35186 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35470 3948
rect 65906 3892 65916 3948
rect 65972 3892 66020 3948
rect 66076 3892 66124 3948
rect 66180 3892 66190 3948
rect 5618 3836 5628 3892
rect 5684 3836 6748 3892
rect 6804 3836 7644 3892
rect 7700 3836 7710 3892
rect 7858 3836 7868 3892
rect 7924 3836 11060 3892
rect 11900 3836 14812 3892
rect 14868 3836 14878 3892
rect 15026 3836 15036 3892
rect 15092 3836 20860 3892
rect 20916 3836 20926 3892
rect 23986 3836 23996 3892
rect 24052 3836 29260 3892
rect 29316 3836 29326 3892
rect 41906 3836 41916 3892
rect 41972 3836 47964 3892
rect 48020 3836 48524 3892
rect 48580 3836 48590 3892
rect 49858 3836 49868 3892
rect 49924 3836 51772 3892
rect 51828 3836 51838 3892
rect 62066 3836 62076 3892
rect 62132 3836 65828 3892
rect 11004 3780 11060 3836
rect 65772 3780 65828 3836
rect 6402 3724 6412 3780
rect 6468 3724 8988 3780
rect 9044 3724 9054 3780
rect 10210 3724 10220 3780
rect 10276 3724 10780 3780
rect 10836 3724 10846 3780
rect 10994 3724 11004 3780
rect 11060 3724 11070 3780
rect 14578 3724 14588 3780
rect 14644 3724 15596 3780
rect 15652 3724 15662 3780
rect 16930 3724 16940 3780
rect 16996 3724 19684 3780
rect 20262 3724 20300 3780
rect 20356 3724 20366 3780
rect 20598 3724 20636 3780
rect 20692 3724 20702 3780
rect 20962 3724 20972 3780
rect 21028 3724 24556 3780
rect 24612 3724 24622 3780
rect 24770 3724 24780 3780
rect 24836 3724 26068 3780
rect 26226 3724 26236 3780
rect 26292 3724 29092 3780
rect 30258 3724 30268 3780
rect 30324 3724 38668 3780
rect 39106 3724 39116 3780
rect 39172 3724 42588 3780
rect 42644 3724 42654 3780
rect 42802 3724 42812 3780
rect 42868 3724 44268 3780
rect 44324 3724 44334 3780
rect 44594 3724 44604 3780
rect 44660 3724 50540 3780
rect 50596 3724 51436 3780
rect 51492 3724 51502 3780
rect 53004 3724 54236 3780
rect 54292 3724 54302 3780
rect 58146 3724 58156 3780
rect 58212 3724 59332 3780
rect 61394 3724 61404 3780
rect 61460 3724 65548 3780
rect 65604 3724 65614 3780
rect 65772 3724 67452 3780
rect 67508 3724 67518 3780
rect 69458 3724 69468 3780
rect 69524 3724 75068 3780
rect 75124 3724 75134 3780
rect 19628 3668 19684 3724
rect 26012 3668 26068 3724
rect 29036 3668 29092 3724
rect 5730 3612 5740 3668
rect 5796 3612 5964 3668
rect 6020 3612 8316 3668
rect 8372 3612 8382 3668
rect 8530 3612 8540 3668
rect 8596 3612 10388 3668
rect 10546 3612 10556 3668
rect 10612 3612 17500 3668
rect 17556 3612 17566 3668
rect 18274 3612 18284 3668
rect 18340 3612 19068 3668
rect 19124 3612 19134 3668
rect 19282 3612 19292 3668
rect 19348 3612 19386 3668
rect 19618 3612 19628 3668
rect 19684 3612 19694 3668
rect 20402 3612 20412 3668
rect 20468 3612 21756 3668
rect 21812 3612 25788 3668
rect 25844 3612 25854 3668
rect 26012 3612 28476 3668
rect 28532 3612 28542 3668
rect 29036 3612 31164 3668
rect 31220 3612 31230 3668
rect 36082 3612 36092 3668
rect 36148 3612 36876 3668
rect 36932 3612 36942 3668
rect 38612 3612 38668 3724
rect 42812 3668 42868 3724
rect 53004 3668 53060 3724
rect 59276 3668 59332 3724
rect 38724 3612 38734 3668
rect 40338 3612 40348 3668
rect 40404 3612 41356 3668
rect 41412 3612 41422 3668
rect 41794 3612 41804 3668
rect 41860 3612 42868 3668
rect 43922 3612 43932 3668
rect 43988 3612 49868 3668
rect 49924 3612 49934 3668
rect 51314 3612 51324 3668
rect 51380 3612 53004 3668
rect 53060 3612 53070 3668
rect 53330 3612 53340 3668
rect 53396 3612 56028 3668
rect 56084 3612 56094 3668
rect 56578 3612 56588 3668
rect 56644 3612 58044 3668
rect 58100 3612 58110 3668
rect 59042 3612 59052 3668
rect 59108 3612 59118 3668
rect 59276 3612 63868 3668
rect 63924 3612 63934 3668
rect 64530 3612 64540 3668
rect 64596 3612 65660 3668
rect 65716 3612 65726 3668
rect 71250 3612 71260 3668
rect 71316 3612 71326 3668
rect 10332 3556 10388 3612
rect 59052 3556 59108 3612
rect 7158 3500 7196 3556
rect 7252 3500 7262 3556
rect 10332 3500 12348 3556
rect 12404 3500 12414 3556
rect 14130 3500 14140 3556
rect 14196 3500 15148 3556
rect 15204 3500 15214 3556
rect 15362 3500 15372 3556
rect 15428 3500 18396 3556
rect 18452 3500 18462 3556
rect 19506 3500 19516 3556
rect 19572 3500 22988 3556
rect 23044 3500 23054 3556
rect 24546 3500 24556 3556
rect 24612 3500 25116 3556
rect 25172 3500 25182 3556
rect 29922 3500 29932 3556
rect 29988 3500 37212 3556
rect 37268 3500 37278 3556
rect 40226 3500 40236 3556
rect 40292 3500 42476 3556
rect 42532 3500 45276 3556
rect 45332 3500 45342 3556
rect 50082 3500 50092 3556
rect 50148 3500 51660 3556
rect 51716 3500 51726 3556
rect 51986 3500 51996 3556
rect 52052 3500 53228 3556
rect 53284 3500 53676 3556
rect 53732 3500 53742 3556
rect 55346 3500 55356 3556
rect 55412 3500 59108 3556
rect 59490 3500 59500 3556
rect 59556 3500 60956 3556
rect 61012 3500 61852 3556
rect 61908 3500 61918 3556
rect 65426 3500 65436 3556
rect 65492 3500 68908 3556
rect 68964 3500 68974 3556
rect 0 3444 800 3472
rect 71260 3444 71316 3612
rect 75282 3500 75292 3556
rect 75348 3500 77868 3556
rect 77924 3500 77934 3556
rect 0 3388 1708 3444
rect 1764 3388 3164 3444
rect 3220 3388 3230 3444
rect 4722 3388 4732 3444
rect 4788 3388 6300 3444
rect 6356 3388 6366 3444
rect 8082 3388 8092 3444
rect 8148 3388 10892 3444
rect 10948 3388 10958 3444
rect 11218 3388 11228 3444
rect 11284 3388 11900 3444
rect 11956 3388 11966 3444
rect 14690 3388 14700 3444
rect 14756 3388 17724 3444
rect 17780 3388 17790 3444
rect 17938 3388 17948 3444
rect 18004 3388 21084 3444
rect 21140 3388 21150 3444
rect 23538 3388 23548 3444
rect 23604 3388 26908 3444
rect 26964 3388 26974 3444
rect 28578 3388 28588 3444
rect 28644 3388 34972 3444
rect 35028 3388 35038 3444
rect 35298 3388 35308 3444
rect 35364 3388 42252 3444
rect 42308 3388 42318 3444
rect 43026 3388 43036 3444
rect 43092 3388 45164 3444
rect 45220 3388 45230 3444
rect 47170 3388 47180 3444
rect 47236 3388 49644 3444
rect 49700 3388 49710 3444
rect 50866 3388 50876 3444
rect 50932 3388 52332 3444
rect 52388 3388 52398 3444
rect 57362 3388 57372 3444
rect 57428 3388 59724 3444
rect 59780 3388 59790 3444
rect 64754 3388 64764 3444
rect 64820 3388 71316 3444
rect 71474 3388 71484 3444
rect 71540 3388 76188 3444
rect 76244 3388 76254 3444
rect 0 3360 800 3388
rect 11890 3276 11900 3332
rect 11956 3276 15484 3332
rect 15540 3276 15550 3332
rect 20066 3276 20076 3332
rect 20132 3276 21028 3332
rect 23650 3276 23660 3332
rect 23716 3276 24220 3332
rect 24276 3276 24286 3332
rect 24994 3276 25004 3332
rect 25060 3276 29260 3332
rect 29316 3276 29326 3332
rect 31602 3276 31612 3332
rect 31668 3276 40460 3332
rect 40516 3276 40526 3332
rect 49186 3276 49196 3332
rect 49252 3276 50204 3332
rect 50260 3276 50270 3332
rect 50428 3276 51212 3332
rect 51268 3276 51278 3332
rect 8754 3164 8764 3220
rect 8820 3164 15148 3220
rect 15204 3164 15214 3220
rect 19826 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20110 3164
rect 20972 2996 21028 3276
rect 50428 3220 50484 3276
rect 21970 3164 21980 3220
rect 22036 3164 26684 3220
rect 26740 3164 26750 3220
rect 30146 3164 30156 3220
rect 30212 3164 50484 3220
rect 50546 3108 50556 3164
rect 50612 3108 50660 3164
rect 50716 3108 50764 3164
rect 50820 3108 50830 3164
rect 21186 3052 21196 3108
rect 21252 3052 29932 3108
rect 29988 3052 29998 3108
rect 79200 2996 80000 3024
rect 20972 2940 27468 2996
rect 27524 2940 27534 2996
rect 28914 2940 28924 2996
rect 28980 2940 37324 2996
rect 37380 2940 37390 2996
rect 74498 2940 74508 2996
rect 74564 2940 80000 2996
rect 79200 2912 80000 2940
rect 27794 2828 27804 2884
rect 27860 2828 36988 2884
rect 37044 2828 37054 2884
rect 24210 2716 24220 2772
rect 24276 2716 30492 2772
rect 30548 2716 30558 2772
rect 26674 2604 26684 2660
rect 26740 2604 32508 2660
rect 32564 2604 32574 2660
rect 21522 2492 21532 2548
rect 21588 2492 28588 2548
rect 28644 2492 28654 2548
rect 40562 2492 40572 2548
rect 40628 2492 49196 2548
rect 49252 2492 49262 2548
rect 11330 2380 11340 2436
rect 11396 2380 28812 2436
rect 28868 2380 28878 2436
rect 0 2324 800 2352
rect 0 2268 2380 2324
rect 2436 2268 2446 2324
rect 14354 2268 14364 2324
rect 14420 2268 23884 2324
rect 23940 2268 23950 2324
rect 29250 2268 29260 2324
rect 29316 2268 36540 2324
rect 36596 2268 36606 2324
rect 0 2240 800 2268
rect 24098 2156 24108 2212
rect 24164 2156 36876 2212
rect 36932 2156 36942 2212
rect 25330 2044 25340 2100
rect 25396 2044 35980 2100
rect 36036 2044 36046 2100
rect 79200 1876 80000 1904
rect 27570 1820 27580 1876
rect 27636 1820 34524 1876
rect 34580 1820 34590 1876
rect 75506 1820 75516 1876
rect 75572 1820 80000 1876
rect 79200 1792 80000 1820
rect 19618 1708 19628 1764
rect 19684 1708 23772 1764
rect 23828 1708 23838 1764
rect 26908 1708 29428 1764
rect 26908 1652 26964 1708
rect 29372 1652 29428 1708
rect 25890 1596 25900 1652
rect 25956 1596 26964 1652
rect 27020 1596 29148 1652
rect 29204 1596 29214 1652
rect 29372 1596 32172 1652
rect 32228 1596 32238 1652
rect 27020 1540 27076 1596
rect 21298 1484 21308 1540
rect 21364 1484 27076 1540
rect 22642 1372 22652 1428
rect 22708 1372 33740 1428
rect 33796 1372 33806 1428
rect 18834 1260 18844 1316
rect 18900 1260 27244 1316
rect 27300 1260 27310 1316
rect 74274 924 74284 980
rect 74340 924 74350 980
rect 74284 756 74340 924
rect 79200 756 80000 784
rect 74284 700 80000 756
rect 79200 672 80000 700
<< via3 >>
rect 19836 76804 19892 76860
rect 19940 76804 19996 76860
rect 20044 76804 20100 76860
rect 50556 76804 50612 76860
rect 50660 76804 50716 76860
rect 50764 76804 50820 76860
rect 73164 76524 73220 76580
rect 47404 76300 47460 76356
rect 4476 76020 4532 76076
rect 4580 76020 4636 76076
rect 4684 76020 4740 76076
rect 35196 76020 35252 76076
rect 35300 76020 35356 76076
rect 35404 76020 35460 76076
rect 65916 76020 65972 76076
rect 66020 76020 66076 76076
rect 66124 76020 66180 76076
rect 47180 75628 47236 75684
rect 76524 75628 76580 75684
rect 19836 75236 19892 75292
rect 19940 75236 19996 75292
rect 20044 75236 20100 75292
rect 50556 75236 50612 75292
rect 50660 75236 50716 75292
rect 50764 75236 50820 75292
rect 4476 74452 4532 74508
rect 4580 74452 4636 74508
rect 4684 74452 4740 74508
rect 35196 74452 35252 74508
rect 35300 74452 35356 74508
rect 35404 74452 35460 74508
rect 65916 74452 65972 74508
rect 66020 74452 66076 74508
rect 66124 74452 66180 74508
rect 19836 73668 19892 73724
rect 19940 73668 19996 73724
rect 20044 73668 20100 73724
rect 50556 73668 50612 73724
rect 50660 73668 50716 73724
rect 50764 73668 50820 73724
rect 4476 72884 4532 72940
rect 4580 72884 4636 72940
rect 4684 72884 4740 72940
rect 35196 72884 35252 72940
rect 35300 72884 35356 72940
rect 35404 72884 35460 72940
rect 65916 72884 65972 72940
rect 66020 72884 66076 72940
rect 66124 72884 66180 72940
rect 19836 72100 19892 72156
rect 19940 72100 19996 72156
rect 20044 72100 20100 72156
rect 50556 72100 50612 72156
rect 50660 72100 50716 72156
rect 50764 72100 50820 72156
rect 4476 71316 4532 71372
rect 4580 71316 4636 71372
rect 4684 71316 4740 71372
rect 35196 71316 35252 71372
rect 35300 71316 35356 71372
rect 35404 71316 35460 71372
rect 65916 71316 65972 71372
rect 66020 71316 66076 71372
rect 66124 71316 66180 71372
rect 19836 70532 19892 70588
rect 19940 70532 19996 70588
rect 20044 70532 20100 70588
rect 50556 70532 50612 70588
rect 50660 70532 50716 70588
rect 50764 70532 50820 70588
rect 4476 69748 4532 69804
rect 4580 69748 4636 69804
rect 4684 69748 4740 69804
rect 35196 69748 35252 69804
rect 35300 69748 35356 69804
rect 35404 69748 35460 69804
rect 65916 69748 65972 69804
rect 66020 69748 66076 69804
rect 66124 69748 66180 69804
rect 76748 69132 76804 69188
rect 19836 68964 19892 69020
rect 19940 68964 19996 69020
rect 20044 68964 20100 69020
rect 50556 68964 50612 69020
rect 50660 68964 50716 69020
rect 50764 68964 50820 69020
rect 76860 68460 76916 68516
rect 4476 68180 4532 68236
rect 4580 68180 4636 68236
rect 4684 68180 4740 68236
rect 35196 68180 35252 68236
rect 35300 68180 35356 68236
rect 35404 68180 35460 68236
rect 65916 68180 65972 68236
rect 66020 68180 66076 68236
rect 66124 68180 66180 68236
rect 19836 67396 19892 67452
rect 19940 67396 19996 67452
rect 20044 67396 20100 67452
rect 50556 67396 50612 67452
rect 50660 67396 50716 67452
rect 50764 67396 50820 67452
rect 4476 66612 4532 66668
rect 4580 66612 4636 66668
rect 4684 66612 4740 66668
rect 35196 66612 35252 66668
rect 35300 66612 35356 66668
rect 35404 66612 35460 66668
rect 65916 66612 65972 66668
rect 66020 66612 66076 66668
rect 66124 66612 66180 66668
rect 76636 65996 76692 66052
rect 19836 65828 19892 65884
rect 19940 65828 19996 65884
rect 20044 65828 20100 65884
rect 50556 65828 50612 65884
rect 50660 65828 50716 65884
rect 50764 65828 50820 65884
rect 4476 65044 4532 65100
rect 4580 65044 4636 65100
rect 4684 65044 4740 65100
rect 35196 65044 35252 65100
rect 35300 65044 35356 65100
rect 35404 65044 35460 65100
rect 65916 65044 65972 65100
rect 66020 65044 66076 65100
rect 66124 65044 66180 65100
rect 77084 64652 77140 64708
rect 19836 64260 19892 64316
rect 19940 64260 19996 64316
rect 20044 64260 20100 64316
rect 50556 64260 50612 64316
rect 50660 64260 50716 64316
rect 50764 64260 50820 64316
rect 76412 63980 76468 64036
rect 4476 63476 4532 63532
rect 4580 63476 4636 63532
rect 4684 63476 4740 63532
rect 35196 63476 35252 63532
rect 35300 63476 35356 63532
rect 35404 63476 35460 63532
rect 65916 63476 65972 63532
rect 66020 63476 66076 63532
rect 66124 63476 66180 63532
rect 19836 62692 19892 62748
rect 19940 62692 19996 62748
rect 20044 62692 20100 62748
rect 50556 62692 50612 62748
rect 50660 62692 50716 62748
rect 50764 62692 50820 62748
rect 76188 62188 76244 62244
rect 4476 61908 4532 61964
rect 4580 61908 4636 61964
rect 4684 61908 4740 61964
rect 35196 61908 35252 61964
rect 35300 61908 35356 61964
rect 35404 61908 35460 61964
rect 65916 61908 65972 61964
rect 66020 61908 66076 61964
rect 66124 61908 66180 61964
rect 75404 61516 75460 61572
rect 19836 61124 19892 61180
rect 19940 61124 19996 61180
rect 20044 61124 20100 61180
rect 50556 61124 50612 61180
rect 50660 61124 50716 61180
rect 50764 61124 50820 61180
rect 76300 60844 76356 60900
rect 4476 60340 4532 60396
rect 4580 60340 4636 60396
rect 4684 60340 4740 60396
rect 35196 60340 35252 60396
rect 35300 60340 35356 60396
rect 35404 60340 35460 60396
rect 65916 60340 65972 60396
rect 66020 60340 66076 60396
rect 66124 60340 66180 60396
rect 19836 59556 19892 59612
rect 19940 59556 19996 59612
rect 20044 59556 20100 59612
rect 50556 59556 50612 59612
rect 50660 59556 50716 59612
rect 50764 59556 50820 59612
rect 74956 59052 75012 59108
rect 4476 58772 4532 58828
rect 4580 58772 4636 58828
rect 4684 58772 4740 58828
rect 35196 58772 35252 58828
rect 35300 58772 35356 58828
rect 35404 58772 35460 58828
rect 65916 58772 65972 58828
rect 66020 58772 66076 58828
rect 66124 58772 66180 58828
rect 19836 57988 19892 58044
rect 19940 57988 19996 58044
rect 20044 57988 20100 58044
rect 50556 57988 50612 58044
rect 50660 57988 50716 58044
rect 50764 57988 50820 58044
rect 4476 57204 4532 57260
rect 4580 57204 4636 57260
rect 4684 57204 4740 57260
rect 35196 57204 35252 57260
rect 35300 57204 35356 57260
rect 35404 57204 35460 57260
rect 65916 57204 65972 57260
rect 66020 57204 66076 57260
rect 66124 57204 66180 57260
rect 19836 56420 19892 56476
rect 19940 56420 19996 56476
rect 20044 56420 20100 56476
rect 50556 56420 50612 56476
rect 50660 56420 50716 56476
rect 50764 56420 50820 56476
rect 4476 55636 4532 55692
rect 4580 55636 4636 55692
rect 4684 55636 4740 55692
rect 35196 55636 35252 55692
rect 35300 55636 35356 55692
rect 35404 55636 35460 55692
rect 65916 55636 65972 55692
rect 66020 55636 66076 55692
rect 66124 55636 66180 55692
rect 19836 54852 19892 54908
rect 19940 54852 19996 54908
rect 20044 54852 20100 54908
rect 50556 54852 50612 54908
rect 50660 54852 50716 54908
rect 50764 54852 50820 54908
rect 4476 54068 4532 54124
rect 4580 54068 4636 54124
rect 4684 54068 4740 54124
rect 35196 54068 35252 54124
rect 35300 54068 35356 54124
rect 35404 54068 35460 54124
rect 65916 54068 65972 54124
rect 66020 54068 66076 54124
rect 66124 54068 66180 54124
rect 72604 54012 72660 54068
rect 19836 53284 19892 53340
rect 19940 53284 19996 53340
rect 20044 53284 20100 53340
rect 50556 53284 50612 53340
rect 50660 53284 50716 53340
rect 50764 53284 50820 53340
rect 4476 52500 4532 52556
rect 4580 52500 4636 52556
rect 4684 52500 4740 52556
rect 35196 52500 35252 52556
rect 35300 52500 35356 52556
rect 35404 52500 35460 52556
rect 65916 52500 65972 52556
rect 66020 52500 66076 52556
rect 66124 52500 66180 52556
rect 19836 51716 19892 51772
rect 19940 51716 19996 51772
rect 20044 51716 20100 51772
rect 50556 51716 50612 51772
rect 50660 51716 50716 51772
rect 50764 51716 50820 51772
rect 4476 50932 4532 50988
rect 4580 50932 4636 50988
rect 4684 50932 4740 50988
rect 35196 50932 35252 50988
rect 35300 50932 35356 50988
rect 35404 50932 35460 50988
rect 65916 50932 65972 50988
rect 66020 50932 66076 50988
rect 66124 50932 66180 50988
rect 19836 50148 19892 50204
rect 19940 50148 19996 50204
rect 20044 50148 20100 50204
rect 50556 50148 50612 50204
rect 50660 50148 50716 50204
rect 50764 50148 50820 50204
rect 4476 49364 4532 49420
rect 4580 49364 4636 49420
rect 4684 49364 4740 49420
rect 35196 49364 35252 49420
rect 35300 49364 35356 49420
rect 35404 49364 35460 49420
rect 65916 49364 65972 49420
rect 66020 49364 66076 49420
rect 66124 49364 66180 49420
rect 19836 48580 19892 48636
rect 19940 48580 19996 48636
rect 20044 48580 20100 48636
rect 50556 48580 50612 48636
rect 50660 48580 50716 48636
rect 50764 48580 50820 48636
rect 4476 47796 4532 47852
rect 4580 47796 4636 47852
rect 4684 47796 4740 47852
rect 35196 47796 35252 47852
rect 35300 47796 35356 47852
rect 35404 47796 35460 47852
rect 65916 47796 65972 47852
rect 66020 47796 66076 47852
rect 66124 47796 66180 47852
rect 19836 47012 19892 47068
rect 19940 47012 19996 47068
rect 20044 47012 20100 47068
rect 50556 47012 50612 47068
rect 50660 47012 50716 47068
rect 50764 47012 50820 47068
rect 74732 46956 74788 47012
rect 74060 46844 74116 46900
rect 4476 46228 4532 46284
rect 4580 46228 4636 46284
rect 4684 46228 4740 46284
rect 35196 46228 35252 46284
rect 35300 46228 35356 46284
rect 35404 46228 35460 46284
rect 65916 46228 65972 46284
rect 66020 46228 66076 46284
rect 66124 46228 66180 46284
rect 19836 45444 19892 45500
rect 19940 45444 19996 45500
rect 20044 45444 20100 45500
rect 50556 45444 50612 45500
rect 50660 45444 50716 45500
rect 50764 45444 50820 45500
rect 4476 44660 4532 44716
rect 4580 44660 4636 44716
rect 4684 44660 4740 44716
rect 35196 44660 35252 44716
rect 35300 44660 35356 44716
rect 35404 44660 35460 44716
rect 65916 44660 65972 44716
rect 66020 44660 66076 44716
rect 66124 44660 66180 44716
rect 19836 43876 19892 43932
rect 19940 43876 19996 43932
rect 20044 43876 20100 43932
rect 50556 43876 50612 43932
rect 50660 43876 50716 43932
rect 50764 43876 50820 43932
rect 4476 43092 4532 43148
rect 4580 43092 4636 43148
rect 4684 43092 4740 43148
rect 35196 43092 35252 43148
rect 35300 43092 35356 43148
rect 35404 43092 35460 43148
rect 65916 43092 65972 43148
rect 66020 43092 66076 43148
rect 66124 43092 66180 43148
rect 77644 42588 77700 42644
rect 19836 42308 19892 42364
rect 19940 42308 19996 42364
rect 20044 42308 20100 42364
rect 50556 42308 50612 42364
rect 50660 42308 50716 42364
rect 50764 42308 50820 42364
rect 74844 41804 74900 41860
rect 4476 41524 4532 41580
rect 4580 41524 4636 41580
rect 4684 41524 4740 41580
rect 35196 41524 35252 41580
rect 35300 41524 35356 41580
rect 35404 41524 35460 41580
rect 65916 41524 65972 41580
rect 66020 41524 66076 41580
rect 66124 41524 66180 41580
rect 72044 41468 72100 41524
rect 72044 40908 72100 40964
rect 77644 40908 77700 40964
rect 72492 40796 72548 40852
rect 19836 40740 19892 40796
rect 19940 40740 19996 40796
rect 20044 40740 20100 40796
rect 50556 40740 50612 40796
rect 50660 40740 50716 40796
rect 50764 40740 50820 40796
rect 74844 40348 74900 40404
rect 4476 39956 4532 40012
rect 4580 39956 4636 40012
rect 4684 39956 4740 40012
rect 35196 39956 35252 40012
rect 35300 39956 35356 40012
rect 35404 39956 35460 40012
rect 65916 39956 65972 40012
rect 66020 39956 66076 40012
rect 66124 39956 66180 40012
rect 19836 39172 19892 39228
rect 19940 39172 19996 39228
rect 20044 39172 20100 39228
rect 50556 39172 50612 39228
rect 50660 39172 50716 39228
rect 50764 39172 50820 39228
rect 69468 39004 69524 39060
rect 74508 39004 74564 39060
rect 74284 38892 74340 38948
rect 76972 38780 77028 38836
rect 4476 38388 4532 38444
rect 4580 38388 4636 38444
rect 4684 38388 4740 38444
rect 35196 38388 35252 38444
rect 35300 38388 35356 38444
rect 35404 38388 35460 38444
rect 65916 38388 65972 38444
rect 66020 38388 66076 38444
rect 66124 38388 66180 38444
rect 69468 38332 69524 38388
rect 75068 38220 75124 38276
rect 73500 37772 73556 37828
rect 74172 37772 74228 37828
rect 77868 37660 77924 37716
rect 19836 37604 19892 37660
rect 19940 37604 19996 37660
rect 20044 37604 20100 37660
rect 50556 37604 50612 37660
rect 50660 37604 50716 37660
rect 50764 37604 50820 37660
rect 74172 37212 74228 37268
rect 76524 37212 76580 37268
rect 74284 36988 74340 37044
rect 76972 36988 77028 37044
rect 72492 36876 72548 36932
rect 4476 36820 4532 36876
rect 4580 36820 4636 36876
rect 4684 36820 4740 36876
rect 35196 36820 35252 36876
rect 35300 36820 35356 36876
rect 35404 36820 35460 36876
rect 65916 36820 65972 36876
rect 66020 36820 66076 36876
rect 66124 36820 66180 36876
rect 73164 36428 73220 36484
rect 19836 36036 19892 36092
rect 19940 36036 19996 36092
rect 20044 36036 20100 36092
rect 50556 36036 50612 36092
rect 50660 36036 50716 36092
rect 50764 36036 50820 36092
rect 75068 35980 75124 36036
rect 74620 35532 74676 35588
rect 74508 35420 74564 35476
rect 4476 35252 4532 35308
rect 4580 35252 4636 35308
rect 4684 35252 4740 35308
rect 35196 35252 35252 35308
rect 35300 35252 35356 35308
rect 35404 35252 35460 35308
rect 65916 35252 65972 35308
rect 66020 35252 66076 35308
rect 66124 35252 66180 35308
rect 77868 35084 77924 35140
rect 75740 34972 75796 35028
rect 73276 34636 73332 34692
rect 19836 34468 19892 34524
rect 19940 34468 19996 34524
rect 20044 34468 20100 34524
rect 50556 34468 50612 34524
rect 50660 34468 50716 34524
rect 50764 34468 50820 34524
rect 4476 33684 4532 33740
rect 4580 33684 4636 33740
rect 4684 33684 4740 33740
rect 35196 33684 35252 33740
rect 35300 33684 35356 33740
rect 35404 33684 35460 33740
rect 65916 33684 65972 33740
rect 66020 33684 66076 33740
rect 66124 33684 66180 33740
rect 75068 33628 75124 33684
rect 76748 33404 76804 33460
rect 19836 32900 19892 32956
rect 19940 32900 19996 32956
rect 20044 32900 20100 32956
rect 50556 32900 50612 32956
rect 50660 32900 50716 32956
rect 50764 32900 50820 32956
rect 75068 32284 75124 32340
rect 4476 32116 4532 32172
rect 4580 32116 4636 32172
rect 4684 32116 4740 32172
rect 35196 32116 35252 32172
rect 35300 32116 35356 32172
rect 35404 32116 35460 32172
rect 65916 32116 65972 32172
rect 66020 32116 66076 32172
rect 66124 32116 66180 32172
rect 71148 32060 71204 32116
rect 75740 31836 75796 31892
rect 76860 31724 76916 31780
rect 74732 31388 74788 31444
rect 19836 31332 19892 31388
rect 19940 31332 19996 31388
rect 20044 31332 20100 31388
rect 50556 31332 50612 31388
rect 50660 31332 50716 31388
rect 50764 31332 50820 31388
rect 73500 30940 73556 30996
rect 74732 30940 74788 30996
rect 77084 30828 77140 30884
rect 51212 30716 51268 30772
rect 70924 30716 70980 30772
rect 4476 30548 4532 30604
rect 4580 30548 4636 30604
rect 4684 30548 4740 30604
rect 35196 30548 35252 30604
rect 35300 30548 35356 30604
rect 35404 30548 35460 30604
rect 65916 30548 65972 30604
rect 66020 30548 66076 30604
rect 66124 30548 66180 30604
rect 71372 30156 71428 30212
rect 76636 30156 76692 30212
rect 72716 30044 72772 30100
rect 72604 29932 72660 29988
rect 19836 29764 19892 29820
rect 19940 29764 19996 29820
rect 20044 29764 20100 29820
rect 50556 29764 50612 29820
rect 50660 29764 50716 29820
rect 50764 29764 50820 29820
rect 76412 29708 76468 29764
rect 76412 29484 76468 29540
rect 18060 29372 18116 29428
rect 69580 29372 69636 29428
rect 75628 29260 75684 29316
rect 4476 28980 4532 29036
rect 4580 28980 4636 29036
rect 4684 28980 4740 29036
rect 35196 28980 35252 29036
rect 35300 28980 35356 29036
rect 35404 28980 35460 29036
rect 65916 28980 65972 29036
rect 66020 28980 66076 29036
rect 66124 28980 66180 29036
rect 75404 28924 75460 28980
rect 76300 28924 76356 28980
rect 74620 28588 74676 28644
rect 72716 28476 72772 28532
rect 74956 28252 75012 28308
rect 19836 28196 19892 28252
rect 19940 28196 19996 28252
rect 20044 28196 20100 28252
rect 50556 28196 50612 28252
rect 50660 28196 50716 28252
rect 50764 28196 50820 28252
rect 74060 27916 74116 27972
rect 74956 27916 75012 27972
rect 76188 27916 76244 27972
rect 76188 27580 76244 27636
rect 4476 27412 4532 27468
rect 4580 27412 4636 27468
rect 4684 27412 4740 27468
rect 35196 27412 35252 27468
rect 35300 27412 35356 27468
rect 35404 27412 35460 27468
rect 65916 27412 65972 27468
rect 66020 27412 66076 27468
rect 66124 27412 66180 27468
rect 75516 27356 75572 27412
rect 73164 27132 73220 27188
rect 72716 26908 72772 26964
rect 74732 26908 74788 26964
rect 56700 26796 56756 26852
rect 75516 26796 75572 26852
rect 46060 26684 46116 26740
rect 51212 26684 51268 26740
rect 19836 26628 19892 26684
rect 19940 26628 19996 26684
rect 20044 26628 20100 26684
rect 50556 26628 50612 26684
rect 50660 26628 50716 26684
rect 50764 26628 50820 26684
rect 73052 26572 73108 26628
rect 56700 26460 56756 26516
rect 70924 26460 70980 26516
rect 69580 26348 69636 26404
rect 75628 26012 75684 26068
rect 4476 25844 4532 25900
rect 4580 25844 4636 25900
rect 4684 25844 4740 25900
rect 35196 25844 35252 25900
rect 35300 25844 35356 25900
rect 35404 25844 35460 25900
rect 65916 25844 65972 25900
rect 66020 25844 66076 25900
rect 66124 25844 66180 25900
rect 71148 25116 71204 25172
rect 19836 25060 19892 25116
rect 19940 25060 19996 25116
rect 20044 25060 20100 25116
rect 50556 25060 50612 25116
rect 50660 25060 50716 25116
rect 50764 25060 50820 25116
rect 18396 24556 18452 24612
rect 4476 24276 4532 24332
rect 4580 24276 4636 24332
rect 4684 24276 4740 24332
rect 43596 24444 43652 24500
rect 71372 24332 71428 24388
rect 35196 24276 35252 24332
rect 35300 24276 35356 24332
rect 35404 24276 35460 24332
rect 65916 24276 65972 24332
rect 66020 24276 66076 24332
rect 66124 24276 66180 24332
rect 18060 23884 18116 23940
rect 73276 23884 73332 23940
rect 18396 23660 18452 23716
rect 19836 23492 19892 23548
rect 19940 23492 19996 23548
rect 20044 23492 20100 23548
rect 40460 23436 40516 23492
rect 50556 23492 50612 23548
rect 50660 23492 50716 23548
rect 50764 23492 50820 23548
rect 40908 23436 40964 23492
rect 50092 23436 50148 23492
rect 46060 23100 46116 23156
rect 43596 22764 43652 22820
rect 4476 22708 4532 22764
rect 4580 22708 4636 22764
rect 4684 22708 4740 22764
rect 35196 22708 35252 22764
rect 35300 22708 35356 22764
rect 35404 22708 35460 22764
rect 65916 22708 65972 22764
rect 66020 22708 66076 22764
rect 66124 22708 66180 22764
rect 76748 22428 76804 22484
rect 47628 22316 47684 22372
rect 75740 22316 75796 22372
rect 77084 22316 77140 22372
rect 47628 21980 47684 22036
rect 19836 21924 19892 21980
rect 19940 21924 19996 21980
rect 20044 21924 20100 21980
rect 50556 21924 50612 21980
rect 50660 21924 50716 21980
rect 50764 21924 50820 21980
rect 74956 21868 75012 21924
rect 34524 21420 34580 21476
rect 4476 21140 4532 21196
rect 4580 21140 4636 21196
rect 4684 21140 4740 21196
rect 35196 21140 35252 21196
rect 35300 21140 35356 21196
rect 35404 21140 35460 21196
rect 65916 21140 65972 21196
rect 66020 21140 66076 21196
rect 66124 21140 66180 21196
rect 47180 20748 47236 20804
rect 19836 20356 19892 20412
rect 19940 20356 19996 20412
rect 20044 20356 20100 20412
rect 50556 20356 50612 20412
rect 50660 20356 50716 20412
rect 50764 20356 50820 20412
rect 34524 19964 34580 20020
rect 50092 19964 50148 20020
rect 4476 19572 4532 19628
rect 4580 19572 4636 19628
rect 4684 19572 4740 19628
rect 35196 19572 35252 19628
rect 35300 19572 35356 19628
rect 35404 19572 35460 19628
rect 65916 19572 65972 19628
rect 66020 19572 66076 19628
rect 66124 19572 66180 19628
rect 28700 19180 28756 19236
rect 19836 18788 19892 18844
rect 19940 18788 19996 18844
rect 20044 18788 20100 18844
rect 50556 18788 50612 18844
rect 50660 18788 50716 18844
rect 50764 18788 50820 18844
rect 28700 18508 28756 18564
rect 4476 18004 4532 18060
rect 4580 18004 4636 18060
rect 4684 18004 4740 18060
rect 35196 18004 35252 18060
rect 35300 18004 35356 18060
rect 35404 18004 35460 18060
rect 65916 18004 65972 18060
rect 66020 18004 66076 18060
rect 66124 18004 66180 18060
rect 19836 17220 19892 17276
rect 19940 17220 19996 17276
rect 20044 17220 20100 17276
rect 50556 17220 50612 17276
rect 50660 17220 50716 17276
rect 50764 17220 50820 17276
rect 47292 16828 47348 16884
rect 4476 16436 4532 16492
rect 4580 16436 4636 16492
rect 4684 16436 4740 16492
rect 35196 16436 35252 16492
rect 35300 16436 35356 16492
rect 35404 16436 35460 16492
rect 65916 16436 65972 16492
rect 66020 16436 66076 16492
rect 66124 16436 66180 16492
rect 19836 15652 19892 15708
rect 19940 15652 19996 15708
rect 20044 15652 20100 15708
rect 50556 15652 50612 15708
rect 50660 15652 50716 15708
rect 50764 15652 50820 15708
rect 77084 15148 77140 15204
rect 4476 14868 4532 14924
rect 4580 14868 4636 14924
rect 4684 14868 4740 14924
rect 35196 14868 35252 14924
rect 35300 14868 35356 14924
rect 35404 14868 35460 14924
rect 65916 14868 65972 14924
rect 66020 14868 66076 14924
rect 66124 14868 66180 14924
rect 19836 14084 19892 14140
rect 19940 14084 19996 14140
rect 20044 14084 20100 14140
rect 50556 14084 50612 14140
rect 50660 14084 50716 14140
rect 50764 14084 50820 14140
rect 76748 13916 76804 13972
rect 4476 13300 4532 13356
rect 4580 13300 4636 13356
rect 4684 13300 4740 13356
rect 35196 13300 35252 13356
rect 35300 13300 35356 13356
rect 35404 13300 35460 13356
rect 65916 13300 65972 13356
rect 66020 13300 66076 13356
rect 66124 13300 66180 13356
rect 75740 13020 75796 13076
rect 19836 12516 19892 12572
rect 19940 12516 19996 12572
rect 20044 12516 20100 12572
rect 50556 12516 50612 12572
rect 50660 12516 50716 12572
rect 50764 12516 50820 12572
rect 4476 11732 4532 11788
rect 4580 11732 4636 11788
rect 4684 11732 4740 11788
rect 35196 11732 35252 11788
rect 35300 11732 35356 11788
rect 35404 11732 35460 11788
rect 65916 11732 65972 11788
rect 66020 11732 66076 11788
rect 66124 11732 66180 11788
rect 44492 11340 44548 11396
rect 19836 10948 19892 11004
rect 19940 10948 19996 11004
rect 20044 10948 20100 11004
rect 50556 10948 50612 11004
rect 50660 10948 50716 11004
rect 50764 10948 50820 11004
rect 17836 10892 17892 10948
rect 44492 10668 44548 10724
rect 4476 10164 4532 10220
rect 4580 10164 4636 10220
rect 4684 10164 4740 10220
rect 35196 10164 35252 10220
rect 35300 10164 35356 10220
rect 35404 10164 35460 10220
rect 65916 10164 65972 10220
rect 66020 10164 66076 10220
rect 66124 10164 66180 10220
rect 19836 9380 19892 9436
rect 19940 9380 19996 9436
rect 20044 9380 20100 9436
rect 50556 9380 50612 9436
rect 50660 9380 50716 9436
rect 50764 9380 50820 9436
rect 4476 8596 4532 8652
rect 4580 8596 4636 8652
rect 4684 8596 4740 8652
rect 35196 8596 35252 8652
rect 35300 8596 35356 8652
rect 35404 8596 35460 8652
rect 65916 8596 65972 8652
rect 66020 8596 66076 8652
rect 66124 8596 66180 8652
rect 19628 8316 19684 8372
rect 20188 8316 20244 8372
rect 14364 7868 14420 7924
rect 19836 7812 19892 7868
rect 19940 7812 19996 7868
rect 20044 7812 20100 7868
rect 17836 7756 17892 7812
rect 50556 7812 50612 7868
rect 50660 7812 50716 7868
rect 50764 7812 50820 7868
rect 19628 7420 19684 7476
rect 20188 7420 20244 7476
rect 4476 7028 4532 7084
rect 4580 7028 4636 7084
rect 4684 7028 4740 7084
rect 35196 7028 35252 7084
rect 35300 7028 35356 7084
rect 35404 7028 35460 7084
rect 65916 7028 65972 7084
rect 66020 7028 66076 7084
rect 66124 7028 66180 7084
rect 23212 6972 23268 7028
rect 17164 6636 17220 6692
rect 30156 6524 30212 6580
rect 14700 6412 14756 6468
rect 21980 6300 22036 6356
rect 19836 6244 19892 6300
rect 19940 6244 19996 6300
rect 20044 6244 20100 6300
rect 50556 6244 50612 6300
rect 50660 6244 50716 6300
rect 50764 6244 50820 6300
rect 17164 5964 17220 6020
rect 4476 5460 4532 5516
rect 4580 5460 4636 5516
rect 4684 5460 4740 5516
rect 35196 5460 35252 5516
rect 35300 5460 35356 5516
rect 35404 5460 35460 5516
rect 65916 5460 65972 5516
rect 66020 5460 66076 5516
rect 66124 5460 66180 5516
rect 22204 5292 22260 5348
rect 14364 5180 14420 5236
rect 14700 5068 14756 5124
rect 20412 4956 20468 5012
rect 23212 4844 23268 4900
rect 15148 4732 15204 4788
rect 19292 4732 19348 4788
rect 19836 4676 19892 4732
rect 19940 4676 19996 4732
rect 20044 4676 20100 4732
rect 50556 4676 50612 4732
rect 50660 4676 50716 4732
rect 50764 4676 50820 4732
rect 7196 4620 7252 4676
rect 20636 4396 20692 4452
rect 20300 4284 20356 4340
rect 15148 4172 15204 4228
rect 22204 4172 22260 4228
rect 4476 3892 4532 3948
rect 4580 3892 4636 3948
rect 4684 3892 4740 3948
rect 35196 3892 35252 3948
rect 35300 3892 35356 3948
rect 35404 3892 35460 3948
rect 65916 3892 65972 3948
rect 66020 3892 66076 3948
rect 66124 3892 66180 3948
rect 20300 3724 20356 3780
rect 20636 3724 20692 3780
rect 19292 3612 19348 3668
rect 20412 3612 20468 3668
rect 7196 3500 7252 3556
rect 15148 3500 15204 3556
rect 19836 3108 19892 3164
rect 19940 3108 19996 3164
rect 20044 3108 20100 3164
rect 21980 3164 22036 3220
rect 30156 3164 30212 3220
rect 50556 3108 50612 3164
rect 50660 3108 50716 3164
rect 50764 3108 50820 3164
<< metal4 >>
rect 4448 76076 4768 76892
rect 4448 76020 4476 76076
rect 4532 76020 4580 76076
rect 4636 76020 4684 76076
rect 4740 76020 4768 76076
rect 4448 74508 4768 76020
rect 4448 74452 4476 74508
rect 4532 74452 4580 74508
rect 4636 74452 4684 74508
rect 4740 74452 4768 74508
rect 4448 72940 4768 74452
rect 4448 72884 4476 72940
rect 4532 72884 4580 72940
rect 4636 72884 4684 72940
rect 4740 72884 4768 72940
rect 4448 71372 4768 72884
rect 4448 71316 4476 71372
rect 4532 71316 4580 71372
rect 4636 71316 4684 71372
rect 4740 71316 4768 71372
rect 4448 69804 4768 71316
rect 4448 69748 4476 69804
rect 4532 69748 4580 69804
rect 4636 69748 4684 69804
rect 4740 69748 4768 69804
rect 4448 68236 4768 69748
rect 4448 68180 4476 68236
rect 4532 68180 4580 68236
rect 4636 68180 4684 68236
rect 4740 68180 4768 68236
rect 4448 66668 4768 68180
rect 4448 66612 4476 66668
rect 4532 66612 4580 66668
rect 4636 66612 4684 66668
rect 4740 66612 4768 66668
rect 4448 65100 4768 66612
rect 4448 65044 4476 65100
rect 4532 65044 4580 65100
rect 4636 65044 4684 65100
rect 4740 65044 4768 65100
rect 4448 63532 4768 65044
rect 4448 63476 4476 63532
rect 4532 63476 4580 63532
rect 4636 63476 4684 63532
rect 4740 63476 4768 63532
rect 4448 61964 4768 63476
rect 4448 61908 4476 61964
rect 4532 61908 4580 61964
rect 4636 61908 4684 61964
rect 4740 61908 4768 61964
rect 4448 60396 4768 61908
rect 4448 60340 4476 60396
rect 4532 60340 4580 60396
rect 4636 60340 4684 60396
rect 4740 60340 4768 60396
rect 4448 58828 4768 60340
rect 4448 58772 4476 58828
rect 4532 58772 4580 58828
rect 4636 58772 4684 58828
rect 4740 58772 4768 58828
rect 4448 57260 4768 58772
rect 4448 57204 4476 57260
rect 4532 57204 4580 57260
rect 4636 57204 4684 57260
rect 4740 57204 4768 57260
rect 4448 55692 4768 57204
rect 4448 55636 4476 55692
rect 4532 55636 4580 55692
rect 4636 55636 4684 55692
rect 4740 55636 4768 55692
rect 4448 54124 4768 55636
rect 4448 54068 4476 54124
rect 4532 54068 4580 54124
rect 4636 54068 4684 54124
rect 4740 54068 4768 54124
rect 4448 52556 4768 54068
rect 4448 52500 4476 52556
rect 4532 52500 4580 52556
rect 4636 52500 4684 52556
rect 4740 52500 4768 52556
rect 4448 50988 4768 52500
rect 4448 50932 4476 50988
rect 4532 50932 4580 50988
rect 4636 50932 4684 50988
rect 4740 50932 4768 50988
rect 4448 49420 4768 50932
rect 4448 49364 4476 49420
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4740 49364 4768 49420
rect 4448 47852 4768 49364
rect 4448 47796 4476 47852
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4740 47796 4768 47852
rect 4448 46284 4768 47796
rect 4448 46228 4476 46284
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4740 46228 4768 46284
rect 4448 44716 4768 46228
rect 4448 44660 4476 44716
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4740 44660 4768 44716
rect 4448 43148 4768 44660
rect 4448 43092 4476 43148
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4740 43092 4768 43148
rect 4448 41580 4768 43092
rect 4448 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4768 41580
rect 4448 40012 4768 41524
rect 4448 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4768 40012
rect 4448 38444 4768 39956
rect 4448 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4768 38444
rect 4448 36876 4768 38388
rect 4448 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4768 36876
rect 4448 35308 4768 36820
rect 4448 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4768 35308
rect 4448 33740 4768 35252
rect 4448 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4768 33740
rect 4448 32172 4768 33684
rect 4448 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4768 32172
rect 4448 30604 4768 32116
rect 4448 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4768 30604
rect 4448 29036 4768 30548
rect 19808 76860 20128 76892
rect 19808 76804 19836 76860
rect 19892 76804 19940 76860
rect 19996 76804 20044 76860
rect 20100 76804 20128 76860
rect 19808 75292 20128 76804
rect 19808 75236 19836 75292
rect 19892 75236 19940 75292
rect 19996 75236 20044 75292
rect 20100 75236 20128 75292
rect 19808 73724 20128 75236
rect 19808 73668 19836 73724
rect 19892 73668 19940 73724
rect 19996 73668 20044 73724
rect 20100 73668 20128 73724
rect 19808 72156 20128 73668
rect 19808 72100 19836 72156
rect 19892 72100 19940 72156
rect 19996 72100 20044 72156
rect 20100 72100 20128 72156
rect 19808 70588 20128 72100
rect 19808 70532 19836 70588
rect 19892 70532 19940 70588
rect 19996 70532 20044 70588
rect 20100 70532 20128 70588
rect 19808 69020 20128 70532
rect 19808 68964 19836 69020
rect 19892 68964 19940 69020
rect 19996 68964 20044 69020
rect 20100 68964 20128 69020
rect 19808 67452 20128 68964
rect 19808 67396 19836 67452
rect 19892 67396 19940 67452
rect 19996 67396 20044 67452
rect 20100 67396 20128 67452
rect 19808 65884 20128 67396
rect 19808 65828 19836 65884
rect 19892 65828 19940 65884
rect 19996 65828 20044 65884
rect 20100 65828 20128 65884
rect 19808 64316 20128 65828
rect 19808 64260 19836 64316
rect 19892 64260 19940 64316
rect 19996 64260 20044 64316
rect 20100 64260 20128 64316
rect 19808 62748 20128 64260
rect 19808 62692 19836 62748
rect 19892 62692 19940 62748
rect 19996 62692 20044 62748
rect 20100 62692 20128 62748
rect 19808 61180 20128 62692
rect 19808 61124 19836 61180
rect 19892 61124 19940 61180
rect 19996 61124 20044 61180
rect 20100 61124 20128 61180
rect 19808 59612 20128 61124
rect 19808 59556 19836 59612
rect 19892 59556 19940 59612
rect 19996 59556 20044 59612
rect 20100 59556 20128 59612
rect 19808 58044 20128 59556
rect 19808 57988 19836 58044
rect 19892 57988 19940 58044
rect 19996 57988 20044 58044
rect 20100 57988 20128 58044
rect 19808 56476 20128 57988
rect 19808 56420 19836 56476
rect 19892 56420 19940 56476
rect 19996 56420 20044 56476
rect 20100 56420 20128 56476
rect 19808 54908 20128 56420
rect 19808 54852 19836 54908
rect 19892 54852 19940 54908
rect 19996 54852 20044 54908
rect 20100 54852 20128 54908
rect 19808 53340 20128 54852
rect 19808 53284 19836 53340
rect 19892 53284 19940 53340
rect 19996 53284 20044 53340
rect 20100 53284 20128 53340
rect 19808 51772 20128 53284
rect 19808 51716 19836 51772
rect 19892 51716 19940 51772
rect 19996 51716 20044 51772
rect 20100 51716 20128 51772
rect 19808 50204 20128 51716
rect 19808 50148 19836 50204
rect 19892 50148 19940 50204
rect 19996 50148 20044 50204
rect 20100 50148 20128 50204
rect 19808 48636 20128 50148
rect 19808 48580 19836 48636
rect 19892 48580 19940 48636
rect 19996 48580 20044 48636
rect 20100 48580 20128 48636
rect 19808 47068 20128 48580
rect 19808 47012 19836 47068
rect 19892 47012 19940 47068
rect 19996 47012 20044 47068
rect 20100 47012 20128 47068
rect 19808 45500 20128 47012
rect 19808 45444 19836 45500
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 20100 45444 20128 45500
rect 19808 43932 20128 45444
rect 19808 43876 19836 43932
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 20100 43876 20128 43932
rect 19808 42364 20128 43876
rect 19808 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20128 42364
rect 19808 40796 20128 42308
rect 19808 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20128 40796
rect 19808 39228 20128 40740
rect 19808 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20128 39228
rect 19808 37660 20128 39172
rect 19808 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20128 37660
rect 19808 36092 20128 37604
rect 19808 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20128 36092
rect 19808 34524 20128 36036
rect 19808 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20128 34524
rect 19808 32956 20128 34468
rect 19808 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20128 32956
rect 19808 31388 20128 32900
rect 19808 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20128 31388
rect 19808 29820 20128 31332
rect 19808 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20128 29820
rect 4448 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4768 29036
rect 4448 27468 4768 28980
rect 4448 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4768 27468
rect 4448 25900 4768 27412
rect 4448 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4768 25900
rect 4448 24332 4768 25844
rect 4448 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4768 24332
rect 4448 22764 4768 24276
rect 18060 29428 18116 29438
rect 18060 23940 18116 29372
rect 19808 28252 20128 29764
rect 19808 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20128 28252
rect 19808 26684 20128 28196
rect 19808 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20128 26684
rect 19808 25116 20128 26628
rect 19808 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20128 25116
rect 18060 23874 18116 23884
rect 18396 24612 18452 24622
rect 18396 23716 18452 24556
rect 18396 23650 18452 23660
rect 4448 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4768 22764
rect 4448 21196 4768 22708
rect 4448 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4768 21196
rect 4448 19628 4768 21140
rect 4448 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4768 19628
rect 4448 18060 4768 19572
rect 4448 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4768 18060
rect 4448 16492 4768 18004
rect 4448 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4768 16492
rect 4448 14924 4768 16436
rect 4448 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4768 14924
rect 4448 13356 4768 14868
rect 4448 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4768 13356
rect 4448 11788 4768 13300
rect 4448 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4768 11788
rect 4448 10220 4768 11732
rect 19808 23548 20128 25060
rect 19808 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20128 23548
rect 19808 21980 20128 23492
rect 19808 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20128 21980
rect 19808 20412 20128 21924
rect 35168 76076 35488 76892
rect 50528 76860 50848 76892
rect 50528 76804 50556 76860
rect 50612 76804 50660 76860
rect 50716 76804 50764 76860
rect 50820 76804 50848 76860
rect 35168 76020 35196 76076
rect 35252 76020 35300 76076
rect 35356 76020 35404 76076
rect 35460 76020 35488 76076
rect 35168 74508 35488 76020
rect 47404 76356 47460 76366
rect 35168 74452 35196 74508
rect 35252 74452 35300 74508
rect 35356 74452 35404 74508
rect 35460 74452 35488 74508
rect 35168 72940 35488 74452
rect 35168 72884 35196 72940
rect 35252 72884 35300 72940
rect 35356 72884 35404 72940
rect 35460 72884 35488 72940
rect 35168 71372 35488 72884
rect 35168 71316 35196 71372
rect 35252 71316 35300 71372
rect 35356 71316 35404 71372
rect 35460 71316 35488 71372
rect 35168 69804 35488 71316
rect 35168 69748 35196 69804
rect 35252 69748 35300 69804
rect 35356 69748 35404 69804
rect 35460 69748 35488 69804
rect 35168 68236 35488 69748
rect 35168 68180 35196 68236
rect 35252 68180 35300 68236
rect 35356 68180 35404 68236
rect 35460 68180 35488 68236
rect 35168 66668 35488 68180
rect 35168 66612 35196 66668
rect 35252 66612 35300 66668
rect 35356 66612 35404 66668
rect 35460 66612 35488 66668
rect 35168 65100 35488 66612
rect 35168 65044 35196 65100
rect 35252 65044 35300 65100
rect 35356 65044 35404 65100
rect 35460 65044 35488 65100
rect 35168 63532 35488 65044
rect 35168 63476 35196 63532
rect 35252 63476 35300 63532
rect 35356 63476 35404 63532
rect 35460 63476 35488 63532
rect 35168 61964 35488 63476
rect 35168 61908 35196 61964
rect 35252 61908 35300 61964
rect 35356 61908 35404 61964
rect 35460 61908 35488 61964
rect 35168 60396 35488 61908
rect 35168 60340 35196 60396
rect 35252 60340 35300 60396
rect 35356 60340 35404 60396
rect 35460 60340 35488 60396
rect 35168 58828 35488 60340
rect 35168 58772 35196 58828
rect 35252 58772 35300 58828
rect 35356 58772 35404 58828
rect 35460 58772 35488 58828
rect 35168 57260 35488 58772
rect 35168 57204 35196 57260
rect 35252 57204 35300 57260
rect 35356 57204 35404 57260
rect 35460 57204 35488 57260
rect 35168 55692 35488 57204
rect 35168 55636 35196 55692
rect 35252 55636 35300 55692
rect 35356 55636 35404 55692
rect 35460 55636 35488 55692
rect 35168 54124 35488 55636
rect 35168 54068 35196 54124
rect 35252 54068 35300 54124
rect 35356 54068 35404 54124
rect 35460 54068 35488 54124
rect 35168 52556 35488 54068
rect 35168 52500 35196 52556
rect 35252 52500 35300 52556
rect 35356 52500 35404 52556
rect 35460 52500 35488 52556
rect 35168 50988 35488 52500
rect 35168 50932 35196 50988
rect 35252 50932 35300 50988
rect 35356 50932 35404 50988
rect 35460 50932 35488 50988
rect 35168 49420 35488 50932
rect 35168 49364 35196 49420
rect 35252 49364 35300 49420
rect 35356 49364 35404 49420
rect 35460 49364 35488 49420
rect 35168 47852 35488 49364
rect 35168 47796 35196 47852
rect 35252 47796 35300 47852
rect 35356 47796 35404 47852
rect 35460 47796 35488 47852
rect 35168 46284 35488 47796
rect 35168 46228 35196 46284
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35460 46228 35488 46284
rect 35168 44716 35488 46228
rect 35168 44660 35196 44716
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35460 44660 35488 44716
rect 35168 43148 35488 44660
rect 35168 43092 35196 43148
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35460 43092 35488 43148
rect 35168 41580 35488 43092
rect 35168 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35488 41580
rect 35168 40012 35488 41524
rect 35168 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35488 40012
rect 35168 38444 35488 39956
rect 35168 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35488 38444
rect 35168 36876 35488 38388
rect 35168 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35488 36876
rect 35168 35308 35488 36820
rect 35168 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35488 35308
rect 35168 33740 35488 35252
rect 35168 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35488 33740
rect 35168 32172 35488 33684
rect 35168 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35488 32172
rect 35168 30604 35488 32116
rect 35168 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35488 30604
rect 35168 29036 35488 30548
rect 35168 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35488 29036
rect 35168 27468 35488 28980
rect 35168 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35488 27468
rect 35168 25900 35488 27412
rect 47180 75684 47236 75694
rect 35168 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35488 25900
rect 35168 24332 35488 25844
rect 46060 26740 46116 26750
rect 35168 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35488 24332
rect 35168 22764 35488 24276
rect 43596 24500 43652 24510
rect 40460 23492 40964 23518
rect 40516 23462 40908 23492
rect 40460 23426 40516 23436
rect 40908 23426 40964 23436
rect 35168 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35488 22764
rect 43596 22820 43652 24444
rect 46060 23156 46116 26684
rect 46060 23090 46116 23100
rect 43596 22754 43652 22764
rect 19808 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20128 20412
rect 19808 18844 20128 20356
rect 34524 21476 34580 21486
rect 34524 20020 34580 21420
rect 34524 19954 34580 19964
rect 35168 21196 35488 22708
rect 35168 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35488 21196
rect 35168 19628 35488 21140
rect 47180 20804 47236 75628
rect 47404 55468 47460 76300
rect 47180 20738 47236 20748
rect 47292 55412 47460 55468
rect 50528 75292 50848 76804
rect 50528 75236 50556 75292
rect 50612 75236 50660 75292
rect 50716 75236 50764 75292
rect 50820 75236 50848 75292
rect 50528 73724 50848 75236
rect 50528 73668 50556 73724
rect 50612 73668 50660 73724
rect 50716 73668 50764 73724
rect 50820 73668 50848 73724
rect 50528 72156 50848 73668
rect 50528 72100 50556 72156
rect 50612 72100 50660 72156
rect 50716 72100 50764 72156
rect 50820 72100 50848 72156
rect 50528 70588 50848 72100
rect 50528 70532 50556 70588
rect 50612 70532 50660 70588
rect 50716 70532 50764 70588
rect 50820 70532 50848 70588
rect 50528 69020 50848 70532
rect 50528 68964 50556 69020
rect 50612 68964 50660 69020
rect 50716 68964 50764 69020
rect 50820 68964 50848 69020
rect 50528 67452 50848 68964
rect 50528 67396 50556 67452
rect 50612 67396 50660 67452
rect 50716 67396 50764 67452
rect 50820 67396 50848 67452
rect 50528 65884 50848 67396
rect 50528 65828 50556 65884
rect 50612 65828 50660 65884
rect 50716 65828 50764 65884
rect 50820 65828 50848 65884
rect 50528 64316 50848 65828
rect 50528 64260 50556 64316
rect 50612 64260 50660 64316
rect 50716 64260 50764 64316
rect 50820 64260 50848 64316
rect 50528 62748 50848 64260
rect 50528 62692 50556 62748
rect 50612 62692 50660 62748
rect 50716 62692 50764 62748
rect 50820 62692 50848 62748
rect 50528 61180 50848 62692
rect 50528 61124 50556 61180
rect 50612 61124 50660 61180
rect 50716 61124 50764 61180
rect 50820 61124 50848 61180
rect 50528 59612 50848 61124
rect 50528 59556 50556 59612
rect 50612 59556 50660 59612
rect 50716 59556 50764 59612
rect 50820 59556 50848 59612
rect 50528 58044 50848 59556
rect 50528 57988 50556 58044
rect 50612 57988 50660 58044
rect 50716 57988 50764 58044
rect 50820 57988 50848 58044
rect 50528 56476 50848 57988
rect 50528 56420 50556 56476
rect 50612 56420 50660 56476
rect 50716 56420 50764 56476
rect 50820 56420 50848 56476
rect 35168 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35488 19628
rect 19808 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20128 18844
rect 19808 17276 20128 18788
rect 28700 19236 28756 19246
rect 28700 18564 28756 19180
rect 28700 18498 28756 18508
rect 19808 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20128 17276
rect 19808 15708 20128 17220
rect 19808 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20128 15708
rect 19808 14140 20128 15652
rect 19808 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20128 14140
rect 19808 12572 20128 14084
rect 19808 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20128 12572
rect 19808 11004 20128 12516
rect 4448 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4768 10220
rect 4448 8652 4768 10164
rect 4448 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4768 8652
rect 4448 7084 4768 8596
rect 17836 10948 17892 10958
rect 4448 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4768 7084
rect 4448 5516 4768 7028
rect 4448 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4768 5516
rect 4448 3948 4768 5460
rect 14364 7924 14420 7934
rect 14364 5236 14420 7868
rect 17836 7812 17892 10892
rect 19808 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20128 11004
rect 19808 9436 20128 10948
rect 19808 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20128 9436
rect 17836 7746 17892 7756
rect 19628 8372 19684 8382
rect 19628 7476 19684 8316
rect 19628 7410 19684 7420
rect 19808 7868 20128 9380
rect 35168 18060 35488 19572
rect 35168 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35488 18060
rect 35168 16492 35488 18004
rect 47292 16884 47348 55412
rect 50528 54908 50848 56420
rect 50528 54852 50556 54908
rect 50612 54852 50660 54908
rect 50716 54852 50764 54908
rect 50820 54852 50848 54908
rect 50528 53340 50848 54852
rect 50528 53284 50556 53340
rect 50612 53284 50660 53340
rect 50716 53284 50764 53340
rect 50820 53284 50848 53340
rect 50528 51772 50848 53284
rect 50528 51716 50556 51772
rect 50612 51716 50660 51772
rect 50716 51716 50764 51772
rect 50820 51716 50848 51772
rect 50528 50204 50848 51716
rect 50528 50148 50556 50204
rect 50612 50148 50660 50204
rect 50716 50148 50764 50204
rect 50820 50148 50848 50204
rect 50528 48636 50848 50148
rect 50528 48580 50556 48636
rect 50612 48580 50660 48636
rect 50716 48580 50764 48636
rect 50820 48580 50848 48636
rect 50528 47068 50848 48580
rect 50528 47012 50556 47068
rect 50612 47012 50660 47068
rect 50716 47012 50764 47068
rect 50820 47012 50848 47068
rect 50528 45500 50848 47012
rect 50528 45444 50556 45500
rect 50612 45444 50660 45500
rect 50716 45444 50764 45500
rect 50820 45444 50848 45500
rect 50528 43932 50848 45444
rect 50528 43876 50556 43932
rect 50612 43876 50660 43932
rect 50716 43876 50764 43932
rect 50820 43876 50848 43932
rect 50528 42364 50848 43876
rect 50528 42308 50556 42364
rect 50612 42308 50660 42364
rect 50716 42308 50764 42364
rect 50820 42308 50848 42364
rect 50528 40796 50848 42308
rect 50528 40740 50556 40796
rect 50612 40740 50660 40796
rect 50716 40740 50764 40796
rect 50820 40740 50848 40796
rect 50528 39228 50848 40740
rect 50528 39172 50556 39228
rect 50612 39172 50660 39228
rect 50716 39172 50764 39228
rect 50820 39172 50848 39228
rect 50528 37660 50848 39172
rect 50528 37604 50556 37660
rect 50612 37604 50660 37660
rect 50716 37604 50764 37660
rect 50820 37604 50848 37660
rect 50528 36092 50848 37604
rect 50528 36036 50556 36092
rect 50612 36036 50660 36092
rect 50716 36036 50764 36092
rect 50820 36036 50848 36092
rect 50528 34524 50848 36036
rect 50528 34468 50556 34524
rect 50612 34468 50660 34524
rect 50716 34468 50764 34524
rect 50820 34468 50848 34524
rect 50528 32956 50848 34468
rect 50528 32900 50556 32956
rect 50612 32900 50660 32956
rect 50716 32900 50764 32956
rect 50820 32900 50848 32956
rect 50528 31388 50848 32900
rect 50528 31332 50556 31388
rect 50612 31332 50660 31388
rect 50716 31332 50764 31388
rect 50820 31332 50848 31388
rect 50528 29820 50848 31332
rect 65888 76076 66208 76892
rect 65888 76020 65916 76076
rect 65972 76020 66020 76076
rect 66076 76020 66124 76076
rect 66180 76020 66208 76076
rect 65888 74508 66208 76020
rect 65888 74452 65916 74508
rect 65972 74452 66020 74508
rect 66076 74452 66124 74508
rect 66180 74452 66208 74508
rect 65888 72940 66208 74452
rect 65888 72884 65916 72940
rect 65972 72884 66020 72940
rect 66076 72884 66124 72940
rect 66180 72884 66208 72940
rect 65888 71372 66208 72884
rect 65888 71316 65916 71372
rect 65972 71316 66020 71372
rect 66076 71316 66124 71372
rect 66180 71316 66208 71372
rect 65888 69804 66208 71316
rect 65888 69748 65916 69804
rect 65972 69748 66020 69804
rect 66076 69748 66124 69804
rect 66180 69748 66208 69804
rect 65888 68236 66208 69748
rect 65888 68180 65916 68236
rect 65972 68180 66020 68236
rect 66076 68180 66124 68236
rect 66180 68180 66208 68236
rect 65888 66668 66208 68180
rect 65888 66612 65916 66668
rect 65972 66612 66020 66668
rect 66076 66612 66124 66668
rect 66180 66612 66208 66668
rect 65888 65100 66208 66612
rect 65888 65044 65916 65100
rect 65972 65044 66020 65100
rect 66076 65044 66124 65100
rect 66180 65044 66208 65100
rect 65888 63532 66208 65044
rect 65888 63476 65916 63532
rect 65972 63476 66020 63532
rect 66076 63476 66124 63532
rect 66180 63476 66208 63532
rect 65888 61964 66208 63476
rect 65888 61908 65916 61964
rect 65972 61908 66020 61964
rect 66076 61908 66124 61964
rect 66180 61908 66208 61964
rect 65888 60396 66208 61908
rect 65888 60340 65916 60396
rect 65972 60340 66020 60396
rect 66076 60340 66124 60396
rect 66180 60340 66208 60396
rect 65888 58828 66208 60340
rect 65888 58772 65916 58828
rect 65972 58772 66020 58828
rect 66076 58772 66124 58828
rect 66180 58772 66208 58828
rect 65888 57260 66208 58772
rect 65888 57204 65916 57260
rect 65972 57204 66020 57260
rect 66076 57204 66124 57260
rect 66180 57204 66208 57260
rect 65888 55692 66208 57204
rect 65888 55636 65916 55692
rect 65972 55636 66020 55692
rect 66076 55636 66124 55692
rect 66180 55636 66208 55692
rect 65888 54124 66208 55636
rect 65888 54068 65916 54124
rect 65972 54068 66020 54124
rect 66076 54068 66124 54124
rect 66180 54068 66208 54124
rect 73164 76580 73220 76590
rect 65888 52556 66208 54068
rect 65888 52500 65916 52556
rect 65972 52500 66020 52556
rect 66076 52500 66124 52556
rect 66180 52500 66208 52556
rect 65888 50988 66208 52500
rect 65888 50932 65916 50988
rect 65972 50932 66020 50988
rect 66076 50932 66124 50988
rect 66180 50932 66208 50988
rect 65888 49420 66208 50932
rect 65888 49364 65916 49420
rect 65972 49364 66020 49420
rect 66076 49364 66124 49420
rect 66180 49364 66208 49420
rect 65888 47852 66208 49364
rect 65888 47796 65916 47852
rect 65972 47796 66020 47852
rect 66076 47796 66124 47852
rect 66180 47796 66208 47852
rect 65888 46284 66208 47796
rect 65888 46228 65916 46284
rect 65972 46228 66020 46284
rect 66076 46228 66124 46284
rect 66180 46228 66208 46284
rect 65888 44716 66208 46228
rect 65888 44660 65916 44716
rect 65972 44660 66020 44716
rect 66076 44660 66124 44716
rect 66180 44660 66208 44716
rect 65888 43148 66208 44660
rect 65888 43092 65916 43148
rect 65972 43092 66020 43148
rect 66076 43092 66124 43148
rect 66180 43092 66208 43148
rect 65888 41580 66208 43092
rect 65888 41524 65916 41580
rect 65972 41524 66020 41580
rect 66076 41524 66124 41580
rect 66180 41524 66208 41580
rect 72604 54068 72660 54078
rect 65888 40012 66208 41524
rect 72044 41524 72100 41534
rect 72044 40964 72100 41468
rect 72044 40898 72100 40908
rect 65888 39956 65916 40012
rect 65972 39956 66020 40012
rect 66076 39956 66124 40012
rect 66180 39956 66208 40012
rect 65888 38444 66208 39956
rect 72492 40852 72548 40862
rect 65888 38388 65916 38444
rect 65972 38388 66020 38444
rect 66076 38388 66124 38444
rect 66180 38388 66208 38444
rect 65888 36876 66208 38388
rect 69468 39060 69524 39070
rect 69468 38388 69524 39004
rect 69468 38322 69524 38332
rect 65888 36820 65916 36876
rect 65972 36820 66020 36876
rect 66076 36820 66124 36876
rect 66180 36820 66208 36876
rect 72492 36932 72548 40796
rect 72492 36866 72548 36876
rect 65888 35308 66208 36820
rect 65888 35252 65916 35308
rect 65972 35252 66020 35308
rect 66076 35252 66124 35308
rect 66180 35252 66208 35308
rect 65888 33740 66208 35252
rect 65888 33684 65916 33740
rect 65972 33684 66020 33740
rect 66076 33684 66124 33740
rect 66180 33684 66208 33740
rect 65888 32172 66208 33684
rect 65888 32116 65916 32172
rect 65972 32116 66020 32172
rect 66076 32116 66124 32172
rect 66180 32116 66208 32172
rect 50528 29764 50556 29820
rect 50612 29764 50660 29820
rect 50716 29764 50764 29820
rect 50820 29764 50848 29820
rect 50528 28252 50848 29764
rect 50528 28196 50556 28252
rect 50612 28196 50660 28252
rect 50716 28196 50764 28252
rect 50820 28196 50848 28252
rect 50528 26684 50848 28196
rect 50528 26628 50556 26684
rect 50612 26628 50660 26684
rect 50716 26628 50764 26684
rect 50820 26628 50848 26684
rect 51212 30772 51268 30782
rect 51212 26740 51268 30716
rect 65888 30604 66208 32116
rect 71148 32116 71204 32126
rect 65888 30548 65916 30604
rect 65972 30548 66020 30604
rect 66076 30548 66124 30604
rect 66180 30548 66208 30604
rect 65888 29036 66208 30548
rect 70924 30772 70980 30782
rect 65888 28980 65916 29036
rect 65972 28980 66020 29036
rect 66076 28980 66124 29036
rect 66180 28980 66208 29036
rect 65888 27468 66208 28980
rect 65888 27412 65916 27468
rect 65972 27412 66020 27468
rect 66076 27412 66124 27468
rect 66180 27412 66208 27468
rect 51212 26674 51268 26684
rect 56700 26852 56756 26862
rect 50528 25116 50848 26628
rect 56700 26516 56756 26796
rect 56700 26450 56756 26460
rect 50528 25060 50556 25116
rect 50612 25060 50660 25116
rect 50716 25060 50764 25116
rect 50820 25060 50848 25116
rect 50528 23548 50848 25060
rect 50092 23492 50148 23502
rect 47628 22372 47684 22382
rect 47628 22036 47684 22316
rect 47628 21970 47684 21980
rect 50092 20020 50148 23436
rect 50092 19954 50148 19964
rect 50528 23492 50556 23548
rect 50612 23492 50660 23548
rect 50716 23492 50764 23548
rect 50820 23492 50848 23548
rect 50528 21980 50848 23492
rect 50528 21924 50556 21980
rect 50612 21924 50660 21980
rect 50716 21924 50764 21980
rect 50820 21924 50848 21980
rect 50528 20412 50848 21924
rect 50528 20356 50556 20412
rect 50612 20356 50660 20412
rect 50716 20356 50764 20412
rect 50820 20356 50848 20412
rect 47292 16818 47348 16828
rect 50528 18844 50848 20356
rect 50528 18788 50556 18844
rect 50612 18788 50660 18844
rect 50716 18788 50764 18844
rect 50820 18788 50848 18844
rect 50528 17276 50848 18788
rect 50528 17220 50556 17276
rect 50612 17220 50660 17276
rect 50716 17220 50764 17276
rect 50820 17220 50848 17276
rect 35168 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35488 16492
rect 35168 14924 35488 16436
rect 35168 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35488 14924
rect 35168 13356 35488 14868
rect 35168 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35488 13356
rect 35168 11788 35488 13300
rect 35168 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35488 11788
rect 35168 10220 35488 11732
rect 50528 15708 50848 17220
rect 50528 15652 50556 15708
rect 50612 15652 50660 15708
rect 50716 15652 50764 15708
rect 50820 15652 50848 15708
rect 50528 14140 50848 15652
rect 50528 14084 50556 14140
rect 50612 14084 50660 14140
rect 50716 14084 50764 14140
rect 50820 14084 50848 14140
rect 50528 12572 50848 14084
rect 50528 12516 50556 12572
rect 50612 12516 50660 12572
rect 50716 12516 50764 12572
rect 50820 12516 50848 12572
rect 44492 11396 44548 11406
rect 44492 10724 44548 11340
rect 44492 10658 44548 10668
rect 50528 11004 50848 12516
rect 50528 10948 50556 11004
rect 50612 10948 50660 11004
rect 50716 10948 50764 11004
rect 50820 10948 50848 11004
rect 35168 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35488 10220
rect 35168 8652 35488 10164
rect 35168 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35488 8652
rect 19808 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20128 7868
rect 17164 6692 17220 6702
rect 14364 5170 14420 5180
rect 14700 6468 14756 6478
rect 14700 5124 14756 6412
rect 17164 6020 17220 6636
rect 17164 5954 17220 5964
rect 19808 6300 20128 7812
rect 20188 8372 20244 8382
rect 20188 7476 20244 8316
rect 20188 7410 20244 7420
rect 35168 7084 35488 8596
rect 23212 7028 23268 7038
rect 19808 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20128 6300
rect 14700 5058 14756 5068
rect 15148 4788 15204 4798
rect 4448 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4768 3948
rect 4448 3076 4768 3892
rect 7196 4676 7252 4686
rect 7196 3556 7252 4620
rect 7196 3490 7252 3500
rect 15148 4228 15204 4732
rect 15148 3556 15204 4172
rect 19292 4788 19348 4798
rect 19292 3668 19348 4732
rect 19292 3602 19348 3612
rect 19808 4732 20128 6244
rect 21980 6356 22036 6366
rect 19808 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20128 4732
rect 15148 3490 15204 3500
rect 19808 3164 20128 4676
rect 20412 5012 20468 5022
rect 20300 4340 20356 4350
rect 20300 3780 20356 4284
rect 20300 3714 20356 3724
rect 20412 3668 20468 4956
rect 20636 4452 20692 4462
rect 20636 3780 20692 4396
rect 20636 3714 20692 3724
rect 20412 3602 20468 3612
rect 19808 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20128 3164
rect 21980 3220 22036 6300
rect 22204 5348 22260 5358
rect 22204 4228 22260 5292
rect 23212 4900 23268 6972
rect 35168 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35488 7084
rect 23212 4834 23268 4844
rect 30156 6580 30212 6590
rect 22204 4162 22260 4172
rect 21980 3154 22036 3164
rect 30156 3220 30212 6524
rect 30156 3154 30212 3164
rect 35168 5516 35488 7028
rect 35168 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35488 5516
rect 35168 3948 35488 5460
rect 35168 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35488 3948
rect 19808 3076 20128 3108
rect 35168 3076 35488 3892
rect 50528 9436 50848 10948
rect 50528 9380 50556 9436
rect 50612 9380 50660 9436
rect 50716 9380 50764 9436
rect 50820 9380 50848 9436
rect 50528 7868 50848 9380
rect 50528 7812 50556 7868
rect 50612 7812 50660 7868
rect 50716 7812 50764 7868
rect 50820 7812 50848 7868
rect 50528 6300 50848 7812
rect 50528 6244 50556 6300
rect 50612 6244 50660 6300
rect 50716 6244 50764 6300
rect 50820 6244 50848 6300
rect 50528 4732 50848 6244
rect 50528 4676 50556 4732
rect 50612 4676 50660 4732
rect 50716 4676 50764 4732
rect 50820 4676 50848 4732
rect 50528 3164 50848 4676
rect 50528 3108 50556 3164
rect 50612 3108 50660 3164
rect 50716 3108 50764 3164
rect 50820 3108 50848 3164
rect 50528 3076 50848 3108
rect 65888 25900 66208 27412
rect 69580 29428 69636 29438
rect 69580 26404 69636 29372
rect 70924 26516 70980 30716
rect 70924 26450 70980 26460
rect 69580 26338 69636 26348
rect 65888 25844 65916 25900
rect 65972 25844 66020 25900
rect 66076 25844 66124 25900
rect 66180 25844 66208 25900
rect 65888 24332 66208 25844
rect 71148 25172 71204 32060
rect 71148 25106 71204 25116
rect 71372 30212 71428 30222
rect 65888 24276 65916 24332
rect 65972 24276 66020 24332
rect 66076 24276 66124 24332
rect 66180 24276 66208 24332
rect 71372 24388 71428 30156
rect 72604 29988 72660 54012
rect 73164 36484 73220 76524
rect 76524 75684 76580 75694
rect 76412 64036 76468 64046
rect 76188 62244 76244 62254
rect 75404 61572 75460 61582
rect 74956 59108 75012 59118
rect 74732 47012 74788 47022
rect 74060 46900 74116 46910
rect 73164 36418 73220 36428
rect 73500 37828 73556 37838
rect 73276 34692 73332 34702
rect 72604 29922 72660 29932
rect 72716 30100 72772 30110
rect 72716 28532 72772 30044
rect 72716 26964 72772 28476
rect 73164 27188 73220 27198
rect 73164 26908 73220 27132
rect 72716 26898 72772 26908
rect 73052 26852 73220 26908
rect 73052 26628 73108 26852
rect 73052 26562 73108 26572
rect 71372 24322 71428 24332
rect 65888 22764 66208 24276
rect 73276 23940 73332 34636
rect 73500 30996 73556 37772
rect 73500 30930 73556 30940
rect 74060 27972 74116 46844
rect 74508 39060 74564 39070
rect 74284 38948 74340 38958
rect 74172 37828 74228 37838
rect 74172 37268 74228 37772
rect 74172 37202 74228 37212
rect 74284 37044 74340 38892
rect 74284 36978 74340 36988
rect 74508 35476 74564 39004
rect 74508 35410 74564 35420
rect 74620 35588 74676 35598
rect 74620 28644 74676 35532
rect 74732 31444 74788 46956
rect 74732 31378 74788 31388
rect 74844 41860 74900 41870
rect 74844 40404 74900 41804
rect 74620 28578 74676 28588
rect 74732 30996 74788 31006
rect 74060 27906 74116 27916
rect 74732 26964 74788 30940
rect 74732 26898 74788 26908
rect 74844 26908 74900 40348
rect 74956 28308 75012 59052
rect 75068 38276 75124 38286
rect 75068 36036 75124 38220
rect 75068 35970 75124 35980
rect 75068 33684 75124 33694
rect 75068 32340 75124 33628
rect 75068 32274 75124 32284
rect 75404 28980 75460 61516
rect 75740 35028 75796 35038
rect 75740 31892 75796 34972
rect 75740 31826 75796 31836
rect 75404 28914 75460 28924
rect 75628 29316 75684 29326
rect 74956 27972 75012 28252
rect 74956 27906 75012 27916
rect 75516 27412 75572 27422
rect 74844 26852 75012 26908
rect 73276 23874 73332 23884
rect 65888 22708 65916 22764
rect 65972 22708 66020 22764
rect 66076 22708 66124 22764
rect 66180 22708 66208 22764
rect 65888 21196 66208 22708
rect 74956 21924 75012 26852
rect 75516 26852 75572 27356
rect 75516 26786 75572 26796
rect 75628 26068 75684 29260
rect 76188 27972 76244 62188
rect 76300 60900 76356 60910
rect 76300 28980 76356 60844
rect 76412 29764 76468 63980
rect 76524 37268 76580 75628
rect 76748 69188 76804 69198
rect 76524 37202 76580 37212
rect 76636 66052 76692 66062
rect 76636 30212 76692 65996
rect 76748 33460 76804 69132
rect 76748 33394 76804 33404
rect 76860 68516 76916 68526
rect 76860 31780 76916 68460
rect 77084 64708 77140 64718
rect 76972 38836 77028 38846
rect 76972 37044 77028 38780
rect 76972 36978 77028 36988
rect 76860 31714 76916 31724
rect 77084 30884 77140 64652
rect 77644 42644 77700 42654
rect 77644 40964 77700 42588
rect 77644 40898 77700 40908
rect 77868 37716 77924 37726
rect 77868 35140 77924 37660
rect 77868 35074 77924 35084
rect 77084 30818 77140 30828
rect 76636 30146 76692 30156
rect 76412 29540 76468 29708
rect 76412 29474 76468 29484
rect 76300 28914 76356 28924
rect 76188 27636 76244 27916
rect 76188 27570 76244 27580
rect 75628 26002 75684 26012
rect 76748 22484 76804 22494
rect 74956 21858 75012 21868
rect 75740 22372 75796 22382
rect 65888 21140 65916 21196
rect 65972 21140 66020 21196
rect 66076 21140 66124 21196
rect 66180 21140 66208 21196
rect 65888 19628 66208 21140
rect 65888 19572 65916 19628
rect 65972 19572 66020 19628
rect 66076 19572 66124 19628
rect 66180 19572 66208 19628
rect 65888 18060 66208 19572
rect 65888 18004 65916 18060
rect 65972 18004 66020 18060
rect 66076 18004 66124 18060
rect 66180 18004 66208 18060
rect 65888 16492 66208 18004
rect 65888 16436 65916 16492
rect 65972 16436 66020 16492
rect 66076 16436 66124 16492
rect 66180 16436 66208 16492
rect 65888 14924 66208 16436
rect 65888 14868 65916 14924
rect 65972 14868 66020 14924
rect 66076 14868 66124 14924
rect 66180 14868 66208 14924
rect 65888 13356 66208 14868
rect 65888 13300 65916 13356
rect 65972 13300 66020 13356
rect 66076 13300 66124 13356
rect 66180 13300 66208 13356
rect 65888 11788 66208 13300
rect 75740 13076 75796 22316
rect 76748 13972 76804 22428
rect 77084 22372 77140 22382
rect 77084 15204 77140 22316
rect 77084 15138 77140 15148
rect 76748 13906 76804 13916
rect 75740 13010 75796 13020
rect 65888 11732 65916 11788
rect 65972 11732 66020 11788
rect 66076 11732 66124 11788
rect 66180 11732 66208 11788
rect 65888 10220 66208 11732
rect 65888 10164 65916 10220
rect 65972 10164 66020 10220
rect 66076 10164 66124 10220
rect 66180 10164 66208 10220
rect 65888 8652 66208 10164
rect 65888 8596 65916 8652
rect 65972 8596 66020 8652
rect 66076 8596 66124 8652
rect 66180 8596 66208 8652
rect 65888 7084 66208 8596
rect 65888 7028 65916 7084
rect 65972 7028 66020 7084
rect 66076 7028 66124 7084
rect 66180 7028 66208 7084
rect 65888 5516 66208 7028
rect 65888 5460 65916 5516
rect 65972 5460 66020 5516
rect 66076 5460 66124 5516
rect 66180 5460 66208 5516
rect 65888 3948 66208 5460
rect 65888 3892 65916 3948
rect 65972 3892 66020 3948
rect 66076 3892 66124 3948
rect 66180 3892 66208 3948
rect 65888 3076 66208 3892
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _0663_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 46480 0 -1 6272
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _0664_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 48832 0 1 6272
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  _0665_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 48048 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _0666_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 32032 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _0667_
timestamp 1698431365
transform 1 0 40320 0 1 4704
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _0668_
timestamp 1698431365
transform 1 0 36400 0 -1 4704
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _0669_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 43232 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _0670_
timestamp 1698431365
transform 1 0 34944 0 -1 6272
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _0671_
timestamp 1698431365
transform -1 0 36624 0 1 4704
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _0672_
timestamp 1698431365
transform 1 0 28560 0 -1 4704
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_4  _0673_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 32704 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _0674_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 41216 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0675_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 35952 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _0676_
timestamp 1698431365
transform 1 0 35840 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _0677_
timestamp 1698431365
transform 1 0 42336 0 -1 6272
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0678_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 43792 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0679_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 40544 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _0680_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 38416 0 1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _0681_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 40096 0 1 4704
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__or4_4  _0682_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 42336 0 1 7840
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _0683_
timestamp 1698431365
transform -1 0 40544 0 -1 6272
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _0684_
timestamp 1698431365
transform 1 0 42112 0 -1 4704
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _0685_
timestamp 1698431365
transform -1 0 44464 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _0686_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 47264 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0687_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 45248 0 -1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _0688_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 43792 0 1 7840
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _0689_
timestamp 1698431365
transform -1 0 46592 0 -1 17248
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _0690_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 46704 0 -1 18816
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _0691_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 41776 0 -1 7840
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _0692_
timestamp 1698431365
transform 1 0 38304 0 1 7840
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _0693_
timestamp 1698431365
transform 1 0 43456 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _0694_
timestamp 1698431365
transform 1 0 41776 0 -1 7840
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0695_
timestamp 1698431365
transform -1 0 42784 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0696_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 70336 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0697_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 72128 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0698_
timestamp 1698431365
transform 1 0 73696 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _0699_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 51856 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _0700_
timestamp 1698431365
transform 1 0 50064 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _0701_
timestamp 1698431365
transform 1 0 44688 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _0702_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 71120 0 1 40768
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _0703_
timestamp 1698431365
transform 1 0 73920 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0704_
timestamp 1698431365
transform 1 0 74816 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _0705_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 40768 0 -1 9408
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _0706_
timestamp 1698431365
transform 1 0 42000 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0707_
timestamp 1698431365
transform 1 0 70224 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0708_
timestamp 1698431365
transform -1 0 68880 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0709_
timestamp 1698431365
transform -1 0 61264 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0710_
timestamp 1698431365
transform -1 0 58912 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _0711_
timestamp 1698431365
transform -1 0 55776 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0712_
timestamp 1698431365
transform 1 0 55104 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _0713_
timestamp 1698431365
transform 1 0 55104 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0714_
timestamp 1698431365
transform 1 0 56000 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _0715_
timestamp 1698431365
transform 1 0 56448 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0716_
timestamp 1698431365
transform 1 0 56896 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _0717_
timestamp 1698431365
transform 1 0 57344 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0718_
timestamp 1698431365
transform 1 0 57792 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _0719_
timestamp 1698431365
transform 1 0 44688 0 1 4704
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0720_
timestamp 1698431365
transform 1 0 72352 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0721_
timestamp 1698431365
transform 1 0 73696 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0722_
timestamp 1698431365
transform 1 0 75152 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _0723_
timestamp 1698431365
transform 1 0 74592 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0724_
timestamp 1698431365
transform -1 0 78064 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _0725_
timestamp 1698431365
transform 1 0 74368 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0726_
timestamp 1698431365
transform 1 0 77728 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _0727_
timestamp 1698431365
transform 1 0 76048 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0728_
timestamp 1698431365
transform -1 0 78064 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _0729_
timestamp 1698431365
transform 1 0 74480 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0730_
timestamp 1698431365
transform 1 0 76832 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _0731_
timestamp 1698431365
transform 1 0 30688 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0732_
timestamp 1698431365
transform -1 0 42672 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0733_
timestamp 1698431365
transform -1 0 40880 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  _0734_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 37968 0 1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0735_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 74704 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0736_
timestamp 1698431365
transform 1 0 75376 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0737_
timestamp 1698431365
transform 1 0 74480 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0738_
timestamp 1698431365
transform 1 0 75152 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0739_
timestamp 1698431365
transform -1 0 44016 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0740_
timestamp 1698431365
transform -1 0 63840 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0741_
timestamp 1698431365
transform -1 0 63840 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _0742_
timestamp 1698431365
transform -1 0 62384 0 -1 40768
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _0743_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 73472 0 -1 26656
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0744_
timestamp 1698431365
transform -1 0 40208 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0745_
timestamp 1698431365
transform -1 0 37520 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0746_
timestamp 1698431365
transform 1 0 33712 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0747_
timestamp 1698431365
transform 1 0 40768 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0748_
timestamp 1698431365
transform -1 0 39536 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0749_
timestamp 1698431365
transform -1 0 36624 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0750_
timestamp 1698431365
transform 1 0 34160 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0751_
timestamp 1698431365
transform -1 0 34832 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0752_
timestamp 1698431365
transform 1 0 39872 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0753_
timestamp 1698431365
transform -1 0 36624 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0754_
timestamp 1698431365
transform -1 0 42336 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0755_
timestamp 1698431365
transform -1 0 37744 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _0756_
timestamp 1698431365
transform 1 0 33712 0 1 26656
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _0757_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 33040 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _0758_
timestamp 1698431365
transform -1 0 27328 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0759_
timestamp 1698431365
transform -1 0 74704 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0760_
timestamp 1698431365
transform -1 0 76496 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _0761_
timestamp 1698431365
transform -1 0 60928 0 -1 40768
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _0762_
timestamp 1698431365
transform 1 0 74144 0 1 25088
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0763_
timestamp 1698431365
transform 1 0 34608 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0764_
timestamp 1698431365
transform 1 0 35952 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0765_
timestamp 1698431365
transform -1 0 35616 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _0766_
timestamp 1698431365
transform -1 0 36400 0 -1 28224
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _0767_
timestamp 1698431365
transform 1 0 35392 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _0768_
timestamp 1698431365
transform 1 0 30240 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0769_
timestamp 1698431365
transform -1 0 73472 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0770_
timestamp 1698431365
transform 1 0 72800 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0771_
timestamp 1698431365
transform 1 0 75152 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _0772_
timestamp 1698431365
transform 1 0 60368 0 1 39200
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _0773_
timestamp 1698431365
transform 1 0 72240 0 1 23520
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0774_
timestamp 1698431365
transform 1 0 34160 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0775_
timestamp 1698431365
transform 1 0 35056 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0776_
timestamp 1698431365
transform 1 0 35728 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _0777_
timestamp 1698431365
transform -1 0 36736 0 -1 26656
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _0778_
timestamp 1698431365
transform 1 0 35616 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _0779_
timestamp 1698431365
transform 1 0 27440 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0780_
timestamp 1698431365
transform 1 0 72464 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0781_
timestamp 1698431365
transform 1 0 73024 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0782_
timestamp 1698431365
transform 1 0 76048 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0783_
timestamp 1698431365
transform 1 0 61488 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _0784_
timestamp 1698431365
transform -1 0 63840 0 -1 40768
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _0785_
timestamp 1698431365
transform 1 0 72128 0 -1 25088
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0786_
timestamp 1698431365
transform 1 0 33264 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0787_
timestamp 1698431365
transform 1 0 35056 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0788_
timestamp 1698431365
transform -1 0 35392 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _0789_
timestamp 1698431365
transform -1 0 36624 0 1 26656
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _0790_
timestamp 1698431365
transform 1 0 35728 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _0791_
timestamp 1698431365
transform -1 0 20272 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  _0792_
timestamp 1698431365
transform -1 0 40096 0 -1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0793_
timestamp 1698431365
transform 1 0 72128 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0794_
timestamp 1698431365
transform 1 0 76720 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0795_
timestamp 1698431365
transform 1 0 77392 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0796_
timestamp 1698431365
transform -1 0 64512 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0797_
timestamp 1698431365
transform -1 0 63392 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0798_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 63616 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0799_
timestamp 1698431365
transform -1 0 36624 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0800_
timestamp 1698431365
transform 1 0 34496 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0801_
timestamp 1698431365
transform -1 0 37520 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0802_
timestamp 1698431365
transform 1 0 35056 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0803_
timestamp 1698431365
transform 1 0 37520 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0804_
timestamp 1698431365
transform 1 0 37072 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0805_
timestamp 1698431365
transform 1 0 37072 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _0806_
timestamp 1698431365
transform 1 0 37632 0 1 28224
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _0807_
timestamp 1698431365
transform 1 0 37968 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _0808_
timestamp 1698431365
transform 1 0 23744 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0809_
timestamp 1698431365
transform 1 0 71008 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0810_
timestamp 1698431365
transform 1 0 76720 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0811_
timestamp 1698431365
transform 1 0 61712 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0812_
timestamp 1698431365
transform -1 0 63616 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0813_
timestamp 1698431365
transform 1 0 33600 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0814_
timestamp 1698431365
transform 1 0 35280 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0815_
timestamp 1698431365
transform 1 0 39200 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _0816_
timestamp 1698431365
transform 1 0 37744 0 -1 28224
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _0817_
timestamp 1698431365
transform 1 0 38080 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _0818_
timestamp 1698431365
transform 1 0 20272 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0819_
timestamp 1698431365
transform 1 0 71232 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0820_
timestamp 1698431365
transform -1 0 72128 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0821_
timestamp 1698431365
transform 1 0 71008 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0822_
timestamp 1698431365
transform 1 0 77392 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _0823_
timestamp 1698431365
transform 1 0 62608 0 1 40768
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _0824_
timestamp 1698431365
transform 1 0 72464 0 1 25088
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0825_
timestamp 1698431365
transform 1 0 34048 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0826_
timestamp 1698431365
transform 1 0 36848 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0827_
timestamp 1698431365
transform 1 0 36960 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _0828_
timestamp 1698431365
transform 1 0 37968 0 -1 26656
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _0829_
timestamp 1698431365
transform 1 0 36960 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _0830_
timestamp 1698431365
transform -1 0 23296 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0831_
timestamp 1698431365
transform -1 0 72912 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0832_
timestamp 1698431365
transform 1 0 70784 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0833_
timestamp 1698431365
transform 1 0 76720 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0834_
timestamp 1698431365
transform 1 0 64176 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _0835_
timestamp 1698431365
transform 1 0 64288 0 -1 40768
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _0836_
timestamp 1698431365
transform 1 0 70784 0 1 25088
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0837_
timestamp 1698431365
transform 1 0 35504 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0838_
timestamp 1698431365
transform 1 0 35616 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0839_
timestamp 1698431365
transform 1 0 41440 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _0840_
timestamp 1698431365
transform 1 0 37968 0 1 26656
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _0841_
timestamp 1698431365
transform -1 0 41888 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _0842_
timestamp 1698431365
transform -1 0 21952 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  _0843_
timestamp 1698431365
transform 1 0 41104 0 -1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0844_
timestamp 1698431365
transform 1 0 71680 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0845_
timestamp 1698431365
transform 1 0 76608 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0846_
timestamp 1698431365
transform 1 0 76608 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0847_
timestamp 1698431365
transform 1 0 65072 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _0848_
timestamp 1698431365
transform -1 0 66976 0 1 40768
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _0849_
timestamp 1698431365
transform 1 0 71008 0 1 20384
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0850_
timestamp 1698431365
transform -1 0 41440 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0851_
timestamp 1698431365
transform 1 0 37520 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0852_
timestamp 1698431365
transform -1 0 40320 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0853_
timestamp 1698431365
transform 1 0 39200 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0854_
timestamp 1698431365
transform 1 0 40096 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0855_
timestamp 1698431365
transform 1 0 42336 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0856_
timestamp 1698431365
transform -1 0 40544 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _0857_
timestamp 1698431365
transform 1 0 40768 0 -1 28224
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _0858_
timestamp 1698431365
transform 1 0 40768 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _0859_
timestamp 1698431365
transform 1 0 23408 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0860_
timestamp 1698431365
transform 1 0 72576 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0861_
timestamp 1698431365
transform -1 0 75824 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _0862_
timestamp 1698431365
transform 1 0 65408 0 1 39200
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _0863_
timestamp 1698431365
transform 1 0 70224 0 -1 21952
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0864_
timestamp 1698431365
transform 1 0 38080 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0865_
timestamp 1698431365
transform 1 0 39200 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0866_
timestamp 1698431365
transform 1 0 41776 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _0867_
timestamp 1698431365
transform 1 0 39424 0 1 26656
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _0868_
timestamp 1698431365
transform 1 0 40880 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _0869_
timestamp 1698431365
transform 1 0 25200 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0870_
timestamp 1698431365
transform 1 0 72240 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0871_
timestamp 1698431365
transform 1 0 72576 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0872_
timestamp 1698431365
transform 1 0 77280 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _0873_
timestamp 1698431365
transform -1 0 67200 0 -1 40768
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _0874_
timestamp 1698431365
transform -1 0 73808 0 -1 21952
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0875_
timestamp 1698431365
transform -1 0 38976 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0876_
timestamp 1698431365
transform 1 0 38304 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0877_
timestamp 1698431365
transform 1 0 41216 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _0878_
timestamp 1698431365
transform 1 0 40880 0 -1 26656
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _0879_
timestamp 1698431365
transform 1 0 40880 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _0880_
timestamp 1698431365
transform 1 0 25088 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0881_
timestamp 1698431365
transform 1 0 74032 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0882_
timestamp 1698431365
transform -1 0 74816 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0883_
timestamp 1698431365
transform 1 0 72912 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0884_
timestamp 1698431365
transform 1 0 75936 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0885_
timestamp 1698431365
transform -1 0 68992 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0886_
timestamp 1698431365
transform -1 0 67984 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _0887_
timestamp 1698431365
transform 1 0 65968 0 -1 39200
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _0888_
timestamp 1698431365
transform 1 0 72688 0 1 20384
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0889_
timestamp 1698431365
transform 1 0 38304 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0890_
timestamp 1698431365
transform 1 0 39200 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0891_
timestamp 1698431365
transform 1 0 40320 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _0892_
timestamp 1698431365
transform 1 0 40880 0 1 26656
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _0893_
timestamp 1698431365
transform 1 0 40880 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _0894_
timestamp 1698431365
transform 1 0 29008 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  _0895_
timestamp 1698431365
transform 1 0 42336 0 -1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0896_
timestamp 1698431365
transform 1 0 73696 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0897_
timestamp 1698431365
transform 1 0 76608 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0898_
timestamp 1698431365
transform 1 0 77056 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0899_
timestamp 1698431365
transform 1 0 65856 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _0900_
timestamp 1698431365
transform -1 0 68880 0 -1 39200
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _0901_
timestamp 1698431365
transform 1 0 72240 0 1 21952
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0902_
timestamp 1698431365
transform 1 0 37184 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0903_
timestamp 1698431365
transform 1 0 37184 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0904_
timestamp 1698431365
transform -1 0 40544 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0905_
timestamp 1698431365
transform 1 0 38752 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0906_
timestamp 1698431365
transform 1 0 41440 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0907_
timestamp 1698431365
transform 1 0 41664 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0908_
timestamp 1698431365
transform 1 0 42560 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _0909_
timestamp 1698431365
transform -1 0 43792 0 1 25088
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _0910_
timestamp 1698431365
transform 1 0 44352 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _0911_
timestamp 1698431365
transform 1 0 33376 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0912_
timestamp 1698431365
transform 1 0 72800 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0913_
timestamp 1698431365
transform 1 0 77280 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _0914_
timestamp 1698431365
transform 1 0 68880 0 -1 39200
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _0915_
timestamp 1698431365
transform 1 0 72128 0 -1 23520
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0916_
timestamp 1698431365
transform 1 0 37520 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0917_
timestamp 1698431365
transform 1 0 39312 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0918_
timestamp 1698431365
transform 1 0 43232 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _0919_
timestamp 1698431365
transform -1 0 44352 0 -1 26656
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _0920_
timestamp 1698431365
transform 1 0 44688 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _0921_
timestamp 1698431365
transform -1 0 30576 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0922_
timestamp 1698431365
transform 1 0 74032 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0923_
timestamp 1698431365
transform -1 0 75488 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0924_
timestamp 1698431365
transform -1 0 77280 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _0925_
timestamp 1698431365
transform 1 0 68208 0 1 37632
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _0926_
timestamp 1698431365
transform 1 0 73920 0 1 21952
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0927_
timestamp 1698431365
transform 1 0 37744 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0928_
timestamp 1698431365
transform 1 0 37856 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0929_
timestamp 1698431365
transform 1 0 43456 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _0930_
timestamp 1698431365
transform -1 0 46144 0 1 25088
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _0931_
timestamp 1698431365
transform -1 0 47040 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _0932_
timestamp 1698431365
transform -1 0 33824 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0933_
timestamp 1698431365
transform -1 0 77280 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0934_
timestamp 1698431365
transform 1 0 76048 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0935_
timestamp 1698431365
transform -1 0 77056 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0936_
timestamp 1698431365
transform -1 0 70336 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _0937_
timestamp 1698431365
transform 1 0 68432 0 1 39200
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _0938_
timestamp 1698431365
transform 1 0 74816 0 -1 23520
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0939_
timestamp 1698431365
transform 1 0 35280 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0940_
timestamp 1698431365
transform 1 0 37856 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0941_
timestamp 1698431365
transform 1 0 44688 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _0942_
timestamp 1698431365
transform 1 0 44016 0 -1 25088
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _0943_
timestamp 1698431365
transform 1 0 43568 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _0944_
timestamp 1698431365
transform 1 0 38752 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0945_
timestamp 1698431365
transform 1 0 46032 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  _0946_
timestamp 1698431365
transform 1 0 47040 0 -1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0947_
timestamp 1698431365
transform 1 0 74928 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0948_
timestamp 1698431365
transform 1 0 75824 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0949_
timestamp 1698431365
transform -1 0 77616 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0950_
timestamp 1698431365
transform 1 0 77616 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0951_
timestamp 1698431365
transform 1 0 68992 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0952_
timestamp 1698431365
transform -1 0 71904 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0953_
timestamp 1698431365
transform 1 0 70112 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0954_
timestamp 1698431365
transform -1 0 71456 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0955_
timestamp 1698431365
transform 1 0 45696 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0956_
timestamp 1698431365
transform 1 0 46144 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0957_
timestamp 1698431365
transform -1 0 48384 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0958_
timestamp 1698431365
transform 1 0 45472 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0959_
timestamp 1698431365
transform 1 0 46816 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0960_
timestamp 1698431365
transform -1 0 48048 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0961_
timestamp 1698431365
transform 1 0 47488 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0962_
timestamp 1698431365
transform 1 0 45136 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0963_
timestamp 1698431365
transform 1 0 45584 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0964_
timestamp 1698431365
transform 1 0 47040 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0965_
timestamp 1698431365
transform -1 0 45584 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _0966_
timestamp 1698431365
transform 1 0 46704 0 -1 18816
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _0967_
timestamp 1698431365
transform 1 0 46368 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _0968_
timestamp 1698431365
transform 1 0 37632 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0969_
timestamp 1698431365
transform 1 0 75712 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0970_
timestamp 1698431365
transform -1 0 75824 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0971_
timestamp 1698431365
transform 1 0 70336 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0972_
timestamp 1698431365
transform -1 0 71120 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0973_
timestamp 1698431365
transform 1 0 44688 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0974_
timestamp 1698431365
transform 1 0 46928 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0975_
timestamp 1698431365
transform 1 0 47824 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _0976_
timestamp 1698431365
transform 1 0 44912 0 1 17248
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _0977_
timestamp 1698431365
transform 1 0 46368 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _0978_
timestamp 1698431365
transform 1 0 34496 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0979_
timestamp 1698431365
transform 1 0 74480 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0980_
timestamp 1698431365
transform 1 0 75936 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0981_
timestamp 1698431365
transform 1 0 77392 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0982_
timestamp 1698431365
transform 1 0 70224 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0983_
timestamp 1698431365
transform -1 0 71568 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0984_
timestamp 1698431365
transform 1 0 44016 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0985_
timestamp 1698431365
transform 1 0 46032 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0986_
timestamp 1698431365
transform 1 0 47712 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _0987_
timestamp 1698431365
transform 1 0 46592 0 -1 17248
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _0988_
timestamp 1698431365
transform 1 0 48608 0 -1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _0989_
timestamp 1698431365
transform 1 0 35504 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0990_
timestamp 1698431365
transform 1 0 74704 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0991_
timestamp 1698431365
transform 1 0 76048 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0992_
timestamp 1698431365
transform -1 0 76720 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0993_
timestamp 1698431365
transform 1 0 70336 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0994_
timestamp 1698431365
transform -1 0 71904 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _0995_
timestamp 1698431365
transform 1 0 73808 0 1 29792
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0996_
timestamp 1698431365
transform 1 0 45248 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0997_
timestamp 1698431365
transform 1 0 46032 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0998_
timestamp 1698431365
transform 1 0 46928 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _0999_
timestamp 1698431365
transform 1 0 46480 0 1 20384
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _1000_
timestamp 1698431365
transform 1 0 46704 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1001_
timestamp 1698431365
transform 1 0 28000 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  _1002_
timestamp 1698431365
transform 1 0 50288 0 1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1003_
timestamp 1698431365
transform 1 0 76160 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1004_
timestamp 1698431365
transform -1 0 78064 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1005_
timestamp 1698431365
transform 1 0 76720 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1006_
timestamp 1698431365
transform -1 0 73696 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1007_
timestamp 1698431365
transform 1 0 72128 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1008_
timestamp 1698431365
transform -1 0 73024 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1009_
timestamp 1698431365
transform 1 0 45584 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1010_
timestamp 1698431365
transform 1 0 46816 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1011_
timestamp 1698431365
transform 1 0 46144 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1012_
timestamp 1698431365
transform 1 0 47152 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1013_
timestamp 1698431365
transform 1 0 49168 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1014_
timestamp 1698431365
transform -1 0 49280 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1015_
timestamp 1698431365
transform -1 0 50176 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1016_
timestamp 1698431365
transform -1 0 49616 0 1 20384
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _1017_
timestamp 1698431365
transform 1 0 48608 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1018_
timestamp 1698431365
transform 1 0 31808 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1019_
timestamp 1698431365
transform 1 0 76944 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1020_
timestamp 1698431365
transform -1 0 75936 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1021_
timestamp 1698431365
transform 1 0 73024 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1022_
timestamp 1698431365
transform -1 0 73920 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1023_
timestamp 1698431365
transform 1 0 44800 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1024_
timestamp 1698431365
transform 1 0 46256 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1025_
timestamp 1698431365
transform 1 0 48608 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1026_
timestamp 1698431365
transform 1 0 48608 0 -1 21952
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _1027_
timestamp 1698431365
transform 1 0 48608 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1028_
timestamp 1698431365
transform 1 0 27552 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1029_
timestamp 1698431365
transform 1 0 76272 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1030_
timestamp 1698431365
transform 1 0 76384 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1031_
timestamp 1698431365
transform 1 0 77056 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1032_
timestamp 1698431365
transform 1 0 72688 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1033_
timestamp 1698431365
transform -1 0 74928 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1034_
timestamp 1698431365
transform 1 0 44688 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1035_
timestamp 1698431365
transform 1 0 47040 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1036_
timestamp 1698431365
transform 1 0 48944 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1037_
timestamp 1698431365
transform 1 0 49616 0 1 20384
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _1038_
timestamp 1698431365
transform 1 0 48720 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1039_
timestamp 1698431365
transform -1 0 32144 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1040_
timestamp 1698431365
transform 1 0 75376 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1041_
timestamp 1698431365
transform 1 0 76384 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1042_
timestamp 1698431365
transform 1 0 77056 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1043_
timestamp 1698431365
transform 1 0 71008 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1044_
timestamp 1698431365
transform -1 0 74816 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1045_
timestamp 1698431365
transform -1 0 74592 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1046_
timestamp 1698431365
transform 1 0 44800 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1047_
timestamp 1698431365
transform 1 0 46144 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1048_
timestamp 1698431365
transform 1 0 49504 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1049_
timestamp 1698431365
transform 1 0 50064 0 -1 21952
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _1050_
timestamp 1698431365
transform 1 0 49056 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1051_
timestamp 1698431365
transform 1 0 43120 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  _1052_
timestamp 1698431365
transform 1 0 51184 0 1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1053_
timestamp 1698431365
transform 1 0 77056 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1054_
timestamp 1698431365
transform -1 0 75152 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1055_
timestamp 1698431365
transform -1 0 74144 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1056_
timestamp 1698431365
transform 1 0 74032 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1057_
timestamp 1698431365
transform 1 0 74368 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1058_
timestamp 1698431365
transform 1 0 74144 0 1 32928
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1059_
timestamp 1698431365
transform 1 0 45248 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1060_
timestamp 1698431365
transform 1 0 44912 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1061_
timestamp 1698431365
transform 1 0 46816 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1062_
timestamp 1698431365
transform 1 0 45920 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1063_
timestamp 1698431365
transform 1 0 50512 0 1 29792
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1064_
timestamp 1698431365
transform -1 0 51968 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1065_
timestamp 1698431365
transform 1 0 52528 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1066_
timestamp 1698431365
transform -1 0 51856 0 1 17248
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _1067_
timestamp 1698431365
transform 1 0 52528 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1068_
timestamp 1698431365
transform 1 0 45136 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1069_
timestamp 1698431365
transform 1 0 76160 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1070_
timestamp 1698431365
transform 1 0 77392 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1071_
timestamp 1698431365
transform 1 0 74704 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1072_
timestamp 1698431365
transform 1 0 74592 0 -1 32928
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1073_
timestamp 1698431365
transform 1 0 44688 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1074_
timestamp 1698431365
transform 1 0 46816 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1075_
timestamp 1698431365
transform 1 0 49952 0 -1 31360
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1076_
timestamp 1698431365
transform 1 0 52640 0 -1 20384
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _1077_
timestamp 1698431365
transform 1 0 52192 0 -1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1078_
timestamp 1698431365
transform 1 0 45248 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1079_
timestamp 1698431365
transform 1 0 75152 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1080_
timestamp 1698431365
transform -1 0 76832 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1081_
timestamp 1698431365
transform 1 0 77392 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1082_
timestamp 1698431365
transform 1 0 74928 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1083_
timestamp 1698431365
transform 1 0 76048 0 1 34496
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1084_
timestamp 1698431365
transform 1 0 44464 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1085_
timestamp 1698431365
transform 1 0 45920 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1086_
timestamp 1698431365
transform 1 0 50960 0 -1 31360
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1087_
timestamp 1698431365
transform -1 0 52976 0 -1 21952
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _1088_
timestamp 1698431365
transform 1 0 52192 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1089_
timestamp 1698431365
transform -1 0 42112 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1090_
timestamp 1698431365
transform 1 0 73696 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1091_
timestamp 1698431365
transform -1 0 77056 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1092_
timestamp 1698431365
transform 1 0 77392 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1093_
timestamp 1698431365
transform 1 0 69104 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1094_
timestamp 1698431365
transform -1 0 76944 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1095_
timestamp 1698431365
transform 1 0 76048 0 1 36064
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1096_
timestamp 1698431365
transform 1 0 44800 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1097_
timestamp 1698431365
transform 1 0 45920 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1098_
timestamp 1698431365
transform 1 0 50960 0 1 31360
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1099_
timestamp 1698431365
transform 1 0 52528 0 1 20384
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _1100_
timestamp 1698431365
transform -1 0 54880 0 -1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1101_
timestamp 1698431365
transform -1 0 40544 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  _1102_
timestamp 1698431365
transform 1 0 52528 0 1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1103_
timestamp 1698431365
transform -1 0 77728 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1104_
timestamp 1698431365
transform -1 0 77952 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1105_
timestamp 1698431365
transform -1 0 75824 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1106_
timestamp 1698431365
transform 1 0 74144 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1107_
timestamp 1698431365
transform 1 0 76944 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1108_
timestamp 1698431365
transform -1 0 78400 0 -1 37632
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1109_
timestamp 1698431365
transform 1 0 45920 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1110_
timestamp 1698431365
transform 1 0 45024 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1111_
timestamp 1698431365
transform 1 0 46592 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1112_
timestamp 1698431365
transform 1 0 45808 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1113_
timestamp 1698431365
transform 1 0 52864 0 1 32928
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1114_
timestamp 1698431365
transform 1 0 52976 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1115_
timestamp 1698431365
transform 1 0 52640 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1116_
timestamp 1698431365
transform 1 0 54096 0 -1 20384
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _1117_
timestamp 1698431365
transform 1 0 52864 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1118_
timestamp 1698431365
transform 1 0 44688 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1119_
timestamp 1698431365
transform -1 0 76720 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1120_
timestamp 1698431365
transform 1 0 77728 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1121_
timestamp 1698431365
transform 1 0 77056 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1122_
timestamp 1698431365
transform 1 0 76720 0 1 37632
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1123_
timestamp 1698431365
transform 1 0 45024 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1124_
timestamp 1698431365
transform 1 0 46592 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1125_
timestamp 1698431365
transform 1 0 53536 0 1 34496
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1126_
timestamp 1698431365
transform 1 0 53984 0 1 20384
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _1127_
timestamp 1698431365
transform 1 0 53536 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1128_
timestamp 1698431365
transform 1 0 40544 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1129_
timestamp 1698431365
transform 1 0 74928 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1130_
timestamp 1698431365
transform 1 0 76048 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1131_
timestamp 1698431365
transform 1 0 76720 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1132_
timestamp 1698431365
transform -1 0 77728 0 1 39200
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1133_
timestamp 1698431365
transform 1 0 44912 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1134_
timestamp 1698431365
transform 1 0 45696 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1135_
timestamp 1698431365
transform 1 0 54880 0 -1 36064
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1136_
timestamp 1698431365
transform -1 0 55328 0 -1 21952
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _1137_
timestamp 1698431365
transform 1 0 56448 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1138_
timestamp 1698431365
transform 1 0 44800 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1139_
timestamp 1698431365
transform -1 0 73472 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1140_
timestamp 1698431365
transform 1 0 77728 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1141_
timestamp 1698431365
transform 1 0 73024 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1142_
timestamp 1698431365
transform -1 0 74144 0 -1 40768
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1143_
timestamp 1698431365
transform 1 0 44912 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1144_
timestamp 1698431365
transform 1 0 45696 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1145_
timestamp 1698431365
transform 1 0 53872 0 -1 36064
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1146_
timestamp 1698431365
transform 1 0 55440 0 1 20384
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _1147_
timestamp 1698431365
transform -1 0 56224 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1148_
timestamp 1698431365
transform -1 0 42448 0 -1 39200
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1149_
timestamp 1698431365
transform -1 0 41440 0 -1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1150_
timestamp 1698431365
transform 1 0 42448 0 -1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1151_
timestamp 1698431365
transform -1 0 43008 0 -1 23520
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1152_
timestamp 1698431365
transform 1 0 74816 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1153_
timestamp 1698431365
transform 1 0 77616 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1154_
timestamp 1698431365
transform 1 0 40320 0 1 6272
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1155_
timestamp 1698431365
transform -1 0 30016 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1156_
timestamp 1698431365
transform -1 0 28448 0 1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1157_
timestamp 1698431365
transform -1 0 16352 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1158_
timestamp 1698431365
transform -1 0 15904 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1159_
timestamp 1698431365
transform 1 0 29568 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1160_
timestamp 1698431365
transform -1 0 28784 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1161_
timestamp 1698431365
transform -1 0 20384 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1162_
timestamp 1698431365
transform 1 0 20944 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1163_
timestamp 1698431365
transform -1 0 20832 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1164_
timestamp 1698431365
transform 1 0 17584 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1165_
timestamp 1698431365
transform -1 0 17920 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1166_
timestamp 1698431365
transform -1 0 11424 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1167_
timestamp 1698431365
transform 1 0 18256 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1168_
timestamp 1698431365
transform -1 0 14896 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1169_
timestamp 1698431365
transform -1 0 12096 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1170_
timestamp 1698431365
transform 1 0 18256 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1171_
timestamp 1698431365
transform -1 0 16016 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1172_
timestamp 1698431365
transform -1 0 15680 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1173_
timestamp 1698431365
transform 1 0 18032 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1174_
timestamp 1698431365
transform -1 0 17920 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1175_
timestamp 1698431365
transform 1 0 15904 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1176_
timestamp 1698431365
transform -1 0 18368 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1177_
timestamp 1698431365
transform -1 0 20384 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1178_
timestamp 1698431365
transform -1 0 21840 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1179_
timestamp 1698431365
transform 1 0 18816 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1180_
timestamp 1698431365
transform -1 0 18256 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1181_
timestamp 1698431365
transform 1 0 18368 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1182_
timestamp 1698431365
transform 1 0 19712 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1183_
timestamp 1698431365
transform 1 0 19936 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1184_
timestamp 1698431365
transform -1 0 17024 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1185_
timestamp 1698431365
transform 1 0 19600 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1186_
timestamp 1698431365
transform -1 0 19600 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1187_
timestamp 1698431365
transform -1 0 18144 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1188_
timestamp 1698431365
transform 1 0 19712 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1189_
timestamp 1698431365
transform -1 0 20160 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1190_
timestamp 1698431365
transform -1 0 28000 0 -1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1191_
timestamp 1698431365
transform -1 0 23072 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1192_
timestamp 1698431365
transform -1 0 20832 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1193_
timestamp 1698431365
transform -1 0 28784 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1194_
timestamp 1698431365
transform -1 0 27440 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1195_
timestamp 1698431365
transform 1 0 26432 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1196_
timestamp 1698431365
transform 1 0 26208 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1197_
timestamp 1698431365
transform -1 0 23520 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1198_
timestamp 1698431365
transform -1 0 22176 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1199_
timestamp 1698431365
transform 1 0 25872 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1200_
timestamp 1698431365
transform -1 0 24304 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1201_
timestamp 1698431365
transform 1 0 23632 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1202_
timestamp 1698431365
transform 1 0 25424 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1203_
timestamp 1698431365
transform -1 0 23632 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1204_
timestamp 1698431365
transform -1 0 21504 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1205_
timestamp 1698431365
transform -1 0 27216 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1206_
timestamp 1698431365
transform 1 0 27216 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1207_
timestamp 1698431365
transform -1 0 22736 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1208_
timestamp 1698431365
transform 1 0 22400 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1209_
timestamp 1698431365
transform -1 0 27440 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1210_
timestamp 1698431365
transform 1 0 14112 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1211_
timestamp 1698431365
transform 1 0 25088 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1212_
timestamp 1698431365
transform 1 0 25088 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1213_
timestamp 1698431365
transform -1 0 23184 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1214_
timestamp 1698431365
transform -1 0 21728 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1215_
timestamp 1698431365
transform -1 0 26880 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1216_
timestamp 1698431365
transform 1 0 26096 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1217_
timestamp 1698431365
transform -1 0 22288 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1218_
timestamp 1698431365
transform 1 0 24640 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1219_
timestamp 1698431365
transform -1 0 22848 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1220_
timestamp 1698431365
transform -1 0 22400 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1221_
timestamp 1698431365
transform 1 0 25088 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1222_
timestamp 1698431365
transform -1 0 23520 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1223_
timestamp 1698431365
transform 1 0 28784 0 -1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1224_
timestamp 1698431365
transform -1 0 28112 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1225_
timestamp 1698431365
transform -1 0 26208 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1226_
timestamp 1698431365
transform 1 0 30688 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1227_
timestamp 1698431365
transform -1 0 32480 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1228_
timestamp 1698431365
transform 1 0 33040 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1229_
timestamp 1698431365
transform 1 0 32032 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1230_
timestamp 1698431365
transform -1 0 30464 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1231_
timestamp 1698431365
transform -1 0 27888 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1232_
timestamp 1698431365
transform -1 0 33376 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1233_
timestamp 1698431365
transform 1 0 33824 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1234_
timestamp 1698431365
transform -1 0 27440 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1235_
timestamp 1698431365
transform 1 0 31584 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1236_
timestamp 1698431365
transform -1 0 30576 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1237_
timestamp 1698431365
transform -1 0 23520 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1238_
timestamp 1698431365
transform 1 0 32928 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1239_
timestamp 1698431365
transform -1 0 29680 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1240_
timestamp 1698431365
transform 1 0 30800 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1241_
timestamp 1698431365
transform 1 0 31920 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1242_
timestamp 1698431365
transform 1 0 32928 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1243_
timestamp 1698431365
transform 1 0 32816 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1244_
timestamp 1698431365
transform 1 0 34384 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1245_
timestamp 1698431365
transform 1 0 34496 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1246_
timestamp 1698431365
transform -1 0 30464 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1247_
timestamp 1698431365
transform 1 0 33600 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1248_
timestamp 1698431365
transform -1 0 31136 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1249_
timestamp 1698431365
transform -1 0 30688 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1250_
timestamp 1698431365
transform 1 0 32928 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1251_
timestamp 1698431365
transform -1 0 32256 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1252_
timestamp 1698431365
transform -1 0 29792 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1253_
timestamp 1698431365
transform 1 0 34496 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1254_
timestamp 1698431365
transform -1 0 34944 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1255_
timestamp 1698431365
transform -1 0 29792 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1256_
timestamp 1698431365
transform -1 0 25984 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1257_
timestamp 1698431365
transform -1 0 26768 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1258_
timestamp 1698431365
transform -1 0 25312 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1259_
timestamp 1698431365
transform 1 0 23296 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1260_
timestamp 1698431365
transform 1 0 23744 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1261_
timestamp 1698431365
transform -1 0 27776 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1262_
timestamp 1698431365
transform 1 0 23856 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1263_
timestamp 1698431365
transform -1 0 25984 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1264_
timestamp 1698431365
transform 1 0 23520 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1265_
timestamp 1698431365
transform -1 0 28336 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1266_
timestamp 1698431365
transform 1 0 23744 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1267_
timestamp 1698431365
transform -1 0 25984 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1268_
timestamp 1698431365
transform -1 0 22848 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1269_
timestamp 1698431365
transform -1 0 20272 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1270_
timestamp 1698431365
transform -1 0 18816 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1271_
timestamp 1698431365
transform 1 0 17360 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1272_
timestamp 1698431365
transform 1 0 20272 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1273_
timestamp 1698431365
transform -1 0 22064 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1274_
timestamp 1698431365
transform -1 0 17808 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1275_
timestamp 1698431365
transform -1 0 18144 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1276_
timestamp 1698431365
transform 1 0 19376 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1277_
timestamp 1698431365
transform -1 0 22064 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1278_
timestamp 1698431365
transform -1 0 22512 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1279_
timestamp 1698431365
transform -1 0 18928 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1280_
timestamp 1698431365
transform 1 0 18816 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1281_
timestamp 1698431365
transform -1 0 20608 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1282_
timestamp 1698431365
transform 1 0 18928 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1283_
timestamp 1698431365
transform -1 0 20944 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1284_
timestamp 1698431365
transform -1 0 18368 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1285_
timestamp 1698431365
transform -1 0 22736 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1286_
timestamp 1698431365
transform 1 0 19040 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1287_
timestamp 1698431365
transform 1 0 22512 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1288_
timestamp 1698431365
transform 1 0 26432 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1289_
timestamp 1698431365
transform 1 0 25200 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1290_
timestamp 1698431365
transform 1 0 26208 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1291_
timestamp 1698431365
transform -1 0 27888 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1292_
timestamp 1698431365
transform 1 0 26096 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1293_
timestamp 1698431365
transform -1 0 31584 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1294_
timestamp 1698431365
transform 1 0 25872 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1295_
timestamp 1698431365
transform -1 0 29904 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1296_
timestamp 1698431365
transform 1 0 27104 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1297_
timestamp 1698431365
transform -1 0 31808 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1298_
timestamp 1698431365
transform 1 0 29344 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1299_
timestamp 1698431365
transform -1 0 35840 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1300_
timestamp 1698431365
transform 1 0 28112 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1301_
timestamp 1698431365
transform 1 0 31360 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1302_
timestamp 1698431365
transform -1 0 31472 0 -1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1303_
timestamp 1698431365
transform -1 0 36176 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1304_
timestamp 1698431365
transform 1 0 32032 0 1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1305_
timestamp 1698431365
transform -1 0 35504 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1306_
timestamp 1698431365
transform 1 0 31472 0 -1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1307_
timestamp 1698431365
transform -1 0 33824 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1308_
timestamp 1698431365
transform 1 0 32032 0 -1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1309_
timestamp 1698431365
transform -1 0 33824 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1310_
timestamp 1698431365
transform -1 0 30576 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1311_
timestamp 1698431365
transform -1 0 29568 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1312_
timestamp 1698431365
transform -1 0 26768 0 -1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1313_
timestamp 1698431365
transform -1 0 26992 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1314_
timestamp 1698431365
transform -1 0 30128 0 -1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1315_
timestamp 1698431365
transform 1 0 27888 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1316_
timestamp 1698431365
transform 1 0 26768 0 -1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1317_
timestamp 1698431365
transform -1 0 27888 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1318_
timestamp 1698431365
transform 1 0 28336 0 -1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1319_
timestamp 1698431365
transform -1 0 29904 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1320_
timestamp 1698431365
transform 1 0 38640 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1321_
timestamp 1698431365
transform 1 0 36960 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1322_
timestamp 1698431365
transform 1 0 37520 0 -1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1323_
timestamp 1698431365
transform -1 0 41664 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1324_
timestamp 1698431365
transform 1 0 40768 0 -1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1325_
timestamp 1698431365
transform -1 0 43456 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1326_
timestamp 1698431365
transform 1 0 38080 0 -1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1327_
timestamp 1698431365
transform -1 0 43120 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1328_
timestamp 1698431365
transform -1 0 39872 0 -1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1329_
timestamp 1698431365
transform -1 0 40320 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1330_
timestamp 1698431365
transform 1 0 38304 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1331_
timestamp 1698431365
transform 1 0 36848 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1332_
timestamp 1698431365
transform 1 0 37184 0 1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1333_
timestamp 1698431365
transform -1 0 39760 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1334_
timestamp 1698431365
transform 1 0 36064 0 1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1335_
timestamp 1698431365
transform -1 0 43792 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1336_
timestamp 1698431365
transform -1 0 39984 0 1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1337_
timestamp 1698431365
transform 1 0 38528 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1338_
timestamp 1698431365
transform -1 0 36064 0 1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1339_
timestamp 1698431365
transform 1 0 43792 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1340_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 37968 0 -1 7840
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1341_
timestamp 1698431365
transform -1 0 38416 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1342_
timestamp 1698431365
transform -1 0 29568 0 1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1343_
timestamp 1698431365
transform -1 0 10640 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1344_
timestamp 1698431365
transform -1 0 9968 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1345_
timestamp 1698431365
transform -1 0 28896 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1346_
timestamp 1698431365
transform -1 0 13552 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1347_
timestamp 1698431365
transform -1 0 14000 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1348_
timestamp 1698431365
transform 1 0 11648 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1349_
timestamp 1698431365
transform -1 0 9632 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1350_
timestamp 1698431365
transform -1 0 8624 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1351_
timestamp 1698431365
transform 1 0 11648 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1352_
timestamp 1698431365
transform -1 0 9744 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1353_
timestamp 1698431365
transform -1 0 9296 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1354_
timestamp 1698431365
transform 1 0 11536 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1355_
timestamp 1698431365
transform -1 0 10080 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1356_
timestamp 1698431365
transform -1 0 9184 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1357_
timestamp 1698431365
transform 1 0 13328 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1358_
timestamp 1698431365
transform -1 0 13552 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1359_
timestamp 1698431365
transform -1 0 9744 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1360_
timestamp 1698431365
transform -1 0 7840 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1361_
timestamp 1698431365
transform -1 0 14000 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1362_
timestamp 1698431365
transform -1 0 15232 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1363_
timestamp 1698431365
transform 1 0 13888 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1364_
timestamp 1698431365
transform -1 0 11424 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1365_
timestamp 1698431365
transform -1 0 8512 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1366_
timestamp 1698431365
transform 1 0 13328 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1367_
timestamp 1698431365
transform -1 0 11088 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1368_
timestamp 1698431365
transform -1 0 9072 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1369_
timestamp 1698431365
transform 1 0 12208 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1370_
timestamp 1698431365
transform -1 0 12096 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1371_
timestamp 1698431365
transform 1 0 9744 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1372_
timestamp 1698431365
transform 1 0 14112 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1373_
timestamp 1698431365
transform -1 0 13888 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _1374_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 15120 0 1 10976
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _1375_
timestamp 1698431365
transform 1 0 13552 0 -1 9408
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _1376_
timestamp 1698431365
transform 1 0 14784 0 1 7840
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _1377_
timestamp 1698431365
transform 1 0 16240 0 1 6272
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _1378_
timestamp 1698431365
transform 1 0 16464 0 1 12544
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _1379_
timestamp 1698431365
transform 1 0 19712 0 -1 14112
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _1380_
timestamp 1698431365
transform 1 0 18480 0 -1 10976
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _1381_
timestamp 1698431365
transform 1 0 19152 0 -1 9408
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1382_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 25088 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1383_
timestamp 1698431365
transform 1 0 23072 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1384_
timestamp 1698431365
transform 1 0 21616 0 -1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1385_
timestamp 1698431365
transform 1 0 25760 0 -1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1386_
timestamp 1698431365
transform 1 0 21952 0 1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1387_
timestamp 1698431365
transform 1 0 25536 0 1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1388_
timestamp 1698431365
transform 1 0 21616 0 -1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1389_
timestamp 1698431365
transform 1 0 22400 0 1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1390_
timestamp 1698431365
transform 1 0 29344 0 -1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1391_
timestamp 1698431365
transform 1 0 33376 0 1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1392_
timestamp 1698431365
transform 1 0 29456 0 -1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1393_
timestamp 1698431365
transform 1 0 28224 0 -1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1394_
timestamp 1698431365
transform 1 0 34048 0 -1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1395_
timestamp 1698431365
transform 1 0 33152 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1396_
timestamp 1698431365
transform 1 0 30240 0 1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1397_
timestamp 1698431365
transform 1 0 34384 0 -1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1398_
timestamp 1698431365
transform 1 0 27776 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1399_
timestamp 1698431365
transform 1 0 24080 0 1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1400_
timestamp 1698431365
transform 1 0 26992 0 -1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1401_
timestamp 1698431365
transform 1 0 24192 0 1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1402_
timestamp 1698431365
transform 1 0 17248 0 -1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1403_
timestamp 1698431365
transform 1 0 20496 0 -1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1404_
timestamp 1698431365
transform 1 0 16352 0 1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1405_
timestamp 1698431365
transform 1 0 20160 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1406_
timestamp 1698431365
transform 1 0 18928 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1407_
timestamp 1698431365
transform 1 0 18368 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1408_
timestamp 1698431365
transform 1 0 21616 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1409_
timestamp 1698431365
transform 1 0 21952 0 1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1410_
timestamp 1698431365
transform 1 0 26208 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1411_
timestamp 1698431365
transform 1 0 29456 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1412_
timestamp 1698431365
transform 1 0 27552 0 -1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1413_
timestamp 1698431365
transform 1 0 30576 0 1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1414_
timestamp 1698431365
transform 1 0 34944 0 -1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1415_
timestamp 1698431365
transform 1 0 33376 0 1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1416_
timestamp 1698431365
transform 1 0 31584 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1417_
timestamp 1698431365
transform 1 0 32256 0 1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1418_
timestamp 1698431365
transform 1 0 25200 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1419_
timestamp 1698431365
transform 1 0 28560 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1420_
timestamp 1698431365
transform 1 0 24752 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1421_
timestamp 1698431365
transform 1 0 29008 0 1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1422_
timestamp 1698431365
transform 1 0 39312 0 1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1423_
timestamp 1698431365
transform 1 0 41888 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1424_
timestamp 1698431365
transform 1 0 42000 0 -1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1425_
timestamp 1698431365
transform 1 0 38864 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1426_
timestamp 1698431365
transform 1 0 37296 0 -1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1427_
timestamp 1698431365
transform 1 0 41216 0 -1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1428_
timestamp 1698431365
transform 1 0 37296 0 -1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1429_
timestamp 1698431365
transform 1 0 41216 0 1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1430_
timestamp 1698431365
transform 1 0 40768 0 -1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1431_
timestamp 1698431365
transform 1 0 37072 0 1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _1432_
timestamp 1698431365
transform 1 0 9408 0 -1 9408
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _1433_
timestamp 1698431365
transform 1 0 9408 0 -1 10976
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _1434_
timestamp 1698431365
transform 1 0 8848 0 1 10976
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _1435_
timestamp 1698431365
transform 1 0 12432 0 -1 12544
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _1436_
timestamp 1698431365
transform 1 0 10416 0 -1 7840
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _1437_
timestamp 1698431365
transform 1 0 9968 0 -1 6272
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _1438_
timestamp 1698431365
transform 1 0 10864 0 -1 4704
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _1439_
timestamp 1698431365
transform 1 0 14224 0 1 4704
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1456_
timestamp 1698431365
transform -1 0 3248 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1457_
timestamp 1698431365
transform -1 0 2576 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1458_
timestamp 1698431365
transform -1 0 2576 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1459_
timestamp 1698431365
transform -1 0 3920 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1460_
timestamp 1698431365
transform -1 0 2576 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1461_
timestamp 1698431365
transform -1 0 3248 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1462_
timestamp 1698431365
transform -1 0 3920 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1463_
timestamp 1698431365
transform -1 0 3360 0 -1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1464_
timestamp 1698431365
transform -1 0 4032 0 -1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1465_
timestamp 1698431365
transform 1 0 2688 0 1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1466_
timestamp 1698431365
transform -1 0 4032 0 1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1467_
timestamp 1698431365
transform -1 0 2576 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1468_
timestamp 1698431365
transform 1 0 3248 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1469_
timestamp 1698431365
transform -1 0 5152 0 1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1470_
timestamp 1698431365
transform -1 0 2576 0 -1 59584
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1471_
timestamp 1698431365
transform -1 0 3248 0 -1 59584
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1472_
timestamp 1698431365
transform -1 0 2576 0 1 61152
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1473_
timestamp 1698431365
transform -1 0 3920 0 1 61152
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1474_
timestamp 1698431365
transform 1 0 2688 0 -1 64288
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1475_
timestamp 1698431365
transform 1 0 3360 0 -1 64288
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1476_
timestamp 1698431365
transform -1 0 5152 0 1 64288
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1477_
timestamp 1698431365
transform -1 0 2576 0 -1 67424
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1478_
timestamp 1698431365
transform -1 0 3920 0 -1 67424
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1479_
timestamp 1698431365
transform -1 0 2576 0 1 68992
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1480_
timestamp 1698431365
transform -1 0 3248 0 1 68992
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1481_
timestamp 1698431365
transform 1 0 2688 0 -1 72128
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1482_
timestamp 1698431365
transform -1 0 4032 0 -1 72128
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1483_
timestamp 1698431365
transform -1 0 5152 0 -1 73696
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1484_
timestamp 1698431365
transform -1 0 5152 0 1 73696
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1485_
timestamp 1698431365
transform -1 0 5152 0 -1 75264
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1486_
timestamp 1698431365
transform -1 0 5152 0 1 75264
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1487_
timestamp 1698431365
transform -1 0 5152 0 -1 76832
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0666__I dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 25984 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0674__I
timestamp 1698431365
transform 1 0 41440 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0678__I
timestamp 1698431365
transform 1 0 44240 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0681__A2
timestamp 1698431365
transform -1 0 34272 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0689__A1
timestamp 1698431365
transform -1 0 45584 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0689__A3
timestamp 1698431365
transform 1 0 46592 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0690__A1
timestamp 1698431365
transform -1 0 46256 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0690__B
timestamp 1698431365
transform 1 0 42784 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0692__A1
timestamp 1698431365
transform 1 0 40992 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0694__A2
timestamp 1698431365
transform 1 0 46816 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0696__I
timestamp 1698431365
transform -1 0 70336 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0697__I
timestamp 1698431365
transform 1 0 71680 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0699__I
timestamp 1698431365
transform 1 0 52080 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0700__I
timestamp 1698431365
transform 1 0 50960 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0701__I
timestamp 1698431365
transform -1 0 46032 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0702__A1
timestamp 1698431365
transform -1 0 71120 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0702__A2
timestamp 1698431365
transform 1 0 70672 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0702__A3
timestamp 1698431365
transform 1 0 70224 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0702__A4
timestamp 1698431365
transform -1 0 70672 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0707__I
timestamp 1698431365
transform 1 0 70000 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0708__I
timestamp 1698431365
transform 1 0 69104 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0711__A1
timestamp 1698431365
transform -1 0 56224 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0713__A1
timestamp 1698431365
transform 1 0 54880 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0715__A1
timestamp 1698431365
transform 1 0 56224 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0717__A1
timestamp 1698431365
transform 1 0 57120 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0720__I
timestamp 1698431365
transform -1 0 72464 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0723__A1
timestamp 1698431365
transform -1 0 74592 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0723__A2
timestamp 1698431365
transform 1 0 76272 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0725__A1
timestamp 1698431365
transform 1 0 75488 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0725__A2
timestamp 1698431365
transform 1 0 75600 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0727__A1
timestamp 1698431365
transform 1 0 76272 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0727__A2
timestamp 1698431365
transform 1 0 77168 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0729__A1
timestamp 1698431365
transform -1 0 73696 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0729__A2
timestamp 1698431365
transform 1 0 78176 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0736__I
timestamp 1698431365
transform 1 0 75152 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0738__A1
timestamp 1698431365
transform 1 0 76272 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0740__I
timestamp 1698431365
transform 1 0 62944 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0742__A1
timestamp 1698431365
transform 1 0 61488 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0743__B
timestamp 1698431365
transform 1 0 73248 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0744__I
timestamp 1698431365
transform -1 0 40544 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0746__I
timestamp 1698431365
transform -1 0 32256 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0747__I
timestamp 1698431365
transform 1 0 44240 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0751__A1
timestamp 1698431365
transform -1 0 33824 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0756__A2
timestamp 1698431365
transform 1 0 34720 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0760__A1
timestamp 1698431365
transform -1 0 71456 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0761__A1
timestamp 1698431365
transform 1 0 60928 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0762__B
timestamp 1698431365
transform -1 0 74256 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0763__I
timestamp 1698431365
transform -1 0 34608 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0765__A1
timestamp 1698431365
transform -1 0 35056 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0766__A2
timestamp 1698431365
transform 1 0 36624 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0772__A1
timestamp 1698431365
transform 1 0 62608 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0773__B
timestamp 1698431365
transform -1 0 72240 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0774__I
timestamp 1698431365
transform -1 0 32704 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0776__A1
timestamp 1698431365
transform -1 0 34384 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0777__A2
timestamp 1698431365
transform -1 0 35280 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0784__A1
timestamp 1698431365
transform -1 0 62384 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0785__B
timestamp 1698431365
transform 1 0 71680 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0786__I
timestamp 1698431365
transform 1 0 33152 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0788__A1
timestamp 1698431365
transform -1 0 34272 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0789__A2
timestamp 1698431365
transform 1 0 37072 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0793__A1
timestamp 1698431365
transform 1 0 72576 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0797__A1
timestamp 1698431365
transform -1 0 62496 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0798__A1
timestamp 1698431365
transform -1 0 64064 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0800__I
timestamp 1698431365
transform 1 0 34272 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0803__A1
timestamp 1698431365
transform -1 0 35728 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0806__A2
timestamp 1698431365
transform -1 0 37632 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0807__A1
timestamp 1698431365
transform 1 0 35504 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0809__A1
timestamp 1698431365
transform -1 0 72128 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0811__A1
timestamp 1698431365
transform 1 0 63616 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0813__I
timestamp 1698431365
transform 1 0 33376 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0815__A1
timestamp 1698431365
transform 1 0 44016 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0816__A2
timestamp 1698431365
transform 1 0 39424 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0817__A1
timestamp 1698431365
transform 1 0 35056 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0819__I
timestamp 1698431365
transform 1 0 71008 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0821__A1
timestamp 1698431365
transform -1 0 71008 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0823__A1
timestamp 1698431365
transform 1 0 64512 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0824__B
timestamp 1698431365
transform 1 0 72352 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0825__I
timestamp 1698431365
transform 1 0 33824 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0827__A1
timestamp 1698431365
transform -1 0 34832 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0828__A2
timestamp 1698431365
transform 1 0 39872 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0829__A1
timestamp 1698431365
transform 1 0 34832 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0832__A1
timestamp 1698431365
transform -1 0 71904 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0835__A1
timestamp 1698431365
transform 1 0 67872 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0836__B
timestamp 1698431365
transform -1 0 70784 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0837__I
timestamp 1698431365
transform 1 0 36176 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0839__A1
timestamp 1698431365
transform -1 0 43456 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0840__A2
timestamp 1698431365
transform -1 0 37744 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0844__A1
timestamp 1698431365
transform -1 0 72800 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0848__A1
timestamp 1698431365
transform 1 0 65296 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0849__B
timestamp 1698431365
transform -1 0 71008 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0851__I
timestamp 1698431365
transform -1 0 37296 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0854__A1
timestamp 1698431365
transform -1 0 41216 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0857__A2
timestamp 1698431365
transform 1 0 40320 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0858__A1
timestamp 1698431365
transform -1 0 40768 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0860__A1
timestamp 1698431365
transform 1 0 73696 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0862__A1
timestamp 1698431365
transform 1 0 67088 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0863__B
timestamp 1698431365
transform 1 0 70000 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0864__I
timestamp 1698431365
transform 1 0 38752 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0866__A1
timestamp 1698431365
transform -1 0 44016 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0867__A2
timestamp 1698431365
transform 1 0 40880 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0868__A1
timestamp 1698431365
transform -1 0 41664 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0871__A1
timestamp 1698431365
transform -1 0 72576 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0873__A1
timestamp 1698431365
transform 1 0 67424 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0874__B
timestamp 1698431365
transform 1 0 74032 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0875__I
timestamp 1698431365
transform 1 0 38304 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0877__A1
timestamp 1698431365
transform -1 0 45136 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0878__A2
timestamp 1698431365
transform 1 0 42560 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0879__A1
timestamp 1698431365
transform -1 0 41664 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0881__I
timestamp 1698431365
transform 1 0 73808 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0883__A1
timestamp 1698431365
transform -1 0 72912 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0885__I
timestamp 1698431365
transform 1 0 68096 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0887__A1
timestamp 1698431365
transform 1 0 67536 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0888__B
timestamp 1698431365
transform -1 0 72688 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0889__I
timestamp 1698431365
transform 1 0 38640 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0891__A1
timestamp 1698431365
transform -1 0 41216 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0892__A2
timestamp 1698431365
transform 1 0 42448 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0893__A1
timestamp 1698431365
transform -1 0 41216 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0896__A1
timestamp 1698431365
transform -1 0 72800 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0900__A1
timestamp 1698431365
transform 1 0 69552 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0901__B
timestamp 1698431365
transform -1 0 72240 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0903__I
timestamp 1698431365
transform -1 0 37296 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0906__A1
timestamp 1698431365
transform -1 0 42560 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0909__A2
timestamp 1698431365
transform 1 0 43792 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0910__A1
timestamp 1698431365
transform 1 0 48832 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0912__A1
timestamp 1698431365
transform 1 0 73696 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0914__A1
timestamp 1698431365
transform 1 0 69888 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0915__B
timestamp 1698431365
transform 1 0 71680 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0916__I
timestamp 1698431365
transform -1 0 36624 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0918__A1
timestamp 1698431365
transform 1 0 45808 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0919__A2
timestamp 1698431365
transform 1 0 44576 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0923__A1
timestamp 1698431365
transform -1 0 71904 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0925__A1
timestamp 1698431365
transform 1 0 69664 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0926__B
timestamp 1698431365
transform -1 0 71792 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0927__I
timestamp 1698431365
transform 1 0 37856 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0929__A1
timestamp 1698431365
transform -1 0 47936 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0930__A2
timestamp 1698431365
transform 1 0 47488 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0934__A1
timestamp 1698431365
transform -1 0 71792 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0937__A1
timestamp 1698431365
transform 1 0 71344 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0938__B
timestamp 1698431365
transform -1 0 74816 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0939__I
timestamp 1698431365
transform 1 0 36400 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0941__A1
timestamp 1698431365
transform -1 0 49392 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0942__A2
timestamp 1698431365
transform 1 0 48160 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0947__A1
timestamp 1698431365
transform -1 0 73472 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0948__I
timestamp 1698431365
transform 1 0 74256 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0951__I
timestamp 1698431365
transform 1 0 68768 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0953__A1
timestamp 1698431365
transform 1 0 72576 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0955__I
timestamp 1698431365
transform 1 0 45472 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0957__I
timestamp 1698431365
transform 1 0 50176 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0961__A1
timestamp 1698431365
transform 1 0 48832 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0966__A2
timestamp 1698431365
transform -1 0 46704 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0969__A1
timestamp 1698431365
transform -1 0 72016 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0971__A1
timestamp 1698431365
transform 1 0 72128 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0973__I
timestamp 1698431365
transform 1 0 49280 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0975__A1
timestamp 1698431365
transform 1 0 50400 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0976__A2
timestamp 1698431365
transform -1 0 46368 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0980__A1
timestamp 1698431365
transform -1 0 72240 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0982__A1
timestamp 1698431365
transform 1 0 71792 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0984__I
timestamp 1698431365
transform 1 0 48272 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0986__A1
timestamp 1698431365
transform -1 0 49952 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0987__A2
timestamp 1698431365
transform 1 0 48048 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0988__A1
timestamp 1698431365
transform 1 0 48832 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0991__A1
timestamp 1698431365
transform -1 0 74480 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0994__A1
timestamp 1698431365
transform 1 0 73024 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0996__I
timestamp 1698431365
transform 1 0 48720 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0998__A1
timestamp 1698431365
transform 1 0 49616 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0999__A2
timestamp 1698431365
transform 1 0 48496 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1003__A1
timestamp 1698431365
transform -1 0 77056 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1007__A1
timestamp 1698431365
transform -1 0 72688 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1010__I
timestamp 1698431365
transform 1 0 47936 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1013__A1
timestamp 1698431365
transform -1 0 50624 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1016__A2
timestamp 1698431365
transform 1 0 50176 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1017__A1
timestamp 1698431365
transform 1 0 51632 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1019__A1
timestamp 1698431365
transform -1 0 71456 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1021__A1
timestamp 1698431365
transform 1 0 73808 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1023__I
timestamp 1698431365
transform -1 0 44464 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1025__A1
timestamp 1698431365
transform -1 0 50176 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1026__A2
timestamp 1698431365
transform 1 0 50848 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1027__A1
timestamp 1698431365
transform 1 0 52080 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1029__I
timestamp 1698431365
transform 1 0 73472 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1030__A1
timestamp 1698431365
transform -1 0 73584 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1032__A1
timestamp 1698431365
transform -1 0 72240 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1034__I
timestamp 1698431365
transform 1 0 45360 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1036__A1
timestamp 1698431365
transform 1 0 50288 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1037__A2
timestamp 1698431365
transform 1 0 51072 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1038__A1
timestamp 1698431365
transform 1 0 52416 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1041__A1
timestamp 1698431365
transform -1 0 71680 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1044__A1
timestamp 1698431365
transform -1 0 71792 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1046__I
timestamp 1698431365
transform 1 0 44576 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1048__A1
timestamp 1698431365
transform 1 0 50736 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1049__A2
timestamp 1698431365
transform 1 0 51744 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1050__A1
timestamp 1698431365
transform -1 0 51520 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1053__A1
timestamp 1698431365
transform -1 0 71904 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1057__A1
timestamp 1698431365
transform 1 0 75264 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1060__I
timestamp 1698431365
transform -1 0 44912 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1063__A1
timestamp 1698431365
transform 1 0 51744 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1066__A2
timestamp 1698431365
transform 1 0 52080 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1069__A1
timestamp 1698431365
transform -1 0 75824 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1071__A1
timestamp 1698431365
transform -1 0 74480 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1073__I
timestamp 1698431365
transform 1 0 45360 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1075__A1
timestamp 1698431365
transform -1 0 52416 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1076__A2
timestamp 1698431365
transform 1 0 55776 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1077__B1
timestamp 1698431365
transform -1 0 51184 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1079__I
timestamp 1698431365
transform 1 0 72128 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1080__A1
timestamp 1698431365
transform -1 0 71456 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1082__A1
timestamp 1698431365
transform 1 0 78176 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1084__I
timestamp 1698431365
transform 1 0 44240 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1086__A1
timestamp 1698431365
transform -1 0 52864 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1087__A2
timestamp 1698431365
transform 1 0 53760 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1090__I
timestamp 1698431365
transform 1 0 73472 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1091__A1
timestamp 1698431365
transform 1 0 77056 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1093__I
timestamp 1698431365
transform -1 0 69104 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1094__A1
timestamp 1698431365
transform 1 0 78064 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1096__I
timestamp 1698431365
transform 1 0 45472 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1098__A1
timestamp 1698431365
transform 1 0 52752 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1099__A2
timestamp 1698431365
transform 1 0 54208 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1100__B1
timestamp 1698431365
transform 1 0 55104 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1103__A1
timestamp 1698431365
transform -1 0 78288 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1107__A1
timestamp 1698431365
transform 1 0 78176 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1110__I
timestamp 1698431365
transform 1 0 45696 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1113__A1
timestamp 1698431365
transform 1 0 54096 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1116__A2
timestamp 1698431365
transform 1 0 56672 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1117__A1
timestamp 1698431365
transform 1 0 56000 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1119__A1
timestamp 1698431365
transform -1 0 77392 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1121__A1
timestamp 1698431365
transform 1 0 77952 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1123__I
timestamp 1698431365
transform -1 0 44464 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1125__A1
timestamp 1698431365
transform 1 0 55328 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1126__A2
timestamp 1698431365
transform 1 0 56000 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1127__A1
timestamp 1698431365
transform 1 0 57344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1129__A1
timestamp 1698431365
transform -1 0 75824 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1131__A1
timestamp 1698431365
transform 1 0 76496 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1133__I
timestamp 1698431365
transform 1 0 44688 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1135__A1
timestamp 1698431365
transform -1 0 56896 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1136__A2
timestamp 1698431365
transform 1 0 55552 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1137__A1
timestamp 1698431365
transform 1 0 57120 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1137__B1
timestamp 1698431365
transform -1 0 56896 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1139__A1
timestamp 1698431365
transform 1 0 74592 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1141__A1
timestamp 1698431365
transform 1 0 73920 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1143__I
timestamp 1698431365
transform 1 0 45584 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1145__A1
timestamp 1698431365
transform -1 0 55104 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1146__A2
timestamp 1698431365
transform 1 0 57120 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1147__A1
timestamp 1698431365
transform 1 0 56672 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1147__B1
timestamp 1698431365
transform 1 0 57120 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1148__A1
timestamp 1698431365
transform 1 0 43232 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1149__A1
timestamp 1698431365
transform 1 0 41440 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1150__A1
timestamp 1698431365
transform 1 0 43680 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1151__A1
timestamp 1698431365
transform 1 0 48832 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1152__A1
timestamp 1698431365
transform -1 0 74816 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1156__A1
timestamp 1698431365
transform -1 0 28672 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1160__A1
timestamp 1698431365
transform -1 0 26432 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1162__I
timestamp 1698431365
transform 1 0 20720 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1163__I
timestamp 1698431365
transform -1 0 18032 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1164__A1
timestamp 1698431365
transform 1 0 18480 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1167__A1
timestamp 1698431365
transform -1 0 17024 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1170__A1
timestamp 1698431365
transform -1 0 16576 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1173__A1
timestamp 1698431365
transform -1 0 18928 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1178__I
timestamp 1698431365
transform -1 0 19712 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1179__A1
timestamp 1698431365
transform 1 0 18592 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1182__A1
timestamp 1698431365
transform 1 0 21392 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1185__A1
timestamp 1698431365
transform 1 0 20720 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1188__A1
timestamp 1698431365
transform -1 0 19488 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1190__A1
timestamp 1698431365
transform 1 0 25760 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1193__A1
timestamp 1698431365
transform -1 0 24864 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1195__I
timestamp 1698431365
transform 1 0 25312 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1210__I
timestamp 1698431365
transform -1 0 13104 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1211__I
timestamp 1698431365
transform 1 0 24640 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1223__A1
timestamp 1698431365
transform -1 0 25536 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1226__A1
timestamp 1698431365
transform -1 0 30912 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1228__I
timestamp 1698431365
transform 1 0 31808 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1243__I
timestamp 1698431365
transform 1 0 31136 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1255__A1
timestamp 1698431365
transform 1 0 29904 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1260__A1
timestamp 1698431365
transform 1 0 24528 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1262__A1
timestamp 1698431365
transform 1 0 23632 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1264__A1
timestamp 1698431365
transform 1 0 23296 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1266__A1
timestamp 1698431365
transform 1 0 23520 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1270__A1
timestamp 1698431365
transform 1 0 17136 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1271__A1
timestamp 1698431365
transform -1 0 18480 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1272__A1
timestamp 1698431365
transform 1 0 19376 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1273__A1
timestamp 1698431365
transform 1 0 22288 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1274__A1
timestamp 1698431365
transform 1 0 16800 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1275__A1
timestamp 1698431365
transform 1 0 18368 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1276__A1
timestamp 1698431365
transform 1 0 19152 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1280__A1
timestamp 1698431365
transform 1 0 18592 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1281__A1
timestamp 1698431365
transform 1 0 20608 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1282__A1
timestamp 1698431365
transform 1 0 18704 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1283__A1
timestamp 1698431365
transform 1 0 21392 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1284__A1
timestamp 1698431365
transform 1 0 17584 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1285__A1
timestamp 1698431365
transform 1 0 22736 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1286__A1
timestamp 1698431365
transform 1 0 18816 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1287__A1
timestamp 1698431365
transform -1 0 21840 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1290__A1
timestamp 1698431365
transform 1 0 24416 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1291__A1
timestamp 1698431365
transform 1 0 28112 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1292__A1
timestamp 1698431365
transform 1 0 26880 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1294__A1
timestamp 1698431365
transform 1 0 25648 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1296__A1
timestamp 1698431365
transform 1 0 27888 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1307__A1
timestamp 1698431365
transform 1 0 34048 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1313__A1
timestamp 1698431365
transform -1 0 25648 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1315__A1
timestamp 1698431365
transform 1 0 29232 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1317__A1
timestamp 1698431365
transform -1 0 26096 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1319__A1
timestamp 1698431365
transform 1 0 30800 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1333__A1
timestamp 1698431365
transform -1 0 40432 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1335__A1
timestamp 1698431365
transform -1 0 45696 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1337__A1
timestamp 1698431365
transform 1 0 41552 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1339__A1
timestamp 1698431365
transform -1 0 46144 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1340__S
timestamp 1698431365
transform -1 0 35952 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1342__A1
timestamp 1698431365
transform 1 0 30352 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1343__I
timestamp 1698431365
transform -1 0 9968 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1345__A1
timestamp 1698431365
transform -1 0 27888 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1347__I
timestamp 1698431365
transform -1 0 14224 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1348__A1
timestamp 1698431365
transform 1 0 10976 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1351__A1
timestamp 1698431365
transform 1 0 12768 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1354__A1
timestamp 1698431365
transform 1 0 12432 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1357__A1
timestamp 1698431365
transform 1 0 14448 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1359__I
timestamp 1698431365
transform -1 0 7504 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1362__I
timestamp 1698431365
transform -1 0 16128 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1363__A1
timestamp 1698431365
transform 1 0 11424 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1366__A1
timestamp 1698431365
transform -1 0 8400 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1369__A1
timestamp 1698431365
transform -1 0 7952 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1372__A1
timestamp 1698431365
transform -1 0 9968 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1411__CLK
timestamp 1698431365
transform 1 0 32704 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1414__CLK
timestamp 1698431365
transform -1 0 38416 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1416__CLK
timestamp 1698431365
transform -1 0 35280 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1417__CLK
timestamp 1698431365
transform 1 0 35392 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1430__CLK
timestamp 1698431365
transform 1 0 40320 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1471__I
timestamp 1698431365
transform 1 0 3472 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_clk_I
timestamp 1698431365
transform 1 0 31248 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_0__f_clk_I
timestamp 1698431365
transform -1 0 20944 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_1__f_clk_I
timestamp 1698431365
transform -1 0 27888 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_2__f_clk_I
timestamp 1698431365
transform -1 0 27552 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_3__f_clk_I
timestamp 1698431365
transform 1 0 28560 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_4__f_clk_I
timestamp 1698431365
transform 1 0 32480 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_5__f_clk_I
timestamp 1698431365
transform 1 0 38304 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_6__f_clk_I
timestamp 1698431365
transform 1 0 28560 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_3_7__f_clk_I
timestamp 1698431365
transform 1 0 33376 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout331_I
timestamp 1698431365
transform -1 0 4368 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout332_I
timestamp 1698431365
transform 1 0 4480 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout334_I
timestamp 1698431365
transform -1 0 2016 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout335_I
timestamp 1698431365
transform 1 0 4928 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout336_I
timestamp 1698431365
transform -1 0 4368 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout338_I
timestamp 1698431365
transform 1 0 2912 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout341_I
timestamp 1698431365
transform -1 0 2016 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout342_I
timestamp 1698431365
transform 1 0 5376 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input1_I
timestamp 1698431365
transform -1 0 24752 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input2_I
timestamp 1698431365
transform -1 0 31808 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input3_I
timestamp 1698431365
transform -1 0 26768 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input4_I
timestamp 1698431365
transform -1 0 21616 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input5_I
timestamp 1698431365
transform -1 0 21056 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input6_I
timestamp 1698431365
transform -1 0 33936 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input7_I
timestamp 1698431365
transform -1 0 25200 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input8_I
timestamp 1698431365
transform -1 0 20944 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input9_I
timestamp 1698431365
transform -1 0 32704 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input10_I
timestamp 1698431365
transform -1 0 31920 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input11_I
timestamp 1698431365
transform -1 0 34384 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input12_I
timestamp 1698431365
transform -1 0 20048 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input13_I
timestamp 1698431365
transform 1 0 40992 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input14_I
timestamp 1698431365
transform 1 0 50176 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input15_I
timestamp 1698431365
transform -1 0 32480 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input16_I
timestamp 1698431365
transform -1 0 48160 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input17_I
timestamp 1698431365
transform 1 0 49056 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input18_I
timestamp 1698431365
transform -1 0 42336 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input19_I
timestamp 1698431365
transform 1 0 51744 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input20_I
timestamp 1698431365
transform 1 0 51408 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input21_I
timestamp 1698431365
transform 1 0 46256 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input22_I
timestamp 1698431365
transform -1 0 47600 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input23_I
timestamp 1698431365
transform -1 0 18480 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input24_I
timestamp 1698431365
transform 1 0 50848 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input25_I
timestamp 1698431365
transform 1 0 51296 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input26_I
timestamp 1698431365
transform -1 0 24416 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input27_I
timestamp 1698431365
transform -1 0 29792 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input28_I
timestamp 1698431365
transform -1 0 23632 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input29_I
timestamp 1698431365
transform -1 0 19600 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input30_I
timestamp 1698431365
transform -1 0 21616 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input31_I
timestamp 1698431365
transform -1 0 23632 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input32_I
timestamp 1698431365
transform -1 0 22064 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input33_I
timestamp 1698431365
transform 1 0 49728 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input34_I
timestamp 1698431365
transform -1 0 3808 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input35_I
timestamp 1698431365
transform -1 0 8512 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input36_I
timestamp 1698431365
transform -1 0 7504 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input37_I
timestamp 1698431365
transform 1 0 14448 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input38_I
timestamp 1698431365
transform -1 0 6272 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input39_I
timestamp 1698431365
transform -1 0 7952 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input40_I
timestamp 1698431365
transform -1 0 10752 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input41_I
timestamp 1698431365
transform -1 0 15680 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input42_I
timestamp 1698431365
transform -1 0 10416 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input43_I
timestamp 1698431365
transform -1 0 15232 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input44_I
timestamp 1698431365
transform -1 0 14112 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input45_I
timestamp 1698431365
transform -1 0 5264 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input46_I
timestamp 1698431365
transform -1 0 12656 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input47_I
timestamp 1698431365
transform -1 0 15344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input48_I
timestamp 1698431365
transform -1 0 12208 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input49_I
timestamp 1698431365
transform -1 0 16576 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input50_I
timestamp 1698431365
transform -1 0 13104 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input51_I
timestamp 1698431365
transform -1 0 15792 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input52_I
timestamp 1698431365
transform -1 0 19376 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input53_I
timestamp 1698431365
transform -1 0 14560 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input54_I
timestamp 1698431365
transform -1 0 17024 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input55_I
timestamp 1698431365
transform -1 0 23072 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input56_I
timestamp 1698431365
transform -1 0 4816 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input57_I
timestamp 1698431365
transform -1 0 16240 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input58_I
timestamp 1698431365
transform -1 0 20496 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input59_I
timestamp 1698431365
transform -1 0 6720 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input60_I
timestamp 1698431365
transform -1 0 5712 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input61_I
timestamp 1698431365
transform -1 0 6272 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input62_I
timestamp 1698431365
transform -1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input63_I
timestamp 1698431365
transform -1 0 7168 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input64_I
timestamp 1698431365
transform -1 0 8064 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input65_I
timestamp 1698431365
transform -1 0 7616 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input66_I
timestamp 1698431365
transform 1 0 52752 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input67_I
timestamp 1698431365
transform 1 0 52528 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input68_I
timestamp 1698431365
transform 1 0 54208 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input69_I
timestamp 1698431365
transform -1 0 53424 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input70_I
timestamp 1698431365
transform -1 0 2240 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input71_I
timestamp 1698431365
transform 1 0 2464 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input72_I
timestamp 1698431365
transform 1 0 2464 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input73_I
timestamp 1698431365
transform 1 0 2464 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input74_I
timestamp 1698431365
transform 1 0 2464 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input75_I
timestamp 1698431365
transform 1 0 2464 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input76_I
timestamp 1698431365
transform 1 0 2464 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input77_I
timestamp 1698431365
transform 1 0 2464 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input78_I
timestamp 1698431365
transform 1 0 2464 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input79_I
timestamp 1698431365
transform 1 0 2464 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input80_I
timestamp 1698431365
transform 1 0 2464 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input81_I
timestamp 1698431365
transform 1 0 3136 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input82_I
timestamp 1698431365
transform 1 0 2464 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input83_I
timestamp 1698431365
transform 1 0 2464 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input84_I
timestamp 1698431365
transform 1 0 2464 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input85_I
timestamp 1698431365
transform 1 0 2464 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input86_I
timestamp 1698431365
transform 1 0 2464 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input87_I
timestamp 1698431365
transform 1 0 2464 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input88_I
timestamp 1698431365
transform 1 0 2464 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input89_I
timestamp 1698431365
transform 1 0 2464 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input90_I
timestamp 1698431365
transform 1 0 2464 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input91_I
timestamp 1698431365
transform 1 0 2464 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input92_I
timestamp 1698431365
transform 1 0 2464 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input93_I
timestamp 1698431365
transform 1 0 2464 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input94_I
timestamp 1698431365
transform 1 0 2464 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input95_I
timestamp 1698431365
transform 1 0 2464 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input96_I
timestamp 1698431365
transform 1 0 2464 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input97_I
timestamp 1698431365
transform 1 0 2464 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input98_I
timestamp 1698431365
transform 1 0 2464 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input99_I
timestamp 1698431365
transform 1 0 2464 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input100_I
timestamp 1698431365
transform 1 0 2464 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input101_I
timestamp 1698431365
transform 1 0 2464 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input102_I
timestamp 1698431365
transform -1 0 75824 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input103_I
timestamp 1698431365
transform -1 0 77728 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input104_I
timestamp 1698431365
transform -1 0 77728 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input105_I
timestamp 1698431365
transform -1 0 77728 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input106_I
timestamp 1698431365
transform -1 0 77728 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input107_I
timestamp 1698431365
transform -1 0 77728 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input108_I
timestamp 1698431365
transform -1 0 77504 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input109_I
timestamp 1698431365
transform -1 0 77728 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input110_I
timestamp 1698431365
transform -1 0 77504 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input111_I
timestamp 1698431365
transform -1 0 77728 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input112_I
timestamp 1698431365
transform -1 0 77504 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input113_I
timestamp 1698431365
transform -1 0 77504 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input114_I
timestamp 1698431365
transform -1 0 77728 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input115_I
timestamp 1698431365
transform -1 0 77728 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input116_I
timestamp 1698431365
transform -1 0 77728 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input117_I
timestamp 1698431365
transform -1 0 77504 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input118_I
timestamp 1698431365
transform -1 0 77728 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input119_I
timestamp 1698431365
transform -1 0 77504 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input120_I
timestamp 1698431365
transform -1 0 77728 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input121_I
timestamp 1698431365
transform -1 0 77728 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input122_I
timestamp 1698431365
transform -1 0 75376 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input123_I
timestamp 1698431365
transform -1 0 77728 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input124_I
timestamp 1698431365
transform -1 0 74144 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input125_I
timestamp 1698431365
transform -1 0 77728 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input126_I
timestamp 1698431365
transform -1 0 77280 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input127_I
timestamp 1698431365
transform 1 0 78176 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input128_I
timestamp 1698431365
transform -1 0 77728 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input129_I
timestamp 1698431365
transform -1 0 77728 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input130_I
timestamp 1698431365
transform -1 0 77728 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input131_I
timestamp 1698431365
transform -1 0 77728 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input132_I
timestamp 1698431365
transform -1 0 77728 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input133_I
timestamp 1698431365
transform -1 0 77728 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input134_I
timestamp 1698431365
transform -1 0 77728 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input135_I
timestamp 1698431365
transform -1 0 74592 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input136_I
timestamp 1698431365
transform -1 0 75376 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input137_I
timestamp 1698431365
transform -1 0 77728 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input138_I
timestamp 1698431365
transform -1 0 77728 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input139_I
timestamp 1698431365
transform -1 0 77056 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input140_I
timestamp 1698431365
transform -1 0 76608 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input141_I
timestamp 1698431365
transform -1 0 74704 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input142_I
timestamp 1698431365
transform -1 0 78400 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input143_I
timestamp 1698431365
transform -1 0 77728 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input144_I
timestamp 1698431365
transform -1 0 74480 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input145_I
timestamp 1698431365
transform -1 0 74704 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input146_I
timestamp 1698431365
transform -1 0 78400 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input147_I
timestamp 1698431365
transform -1 0 78400 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input148_I
timestamp 1698431365
transform -1 0 72464 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input149_I
timestamp 1698431365
transform -1 0 73024 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input150_I
timestamp 1698431365
transform -1 0 76608 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input151_I
timestamp 1698431365
transform -1 0 71344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input152_I
timestamp 1698431365
transform -1 0 71008 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input153_I
timestamp 1698431365
transform -1 0 75376 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input154_I
timestamp 1698431365
transform -1 0 71008 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input155_I
timestamp 1698431365
transform -1 0 77728 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input156_I
timestamp 1698431365
transform -1 0 71344 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input157_I
timestamp 1698431365
transform -1 0 71232 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input158_I
timestamp 1698431365
transform -1 0 77056 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input159_I
timestamp 1698431365
transform -1 0 78400 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input160_I
timestamp 1698431365
transform -1 0 76048 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input161_I
timestamp 1698431365
transform -1 0 76944 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input162_I
timestamp 1698431365
transform -1 0 77728 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input163_I
timestamp 1698431365
transform -1 0 77056 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input164_I
timestamp 1698431365
transform -1 0 76608 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input165_I
timestamp 1698431365
transform -1 0 77728 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input166_I
timestamp 1698431365
transform -1 0 77728 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input167_I
timestamp 1698431365
transform -1 0 77728 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input168_I
timestamp 1698431365
transform 1 0 34608 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input169_I
timestamp 1698431365
transform 1 0 42000 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input170_I
timestamp 1698431365
transform -1 0 41552 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input171_I
timestamp 1698431365
transform 1 0 42448 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input172_I
timestamp 1698431365
transform -1 0 43456 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input173_I
timestamp 1698431365
transform -1 0 44016 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input174_I
timestamp 1698431365
transform 1 0 46032 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input175_I
timestamp 1698431365
transform -1 0 44464 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input176_I
timestamp 1698431365
transform -1 0 46704 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input177_I
timestamp 1698431365
transform 1 0 48048 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input178_I
timestamp 1698431365
transform -1 0 46928 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input179_I
timestamp 1698431365
transform 1 0 35504 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input180_I
timestamp 1698431365
transform 1 0 48496 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input181_I
timestamp 1698431365
transform -1 0 49168 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input182_I
timestamp 1698431365
transform 1 0 50736 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input183_I
timestamp 1698431365
transform -1 0 49616 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input184_I
timestamp 1698431365
transform 1 0 51184 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input185_I
timestamp 1698431365
transform -1 0 51856 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input186_I
timestamp 1698431365
transform -1 0 52864 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input187_I
timestamp 1698431365
transform -1 0 52304 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input188_I
timestamp 1698431365
transform 1 0 55104 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input189_I
timestamp 1698431365
transform -1 0 53648 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input190_I
timestamp 1698431365
transform 1 0 35952 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input191_I
timestamp 1698431365
transform -1 0 54544 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input192_I
timestamp 1698431365
transform -1 0 55440 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input193_I
timestamp 1698431365
transform 1 0 36736 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input194_I
timestamp 1698431365
transform 1 0 37632 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input195_I
timestamp 1698431365
transform 1 0 38192 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input196_I
timestamp 1698431365
transform -1 0 37296 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input197_I
timestamp 1698431365
transform -1 0 38864 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input198_I
timestamp 1698431365
transform 1 0 39424 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input199_I
timestamp 1698431365
transform 1 0 40880 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input200_I
timestamp 1698431365
transform -1 0 32816 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input201_I
timestamp 1698431365
transform -1 0 59248 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input202_I
timestamp 1698431365
transform -1 0 65072 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input203_I
timestamp 1698431365
transform 1 0 66416 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input204_I
timestamp 1698431365
transform -1 0 67088 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input205_I
timestamp 1698431365
transform -1 0 67648 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input206_I
timestamp 1698431365
transform 1 0 68432 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input207_I
timestamp 1698431365
transform -1 0 69216 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input208_I
timestamp 1698431365
transform -1 0 70112 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input209_I
timestamp 1698431365
transform -1 0 70784 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input210_I
timestamp 1698431365
transform -1 0 71456 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input211_I
timestamp 1698431365
transform -1 0 72016 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input212_I
timestamp 1698431365
transform 1 0 61264 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input213_I
timestamp 1698431365
transform 1 0 73360 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input214_I
timestamp 1698431365
transform -1 0 72464 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input215_I
timestamp 1698431365
transform -1 0 74032 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input216_I
timestamp 1698431365
transform -1 0 74592 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input217_I
timestamp 1698431365
transform -1 0 75152 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input218_I
timestamp 1698431365
transform -1 0 75824 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input219_I
timestamp 1698431365
transform -1 0 75040 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input220_I
timestamp 1698431365
transform -1 0 76720 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input221_I
timestamp 1698431365
transform -1 0 76272 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input222_I
timestamp 1698431365
transform -1 0 77280 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input223_I
timestamp 1698431365
transform 1 0 62832 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input224_I
timestamp 1698431365
transform -1 0 76496 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input225_I
timestamp 1698431365
transform -1 0 75488 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input226_I
timestamp 1698431365
transform 1 0 61712 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input227_I
timestamp 1698431365
transform 1 0 62160 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input228_I
timestamp 1698431365
transform 1 0 63280 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input229_I
timestamp 1698431365
transform 1 0 63728 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input230_I
timestamp 1698431365
transform 1 0 64176 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input231_I
timestamp 1698431365
transform -1 0 64736 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input232_I
timestamp 1698431365
transform 1 0 65968 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output233_I
timestamp 1698431365
transform 1 0 14336 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output234_I
timestamp 1698431365
transform -1 0 18032 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output235_I
timestamp 1698431365
transform 1 0 19824 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output236_I
timestamp 1698431365
transform 1 0 19376 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output237_I
timestamp 1698431365
transform 1 0 22960 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output238_I
timestamp 1698431365
transform 1 0 24752 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output239_I
timestamp 1698431365
transform 1 0 25200 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output240_I
timestamp 1698431365
transform 1 0 14112 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output241_I
timestamp 1698431365
transform 1 0 13552 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output242_I
timestamp 1698431365
transform -1 0 14336 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output243_I
timestamp 1698431365
transform -1 0 13440 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output244_I
timestamp 1698431365
transform -1 0 14112 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output245_I
timestamp 1698431365
transform -1 0 14784 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output246_I
timestamp 1698431365
transform 1 0 18032 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output247_I
timestamp 1698431365
transform -1 0 17248 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output248_I
timestamp 1698431365
transform 1 0 18256 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output249_I
timestamp 1698431365
transform 1 0 52528 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output250_I
timestamp 1698431365
transform 1 0 59472 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output251_I
timestamp 1698431365
transform -1 0 60144 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output252_I
timestamp 1698431365
transform -1 0 63280 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output253_I
timestamp 1698431365
transform 1 0 65632 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output254_I
timestamp 1698431365
transform 1 0 66416 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output255_I
timestamp 1698431365
transform -1 0 63280 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output256_I
timestamp 1698431365
transform 1 0 63840 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output257_I
timestamp 1698431365
transform 1 0 67424 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output258_I
timestamp 1698431365
transform -1 0 69888 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output259_I
timestamp 1698431365
transform -1 0 67200 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output260_I
timestamp 1698431365
transform 1 0 55888 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output261_I
timestamp 1698431365
transform 1 0 67312 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output262_I
timestamp 1698431365
transform 1 0 66640 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output263_I
timestamp 1698431365
transform -1 0 67984 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output264_I
timestamp 1698431365
transform -1 0 71120 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output265_I
timestamp 1698431365
transform 1 0 71680 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output266_I
timestamp 1698431365
transform 1 0 70448 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output267_I
timestamp 1698431365
transform -1 0 71120 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output268_I
timestamp 1698431365
transform 1 0 71680 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output269_I
timestamp 1698431365
transform 1 0 70448 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output270_I
timestamp 1698431365
transform 1 0 71680 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output271_I
timestamp 1698431365
transform -1 0 54096 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output272_I
timestamp 1698431365
transform -1 0 74480 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output273_I
timestamp 1698431365
transform 1 0 76272 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output274_I
timestamp 1698431365
transform 1 0 58016 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output275_I
timestamp 1698431365
transform 1 0 61824 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output276_I
timestamp 1698431365
transform 1 0 56784 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output277_I
timestamp 1698431365
transform 1 0 56000 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output278_I
timestamp 1698431365
transform 1 0 62496 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output279_I
timestamp 1698431365
transform 1 0 63504 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output280_I
timestamp 1698431365
transform 1 0 60144 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output281_I
timestamp 1698431365
transform 1 0 50400 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output283_I
timestamp 1698431365
transform 1 0 4704 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output284_I
timestamp 1698431365
transform 1 0 4704 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output285_I
timestamp 1698431365
transform 1 0 4704 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output324_I
timestamp 1698431365
transform 1 0 35056 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output325_I
timestamp 1698431365
transform 1 0 58464 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output326_I
timestamp 1698431365
transform 1 0 59472 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output327_I
timestamp 1698431365
transform -1 0 57680 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output328_I
timestamp 1698431365
transform 1 0 60816 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_clk dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 31248 0 -1 15680
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_0__f_clk
timestamp 1698431365
transform -1 0 20496 0 1 9408
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_1__f_clk
timestamp 1698431365
transform 1 0 21168 0 1 9408
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_2__f_clk
timestamp 1698431365
transform -1 0 24864 0 -1 20384
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_3__f_clk
timestamp 1698431365
transform -1 0 28336 0 1 17248
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_4__f_clk
timestamp 1698431365
transform -1 0 38528 0 -1 10976
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_5__f_clk
timestamp 1698431365
transform 1 0 38528 0 1 10976
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_6__f_clk
timestamp 1698431365
transform -1 0 35280 0 1 18816
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_3_7__f_clk
timestamp 1698431365
transform 1 0 34272 0 -1 18816
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout329
timestamp 1698431365
transform 1 0 2016 0 -1 64288
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout330
timestamp 1698431365
transform 1 0 2576 0 -1 67424
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout331
timestamp 1698431365
transform -1 0 3248 0 1 61152
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  fanout332
timestamp 1698431365
transform -1 0 4256 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout333
timestamp 1698431365
transform -1 0 3248 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout334
timestamp 1698431365
transform 1 0 2016 0 1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  fanout335
timestamp 1698431365
transform -1 0 3360 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout336
timestamp 1698431365
transform 1 0 2576 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout337
timestamp 1698431365
transform 1 0 2016 0 -1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  fanout338
timestamp 1698431365
transform -1 0 2688 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout339
timestamp 1698431365
transform -1 0 4704 0 -1 72128
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout340
timestamp 1698431365
transform -1 0 6048 0 -1 76832
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout341
timestamp 1698431365
transform 1 0 2016 0 -1 72128
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  fanout342
timestamp 1698431365
transform -1 0 2464 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_14 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 2912 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_18
timestamp 1698431365
transform 1 0 3360 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_36
timestamp 1698431365
transform 1 0 5376 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_70
timestamp 1698431365
transform 1 0 9184 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_104
timestamp 1698431365
transform 1 0 12992 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_138
timestamp 1698431365
transform 1 0 16800 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_172
timestamp 1698431365
transform 1 0 20608 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_206
timestamp 1698431365
transform 1 0 24416 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_216
timestamp 1698431365
transform 1 0 25536 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_240
timestamp 1698431365
transform 1 0 28224 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_470
timestamp 1698431365
transform 1 0 53984 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_474
timestamp 1698431365
transform 1 0 54432 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_504
timestamp 1698431365
transform 1 0 57792 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_508
timestamp 1698431365
transform 1 0 58240 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_538
timestamp 1698431365
transform 1 0 61600 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_542
timestamp 1698431365
transform 1 0 62048 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_572
timestamp 1698431365
transform 1 0 65408 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_576
timestamp 1698431365
transform 1 0 65856 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_606 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 69216 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_640
timestamp 1698431365
transform 1 0 73024 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_2
timestamp 1698431365
transform 1 0 1568 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_8 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 2240 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_24
timestamp 1698431365
transform 1 0 4032 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_28 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 4480 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_31
timestamp 1698431365
transform 1 0 4816 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_35
timestamp 1698431365
transform 1 0 5264 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_45
timestamp 1698431365
transform 1 0 6384 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_72
timestamp 1698431365
transform 1 0 9408 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_142
timestamp 1698431365
transform 1 0 17248 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_241
timestamp 1698431365
transform 1 0 28336 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_282
timestamp 1698431365
transform 1 0 32928 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_417
timestamp 1698431365
transform 1 0 48048 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_419
timestamp 1698431365
transform 1 0 48272 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_428
timestamp 1698431365
transform 1 0 49280 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_455
timestamp 1698431365
transform 1 0 52304 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_485
timestamp 1698431365
transform 1 0 55664 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_489
timestamp 1698431365
transform 1 0 56112 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_544
timestamp 1698431365
transform 1 0 62272 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_548
timestamp 1698431365
transform 1 0 62720 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_550
timestamp 1698431365
transform 1 0 62944 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_553
timestamp 1698431365
transform 1 0 63280 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_557
timestamp 1698431365
transform 1 0 63728 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_559
timestamp 1698431365
transform 1 0 63952 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_614
timestamp 1698431365
transform 1 0 70112 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_616
timestamp 1698431365
transform 1 0 70336 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_619
timestamp 1698431365
transform 1 0 70672 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_623
timestamp 1698431365
transform 1 0 71120 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_627
timestamp 1698431365
transform 1 0 71568 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_684
timestamp 1698431365
transform 1 0 77952 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_8
timestamp 1698431365
transform 1 0 2240 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_12
timestamp 1698431365
transform 1 0 2688 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_28
timestamp 1698431365
transform 1 0 4480 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_32
timestamp 1698431365
transform 1 0 4928 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_37
timestamp 1698431365
transform 1 0 5488 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_41
timestamp 1698431365
transform 1 0 5936 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_50
timestamp 1698431365
transform 1 0 6944 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_52
timestamp 1698431365
transform 1 0 7168 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_55
timestamp 1698431365
transform 1 0 7504 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_59
timestamp 1698431365
transform 1 0 7952 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_87
timestamp 1698431365
transform 1 0 11088 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_89
timestamp 1698431365
transform 1 0 11312 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_96
timestamp 1698431365
transform 1 0 12096 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_158
timestamp 1698431365
transform 1 0 19040 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_160
timestamp 1698431365
transform 1 0 19264 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_163
timestamp 1698431365
transform 1 0 19600 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_167
timestamp 1698431365
transform 1 0 20048 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_171
timestamp 1698431365
transform 1 0 20496 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_177
timestamp 1698431365
transform 1 0 21168 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_187
timestamp 1698431365
transform 1 0 22288 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_223
timestamp 1698431365
transform 1 0 26320 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_247
timestamp 1698431365
transform 1 0 29008 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_274
timestamp 1698431365
transform 1 0 32032 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_331
timestamp 1698431365
transform 1 0 38416 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_346
timestamp 1698431365
transform 1 0 40096 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_436
timestamp 1698431365
transform 1 0 50176 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_440
timestamp 1698431365
transform 1 0 50624 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_444
timestamp 1698431365
transform 1 0 51072 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_448
timestamp 1698431365
transform 1 0 51520 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_452
timestamp 1698431365
transform 1 0 51968 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_454
timestamp 1698431365
transform 1 0 52192 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_457
timestamp 1698431365
transform 1 0 52528 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_461
timestamp 1698431365
transform 1 0 52976 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_465
timestamp 1698431365
transform 1 0 53424 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_523
timestamp 1698431365
transform 1 0 59920 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_579
timestamp 1698431365
transform 1 0 66192 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_583
timestamp 1698431365
transform 1 0 66640 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_585
timestamp 1698431365
transform 1 0 66864 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_588
timestamp 1698431365
transform 1 0 67200 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_592
timestamp 1698431365
transform 1 0 67648 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_594
timestamp 1698431365
transform 1 0 67872 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_649
timestamp 1698431365
transform 1 0 74032 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_661
timestamp 1698431365
transform 1 0 75376 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_675
timestamp 1698431365
transform 1 0 76944 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_685
timestamp 1698431365
transform 1 0 78064 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_687
timestamp 1698431365
transform 1 0 78288 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_8
timestamp 1698431365
transform 1 0 2240 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_12
timestamp 1698431365
transform 1 0 2688 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_28 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 4480 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_36
timestamp 1698431365
transform 1 0 5376 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_40
timestamp 1698431365
transform 1 0 5824 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_44
timestamp 1698431365
transform 1 0 6272 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_48
timestamp 1698431365
transform 1 0 6720 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_52
timestamp 1698431365
transform 1 0 7168 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_56
timestamp 1698431365
transform 1 0 7616 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_60
timestamp 1698431365
transform 1 0 8064 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_72
timestamp 1698431365
transform 1 0 9408 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_74
timestamp 1698431365
transform 1 0 9632 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_122
timestamp 1698431365
transform 1 0 15008 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_130
timestamp 1698431365
transform 1 0 15904 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_136
timestamp 1698431365
transform 1 0 16576 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_148
timestamp 1698431365
transform 1 0 17920 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_150
timestamp 1698431365
transform 1 0 18144 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_153
timestamp 1698431365
transform 1 0 18480 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_157
timestamp 1698431365
transform 1 0 18928 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_161
timestamp 1698431365
transform 1 0 19376 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_163
timestamp 1698431365
transform 1 0 19600 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_170
timestamp 1698431365
transform 1 0 20384 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_194
timestamp 1698431365
transform 1 0 23072 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_196
timestamp 1698431365
transform 1 0 23296 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_205
timestamp 1698431365
transform 1 0 24304 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_207
timestamp 1698431365
transform 1 0 24528 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_212
timestamp 1698431365
transform 1 0 25088 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_230
timestamp 1698431365
transform 1 0 27104 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_276
timestamp 1698431365
transform 1 0 32256 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_290
timestamp 1698431365
transform 1 0 33824 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_352
timestamp 1698431365
transform 1 0 40768 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_356
timestamp 1698431365
transform 1 0 41216 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_360
timestamp 1698431365
transform 1 0 41664 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_419
timestamp 1698431365
transform 1 0 48272 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_430
timestamp 1698431365
transform 1 0 49504 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_434
timestamp 1698431365
transform 1 0 49952 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_438
timestamp 1698431365
transform 1 0 50400 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_442
timestamp 1698431365
transform 1 0 50848 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_445
timestamp 1698431365
transform 1 0 51184 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_449
timestamp 1698431365
transform 1 0 51632 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_459
timestamp 1698431365
transform 1 0 52752 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_475
timestamp 1698431365
transform 1 0 54544 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_483
timestamp 1698431365
transform 1 0 55440 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_487
timestamp 1698431365
transform 1 0 55888 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_492
timestamp 1698431365
transform 1 0 56448 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_494
timestamp 1698431365
transform 1 0 56672 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_547
timestamp 1698431365
transform 1 0 62608 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_553
timestamp 1698431365
transform 1 0 63280 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_557
timestamp 1698431365
transform 1 0 63728 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_614
timestamp 1698431365
transform 1 0 70112 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_616
timestamp 1698431365
transform 1 0 70336 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_619
timestamp 1698431365
transform 1 0 70672 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_623
timestamp 1698431365
transform 1 0 71120 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_627
timestamp 1698431365
transform 1 0 71568 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_684
timestamp 1698431365
transform 1 0 77952 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1568 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_34
timestamp 1698431365
transform 1 0 5152 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_4_37
timestamp 1698431365
transform 1 0 5488 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_55
timestamp 1698431365
transform 1 0 7504 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_83
timestamp 1698431365
transform 1 0 10640 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_90
timestamp 1698431365
transform 1 0 11424 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_94
timestamp 1698431365
transform 1 0 11872 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_97
timestamp 1698431365
transform 1 0 12208 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_101
timestamp 1698431365
transform 1 0 12656 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_113
timestamp 1698431365
transform 1 0 14000 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_115
timestamp 1698431365
transform 1 0 14224 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_124
timestamp 1698431365
transform 1 0 15232 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_126
timestamp 1698431365
transform 1 0 15456 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_129
timestamp 1698431365
transform 1 0 15792 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_170
timestamp 1698431365
transform 1 0 20384 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_172
timestamp 1698431365
transform 1 0 20608 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_177
timestamp 1698431365
transform 1 0 21168 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_181
timestamp 1698431365
transform 1 0 21616 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_191
timestamp 1698431365
transform 1 0 22736 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_205
timestamp 1698431365
transform 1 0 24304 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_209
timestamp 1698431365
transform 1 0 24752 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_233
timestamp 1698431365
transform 1 0 27440 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_287
timestamp 1698431365
transform 1 0 33488 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_304
timestamp 1698431365
transform 1 0 35392 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_306
timestamp 1698431365
transform 1 0 35616 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_317
timestamp 1698431365
transform 1 0 36848 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_424
timestamp 1698431365
transform 1 0 48832 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_428
timestamp 1698431365
transform 1 0 49280 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_432
timestamp 1698431365
transform 1 0 49728 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_434
timestamp 1698431365
transform 1 0 49952 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_451
timestamp 1698431365
transform 1 0 51856 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_457
timestamp 1698431365
transform 1 0 52528 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_489
timestamp 1698431365
transform 1 0 56112 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_493
timestamp 1698431365
transform 1 0 56560 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_4_497
timestamp 1698431365
transform 1 0 57008 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_513
timestamp 1698431365
transform 1 0 58800 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_517
timestamp 1698431365
transform 1 0 59248 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_521
timestamp 1698431365
transform 1 0 59696 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_579
timestamp 1698431365
transform 1 0 66192 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_587
timestamp 1698431365
transform 1 0 67088 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_591
timestamp 1698431365
transform 1 0 67536 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_649
timestamp 1698431365
transform 1 0 74032 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_651
timestamp 1698431365
transform 1 0 74256 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_660
timestamp 1698431365
transform 1 0 75264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_664
timestamp 1698431365
transform 1 0 75712 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_675
timestamp 1698431365
transform 1 0 76944 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_8
timestamp 1698431365
transform 1 0 2240 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_5_12
timestamp 1698431365
transform 1 0 2688 0 -1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_5_44
timestamp 1698431365
transform 1 0 6272 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_60
timestamp 1698431365
transform 1 0 8064 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_68
timestamp 1698431365
transform 1 0 8960 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_72
timestamp 1698431365
transform 1 0 9408 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_74
timestamp 1698431365
transform 1 0 9632 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_77
timestamp 1698431365
transform 1 0 9968 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_120
timestamp 1698431365
transform 1 0 14784 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_122
timestamp 1698431365
transform 1 0 15008 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_131
timestamp 1698431365
transform 1 0 16016 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_133
timestamp 1698431365
transform 1 0 16240 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_136
timestamp 1698431365
transform 1 0 16576 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_142
timestamp 1698431365
transform 1 0 17248 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_146
timestamp 1698431365
transform 1 0 17696 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_157
timestamp 1698431365
transform 1 0 18928 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_159
timestamp 1698431365
transform 1 0 19152 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_174
timestamp 1698431365
transform 1 0 20832 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_212
timestamp 1698431365
transform 1 0 25088 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_216
timestamp 1698431365
transform 1 0 25536 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_220
timestamp 1698431365
transform 1 0 25984 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_230
timestamp 1698431365
transform 1 0 27104 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_232
timestamp 1698431365
transform 1 0 27328 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_260
timestamp 1698431365
transform 1 0 30464 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_262
timestamp 1698431365
transform 1 0 30688 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_269
timestamp 1698431365
transform 1 0 31472 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_279
timestamp 1698431365
transform 1 0 32592 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_294
timestamp 1698431365
transform 1 0 34272 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_324
timestamp 1698431365
transform 1 0 37632 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_326
timestamp 1698431365
transform 1 0 37856 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_404
timestamp 1698431365
transform 1 0 46592 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_408
timestamp 1698431365
transform 1 0 47040 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_410
timestamp 1698431365
transform 1 0 47264 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_413
timestamp 1698431365
transform 1 0 47600 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_415
timestamp 1698431365
transform 1 0 47824 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_418
timestamp 1698431365
transform 1 0 48160 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_422 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 48608 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_486
timestamp 1698431365
transform 1 0 55776 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_5_492
timestamp 1698431365
transform 1 0 56448 0 -1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_524
timestamp 1698431365
transform 1 0 60032 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_5_527
timestamp 1698431365
transform 1 0 60368 0 -1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_559
timestamp 1698431365
transform 1 0 63952 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_5_562
timestamp 1698431365
transform 1 0 64288 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_578
timestamp 1698431365
transform 1 0 66080 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_582
timestamp 1698431365
transform 1 0 66528 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_5_611
timestamp 1698431365
transform 1 0 69776 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_627
timestamp 1698431365
transform 1 0 71568 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_632
timestamp 1698431365
transform 1 0 72128 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_685
timestamp 1698431365
transform 1 0 78064 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_687
timestamp 1698431365
transform 1 0 78288 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_8
timestamp 1698431365
transform 1 0 2240 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_12
timestamp 1698431365
transform 1 0 2688 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_28
timestamp 1698431365
transform 1 0 4480 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_32
timestamp 1698431365
transform 1 0 4928 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_34
timestamp 1698431365
transform 1 0 5152 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_37
timestamp 1698431365
transform 1 0 5488 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_53
timestamp 1698431365
transform 1 0 7280 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_61
timestamp 1698431365
transform 1 0 8176 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_65
timestamp 1698431365
transform 1 0 8624 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_67
timestamp 1698431365
transform 1 0 8848 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_74
timestamp 1698431365
transform 1 0 9632 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_84
timestamp 1698431365
transform 1 0 10752 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_88
timestamp 1698431365
transform 1 0 11200 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_100
timestamp 1698431365
transform 1 0 12544 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_102
timestamp 1698431365
transform 1 0 12768 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_107
timestamp 1698431365
transform 1 0 13328 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_111
timestamp 1698431365
transform 1 0 13776 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_159
timestamp 1698431365
transform 1 0 19152 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_161
timestamp 1698431365
transform 1 0 19376 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_172
timestamp 1698431365
transform 1 0 20608 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_174
timestamp 1698431365
transform 1 0 20832 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_183
timestamp 1698431365
transform 1 0 21840 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_213
timestamp 1698431365
transform 1 0 25200 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_242
timestamp 1698431365
transform 1 0 28448 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_244
timestamp 1698431365
transform 1 0 28672 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_247
timestamp 1698431365
transform 1 0 29008 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_251
timestamp 1698431365
transform 1 0 29456 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_260
timestamp 1698431365
transform 1 0 30464 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_264
timestamp 1698431365
transform 1 0 30912 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_268
timestamp 1698431365
transform 1 0 31360 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_278
timestamp 1698431365
transform 1 0 32480 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_280
timestamp 1698431365
transform 1 0 32704 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_287
timestamp 1698431365
transform 1 0 33488 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_291
timestamp 1698431365
transform 1 0 33936 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_317
timestamp 1698431365
transform 1 0 36848 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_395
timestamp 1698431365
transform 1 0 45584 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_399
timestamp 1698431365
transform 1 0 46032 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_403
timestamp 1698431365
transform 1 0 46480 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_435
timestamp 1698431365
transform 1 0 50064 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_451
timestamp 1698431365
transform 1 0 51856 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_457
timestamp 1698431365
transform 1 0 52528 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_521
timestamp 1698431365
transform 1 0 59696 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_527
timestamp 1698431365
transform 1 0 60368 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_591
timestamp 1698431365
transform 1 0 67536 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_597
timestamp 1698431365
transform 1 0 68208 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_629
timestamp 1698431365
transform 1 0 71792 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_637
timestamp 1698431365
transform 1 0 72688 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_667
timestamp 1698431365
transform 1 0 76048 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_671
timestamp 1698431365
transform 1 0 76496 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_675
timestamp 1698431365
transform 1 0 76944 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_2
timestamp 1698431365
transform 1 0 1568 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_66
timestamp 1698431365
transform 1 0 8736 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_148
timestamp 1698431365
transform 1 0 17920 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_150
timestamp 1698431365
transform 1 0 18144 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_190
timestamp 1698431365
transform 1 0 22624 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_194
timestamp 1698431365
transform 1 0 23072 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_196
timestamp 1698431365
transform 1 0 23296 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_199
timestamp 1698431365
transform 1 0 23632 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_203
timestamp 1698431365
transform 1 0 24080 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_206
timestamp 1698431365
transform 1 0 24416 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_247
timestamp 1698431365
transform 1 0 29008 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_249
timestamp 1698431365
transform 1 0 29232 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_279
timestamp 1698431365
transform 1 0 32592 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_282
timestamp 1698431365
transform 1 0 32928 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_289
timestamp 1698431365
transform 1 0 33712 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_291
timestamp 1698431365
transform 1 0 33936 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_392
timestamp 1698431365
transform 1 0 45248 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_396
timestamp 1698431365
transform 1 0 45696 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_400
timestamp 1698431365
transform 1 0 46144 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_416
timestamp 1698431365
transform 1 0 47936 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_422
timestamp 1698431365
transform 1 0 48608 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_486
timestamp 1698431365
transform 1 0 55776 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_492
timestamp 1698431365
transform 1 0 56448 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_556
timestamp 1698431365
transform 1 0 63616 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_562
timestamp 1698431365
transform 1 0 64288 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_626
timestamp 1698431365
transform 1 0 71456 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_632
timestamp 1698431365
transform 1 0 72128 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_8
timestamp 1698431365
transform 1 0 2240 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_12
timestamp 1698431365
transform 1 0 2688 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_28
timestamp 1698431365
transform 1 0 4480 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_32
timestamp 1698431365
transform 1 0 4928 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_34
timestamp 1698431365
transform 1 0 5152 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_37
timestamp 1698431365
transform 1 0 5488 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_75
timestamp 1698431365
transform 1 0 9744 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_91
timestamp 1698431365
transform 1 0 11536 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_100
timestamp 1698431365
transform 1 0 12544 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_104
timestamp 1698431365
transform 1 0 12992 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_113
timestamp 1698431365
transform 1 0 14000 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_171
timestamp 1698431365
transform 1 0 20496 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_233
timestamp 1698431365
transform 1 0 27440 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_237
timestamp 1698431365
transform 1 0 27888 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_241
timestamp 1698431365
transform 1 0 28336 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_244
timestamp 1698431365
transform 1 0 28672 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_253
timestamp 1698431365
transform 1 0 29680 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_257
timestamp 1698431365
transform 1 0 30128 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_261
timestamp 1698431365
transform 1 0 30576 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_269
timestamp 1698431365
transform 1 0 31472 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_271
timestamp 1698431365
transform 1 0 31696 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_302
timestamp 1698431365
transform 1 0 35168 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_304
timestamp 1698431365
transform 1 0 35392 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_317
timestamp 1698431365
transform 1 0 36848 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_319
timestamp 1698431365
transform 1 0 37072 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_331
timestamp 1698431365
transform 1 0 38416 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_345
timestamp 1698431365
transform 1 0 39984 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_349
timestamp 1698431365
transform 1 0 40432 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_387
timestamp 1698431365
transform 1 0 44688 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_394
timestamp 1698431365
transform 1 0 45472 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_426
timestamp 1698431365
transform 1 0 49056 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_442
timestamp 1698431365
transform 1 0 50848 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_450
timestamp 1698431365
transform 1 0 51744 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_454
timestamp 1698431365
transform 1 0 52192 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_457
timestamp 1698431365
transform 1 0 52528 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_521
timestamp 1698431365
transform 1 0 59696 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_527
timestamp 1698431365
transform 1 0 60368 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_591
timestamp 1698431365
transform 1 0 67536 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_597
timestamp 1698431365
transform 1 0 68208 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_629
timestamp 1698431365
transform 1 0 71792 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_645
timestamp 1698431365
transform 1 0 73584 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_653
timestamp 1698431365
transform 1 0 74480 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_657
timestamp 1698431365
transform 1 0 74928 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_661
timestamp 1698431365
transform 1 0 75376 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_667
timestamp 1698431365
transform 1 0 76048 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_671
timestamp 1698431365
transform 1 0 76496 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_673
timestamp 1698431365
transform 1 0 76720 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_676
timestamp 1698431365
transform 1 0 77056 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_8
timestamp 1698431365
transform 1 0 2240 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_9_12
timestamp 1698431365
transform 1 0 2688 0 -1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_9_44
timestamp 1698431365
transform 1 0 6272 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_60
timestamp 1698431365
transform 1 0 8064 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_68
timestamp 1698431365
transform 1 0 8960 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_109
timestamp 1698431365
transform 1 0 13552 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_115
timestamp 1698431365
transform 1 0 14224 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_119
timestamp 1698431365
transform 1 0 14672 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_121
timestamp 1698431365
transform 1 0 14896 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_124
timestamp 1698431365
transform 1 0 15232 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_128
timestamp 1698431365
transform 1 0 15680 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_132
timestamp 1698431365
transform 1 0 16128 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_142
timestamp 1698431365
transform 1 0 17248 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_144
timestamp 1698431365
transform 1 0 17472 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_184
timestamp 1698431365
transform 1 0 21952 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_188
timestamp 1698431365
transform 1 0 22400 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_195
timestamp 1698431365
transform 1 0 23184 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_203
timestamp 1698431365
transform 1 0 24080 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_207
timestamp 1698431365
transform 1 0 24528 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_209
timestamp 1698431365
transform 1 0 24752 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_228
timestamp 1698431365
transform 1 0 26880 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_236
timestamp 1698431365
transform 1 0 27776 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_269
timestamp 1698431365
transform 1 0 31472 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_277
timestamp 1698431365
transform 1 0 32368 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_332
timestamp 1698431365
transform 1 0 38528 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_334
timestamp 1698431365
transform 1 0 38752 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_343
timestamp 1698431365
transform 1 0 39760 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_352
timestamp 1698431365
transform 1 0 40768 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_9_385
timestamp 1698431365
transform 1 0 44464 0 -1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_417
timestamp 1698431365
transform 1 0 48048 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_419
timestamp 1698431365
transform 1 0 48272 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_422
timestamp 1698431365
transform 1 0 48608 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_486
timestamp 1698431365
transform 1 0 55776 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_492
timestamp 1698431365
transform 1 0 56448 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_556
timestamp 1698431365
transform 1 0 63616 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_562
timestamp 1698431365
transform 1 0 64288 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_626
timestamp 1698431365
transform 1 0 71456 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_9_632
timestamp 1698431365
transform 1 0 72128 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_648
timestamp 1698431365
transform 1 0 73920 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_656
timestamp 1698431365
transform 1 0 74816 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_660
timestamp 1698431365
transform 1 0 75264 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_8
timestamp 1698431365
transform 1 0 2240 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_12
timestamp 1698431365
transform 1 0 2688 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_28
timestamp 1698431365
transform 1 0 4480 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_32
timestamp 1698431365
transform 1 0 4928 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_34
timestamp 1698431365
transform 1 0 5152 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_37
timestamp 1698431365
transform 1 0 5488 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_53
timestamp 1698431365
transform 1 0 7280 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_61
timestamp 1698431365
transform 1 0 8176 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_65
timestamp 1698431365
transform 1 0 8624 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_98
timestamp 1698431365
transform 1 0 12320 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_102
timestamp 1698431365
transform 1 0 12768 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_104
timestamp 1698431365
transform 1 0 12992 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_115
timestamp 1698431365
transform 1 0 14224 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_119
timestamp 1698431365
transform 1 0 14672 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_154
timestamp 1698431365
transform 1 0 18592 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_156
timestamp 1698431365
transform 1 0 18816 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_171
timestamp 1698431365
transform 1 0 20496 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_177
timestamp 1698431365
transform 1 0 21168 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_185
timestamp 1698431365
transform 1 0 22064 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_198
timestamp 1698431365
transform 1 0 23520 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_206
timestamp 1698431365
transform 1 0 24416 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_247
timestamp 1698431365
transform 1 0 29008 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_261
timestamp 1698431365
transform 1 0 30576 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_269
timestamp 1698431365
transform 1 0 31472 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_327
timestamp 1698431365
transform 1 0 37968 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_329
timestamp 1698431365
transform 1 0 38192 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_382
timestamp 1698431365
transform 1 0 44128 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_384
timestamp 1698431365
transform 1 0 44352 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_393
timestamp 1698431365
transform 1 0 45360 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_425
timestamp 1698431365
transform 1 0 48944 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_441
timestamp 1698431365
transform 1 0 50736 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_449
timestamp 1698431365
transform 1 0 51632 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_453
timestamp 1698431365
transform 1 0 52080 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_457
timestamp 1698431365
transform 1 0 52528 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_521
timestamp 1698431365
transform 1 0 59696 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_527
timestamp 1698431365
transform 1 0 60368 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_591
timestamp 1698431365
transform 1 0 67536 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_597
timestamp 1698431365
transform 1 0 68208 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_661
timestamp 1698431365
transform 1 0 75376 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_667
timestamp 1698431365
transform 1 0 76048 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_669
timestamp 1698431365
transform 1 0 76272 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_672
timestamp 1698431365
transform 1 0 76608 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_2
timestamp 1698431365
transform 1 0 1568 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_66
timestamp 1698431365
transform 1 0 8736 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_78
timestamp 1698431365
transform 1 0 10080 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_86
timestamp 1698431365
transform 1 0 10976 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_90
timestamp 1698431365
transform 1 0 11424 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_130
timestamp 1698431365
transform 1 0 15904 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_138
timestamp 1698431365
transform 1 0 16800 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_142
timestamp 1698431365
transform 1 0 17248 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_144
timestamp 1698431365
transform 1 0 17472 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_151
timestamp 1698431365
transform 1 0 18256 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_155
timestamp 1698431365
transform 1 0 18704 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_171
timestamp 1698431365
transform 1 0 20496 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_179
timestamp 1698431365
transform 1 0 21392 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_220
timestamp 1698431365
transform 1 0 25984 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_227
timestamp 1698431365
transform 1 0 26768 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_243
timestamp 1698431365
transform 1 0 28560 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_282
timestamp 1698431365
transform 1 0 32928 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_290
timestamp 1698431365
transform 1 0 33824 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_294
timestamp 1698431365
transform 1 0 34272 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_296
timestamp 1698431365
transform 1 0 34496 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_309
timestamp 1698431365
transform 1 0 35952 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_313
timestamp 1698431365
transform 1 0 36400 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_317
timestamp 1698431365
transform 1 0 36848 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_357
timestamp 1698431365
transform 1 0 41328 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_11_361
timestamp 1698431365
transform 1 0 41776 0 -1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_393
timestamp 1698431365
transform 1 0 45360 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_409
timestamp 1698431365
transform 1 0 47152 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_417
timestamp 1698431365
transform 1 0 48048 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_419
timestamp 1698431365
transform 1 0 48272 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_422
timestamp 1698431365
transform 1 0 48608 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_486
timestamp 1698431365
transform 1 0 55776 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_492
timestamp 1698431365
transform 1 0 56448 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_556
timestamp 1698431365
transform 1 0 63616 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_562
timestamp 1698431365
transform 1 0 64288 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_626
timestamp 1698431365
transform 1 0 71456 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_11_632
timestamp 1698431365
transform 1 0 72128 0 -1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_664
timestamp 1698431365
transform 1 0 75712 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_672
timestamp 1698431365
transform 1 0 76608 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_676
timestamp 1698431365
transform 1 0 77056 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_678
timestamp 1698431365
transform 1 0 77280 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_685
timestamp 1698431365
transform 1 0 78064 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_687
timestamp 1698431365
transform 1 0 78288 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_8
timestamp 1698431365
transform 1 0 2240 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_12
timestamp 1698431365
transform 1 0 2688 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_28
timestamp 1698431365
transform 1 0 4480 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_32
timestamp 1698431365
transform 1 0 4928 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_34
timestamp 1698431365
transform 1 0 5152 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_37
timestamp 1698431365
transform 1 0 5488 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_69
timestamp 1698431365
transform 1 0 9072 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_85
timestamp 1698431365
transform 1 0 10864 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_93
timestamp 1698431365
transform 1 0 11760 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_97
timestamp 1698431365
transform 1 0 12208 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_101
timestamp 1698431365
transform 1 0 12656 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_107
timestamp 1698431365
transform 1 0 13328 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_123
timestamp 1698431365
transform 1 0 15120 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_131
timestamp 1698431365
transform 1 0 16016 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_172
timestamp 1698431365
transform 1 0 20608 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_174
timestamp 1698431365
transform 1 0 20832 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_177
timestamp 1698431365
transform 1 0 21168 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_185
timestamp 1698431365
transform 1 0 22064 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_187
timestamp 1698431365
transform 1 0 22288 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_217
timestamp 1698431365
transform 1 0 25648 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_233
timestamp 1698431365
transform 1 0 27440 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_237
timestamp 1698431365
transform 1 0 27888 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_247
timestamp 1698431365
transform 1 0 29008 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_249
timestamp 1698431365
transform 1 0 29232 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_256
timestamp 1698431365
transform 1 0 30016 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_264
timestamp 1698431365
transform 1 0 30912 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_279
timestamp 1698431365
transform 1 0 32592 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_283
timestamp 1698431365
transform 1 0 33040 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_285
timestamp 1698431365
transform 1 0 33264 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_317
timestamp 1698431365
transform 1 0 36848 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_336
timestamp 1698431365
transform 1 0 38976 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_338
timestamp 1698431365
transform 1 0 39200 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_376
timestamp 1698431365
transform 1 0 43456 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_384
timestamp 1698431365
transform 1 0 44352 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_387
timestamp 1698431365
transform 1 0 44688 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_451
timestamp 1698431365
transform 1 0 51856 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_457
timestamp 1698431365
transform 1 0 52528 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_521
timestamp 1698431365
transform 1 0 59696 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_527
timestamp 1698431365
transform 1 0 60368 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_591
timestamp 1698431365
transform 1 0 67536 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_597
timestamp 1698431365
transform 1 0 68208 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_629
timestamp 1698431365
transform 1 0 71792 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_645
timestamp 1698431365
transform 1 0 73584 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_649
timestamp 1698431365
transform 1 0 74032 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_651
timestamp 1698431365
transform 1 0 74256 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_662
timestamp 1698431365
transform 1 0 75488 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_664
timestamp 1698431365
transform 1 0 75712 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_667
timestamp 1698431365
transform 1 0 76048 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_671
timestamp 1698431365
transform 1 0 76496 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_687
timestamp 1698431365
transform 1 0 78288 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_8
timestamp 1698431365
transform 1 0 2240 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_13_12
timestamp 1698431365
transform 1 0 2688 0 -1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_44
timestamp 1698431365
transform 1 0 6272 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_60
timestamp 1698431365
transform 1 0 8064 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_68
timestamp 1698431365
transform 1 0 8960 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_72
timestamp 1698431365
transform 1 0 9408 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_136
timestamp 1698431365
transform 1 0 16576 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_142
timestamp 1698431365
transform 1 0 17248 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_150
timestamp 1698431365
transform 1 0 18144 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_195
timestamp 1698431365
transform 1 0 23184 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_203
timestamp 1698431365
transform 1 0 24080 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_207
timestamp 1698431365
transform 1 0 24528 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_209
timestamp 1698431365
transform 1 0 24752 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_212
timestamp 1698431365
transform 1 0 25088 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_220
timestamp 1698431365
transform 1 0 25984 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_232
timestamp 1698431365
transform 1 0 27328 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_240
timestamp 1698431365
transform 1 0 28224 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_257
timestamp 1698431365
transform 1 0 30128 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_261
timestamp 1698431365
transform 1 0 30576 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_263
timestamp 1698431365
transform 1 0 30800 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_279
timestamp 1698431365
transform 1 0 32592 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_290
timestamp 1698431365
transform 1 0 33824 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_294
timestamp 1698431365
transform 1 0 34272 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_308
timestamp 1698431365
transform 1 0 35840 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_316
timestamp 1698431365
transform 1 0 36736 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_320
timestamp 1698431365
transform 1 0 37184 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_322
timestamp 1698431365
transform 1 0 37408 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_344
timestamp 1698431365
transform 1 0 39872 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_348
timestamp 1698431365
transform 1 0 40320 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_360
timestamp 1698431365
transform 1 0 41664 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_395
timestamp 1698431365
transform 1 0 45584 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_403
timestamp 1698431365
transform 1 0 46480 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_406
timestamp 1698431365
transform 1 0 46816 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_414
timestamp 1698431365
transform 1 0 47712 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_416
timestamp 1698431365
transform 1 0 47936 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_419
timestamp 1698431365
transform 1 0 48272 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_422
timestamp 1698431365
transform 1 0 48608 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_426
timestamp 1698431365
transform 1 0 49056 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_442
timestamp 1698431365
transform 1 0 50848 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_478
timestamp 1698431365
transform 1 0 54880 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_482
timestamp 1698431365
transform 1 0 55328 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_492
timestamp 1698431365
transform 1 0 56448 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_556
timestamp 1698431365
transform 1 0 63616 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_562
timestamp 1698431365
transform 1 0 64288 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_626
timestamp 1698431365
transform 1 0 71456 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_13_632
timestamp 1698431365
transform 1 0 72128 0 -1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_664
timestamp 1698431365
transform 1 0 75712 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_2
timestamp 1698431365
transform 1 0 1568 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_34
timestamp 1698431365
transform 1 0 5152 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_37
timestamp 1698431365
transform 1 0 5488 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_101
timestamp 1698431365
transform 1 0 12656 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_107
timestamp 1698431365
transform 1 0 13328 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_139
timestamp 1698431365
transform 1 0 16912 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_155
timestamp 1698431365
transform 1 0 18704 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_163
timestamp 1698431365
transform 1 0 19600 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_172
timestamp 1698431365
transform 1 0 20608 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_174
timestamp 1698431365
transform 1 0 20832 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_177
timestamp 1698431365
transform 1 0 21168 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_181
timestamp 1698431365
transform 1 0 21616 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_197
timestamp 1698431365
transform 1 0 23408 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_205
timestamp 1698431365
transform 1 0 24304 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_244
timestamp 1698431365
transform 1 0 28672 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_261
timestamp 1698431365
transform 1 0 30576 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_265
timestamp 1698431365
transform 1 0 31024 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_269
timestamp 1698431365
transform 1 0 31472 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_299
timestamp 1698431365
transform 1 0 34832 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_311
timestamp 1698431365
transform 1 0 36176 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_317
timestamp 1698431365
transform 1 0 36848 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_321
timestamp 1698431365
transform 1 0 37296 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_331
timestamp 1698431365
transform 1 0 38416 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_364
timestamp 1698431365
transform 1 0 42112 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_377
timestamp 1698431365
transform 1 0 43568 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_381
timestamp 1698431365
transform 1 0 44016 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_387
timestamp 1698431365
transform 1 0 44688 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_395
timestamp 1698431365
transform 1 0 45584 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_399
timestamp 1698431365
transform 1 0 46032 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_434
timestamp 1698431365
transform 1 0 49952 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_442
timestamp 1698431365
transform 1 0 50848 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_467
timestamp 1698431365
transform 1 0 53648 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_499
timestamp 1698431365
transform 1 0 57232 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_515
timestamp 1698431365
transform 1 0 59024 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_523
timestamp 1698431365
transform 1 0 59920 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_527
timestamp 1698431365
transform 1 0 60368 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_591
timestamp 1698431365
transform 1 0 67536 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_597
timestamp 1698431365
transform 1 0 68208 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_661
timestamp 1698431365
transform 1 0 75376 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_667
timestamp 1698431365
transform 1 0 76048 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_675
timestamp 1698431365
transform 1 0 76944 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_679
timestamp 1698431365
transform 1 0 77392 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_8
timestamp 1698431365
transform 1 0 2240 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_15_12
timestamp 1698431365
transform 1 0 2688 0 -1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_44
timestamp 1698431365
transform 1 0 6272 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_60
timestamp 1698431365
transform 1 0 8064 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_68
timestamp 1698431365
transform 1 0 8960 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_72
timestamp 1698431365
transform 1 0 9408 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_136
timestamp 1698431365
transform 1 0 16576 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_142
timestamp 1698431365
transform 1 0 17248 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_206
timestamp 1698431365
transform 1 0 24416 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_212
timestamp 1698431365
transform 1 0 25088 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_216
timestamp 1698431365
transform 1 0 25536 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_267
timestamp 1698431365
transform 1 0 31248 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_275
timestamp 1698431365
transform 1 0 32144 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_279
timestamp 1698431365
transform 1 0 32592 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_290
timestamp 1698431365
transform 1 0 33824 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_298
timestamp 1698431365
transform 1 0 34720 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_329
timestamp 1698431365
transform 1 0 38192 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_348
timestamp 1698431365
transform 1 0 40320 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_352
timestamp 1698431365
transform 1 0 40768 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_356
timestamp 1698431365
transform 1 0 41216 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_360
timestamp 1698431365
transform 1 0 41664 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_362
timestamp 1698431365
transform 1 0 41888 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_396
timestamp 1698431365
transform 1 0 45696 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_398
timestamp 1698431365
transform 1 0 45920 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_401
timestamp 1698431365
transform 1 0 46256 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_405
timestamp 1698431365
transform 1 0 46704 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_407
timestamp 1698431365
transform 1 0 46928 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_418
timestamp 1698431365
transform 1 0 48160 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_486
timestamp 1698431365
transform 1 0 55776 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_492
timestamp 1698431365
transform 1 0 56448 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_556
timestamp 1698431365
transform 1 0 63616 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_562
timestamp 1698431365
transform 1 0 64288 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_626
timestamp 1698431365
transform 1 0 71456 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_15_632
timestamp 1698431365
transform 1 0 72128 0 -1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_664
timestamp 1698431365
transform 1 0 75712 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_680
timestamp 1698431365
transform 1 0 77504 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_8
timestamp 1698431365
transform 1 0 2240 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_12
timestamp 1698431365
transform 1 0 2688 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_28
timestamp 1698431365
transform 1 0 4480 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_32
timestamp 1698431365
transform 1 0 4928 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_34
timestamp 1698431365
transform 1 0 5152 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_37
timestamp 1698431365
transform 1 0 5488 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_101
timestamp 1698431365
transform 1 0 12656 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_107
timestamp 1698431365
transform 1 0 13328 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_171
timestamp 1698431365
transform 1 0 20496 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_177
timestamp 1698431365
transform 1 0 21168 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_209
timestamp 1698431365
transform 1 0 24752 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_213
timestamp 1698431365
transform 1 0 25200 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_217
timestamp 1698431365
transform 1 0 25648 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_311
timestamp 1698431365
transform 1 0 36176 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_317
timestamp 1698431365
transform 1 0 36848 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_319
timestamp 1698431365
transform 1 0 37072 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_324
timestamp 1698431365
transform 1 0 37632 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_328
timestamp 1698431365
transform 1 0 38080 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_332
timestamp 1698431365
transform 1 0 38528 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_336
timestamp 1698431365
transform 1 0 38976 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_346
timestamp 1698431365
transform 1 0 40096 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_352
timestamp 1698431365
transform 1 0 40768 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_356
timestamp 1698431365
transform 1 0 41216 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_364
timestamp 1698431365
transform 1 0 42112 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_368
timestamp 1698431365
transform 1 0 42560 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_372
timestamp 1698431365
transform 1 0 43008 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_383
timestamp 1698431365
transform 1 0 44240 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_387
timestamp 1698431365
transform 1 0 44688 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_391
timestamp 1698431365
transform 1 0 45136 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_395
timestamp 1698431365
transform 1 0 45584 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_447
timestamp 1698431365
transform 1 0 51408 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_451
timestamp 1698431365
transform 1 0 51856 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_489
timestamp 1698431365
transform 1 0 56112 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_521
timestamp 1698431365
transform 1 0 59696 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_527
timestamp 1698431365
transform 1 0 60368 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_591
timestamp 1698431365
transform 1 0 67536 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_597
timestamp 1698431365
transform 1 0 68208 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_661
timestamp 1698431365
transform 1 0 75376 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_667
timestamp 1698431365
transform 1 0 76048 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_675
timestamp 1698431365
transform 1 0 76944 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_679
timestamp 1698431365
transform 1 0 77392 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_2
timestamp 1698431365
transform 1 0 1568 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_66
timestamp 1698431365
transform 1 0 8736 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_72
timestamp 1698431365
transform 1 0 9408 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_136
timestamp 1698431365
transform 1 0 16576 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_142
timestamp 1698431365
transform 1 0 17248 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_174
timestamp 1698431365
transform 1 0 20832 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_190
timestamp 1698431365
transform 1 0 22624 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_193
timestamp 1698431365
transform 1 0 22960 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_209
timestamp 1698431365
transform 1 0 24752 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_212
timestamp 1698431365
transform 1 0 25088 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_242
timestamp 1698431365
transform 1 0 28448 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_278
timestamp 1698431365
transform 1 0 32480 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_282
timestamp 1698431365
transform 1 0 32928 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_288
timestamp 1698431365
transform 1 0 33600 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_292
timestamp 1698431365
transform 1 0 34048 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_296
timestamp 1698431365
transform 1 0 34496 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_314
timestamp 1698431365
transform 1 0 36512 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_316
timestamp 1698431365
transform 1 0 36736 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_327
timestamp 1698431365
transform 1 0 37968 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_336
timestamp 1698431365
transform 1 0 38976 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_346
timestamp 1698431365
transform 1 0 40096 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_352
timestamp 1698431365
transform 1 0 40768 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_366
timestamp 1698431365
transform 1 0 42336 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_417
timestamp 1698431365
transform 1 0 48048 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_419
timestamp 1698431365
transform 1 0 48272 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_486
timestamp 1698431365
transform 1 0 55776 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_492
timestamp 1698431365
transform 1 0 56448 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_496
timestamp 1698431365
transform 1 0 56896 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_500
timestamp 1698431365
transform 1 0 57344 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_532
timestamp 1698431365
transform 1 0 60928 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_548
timestamp 1698431365
transform 1 0 62720 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_556
timestamp 1698431365
transform 1 0 63616 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_562
timestamp 1698431365
transform 1 0 64288 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_626
timestamp 1698431365
transform 1 0 71456 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_632
timestamp 1698431365
transform 1 0 72128 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_664
timestamp 1698431365
transform 1 0 75712 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_8
timestamp 1698431365
transform 1 0 2240 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_12
timestamp 1698431365
transform 1 0 2688 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_28
timestamp 1698431365
transform 1 0 4480 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_32
timestamp 1698431365
transform 1 0 4928 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_34
timestamp 1698431365
transform 1 0 5152 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_37
timestamp 1698431365
transform 1 0 5488 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_101
timestamp 1698431365
transform 1 0 12656 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_107
timestamp 1698431365
transform 1 0 13328 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_139
timestamp 1698431365
transform 1 0 16912 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_162
timestamp 1698431365
transform 1 0 19488 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_166
timestamp 1698431365
transform 1 0 19936 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_177
timestamp 1698431365
transform 1 0 21168 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_181
timestamp 1698431365
transform 1 0 21616 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_241
timestamp 1698431365
transform 1 0 28336 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_247
timestamp 1698431365
transform 1 0 29008 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_251
timestamp 1698431365
transform 1 0 29456 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_259
timestamp 1698431365
transform 1 0 30352 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_261
timestamp 1698431365
transform 1 0 30576 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_270
timestamp 1698431365
transform 1 0 31584 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_278
timestamp 1698431365
transform 1 0 32480 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_282
timestamp 1698431365
transform 1 0 32928 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_300
timestamp 1698431365
transform 1 0 34944 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_329
timestamp 1698431365
transform 1 0 38192 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_351
timestamp 1698431365
transform 1 0 40656 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_387
timestamp 1698431365
transform 1 0 44688 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_434
timestamp 1698431365
transform 1 0 49952 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_451
timestamp 1698431365
transform 1 0 51856 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_457
timestamp 1698431365
transform 1 0 52528 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_459
timestamp 1698431365
transform 1 0 52752 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_524
timestamp 1698431365
transform 1 0 60032 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_527
timestamp 1698431365
transform 1 0 60368 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_591
timestamp 1698431365
transform 1 0 67536 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_597
timestamp 1698431365
transform 1 0 68208 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_613
timestamp 1698431365
transform 1 0 70000 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_622
timestamp 1698431365
transform 1 0 71008 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_654
timestamp 1698431365
transform 1 0 74592 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_662
timestamp 1698431365
transform 1 0 75488 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_664
timestamp 1698431365
transform 1 0 75712 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_667
timestamp 1698431365
transform 1 0 76048 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_675
timestamp 1698431365
transform 1 0 76944 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_679
timestamp 1698431365
transform 1 0 77392 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_8
timestamp 1698431365
transform 1 0 2240 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_12
timestamp 1698431365
transform 1 0 2688 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_44
timestamp 1698431365
transform 1 0 6272 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_60
timestamp 1698431365
transform 1 0 8064 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_68
timestamp 1698431365
transform 1 0 8960 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_72
timestamp 1698431365
transform 1 0 9408 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_136
timestamp 1698431365
transform 1 0 16576 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_142
timestamp 1698431365
transform 1 0 17248 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_144
timestamp 1698431365
transform 1 0 17472 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_212
timestamp 1698431365
transform 1 0 25088 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_219
timestamp 1698431365
transform 1 0 25872 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_221
timestamp 1698431365
transform 1 0 26096 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_282
timestamp 1698431365
transform 1 0 32928 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_292
timestamp 1698431365
transform 1 0 34048 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_369
timestamp 1698431365
transform 1 0 42672 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_371
timestamp 1698431365
transform 1 0 42896 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_418
timestamp 1698431365
transform 1 0 48160 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_454
timestamp 1698431365
transform 1 0 52192 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_492
timestamp 1698431365
transform 1 0 56448 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_496
timestamp 1698431365
transform 1 0 56896 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_500
timestamp 1698431365
transform 1 0 57344 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_532
timestamp 1698431365
transform 1 0 60928 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_548
timestamp 1698431365
transform 1 0 62720 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_556
timestamp 1698431365
transform 1 0 63616 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_562
timestamp 1698431365
transform 1 0 64288 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_626
timestamp 1698431365
transform 1 0 71456 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_632
timestamp 1698431365
transform 1 0 72128 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_664
timestamp 1698431365
transform 1 0 75712 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_672
timestamp 1698431365
transform 1 0 76608 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_8
timestamp 1698431365
transform 1 0 2240 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_12
timestamp 1698431365
transform 1 0 2688 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_28
timestamp 1698431365
transform 1 0 4480 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_32
timestamp 1698431365
transform 1 0 4928 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_34
timestamp 1698431365
transform 1 0 5152 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_37
timestamp 1698431365
transform 1 0 5488 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_101
timestamp 1698431365
transform 1 0 12656 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_107
timestamp 1698431365
transform 1 0 13328 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_139
timestamp 1698431365
transform 1 0 16912 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_155
timestamp 1698431365
transform 1 0 18704 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_163
timestamp 1698431365
transform 1 0 19600 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_172
timestamp 1698431365
transform 1 0 20608 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_174
timestamp 1698431365
transform 1 0 20832 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_177
timestamp 1698431365
transform 1 0 21168 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_203
timestamp 1698431365
transform 1 0 24080 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_205
timestamp 1698431365
transform 1 0 24304 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_220
timestamp 1698431365
transform 1 0 25984 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_227
timestamp 1698431365
transform 1 0 26768 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_237
timestamp 1698431365
transform 1 0 27888 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_241
timestamp 1698431365
transform 1 0 28336 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_311
timestamp 1698431365
transform 1 0 36176 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_317
timestamp 1698431365
transform 1 0 36848 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_319
timestamp 1698431365
transform 1 0 37072 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_419
timestamp 1698431365
transform 1 0 48272 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_465
timestamp 1698431365
transform 1 0 53424 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_498
timestamp 1698431365
transform 1 0 57120 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_502
timestamp 1698431365
transform 1 0 57568 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_518
timestamp 1698431365
transform 1 0 59360 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_522
timestamp 1698431365
transform 1 0 59808 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_524
timestamp 1698431365
transform 1 0 60032 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_527
timestamp 1698431365
transform 1 0 60368 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_591
timestamp 1698431365
transform 1 0 67536 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_597
timestamp 1698431365
transform 1 0 68208 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_661
timestamp 1698431365
transform 1 0 75376 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_667
timestamp 1698431365
transform 1 0 76048 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_669
timestamp 1698431365
transform 1 0 76272 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_684
timestamp 1698431365
transform 1 0 77952 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_2
timestamp 1698431365
transform 1 0 1568 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_66
timestamp 1698431365
transform 1 0 8736 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_72
timestamp 1698431365
transform 1 0 9408 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_136
timestamp 1698431365
transform 1 0 16576 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_142
timestamp 1698431365
transform 1 0 17248 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_150
timestamp 1698431365
transform 1 0 18144 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_157
timestamp 1698431365
transform 1 0 18928 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_159
timestamp 1698431365
transform 1 0 19152 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_218
timestamp 1698431365
transform 1 0 25760 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_220
timestamp 1698431365
transform 1 0 25984 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_226
timestamp 1698431365
transform 1 0 26656 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_230
timestamp 1698431365
transform 1 0 27104 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_263
timestamp 1698431365
transform 1 0 30800 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_272
timestamp 1698431365
transform 1 0 31808 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_276
timestamp 1698431365
transform 1 0 32256 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_282
timestamp 1698431365
transform 1 0 32928 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_284
timestamp 1698431365
transform 1 0 33152 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_301
timestamp 1698431365
transform 1 0 35056 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_347
timestamp 1698431365
transform 1 0 40208 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_349
timestamp 1698431365
transform 1 0 40432 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_422
timestamp 1698431365
transform 1 0 48608 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_484
timestamp 1698431365
transform 1 0 55552 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_488
timestamp 1698431365
transform 1 0 56000 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_492
timestamp 1698431365
transform 1 0 56448 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_496
timestamp 1698431365
transform 1 0 56896 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_562
timestamp 1698431365
transform 1 0 64288 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_626
timestamp 1698431365
transform 1 0 71456 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_632
timestamp 1698431365
transform 1 0 72128 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_634
timestamp 1698431365
transform 1 0 72352 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_637
timestamp 1698431365
transform 1 0 72688 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_655
timestamp 1698431365
transform 1 0 74704 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_661
timestamp 1698431365
transform 1 0 75376 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_665
timestamp 1698431365
transform 1 0 75824 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_678
timestamp 1698431365
transform 1 0 77280 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_8
timestamp 1698431365
transform 1 0 2240 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_12
timestamp 1698431365
transform 1 0 2688 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_28
timestamp 1698431365
transform 1 0 4480 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_32
timestamp 1698431365
transform 1 0 4928 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_34
timestamp 1698431365
transform 1 0 5152 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_37
timestamp 1698431365
transform 1 0 5488 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_101
timestamp 1698431365
transform 1 0 12656 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_107
timestamp 1698431365
transform 1 0 13328 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_139
timestamp 1698431365
transform 1 0 16912 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_147
timestamp 1698431365
transform 1 0 17808 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_151
timestamp 1698431365
transform 1 0 18256 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_153
timestamp 1698431365
transform 1 0 18480 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_161
timestamp 1698431365
transform 1 0 19376 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_169
timestamp 1698431365
transform 1 0 20272 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_171
timestamp 1698431365
transform 1 0 20496 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_174
timestamp 1698431365
transform 1 0 20832 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_177
timestamp 1698431365
transform 1 0 21168 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_235
timestamp 1698431365
transform 1 0 27664 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_239
timestamp 1698431365
transform 1 0 28112 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_243
timestamp 1698431365
transform 1 0 28560 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_290
timestamp 1698431365
transform 1 0 33824 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_292
timestamp 1698431365
transform 1 0 34048 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_323
timestamp 1698431365
transform 1 0 37520 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_325
timestamp 1698431365
transform 1 0 37744 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_334
timestamp 1698431365
transform 1 0 38752 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_416
timestamp 1698431365
transform 1 0 47936 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_452
timestamp 1698431365
transform 1 0 51968 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_454
timestamp 1698431365
transform 1 0 52192 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_496
timestamp 1698431365
transform 1 0 56896 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_500
timestamp 1698431365
transform 1 0 57344 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_516
timestamp 1698431365
transform 1 0 59136 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_524
timestamp 1698431365
transform 1 0 60032 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_527
timestamp 1698431365
transform 1 0 60368 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_591
timestamp 1698431365
transform 1 0 67536 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_597
timestamp 1698431365
transform 1 0 68208 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_613
timestamp 1698431365
transform 1 0 70000 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_617
timestamp 1698431365
transform 1 0 70448 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_619
timestamp 1698431365
transform 1 0 70672 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_652
timestamp 1698431365
transform 1 0 74368 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_656
timestamp 1698431365
transform 1 0 74816 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_658
timestamp 1698431365
transform 1 0 75040 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_667
timestamp 1698431365
transform 1 0 76048 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_671
timestamp 1698431365
transform 1 0 76496 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_684
timestamp 1698431365
transform 1 0 77952 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_8
timestamp 1698431365
transform 1 0 2240 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_12
timestamp 1698431365
transform 1 0 2688 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_44
timestamp 1698431365
transform 1 0 6272 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_60
timestamp 1698431365
transform 1 0 8064 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_68
timestamp 1698431365
transform 1 0 8960 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_72
timestamp 1698431365
transform 1 0 9408 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_136
timestamp 1698431365
transform 1 0 16576 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_150
timestamp 1698431365
transform 1 0 18144 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_154
timestamp 1698431365
transform 1 0 18592 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_156
timestamp 1698431365
transform 1 0 18816 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_192
timestamp 1698431365
transform 1 0 22848 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_196
timestamp 1698431365
transform 1 0 23296 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_205
timestamp 1698431365
transform 1 0 24304 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_209
timestamp 1698431365
transform 1 0 24752 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_212
timestamp 1698431365
transform 1 0 25088 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_216
timestamp 1698431365
transform 1 0 25536 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_219
timestamp 1698431365
transform 1 0 25872 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_227
timestamp 1698431365
transform 1 0 26768 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_259
timestamp 1698431365
transform 1 0 30352 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_275
timestamp 1698431365
transform 1 0 32144 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_279
timestamp 1698431365
transform 1 0 32592 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_282
timestamp 1698431365
transform 1 0 32928 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_290
timestamp 1698431365
transform 1 0 33824 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_294
timestamp 1698431365
transform 1 0 34272 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_297
timestamp 1698431365
transform 1 0 34608 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_317
timestamp 1698431365
transform 1 0 36848 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_352
timestamp 1698431365
transform 1 0 40768 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_354
timestamp 1698431365
transform 1 0 40992 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_365
timestamp 1698431365
transform 1 0 42224 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_376
timestamp 1698431365
transform 1 0 43456 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_417
timestamp 1698431365
transform 1 0 48048 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_419
timestamp 1698431365
transform 1 0 48272 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_482
timestamp 1698431365
transform 1 0 55328 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_486
timestamp 1698431365
transform 1 0 55776 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_492
timestamp 1698431365
transform 1 0 56448 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_556
timestamp 1698431365
transform 1 0 63616 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_562
timestamp 1698431365
transform 1 0 64288 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_594
timestamp 1698431365
transform 1 0 67872 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_610
timestamp 1698431365
transform 1 0 69664 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_612
timestamp 1698431365
transform 1 0 69888 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_647
timestamp 1698431365
transform 1 0 73808 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_651
timestamp 1698431365
transform 1 0 74256 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_667
timestamp 1698431365
transform 1 0 76048 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_669
timestamp 1698431365
transform 1 0 76272 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_2
timestamp 1698431365
transform 1 0 1568 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_34
timestamp 1698431365
transform 1 0 5152 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_37
timestamp 1698431365
transform 1 0 5488 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_101
timestamp 1698431365
transform 1 0 12656 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_107
timestamp 1698431365
transform 1 0 13328 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_123
timestamp 1698431365
transform 1 0 15120 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_131
timestamp 1698431365
transform 1 0 16016 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_133
timestamp 1698431365
transform 1 0 16240 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_185
timestamp 1698431365
transform 1 0 22064 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_189
timestamp 1698431365
transform 1 0 22512 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_202
timestamp 1698431365
transform 1 0 23968 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_237
timestamp 1698431365
transform 1 0 27888 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_247
timestamp 1698431365
transform 1 0 29008 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_255
timestamp 1698431365
transform 1 0 29904 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_259
timestamp 1698431365
transform 1 0 30352 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_261
timestamp 1698431365
transform 1 0 30576 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_266
timestamp 1698431365
transform 1 0 31136 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_282
timestamp 1698431365
transform 1 0 32928 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_327
timestamp 1698431365
transform 1 0 37968 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_329
timestamp 1698431365
transform 1 0 38192 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_370
timestamp 1698431365
transform 1 0 42784 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_372
timestamp 1698431365
transform 1 0 43008 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_381
timestamp 1698431365
transform 1 0 44016 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_397
timestamp 1698431365
transform 1 0 45808 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_436
timestamp 1698431365
transform 1 0 50176 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_440
timestamp 1698431365
transform 1 0 50624 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_444
timestamp 1698431365
transform 1 0 51072 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_448
timestamp 1698431365
transform 1 0 51520 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_452
timestamp 1698431365
transform 1 0 51968 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_454
timestamp 1698431365
transform 1 0 52192 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_457
timestamp 1698431365
transform 1 0 52528 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_466
timestamp 1698431365
transform 1 0 53536 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_470
timestamp 1698431365
transform 1 0 53984 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_474
timestamp 1698431365
transform 1 0 54432 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_506
timestamp 1698431365
transform 1 0 58016 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_522
timestamp 1698431365
transform 1 0 59808 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_524
timestamp 1698431365
transform 1 0 60032 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_527
timestamp 1698431365
transform 1 0 60368 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_591
timestamp 1698431365
transform 1 0 67536 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_597
timestamp 1698431365
transform 1 0 68208 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_613
timestamp 1698431365
transform 1 0 70000 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_621
timestamp 1698431365
transform 1 0 70896 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_625
timestamp 1698431365
transform 1 0 71344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_629
timestamp 1698431365
transform 1 0 71792 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_663
timestamp 1698431365
transform 1 0 75600 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_667
timestamp 1698431365
transform 1 0 76048 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_669
timestamp 1698431365
transform 1 0 76272 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_678
timestamp 1698431365
transform 1 0 77280 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_685
timestamp 1698431365
transform 1 0 78064 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_687
timestamp 1698431365
transform 1 0 78288 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_8
timestamp 1698431365
transform 1 0 2240 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_12
timestamp 1698431365
transform 1 0 2688 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_44
timestamp 1698431365
transform 1 0 6272 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_60
timestamp 1698431365
transform 1 0 8064 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_68
timestamp 1698431365
transform 1 0 8960 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_72
timestamp 1698431365
transform 1 0 9408 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_136
timestamp 1698431365
transform 1 0 16576 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_147
timestamp 1698431365
transform 1 0 17808 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_153
timestamp 1698431365
transform 1 0 18480 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_157
timestamp 1698431365
transform 1 0 18928 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_166
timestamp 1698431365
transform 1 0 19936 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_197
timestamp 1698431365
transform 1 0 23408 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_199
timestamp 1698431365
transform 1 0 23632 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_205
timestamp 1698431365
transform 1 0 24304 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_209
timestamp 1698431365
transform 1 0 24752 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_220
timestamp 1698431365
transform 1 0 25984 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_265
timestamp 1698431365
transform 1 0 31024 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_273
timestamp 1698431365
transform 1 0 31920 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_277
timestamp 1698431365
transform 1 0 32368 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_279
timestamp 1698431365
transform 1 0 32592 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_282
timestamp 1698431365
transform 1 0 32928 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_286
timestamp 1698431365
transform 1 0 33376 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_290
timestamp 1698431365
transform 1 0 33824 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_346
timestamp 1698431365
transform 1 0 40096 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_372
timestamp 1698431365
transform 1 0 43008 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_419
timestamp 1698431365
transform 1 0 48272 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_422
timestamp 1698431365
transform 1 0 48608 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_426
timestamp 1698431365
transform 1 0 49056 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_430
timestamp 1698431365
transform 1 0 49504 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_434
timestamp 1698431365
transform 1 0 49952 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_438
timestamp 1698431365
transform 1 0 50400 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_442
timestamp 1698431365
transform 1 0 50848 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_446
timestamp 1698431365
transform 1 0 51296 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_478
timestamp 1698431365
transform 1 0 54880 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_486
timestamp 1698431365
transform 1 0 55776 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_492
timestamp 1698431365
transform 1 0 56448 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_556
timestamp 1698431365
transform 1 0 63616 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_562
timestamp 1698431365
transform 1 0 64288 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_626
timestamp 1698431365
transform 1 0 71456 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_647
timestamp 1698431365
transform 1 0 73808 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_653
timestamp 1698431365
transform 1 0 74480 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_655
timestamp 1698431365
transform 1 0 74704 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_671
timestamp 1698431365
transform 1 0 76496 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_685
timestamp 1698431365
transform 1 0 78064 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_687
timestamp 1698431365
transform 1 0 78288 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_8
timestamp 1698431365
transform 1 0 2240 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_12
timestamp 1698431365
transform 1 0 2688 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_28
timestamp 1698431365
transform 1 0 4480 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_32
timestamp 1698431365
transform 1 0 4928 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_34
timestamp 1698431365
transform 1 0 5152 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_37
timestamp 1698431365
transform 1 0 5488 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_101
timestamp 1698431365
transform 1 0 12656 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_107
timestamp 1698431365
transform 1 0 13328 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_139
timestamp 1698431365
transform 1 0 16912 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_156
timestamp 1698431365
transform 1 0 18816 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_160
timestamp 1698431365
transform 1 0 19264 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_174
timestamp 1698431365
transform 1 0 20832 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_185
timestamp 1698431365
transform 1 0 22064 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_189
timestamp 1698431365
transform 1 0 22512 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_193
timestamp 1698431365
transform 1 0 22960 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_195
timestamp 1698431365
transform 1 0 23184 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_232
timestamp 1698431365
transform 1 0 27328 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_241
timestamp 1698431365
transform 1 0 28336 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_247
timestamp 1698431365
transform 1 0 29008 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_279
timestamp 1698431365
transform 1 0 32592 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_287
timestamp 1698431365
transform 1 0 33488 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_291
timestamp 1698431365
transform 1 0 33936 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_295
timestamp 1698431365
transform 1 0 34384 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_299
timestamp 1698431365
transform 1 0 34832 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_303
timestamp 1698431365
transform 1 0 35280 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_312
timestamp 1698431365
transform 1 0 36288 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_314
timestamp 1698431365
transform 1 0 36512 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_317
timestamp 1698431365
transform 1 0 36848 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_396
timestamp 1698431365
transform 1 0 45696 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_398
timestamp 1698431365
transform 1 0 45920 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_417
timestamp 1698431365
transform 1 0 48048 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_421
timestamp 1698431365
transform 1 0 48496 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_425
timestamp 1698431365
transform 1 0 48944 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_429
timestamp 1698431365
transform 1 0 49392 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_433
timestamp 1698431365
transform 1 0 49840 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_449
timestamp 1698431365
transform 1 0 51632 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_453
timestamp 1698431365
transform 1 0 52080 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_457
timestamp 1698431365
transform 1 0 52528 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_521
timestamp 1698431365
transform 1 0 59696 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_527
timestamp 1698431365
transform 1 0 60368 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_591
timestamp 1698431365
transform 1 0 67536 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_597
timestamp 1698431365
transform 1 0 68208 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_629
timestamp 1698431365
transform 1 0 71792 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_648
timestamp 1698431365
transform 1 0 73920 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_650
timestamp 1698431365
transform 1 0 74144 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_679
timestamp 1698431365
transform 1 0 77392 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_681
timestamp 1698431365
transform 1 0 77616 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_2
timestamp 1698431365
transform 1 0 1568 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_66
timestamp 1698431365
transform 1 0 8736 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_72
timestamp 1698431365
transform 1 0 9408 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_136
timestamp 1698431365
transform 1 0 16576 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_206
timestamp 1698431365
transform 1 0 24416 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_220
timestamp 1698431365
transform 1 0 25984 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_228
timestamp 1698431365
transform 1 0 26880 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_262
timestamp 1698431365
transform 1 0 30688 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_278
timestamp 1698431365
transform 1 0 32480 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_282
timestamp 1698431365
transform 1 0 32928 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_298
timestamp 1698431365
transform 1 0 34720 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_343
timestamp 1698431365
transform 1 0 39760 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_412
timestamp 1698431365
transform 1 0 47488 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_416
timestamp 1698431365
transform 1 0 47936 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_422
timestamp 1698431365
transform 1 0 48608 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_426
timestamp 1698431365
transform 1 0 49056 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_492
timestamp 1698431365
transform 1 0 56448 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_524
timestamp 1698431365
transform 1 0 60032 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_540
timestamp 1698431365
transform 1 0 61824 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_556
timestamp 1698431365
transform 1 0 63616 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_562
timestamp 1698431365
transform 1 0 64288 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_594
timestamp 1698431365
transform 1 0 67872 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_610
timestamp 1698431365
transform 1 0 69664 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_618
timestamp 1698431365
transform 1 0 70560 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_622
timestamp 1698431365
transform 1 0 71008 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_626
timestamp 1698431365
transform 1 0 71456 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_647
timestamp 1698431365
transform 1 0 73808 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_651
timestamp 1698431365
transform 1 0 74256 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_671
timestamp 1698431365
transform 1 0 76496 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_685
timestamp 1698431365
transform 1 0 78064 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_687
timestamp 1698431365
transform 1 0 78288 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_8
timestamp 1698431365
transform 1 0 2240 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_12
timestamp 1698431365
transform 1 0 2688 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_28
timestamp 1698431365
transform 1 0 4480 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_32
timestamp 1698431365
transform 1 0 4928 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_34
timestamp 1698431365
transform 1 0 5152 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_37
timestamp 1698431365
transform 1 0 5488 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_101
timestamp 1698431365
transform 1 0 12656 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_107
timestamp 1698431365
transform 1 0 13328 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_171
timestamp 1698431365
transform 1 0 20496 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_177
timestamp 1698431365
transform 1 0 21168 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_193
timestamp 1698431365
transform 1 0 22960 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_197
timestamp 1698431365
transform 1 0 23408 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_206
timestamp 1698431365
transform 1 0 24416 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_222
timestamp 1698431365
transform 1 0 26208 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_226
timestamp 1698431365
transform 1 0 26656 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_232
timestamp 1698431365
transform 1 0 27328 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_240
timestamp 1698431365
transform 1 0 28224 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_244
timestamp 1698431365
transform 1 0 28672 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_247
timestamp 1698431365
transform 1 0 29008 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_279
timestamp 1698431365
transform 1 0 32592 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_295
timestamp 1698431365
transform 1 0 34384 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_303
timestamp 1698431365
transform 1 0 35280 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_317
timestamp 1698431365
transform 1 0 36848 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_359
timestamp 1698431365
transform 1 0 41552 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_379
timestamp 1698431365
transform 1 0 43792 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_383
timestamp 1698431365
transform 1 0 44240 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_410
timestamp 1698431365
transform 1 0 47264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_414
timestamp 1698431365
transform 1 0 47712 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_418
timestamp 1698431365
transform 1 0 48160 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_450
timestamp 1698431365
transform 1 0 51744 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_454
timestamp 1698431365
transform 1 0 52192 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_457
timestamp 1698431365
transform 1 0 52528 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_521
timestamp 1698431365
transform 1 0 59696 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_527
timestamp 1698431365
transform 1 0 60368 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_543
timestamp 1698431365
transform 1 0 62160 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_547
timestamp 1698431365
transform 1 0 62608 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_556
timestamp 1698431365
transform 1 0 63616 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_588
timestamp 1698431365
transform 1 0 67200 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_592
timestamp 1698431365
transform 1 0 67648 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_594
timestamp 1698431365
transform 1 0 67872 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_597
timestamp 1698431365
transform 1 0 68208 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_613
timestamp 1698431365
transform 1 0 70000 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_617
timestamp 1698431365
transform 1 0 70448 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_667
timestamp 1698431365
transform 1 0 76048 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_687
timestamp 1698431365
transform 1 0 78288 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_8
timestamp 1698431365
transform 1 0 2240 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_12
timestamp 1698431365
transform 1 0 2688 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_44
timestamp 1698431365
transform 1 0 6272 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_60
timestamp 1698431365
transform 1 0 8064 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_68
timestamp 1698431365
transform 1 0 8960 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_72
timestamp 1698431365
transform 1 0 9408 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_136
timestamp 1698431365
transform 1 0 16576 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_142
timestamp 1698431365
transform 1 0 17248 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_206
timestamp 1698431365
transform 1 0 24416 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_212
timestamp 1698431365
transform 1 0 25088 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_276
timestamp 1698431365
transform 1 0 32256 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_282
timestamp 1698431365
transform 1 0 32928 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_298
timestamp 1698431365
transform 1 0 34720 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_300
timestamp 1698431365
transform 1 0 34944 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_316
timestamp 1698431365
transform 1 0 36736 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_318
timestamp 1698431365
transform 1 0 36960 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_340
timestamp 1698431365
transform 1 0 39424 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_352
timestamp 1698431365
transform 1 0 40768 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_366
timestamp 1698431365
transform 1 0 42336 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_370
timestamp 1698431365
transform 1 0 42784 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_384
timestamp 1698431365
transform 1 0 44352 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_392
timestamp 1698431365
transform 1 0 45248 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_394
timestamp 1698431365
transform 1 0 45472 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_417
timestamp 1698431365
transform 1 0 48048 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_419
timestamp 1698431365
transform 1 0 48272 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_432
timestamp 1698431365
transform 1 0 49728 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_436
timestamp 1698431365
transform 1 0 50176 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_440
timestamp 1698431365
transform 1 0 50624 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_472
timestamp 1698431365
transform 1 0 54208 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_488
timestamp 1698431365
transform 1 0 56000 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_492
timestamp 1698431365
transform 1 0 56448 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_556
timestamp 1698431365
transform 1 0 63616 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_562
timestamp 1698431365
transform 1 0 64288 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_594
timestamp 1698431365
transform 1 0 67872 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_610
timestamp 1698431365
transform 1 0 69664 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_618
timestamp 1698431365
transform 1 0 70560 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_627
timestamp 1698431365
transform 1 0 71568 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_629
timestamp 1698431365
transform 1 0 71792 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_632
timestamp 1698431365
transform 1 0 72128 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_636
timestamp 1698431365
transform 1 0 72576 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_640
timestamp 1698431365
transform 1 0 73024 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_671
timestamp 1698431365
transform 1 0 76496 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_673
timestamp 1698431365
transform 1 0 76720 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_8
timestamp 1698431365
transform 1 0 2240 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_12
timestamp 1698431365
transform 1 0 2688 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_28
timestamp 1698431365
transform 1 0 4480 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_32
timestamp 1698431365
transform 1 0 4928 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_34
timestamp 1698431365
transform 1 0 5152 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_37
timestamp 1698431365
transform 1 0 5488 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_101
timestamp 1698431365
transform 1 0 12656 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_107
timestamp 1698431365
transform 1 0 13328 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_171
timestamp 1698431365
transform 1 0 20496 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_177
timestamp 1698431365
transform 1 0 21168 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_241
timestamp 1698431365
transform 1 0 28336 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_247
timestamp 1698431365
transform 1 0 29008 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_279
timestamp 1698431365
transform 1 0 32592 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_287
timestamp 1698431365
transform 1 0 33488 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_325
timestamp 1698431365
transform 1 0 37744 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_374
timestamp 1698431365
transform 1 0 43232 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_378
timestamp 1698431365
transform 1 0 43680 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_381
timestamp 1698431365
transform 1 0 44016 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_391
timestamp 1698431365
transform 1 0 45136 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_395
timestamp 1698431365
transform 1 0 45584 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_399
timestamp 1698431365
transform 1 0 46032 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_416
timestamp 1698431365
transform 1 0 47936 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_424
timestamp 1698431365
transform 1 0 48832 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_435
timestamp 1698431365
transform 1 0 50064 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_439
timestamp 1698431365
transform 1 0 50512 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_443
timestamp 1698431365
transform 1 0 50960 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_451
timestamp 1698431365
transform 1 0 51856 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_457
timestamp 1698431365
transform 1 0 52528 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_521
timestamp 1698431365
transform 1 0 59696 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_527
timestamp 1698431365
transform 1 0 60368 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_591
timestamp 1698431365
transform 1 0 67536 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_597
timestamp 1698431365
transform 1 0 68208 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_613
timestamp 1698431365
transform 1 0 70000 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_617
timestamp 1698431365
transform 1 0 70448 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_626
timestamp 1698431365
transform 1 0 71456 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_628
timestamp 1698431365
transform 1 0 71680 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_631
timestamp 1698431365
transform 1 0 72016 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_635
timestamp 1698431365
transform 1 0 72464 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_647
timestamp 1698431365
transform 1 0 73808 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_649
timestamp 1698431365
transform 1 0 74032 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_656
timestamp 1698431365
transform 1 0 74816 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_658
timestamp 1698431365
transform 1 0 75040 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_685
timestamp 1698431365
transform 1 0 78064 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_687
timestamp 1698431365
transform 1 0 78288 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_2
timestamp 1698431365
transform 1 0 1568 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_66
timestamp 1698431365
transform 1 0 8736 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_72
timestamp 1698431365
transform 1 0 9408 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_136
timestamp 1698431365
transform 1 0 16576 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_142
timestamp 1698431365
transform 1 0 17248 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_206
timestamp 1698431365
transform 1 0 24416 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_212
timestamp 1698431365
transform 1 0 25088 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_276
timestamp 1698431365
transform 1 0 32256 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_282
timestamp 1698431365
transform 1 0 32928 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_313
timestamp 1698431365
transform 1 0 36400 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_317
timestamp 1698431365
transform 1 0 36848 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_321
timestamp 1698431365
transform 1 0 37296 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_338
timestamp 1698431365
transform 1 0 39200 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_342
timestamp 1698431365
transform 1 0 39648 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_346
timestamp 1698431365
transform 1 0 40096 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_365
timestamp 1698431365
transform 1 0 42224 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_369
timestamp 1698431365
transform 1 0 42672 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_385
timestamp 1698431365
transform 1 0 44464 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_392
timestamp 1698431365
transform 1 0 45248 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_408
timestamp 1698431365
transform 1 0 47040 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_416
timestamp 1698431365
transform 1 0 47936 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_422
timestamp 1698431365
transform 1 0 48608 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_486
timestamp 1698431365
transform 1 0 55776 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_492
timestamp 1698431365
transform 1 0 56448 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_556
timestamp 1698431365
transform 1 0 63616 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_31_562
timestamp 1698431365
transform 1 0 64288 0 -1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_594
timestamp 1698431365
transform 1 0 67872 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_610
timestamp 1698431365
transform 1 0 69664 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_614
timestamp 1698431365
transform 1 0 70112 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_623
timestamp 1698431365
transform 1 0 71120 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_627
timestamp 1698431365
transform 1 0 71568 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_632
timestamp 1698431365
transform 1 0 72128 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_662
timestamp 1698431365
transform 1 0 75488 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_678
timestamp 1698431365
transform 1 0 77280 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_8
timestamp 1698431365
transform 1 0 2240 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_12
timestamp 1698431365
transform 1 0 2688 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_28
timestamp 1698431365
transform 1 0 4480 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_32
timestamp 1698431365
transform 1 0 4928 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_34
timestamp 1698431365
transform 1 0 5152 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_37
timestamp 1698431365
transform 1 0 5488 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_101
timestamp 1698431365
transform 1 0 12656 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_107
timestamp 1698431365
transform 1 0 13328 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_171
timestamp 1698431365
transform 1 0 20496 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_177
timestamp 1698431365
transform 1 0 21168 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_241
timestamp 1698431365
transform 1 0 28336 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_247
timestamp 1698431365
transform 1 0 29008 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_311
timestamp 1698431365
transform 1 0 36176 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_317
timestamp 1698431365
transform 1 0 36848 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_321
timestamp 1698431365
transform 1 0 37296 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_337
timestamp 1698431365
transform 1 0 39088 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_355
timestamp 1698431365
transform 1 0 41104 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_371
timestamp 1698431365
transform 1 0 42896 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_379
timestamp 1698431365
transform 1 0 43792 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_383
timestamp 1698431365
transform 1 0 44240 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_387
timestamp 1698431365
transform 1 0 44688 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_451
timestamp 1698431365
transform 1 0 51856 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_457
timestamp 1698431365
transform 1 0 52528 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_521
timestamp 1698431365
transform 1 0 59696 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_527
timestamp 1698431365
transform 1 0 60368 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_591
timestamp 1698431365
transform 1 0 67536 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_597
timestamp 1698431365
transform 1 0 68208 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_613
timestamp 1698431365
transform 1 0 70000 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_621
timestamp 1698431365
transform 1 0 70896 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_625
timestamp 1698431365
transform 1 0 71344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_629
timestamp 1698431365
transform 1 0 71792 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_639
timestamp 1698431365
transform 1 0 72912 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_641
timestamp 1698431365
transform 1 0 73136 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_644
timestamp 1698431365
transform 1 0 73472 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_648
timestamp 1698431365
transform 1 0 73920 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_655
timestamp 1698431365
transform 1 0 74704 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_675
timestamp 1698431365
transform 1 0 76944 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_8
timestamp 1698431365
transform 1 0 2240 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_33_12
timestamp 1698431365
transform 1 0 2688 0 -1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_33_44
timestamp 1698431365
transform 1 0 6272 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_60
timestamp 1698431365
transform 1 0 8064 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_68
timestamp 1698431365
transform 1 0 8960 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_72
timestamp 1698431365
transform 1 0 9408 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_136
timestamp 1698431365
transform 1 0 16576 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_142
timestamp 1698431365
transform 1 0 17248 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_206
timestamp 1698431365
transform 1 0 24416 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_212
timestamp 1698431365
transform 1 0 25088 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_276
timestamp 1698431365
transform 1 0 32256 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_282
timestamp 1698431365
transform 1 0 32928 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_346
timestamp 1698431365
transform 1 0 40096 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_33_352
timestamp 1698431365
transform 1 0 40768 0 -1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_384
timestamp 1698431365
transform 1 0 44352 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_386
timestamp 1698431365
transform 1 0 44576 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_33_393
timestamp 1698431365
transform 1 0 45360 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_409
timestamp 1698431365
transform 1 0 47152 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_417
timestamp 1698431365
transform 1 0 48048 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_419
timestamp 1698431365
transform 1 0 48272 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_422
timestamp 1698431365
transform 1 0 48608 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_486
timestamp 1698431365
transform 1 0 55776 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_492
timestamp 1698431365
transform 1 0 56448 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_556
timestamp 1698431365
transform 1 0 63616 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_33_562
timestamp 1698431365
transform 1 0 64288 0 -1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_33_594
timestamp 1698431365
transform 1 0 67872 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_610
timestamp 1698431365
transform 1 0 69664 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_618
timestamp 1698431365
transform 1 0 70560 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_648
timestamp 1698431365
transform 1 0 73920 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_650
timestamp 1698431365
transform 1 0 74144 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_659
timestamp 1698431365
transform 1 0 75152 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_674
timestamp 1698431365
transform 1 0 76832 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_2
timestamp 1698431365
transform 1 0 1568 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_34
timestamp 1698431365
transform 1 0 5152 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_37
timestamp 1698431365
transform 1 0 5488 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_101
timestamp 1698431365
transform 1 0 12656 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_107
timestamp 1698431365
transform 1 0 13328 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_171
timestamp 1698431365
transform 1 0 20496 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_177
timestamp 1698431365
transform 1 0 21168 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_241
timestamp 1698431365
transform 1 0 28336 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_247
timestamp 1698431365
transform 1 0 29008 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_311
timestamp 1698431365
transform 1 0 36176 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_317
timestamp 1698431365
transform 1 0 36848 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_381
timestamp 1698431365
transform 1 0 44016 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_391
timestamp 1698431365
transform 1 0 45136 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_395
timestamp 1698431365
transform 1 0 45584 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_397
timestamp 1698431365
transform 1 0 45808 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_34_412
timestamp 1698431365
transform 1 0 47488 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_428
timestamp 1698431365
transform 1 0 49280 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_436
timestamp 1698431365
transform 1 0 50176 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_438
timestamp 1698431365
transform 1 0 50400 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_448
timestamp 1698431365
transform 1 0 51520 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_452
timestamp 1698431365
transform 1 0 51968 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_454
timestamp 1698431365
transform 1 0 52192 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_457
timestamp 1698431365
transform 1 0 52528 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_521
timestamp 1698431365
transform 1 0 59696 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_527
timestamp 1698431365
transform 1 0 60368 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_591
timestamp 1698431365
transform 1 0 67536 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_34_597
timestamp 1698431365
transform 1 0 68208 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_613
timestamp 1698431365
transform 1 0 70000 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_621
timestamp 1698431365
transform 1 0 70896 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_625
timestamp 1698431365
transform 1 0 71344 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_632
timestamp 1698431365
transform 1 0 72128 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_644
timestamp 1698431365
transform 1 0 73472 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_646
timestamp 1698431365
transform 1 0 73696 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_662
timestamp 1698431365
transform 1 0 75488 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_664
timestamp 1698431365
transform 1 0 75712 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_667
timestamp 1698431365
transform 1 0 76048 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_676
timestamp 1698431365
transform 1 0 77056 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_678
timestamp 1698431365
transform 1 0 77280 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_685
timestamp 1698431365
transform 1 0 78064 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_687
timestamp 1698431365
transform 1 0 78288 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_8
timestamp 1698431365
transform 1 0 2240 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_35_12
timestamp 1698431365
transform 1 0 2688 0 -1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_35_44
timestamp 1698431365
transform 1 0 6272 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_60
timestamp 1698431365
transform 1 0 8064 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_68
timestamp 1698431365
transform 1 0 8960 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_72
timestamp 1698431365
transform 1 0 9408 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_136
timestamp 1698431365
transform 1 0 16576 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_142
timestamp 1698431365
transform 1 0 17248 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_206
timestamp 1698431365
transform 1 0 24416 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_212
timestamp 1698431365
transform 1 0 25088 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_276
timestamp 1698431365
transform 1 0 32256 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_282
timestamp 1698431365
transform 1 0 32928 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_346
timestamp 1698431365
transform 1 0 40096 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_35_352
timestamp 1698431365
transform 1 0 40768 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_368
timestamp 1698431365
transform 1 0 42560 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_376
timestamp 1698431365
transform 1 0 43456 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_380
timestamp 1698431365
transform 1 0 43904 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_382
timestamp 1698431365
transform 1 0 44128 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_389
timestamp 1698431365
transform 1 0 44912 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_391
timestamp 1698431365
transform 1 0 45136 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_414
timestamp 1698431365
transform 1 0 47712 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_418
timestamp 1698431365
transform 1 0 48160 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_422
timestamp 1698431365
transform 1 0 48608 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_430
timestamp 1698431365
transform 1 0 49504 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_452
timestamp 1698431365
transform 1 0 51968 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_456
timestamp 1698431365
transform 1 0 52416 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_35_460
timestamp 1698431365
transform 1 0 52864 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_476
timestamp 1698431365
transform 1 0 54656 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_484
timestamp 1698431365
transform 1 0 55552 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_488
timestamp 1698431365
transform 1 0 56000 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_492
timestamp 1698431365
transform 1 0 56448 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_556
timestamp 1698431365
transform 1 0 63616 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_35_562
timestamp 1698431365
transform 1 0 64288 0 -1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_35_594
timestamp 1698431365
transform 1 0 67872 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_610
timestamp 1698431365
transform 1 0 69664 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_618
timestamp 1698431365
transform 1 0 70560 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_622
timestamp 1698431365
transform 1 0 71008 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_626
timestamp 1698431365
transform 1 0 71456 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_632
timestamp 1698431365
transform 1 0 72128 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_638
timestamp 1698431365
transform 1 0 72800 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_642
timestamp 1698431365
transform 1 0 73248 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_645
timestamp 1698431365
transform 1 0 73584 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_683
timestamp 1698431365
transform 1 0 77840 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_687
timestamp 1698431365
transform 1 0 78288 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_8
timestamp 1698431365
transform 1 0 2240 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_36_12
timestamp 1698431365
transform 1 0 2688 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_28
timestamp 1698431365
transform 1 0 4480 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_32
timestamp 1698431365
transform 1 0 4928 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_34
timestamp 1698431365
transform 1 0 5152 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_37
timestamp 1698431365
transform 1 0 5488 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_101
timestamp 1698431365
transform 1 0 12656 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_107
timestamp 1698431365
transform 1 0 13328 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_171
timestamp 1698431365
transform 1 0 20496 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_177
timestamp 1698431365
transform 1 0 21168 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_241
timestamp 1698431365
transform 1 0 28336 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_247
timestamp 1698431365
transform 1 0 29008 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_311
timestamp 1698431365
transform 1 0 36176 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_317
timestamp 1698431365
transform 1 0 36848 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_381
timestamp 1698431365
transform 1 0 44016 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_387
timestamp 1698431365
transform 1 0 44688 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_392
timestamp 1698431365
transform 1 0 45248 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_396
timestamp 1698431365
transform 1 0 45696 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_406
timestamp 1698431365
transform 1 0 46816 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_438
timestamp 1698431365
transform 1 0 50400 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_442
timestamp 1698431365
transform 1 0 50848 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_452
timestamp 1698431365
transform 1 0 51968 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_454
timestamp 1698431365
transform 1 0 52192 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_457
timestamp 1698431365
transform 1 0 52528 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_461
timestamp 1698431365
transform 1 0 52976 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_527
timestamp 1698431365
transform 1 0 60368 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_591
timestamp 1698431365
transform 1 0 67536 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_36_597
timestamp 1698431365
transform 1 0 68208 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_613
timestamp 1698431365
transform 1 0 70000 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_617
timestamp 1698431365
transform 1 0 70448 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_619
timestamp 1698431365
transform 1 0 70672 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_644
timestamp 1698431365
transform 1 0 73472 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_648
timestamp 1698431365
transform 1 0 73920 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_657
timestamp 1698431365
transform 1 0 74928 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_661
timestamp 1698431365
transform 1 0 75376 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_667
timestamp 1698431365
transform 1 0 76048 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_669
timestamp 1698431365
transform 1 0 76272 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_678
timestamp 1698431365
transform 1 0 77280 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_685
timestamp 1698431365
transform 1 0 78064 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_687
timestamp 1698431365
transform 1 0 78288 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_2
timestamp 1698431365
transform 1 0 1568 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_66
timestamp 1698431365
transform 1 0 8736 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_72
timestamp 1698431365
transform 1 0 9408 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_136
timestamp 1698431365
transform 1 0 16576 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_142
timestamp 1698431365
transform 1 0 17248 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_206
timestamp 1698431365
transform 1 0 24416 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_212
timestamp 1698431365
transform 1 0 25088 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_276
timestamp 1698431365
transform 1 0 32256 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_282
timestamp 1698431365
transform 1 0 32928 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_346
timestamp 1698431365
transform 1 0 40096 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_37_352
timestamp 1698431365
transform 1 0 40768 0 -1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_384
timestamp 1698431365
transform 1 0 44352 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_392
timestamp 1698431365
transform 1 0 45248 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_37_402
timestamp 1698431365
transform 1 0 46368 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_418
timestamp 1698431365
transform 1 0 48160 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_422
timestamp 1698431365
transform 1 0 48608 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_486
timestamp 1698431365
transform 1 0 55776 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_492
timestamp 1698431365
transform 1 0 56448 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_556
timestamp 1698431365
transform 1 0 63616 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_37_562
timestamp 1698431365
transform 1 0 64288 0 -1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_37_594
timestamp 1698431365
transform 1 0 67872 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_610
timestamp 1698431365
transform 1 0 69664 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_618
timestamp 1698431365
transform 1 0 70560 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_632
timestamp 1698431365
transform 1 0 72128 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_639
timestamp 1698431365
transform 1 0 72912 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_643
timestamp 1698431365
transform 1 0 73360 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_675
timestamp 1698431365
transform 1 0 76944 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_685
timestamp 1698431365
transform 1 0 78064 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_687
timestamp 1698431365
transform 1 0 78288 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_8
timestamp 1698431365
transform 1 0 2240 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_38_12
timestamp 1698431365
transform 1 0 2688 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_28
timestamp 1698431365
transform 1 0 4480 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_32
timestamp 1698431365
transform 1 0 4928 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_34
timestamp 1698431365
transform 1 0 5152 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_37
timestamp 1698431365
transform 1 0 5488 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_101
timestamp 1698431365
transform 1 0 12656 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_107
timestamp 1698431365
transform 1 0 13328 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_171
timestamp 1698431365
transform 1 0 20496 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_177
timestamp 1698431365
transform 1 0 21168 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_241
timestamp 1698431365
transform 1 0 28336 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_247
timestamp 1698431365
transform 1 0 29008 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_311
timestamp 1698431365
transform 1 0 36176 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_317
timestamp 1698431365
transform 1 0 36848 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_381
timestamp 1698431365
transform 1 0 44016 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_387
timestamp 1698431365
transform 1 0 44688 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_389
timestamp 1698431365
transform 1 0 44912 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_394
timestamp 1698431365
transform 1 0 45472 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_410
timestamp 1698431365
transform 1 0 47264 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_442
timestamp 1698431365
transform 1 0 50848 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_450
timestamp 1698431365
transform 1 0 51744 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_454
timestamp 1698431365
transform 1 0 52192 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_457
timestamp 1698431365
transform 1 0 52528 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_459
timestamp 1698431365
transform 1 0 52752 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_469
timestamp 1698431365
transform 1 0 53872 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_473
timestamp 1698431365
transform 1 0 54320 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_38_505
timestamp 1698431365
transform 1 0 57904 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_521
timestamp 1698431365
transform 1 0 59696 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_527
timestamp 1698431365
transform 1 0 60368 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_591
timestamp 1698431365
transform 1 0 67536 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_38_597
timestamp 1698431365
transform 1 0 68208 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_613
timestamp 1698431365
transform 1 0 70000 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_621
timestamp 1698431365
transform 1 0 70896 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_624
timestamp 1698431365
transform 1 0 71232 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_628
timestamp 1698431365
transform 1 0 71680 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_632
timestamp 1698431365
transform 1 0 72128 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_634
timestamp 1698431365
transform 1 0 72352 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_641
timestamp 1698431365
transform 1 0 73136 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_643
timestamp 1698431365
transform 1 0 73360 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_667
timestamp 1698431365
transform 1 0 76048 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_669
timestamp 1698431365
transform 1 0 76272 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_684
timestamp 1698431365
transform 1 0 77952 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_8
timestamp 1698431365
transform 1 0 2240 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_39_12
timestamp 1698431365
transform 1 0 2688 0 -1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_39_44
timestamp 1698431365
transform 1 0 6272 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_60
timestamp 1698431365
transform 1 0 8064 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_68
timestamp 1698431365
transform 1 0 8960 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_72
timestamp 1698431365
transform 1 0 9408 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_136
timestamp 1698431365
transform 1 0 16576 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_142
timestamp 1698431365
transform 1 0 17248 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_206
timestamp 1698431365
transform 1 0 24416 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_212
timestamp 1698431365
transform 1 0 25088 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_276
timestamp 1698431365
transform 1 0 32256 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_282
timestamp 1698431365
transform 1 0 32928 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_346
timestamp 1698431365
transform 1 0 40096 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_39_352
timestamp 1698431365
transform 1 0 40768 0 -1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_384
timestamp 1698431365
transform 1 0 44352 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_392
timestamp 1698431365
transform 1 0 45248 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_396
timestamp 1698431365
transform 1 0 45696 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_405
timestamp 1698431365
transform 1 0 46704 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_413
timestamp 1698431365
transform 1 0 47600 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_417
timestamp 1698431365
transform 1 0 48048 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_419
timestamp 1698431365
transform 1 0 48272 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_422
timestamp 1698431365
transform 1 0 48608 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_486
timestamp 1698431365
transform 1 0 55776 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_492
timestamp 1698431365
transform 1 0 56448 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_556
timestamp 1698431365
transform 1 0 63616 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_39_562
timestamp 1698431365
transform 1 0 64288 0 -1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_39_594
timestamp 1698431365
transform 1 0 67872 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_610
timestamp 1698431365
transform 1 0 69664 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_618
timestamp 1698431365
transform 1 0 70560 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_648
timestamp 1698431365
transform 1 0 73920 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_684
timestamp 1698431365
transform 1 0 77952 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_8
timestamp 1698431365
transform 1 0 2240 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_40_12
timestamp 1698431365
transform 1 0 2688 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_28
timestamp 1698431365
transform 1 0 4480 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_32
timestamp 1698431365
transform 1 0 4928 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_34
timestamp 1698431365
transform 1 0 5152 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_37
timestamp 1698431365
transform 1 0 5488 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_101
timestamp 1698431365
transform 1 0 12656 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_107
timestamp 1698431365
transform 1 0 13328 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_171
timestamp 1698431365
transform 1 0 20496 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_177
timestamp 1698431365
transform 1 0 21168 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_241
timestamp 1698431365
transform 1 0 28336 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_247
timestamp 1698431365
transform 1 0 29008 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_311
timestamp 1698431365
transform 1 0 36176 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_317
timestamp 1698431365
transform 1 0 36848 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_381
timestamp 1698431365
transform 1 0 44016 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_387
timestamp 1698431365
transform 1 0 44688 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_389
timestamp 1698431365
transform 1 0 44912 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_394
timestamp 1698431365
transform 1 0 45472 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_412
timestamp 1698431365
transform 1 0 47488 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_444
timestamp 1698431365
transform 1 0 51072 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_452
timestamp 1698431365
transform 1 0 51968 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_454
timestamp 1698431365
transform 1 0 52192 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_457
timestamp 1698431365
transform 1 0 52528 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_465
timestamp 1698431365
transform 1 0 53424 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_475
timestamp 1698431365
transform 1 0 54544 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_477
timestamp 1698431365
transform 1 0 54768 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_480
timestamp 1698431365
transform 1 0 55104 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_484
timestamp 1698431365
transform 1 0 55552 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_516
timestamp 1698431365
transform 1 0 59136 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_524
timestamp 1698431365
transform 1 0 60032 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_527
timestamp 1698431365
transform 1 0 60368 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_591
timestamp 1698431365
transform 1 0 67536 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_40_597
timestamp 1698431365
transform 1 0 68208 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_613
timestamp 1698431365
transform 1 0 70000 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_621
timestamp 1698431365
transform 1 0 70896 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_625
timestamp 1698431365
transform 1 0 71344 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_627
timestamp 1698431365
transform 1 0 71568 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_630
timestamp 1698431365
transform 1 0 71904 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_634
timestamp 1698431365
transform 1 0 72352 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_652
timestamp 1698431365
transform 1 0 74368 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_2
timestamp 1698431365
transform 1 0 1568 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_66
timestamp 1698431365
transform 1 0 8736 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_72
timestamp 1698431365
transform 1 0 9408 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_136
timestamp 1698431365
transform 1 0 16576 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_142
timestamp 1698431365
transform 1 0 17248 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_206
timestamp 1698431365
transform 1 0 24416 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_212
timestamp 1698431365
transform 1 0 25088 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_276
timestamp 1698431365
transform 1 0 32256 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_282
timestamp 1698431365
transform 1 0 32928 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_346
timestamp 1698431365
transform 1 0 40096 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_41_352
timestamp 1698431365
transform 1 0 40768 0 -1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_384
timestamp 1698431365
transform 1 0 44352 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_386
timestamp 1698431365
transform 1 0 44576 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_393
timestamp 1698431365
transform 1 0 45360 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_395
timestamp 1698431365
transform 1 0 45584 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_41_404
timestamp 1698431365
transform 1 0 46592 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_41_422
timestamp 1698431365
transform 1 0 48608 0 -1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_454
timestamp 1698431365
transform 1 0 52192 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_462
timestamp 1698431365
transform 1 0 53088 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_466
timestamp 1698431365
transform 1 0 53536 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_468
timestamp 1698431365
transform 1 0 53760 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_487
timestamp 1698431365
transform 1 0 55888 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_489
timestamp 1698431365
transform 1 0 56112 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_492
timestamp 1698431365
transform 1 0 56448 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_496
timestamp 1698431365
transform 1 0 56896 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_41_562
timestamp 1698431365
transform 1 0 64288 0 -1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_41_594
timestamp 1698431365
transform 1 0 67872 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_610
timestamp 1698431365
transform 1 0 69664 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_618
timestamp 1698431365
transform 1 0 70560 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_622
timestamp 1698431365
transform 1 0 71008 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_626
timestamp 1698431365
transform 1 0 71456 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_644
timestamp 1698431365
transform 1 0 73472 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_646
timestamp 1698431365
transform 1 0 73696 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_663
timestamp 1698431365
transform 1 0 75600 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_665
timestamp 1698431365
transform 1 0 75824 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_8
timestamp 1698431365
transform 1 0 2240 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_12
timestamp 1698431365
transform 1 0 2688 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_28
timestamp 1698431365
transform 1 0 4480 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_32
timestamp 1698431365
transform 1 0 4928 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_34
timestamp 1698431365
transform 1 0 5152 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_37
timestamp 1698431365
transform 1 0 5488 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_101
timestamp 1698431365
transform 1 0 12656 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_107
timestamp 1698431365
transform 1 0 13328 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_171
timestamp 1698431365
transform 1 0 20496 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_177
timestamp 1698431365
transform 1 0 21168 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_241
timestamp 1698431365
transform 1 0 28336 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_247
timestamp 1698431365
transform 1 0 29008 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_311
timestamp 1698431365
transform 1 0 36176 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_317
timestamp 1698431365
transform 1 0 36848 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_381
timestamp 1698431365
transform 1 0 44016 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_387
timestamp 1698431365
transform 1 0 44688 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_393
timestamp 1698431365
transform 1 0 45360 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_397
timestamp 1698431365
transform 1 0 45808 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_429
timestamp 1698431365
transform 1 0 49392 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_445
timestamp 1698431365
transform 1 0 51184 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_453
timestamp 1698431365
transform 1 0 52080 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_457
timestamp 1698431365
transform 1 0 52528 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_521
timestamp 1698431365
transform 1 0 59696 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_527
timestamp 1698431365
transform 1 0 60368 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_591
timestamp 1698431365
transform 1 0 67536 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_597
timestamp 1698431365
transform 1 0 68208 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_601
timestamp 1698431365
transform 1 0 68656 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_604
timestamp 1698431365
transform 1 0 68992 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_608
timestamp 1698431365
transform 1 0 69440 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_612
timestamp 1698431365
transform 1 0 69888 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_620
timestamp 1698431365
transform 1 0 70784 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_622
timestamp 1698431365
transform 1 0 71008 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_625
timestamp 1698431365
transform 1 0 71344 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_629
timestamp 1698431365
transform 1 0 71792 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_633
timestamp 1698431365
transform 1 0 72240 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_645
timestamp 1698431365
transform 1 0 73584 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_649
timestamp 1698431365
transform 1 0 74032 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_8
timestamp 1698431365
transform 1 0 2240 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_43_12
timestamp 1698431365
transform 1 0 2688 0 -1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_44
timestamp 1698431365
transform 1 0 6272 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_60
timestamp 1698431365
transform 1 0 8064 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_68
timestamp 1698431365
transform 1 0 8960 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_72
timestamp 1698431365
transform 1 0 9408 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_136
timestamp 1698431365
transform 1 0 16576 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_142
timestamp 1698431365
transform 1 0 17248 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_206
timestamp 1698431365
transform 1 0 24416 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_212
timestamp 1698431365
transform 1 0 25088 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_276
timestamp 1698431365
transform 1 0 32256 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_282
timestamp 1698431365
transform 1 0 32928 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_346
timestamp 1698431365
transform 1 0 40096 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_352
timestamp 1698431365
transform 1 0 40768 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_416
timestamp 1698431365
transform 1 0 47936 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_422
timestamp 1698431365
transform 1 0 48608 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_486
timestamp 1698431365
transform 1 0 55776 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_492
timestamp 1698431365
transform 1 0 56448 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_556
timestamp 1698431365
transform 1 0 63616 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_43_562
timestamp 1698431365
transform 1 0 64288 0 -1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_594
timestamp 1698431365
transform 1 0 67872 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_628
timestamp 1698431365
transform 1 0 71680 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_656
timestamp 1698431365
transform 1 0 74816 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_2
timestamp 1698431365
transform 1 0 1568 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_12
timestamp 1698431365
transform 1 0 2688 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_44_16
timestamp 1698431365
transform 1 0 3136 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_32
timestamp 1698431365
transform 1 0 4928 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_34
timestamp 1698431365
transform 1 0 5152 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_37
timestamp 1698431365
transform 1 0 5488 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_101
timestamp 1698431365
transform 1 0 12656 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_107
timestamp 1698431365
transform 1 0 13328 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_171
timestamp 1698431365
transform 1 0 20496 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_177
timestamp 1698431365
transform 1 0 21168 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_241
timestamp 1698431365
transform 1 0 28336 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_247
timestamp 1698431365
transform 1 0 29008 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_311
timestamp 1698431365
transform 1 0 36176 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_317
timestamp 1698431365
transform 1 0 36848 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_349
timestamp 1698431365
transform 1 0 40432 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_357
timestamp 1698431365
transform 1 0 41328 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_44_360
timestamp 1698431365
transform 1 0 41664 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_376
timestamp 1698431365
transform 1 0 43456 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_384
timestamp 1698431365
transform 1 0 44352 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_387
timestamp 1698431365
transform 1 0 44688 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_451
timestamp 1698431365
transform 1 0 51856 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_457
timestamp 1698431365
transform 1 0 52528 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_521
timestamp 1698431365
transform 1 0 59696 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_527
timestamp 1698431365
transform 1 0 60368 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_44_559
timestamp 1698431365
transform 1 0 63952 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_575
timestamp 1698431365
transform 1 0 65744 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_584
timestamp 1698431365
transform 1 0 66752 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_586
timestamp 1698431365
transform 1 0 66976 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_610
timestamp 1698431365
transform 1 0 69664 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_630
timestamp 1698431365
transform 1 0 71904 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_634
timestamp 1698431365
transform 1 0 72352 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_638
timestamp 1698431365
transform 1 0 72800 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_642
timestamp 1698431365
transform 1 0 73248 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_660
timestamp 1698431365
transform 1 0 75264 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_662
timestamp 1698431365
transform 1 0 75488 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_45_28
timestamp 1698431365
transform 1 0 4480 0 -1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_60
timestamp 1698431365
transform 1 0 8064 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_68
timestamp 1698431365
transform 1 0 8960 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_72
timestamp 1698431365
transform 1 0 9408 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_136
timestamp 1698431365
transform 1 0 16576 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_142
timestamp 1698431365
transform 1 0 17248 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_206
timestamp 1698431365
transform 1 0 24416 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_212
timestamp 1698431365
transform 1 0 25088 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_276
timestamp 1698431365
transform 1 0 32256 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_282
timestamp 1698431365
transform 1 0 32928 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_346
timestamp 1698431365
transform 1 0 40096 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_352
timestamp 1698431365
transform 1 0 40768 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_372
timestamp 1698431365
transform 1 0 43008 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_376
timestamp 1698431365
transform 1 0 43456 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_45_380
timestamp 1698431365
transform 1 0 43904 0 -1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_412
timestamp 1698431365
transform 1 0 47488 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_422
timestamp 1698431365
transform 1 0 48608 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_486
timestamp 1698431365
transform 1 0 55776 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_45_492
timestamp 1698431365
transform 1 0 56448 0 -1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_524
timestamp 1698431365
transform 1 0 60032 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_45_534
timestamp 1698431365
transform 1 0 61152 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_558
timestamp 1698431365
transform 1 0 63840 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_562
timestamp 1698431365
transform 1 0 64288 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_566
timestamp 1698431365
transform 1 0 64736 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_568
timestamp 1698431365
transform 1 0 64960 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_632
timestamp 1698431365
transform 1 0 72128 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_646
timestamp 1698431365
transform 1 0 73696 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_648
timestamp 1698431365
transform 1 0 73920 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_663
timestamp 1698431365
transform 1 0 75600 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_667
timestamp 1698431365
transform 1 0 76048 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_684
timestamp 1698431365
transform 1 0 77952 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_28
timestamp 1698431365
transform 1 0 4480 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_32
timestamp 1698431365
transform 1 0 4928 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_34
timestamp 1698431365
transform 1 0 5152 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_46_37
timestamp 1698431365
transform 1 0 5488 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_101
timestamp 1698431365
transform 1 0 12656 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_46_107
timestamp 1698431365
transform 1 0 13328 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_171
timestamp 1698431365
transform 1 0 20496 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_46_177
timestamp 1698431365
transform 1 0 21168 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_241
timestamp 1698431365
transform 1 0 28336 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_46_247
timestamp 1698431365
transform 1 0 29008 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_311
timestamp 1698431365
transform 1 0 36176 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_46_317
timestamp 1698431365
transform 1 0 36848 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_381
timestamp 1698431365
transform 1 0 44016 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_46_387
timestamp 1698431365
transform 1 0 44688 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_451
timestamp 1698431365
transform 1 0 51856 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_46_457
timestamp 1698431365
transform 1 0 52528 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_521
timestamp 1698431365
transform 1 0 59696 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_540
timestamp 1698431365
transform 1 0 61824 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_542
timestamp 1698431365
transform 1 0 62048 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_545
timestamp 1698431365
transform 1 0 62384 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_549
timestamp 1698431365
transform 1 0 62832 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_564
timestamp 1698431365
transform 1 0 64512 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_585
timestamp 1698431365
transform 1 0 66864 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_589
timestamp 1698431365
transform 1 0 67312 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_593
timestamp 1698431365
transform 1 0 67760 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_597
timestamp 1698431365
transform 1 0 68208 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_612
timestamp 1698431365
transform 1 0 69888 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_614
timestamp 1698431365
transform 1 0 70112 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_623
timestamp 1698431365
transform 1 0 71120 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_627
timestamp 1698431365
transform 1 0 71568 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_631
timestamp 1698431365
transform 1 0 72016 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_635
timestamp 1698431365
transform 1 0 72464 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_644
timestamp 1698431365
transform 1 0 73472 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_652
timestamp 1698431365
transform 1 0 74368 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_656
timestamp 1698431365
transform 1 0 74816 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_26
timestamp 1698431365
transform 1 0 4256 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_30
timestamp 1698431365
transform 1 0 4704 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_34
timestamp 1698431365
transform 1 0 5152 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_47_38
timestamp 1698431365
transform 1 0 5600 0 -1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_72
timestamp 1698431365
transform 1 0 9408 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_136
timestamp 1698431365
transform 1 0 16576 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_142
timestamp 1698431365
transform 1 0 17248 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_206
timestamp 1698431365
transform 1 0 24416 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_212
timestamp 1698431365
transform 1 0 25088 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_276
timestamp 1698431365
transform 1 0 32256 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_282
timestamp 1698431365
transform 1 0 32928 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_346
timestamp 1698431365
transform 1 0 40096 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_352
timestamp 1698431365
transform 1 0 40768 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_416
timestamp 1698431365
transform 1 0 47936 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_422
timestamp 1698431365
transform 1 0 48608 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_486
timestamp 1698431365
transform 1 0 55776 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_47_492
timestamp 1698431365
transform 1 0 56448 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_508
timestamp 1698431365
transform 1 0 58240 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_516
timestamp 1698431365
transform 1 0 59136 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_518
timestamp 1698431365
transform 1 0 59360 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_558
timestamp 1698431365
transform 1 0 63840 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_588
timestamp 1698431365
transform 1 0 67200 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_592
timestamp 1698431365
transform 1 0 67648 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_596
timestamp 1698431365
transform 1 0 68096 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_603
timestamp 1698431365
transform 1 0 68880 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_607
timestamp 1698431365
transform 1 0 69328 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_611
timestamp 1698431365
transform 1 0 69776 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_617
timestamp 1698431365
transform 1 0 70448 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_621
timestamp 1698431365
transform 1 0 70896 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_629
timestamp 1698431365
transform 1 0 71792 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_632
timestamp 1698431365
transform 1 0 72128 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_634
timestamp 1698431365
transform 1 0 72352 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_28
timestamp 1698431365
transform 1 0 4480 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_32
timestamp 1698431365
transform 1 0 4928 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_34
timestamp 1698431365
transform 1 0 5152 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_37
timestamp 1698431365
transform 1 0 5488 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_101
timestamp 1698431365
transform 1 0 12656 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_107
timestamp 1698431365
transform 1 0 13328 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_171
timestamp 1698431365
transform 1 0 20496 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_177
timestamp 1698431365
transform 1 0 21168 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_241
timestamp 1698431365
transform 1 0 28336 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_247
timestamp 1698431365
transform 1 0 29008 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_311
timestamp 1698431365
transform 1 0 36176 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_317
timestamp 1698431365
transform 1 0 36848 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_381
timestamp 1698431365
transform 1 0 44016 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_387
timestamp 1698431365
transform 1 0 44688 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_451
timestamp 1698431365
transform 1 0 51856 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_48_457
timestamp 1698431365
transform 1 0 52528 0 1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_473
timestamp 1698431365
transform 1 0 54320 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_477
timestamp 1698431365
transform 1 0 54768 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_488
timestamp 1698431365
transform 1 0 56000 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_492
timestamp 1698431365
transform 1 0 56448 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_496
timestamp 1698431365
transform 1 0 56896 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_48_500
timestamp 1698431365
transform 1 0 57344 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_48_514
timestamp 1698431365
transform 1 0 58912 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_522
timestamp 1698431365
transform 1 0 59808 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_524
timestamp 1698431365
transform 1 0 60032 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_535
timestamp 1698431365
transform 1 0 61264 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_560
timestamp 1698431365
transform 1 0 64064 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_569
timestamp 1698431365
transform 1 0 65072 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_48_586
timestamp 1698431365
transform 1 0 66976 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_594
timestamp 1698431365
transform 1 0 67872 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_597
timestamp 1698431365
transform 1 0 68208 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_601
timestamp 1698431365
transform 1 0 68656 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_611
timestamp 1698431365
transform 1 0 69776 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_633
timestamp 1698431365
transform 1 0 72240 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_637
timestamp 1698431365
transform 1 0 72688 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_639
timestamp 1698431365
transform 1 0 72912 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_664
timestamp 1698431365
transform 1 0 75712 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_683
timestamp 1698431365
transform 1 0 77840 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_687
timestamp 1698431365
transform 1 0 78288 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_28
timestamp 1698431365
transform 1 0 4480 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_49_32
timestamp 1698431365
transform 1 0 4928 0 -1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_64
timestamp 1698431365
transform 1 0 8512 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_68
timestamp 1698431365
transform 1 0 8960 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_49_72
timestamp 1698431365
transform 1 0 9408 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_136
timestamp 1698431365
transform 1 0 16576 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_49_142
timestamp 1698431365
transform 1 0 17248 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_206
timestamp 1698431365
transform 1 0 24416 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_49_212
timestamp 1698431365
transform 1 0 25088 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_276
timestamp 1698431365
transform 1 0 32256 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_49_282
timestamp 1698431365
transform 1 0 32928 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_346
timestamp 1698431365
transform 1 0 40096 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_49_352
timestamp 1698431365
transform 1 0 40768 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_416
timestamp 1698431365
transform 1 0 47936 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_49_422
timestamp 1698431365
transform 1 0 48608 0 -1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_49_454
timestamp 1698431365
transform 1 0 52192 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_470
timestamp 1698431365
transform 1 0 53984 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_486
timestamp 1698431365
transform 1 0 55776 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_49_508
timestamp 1698431365
transform 1 0 58240 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_524
timestamp 1698431365
transform 1 0 60032 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_532
timestamp 1698431365
transform 1 0 60928 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_536
timestamp 1698431365
transform 1 0 61376 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_545
timestamp 1698431365
transform 1 0 62384 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_554
timestamp 1698431365
transform 1 0 63392 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_558
timestamp 1698431365
transform 1 0 63840 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_562
timestamp 1698431365
transform 1 0 64288 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_49_566
timestamp 1698431365
transform 1 0 64736 0 -1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_49_598
timestamp 1698431365
transform 1 0 68320 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_614
timestamp 1698431365
transform 1 0 70112 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_616
timestamp 1698431365
transform 1 0 70336 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_619
timestamp 1698431365
transform 1 0 70672 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_623
timestamp 1698431365
transform 1 0 71120 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_627
timestamp 1698431365
transform 1 0 71568 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_629
timestamp 1698431365
transform 1 0 71792 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_49_632
timestamp 1698431365
transform 1 0 72128 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_650
timestamp 1698431365
transform 1 0 74144 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_28
timestamp 1698431365
transform 1 0 4480 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_32
timestamp 1698431365
transform 1 0 4928 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_34
timestamp 1698431365
transform 1 0 5152 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_50_37
timestamp 1698431365
transform 1 0 5488 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_101
timestamp 1698431365
transform 1 0 12656 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_50_107
timestamp 1698431365
transform 1 0 13328 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_171
timestamp 1698431365
transform 1 0 20496 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_50_177
timestamp 1698431365
transform 1 0 21168 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_241
timestamp 1698431365
transform 1 0 28336 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_50_247
timestamp 1698431365
transform 1 0 29008 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_311
timestamp 1698431365
transform 1 0 36176 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_50_317
timestamp 1698431365
transform 1 0 36848 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_381
timestamp 1698431365
transform 1 0 44016 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_50_387
timestamp 1698431365
transform 1 0 44688 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_451
timestamp 1698431365
transform 1 0 51856 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_50_457
timestamp 1698431365
transform 1 0 52528 0 1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_473
timestamp 1698431365
transform 1 0 54320 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_477
timestamp 1698431365
transform 1 0 54768 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_479
timestamp 1698431365
transform 1 0 54992 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_512
timestamp 1698431365
transform 1 0 58688 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_520
timestamp 1698431365
transform 1 0 59584 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_524
timestamp 1698431365
transform 1 0 60032 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_50_527
timestamp 1698431365
transform 1 0 60368 0 1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_543
timestamp 1698431365
transform 1 0 62160 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_50_546
timestamp 1698431365
transform 1 0 62496 0 1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_50_578
timestamp 1698431365
transform 1 0 66080 0 1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_594
timestamp 1698431365
transform 1 0 67872 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_50_597
timestamp 1698431365
transform 1 0 68208 0 1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_50_629
timestamp 1698431365
transform 1 0 71792 0 1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_645
timestamp 1698431365
transform 1 0 73584 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_653
timestamp 1698431365
transform 1 0 74480 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_657
timestamp 1698431365
transform 1 0 74928 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_659
timestamp 1698431365
transform 1 0 75152 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_662
timestamp 1698431365
transform 1 0 75488 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_664
timestamp 1698431365
transform 1 0 75712 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_667
timestamp 1698431365
transform 1 0 76048 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_687
timestamp 1698431365
transform 1 0 78288 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_2
timestamp 1698431365
transform 1 0 1568 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_4
timestamp 1698431365
transform 1 0 1792 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_51_17
timestamp 1698431365
transform 1 0 3248 0 -1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_51_49
timestamp 1698431365
transform 1 0 6832 0 -1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_65
timestamp 1698431365
transform 1 0 8624 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_69
timestamp 1698431365
transform 1 0 9072 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_51_72
timestamp 1698431365
transform 1 0 9408 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_136
timestamp 1698431365
transform 1 0 16576 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_51_142
timestamp 1698431365
transform 1 0 17248 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_206
timestamp 1698431365
transform 1 0 24416 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_51_212
timestamp 1698431365
transform 1 0 25088 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_276
timestamp 1698431365
transform 1 0 32256 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_51_282
timestamp 1698431365
transform 1 0 32928 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_346
timestamp 1698431365
transform 1 0 40096 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_51_352
timestamp 1698431365
transform 1 0 40768 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_416
timestamp 1698431365
transform 1 0 47936 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_51_422
timestamp 1698431365
transform 1 0 48608 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_486
timestamp 1698431365
transform 1 0 55776 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_51_492
timestamp 1698431365
transform 1 0 56448 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_556
timestamp 1698431365
transform 1 0 63616 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_51_562
timestamp 1698431365
transform 1 0 64288 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_626
timestamp 1698431365
transform 1 0 71456 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_51_632
timestamp 1698431365
transform 1 0 72128 0 -1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_51_664
timestamp 1698431365
transform 1 0 75712 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_672
timestamp 1698431365
transform 1 0 76608 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_678
timestamp 1698431365
transform 1 0 77280 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_28
timestamp 1698431365
transform 1 0 4480 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_32
timestamp 1698431365
transform 1 0 4928 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_34
timestamp 1698431365
transform 1 0 5152 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_52_37
timestamp 1698431365
transform 1 0 5488 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_101
timestamp 1698431365
transform 1 0 12656 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_52_107
timestamp 1698431365
transform 1 0 13328 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_171
timestamp 1698431365
transform 1 0 20496 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_52_177
timestamp 1698431365
transform 1 0 21168 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_241
timestamp 1698431365
transform 1 0 28336 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_52_247
timestamp 1698431365
transform 1 0 29008 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_311
timestamp 1698431365
transform 1 0 36176 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_52_317
timestamp 1698431365
transform 1 0 36848 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_381
timestamp 1698431365
transform 1 0 44016 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_52_387
timestamp 1698431365
transform 1 0 44688 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_451
timestamp 1698431365
transform 1 0 51856 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_52_457
timestamp 1698431365
transform 1 0 52528 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_521
timestamp 1698431365
transform 1 0 59696 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_52_527
timestamp 1698431365
transform 1 0 60368 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_591
timestamp 1698431365
transform 1 0 67536 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_52_597
timestamp 1698431365
transform 1 0 68208 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_661
timestamp 1698431365
transform 1 0 75376 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_52_667
timestamp 1698431365
transform 1 0 76048 0 1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_683
timestamp 1698431365
transform 1 0 77840 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_686
timestamp 1698431365
transform 1 0 78176 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_53_28
timestamp 1698431365
transform 1 0 4480 0 -1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_53_60
timestamp 1698431365
transform 1 0 8064 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_68
timestamp 1698431365
transform 1 0 8960 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_53_72
timestamp 1698431365
transform 1 0 9408 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_136
timestamp 1698431365
transform 1 0 16576 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_53_142
timestamp 1698431365
transform 1 0 17248 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_206
timestamp 1698431365
transform 1 0 24416 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_53_212
timestamp 1698431365
transform 1 0 25088 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_276
timestamp 1698431365
transform 1 0 32256 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_53_282
timestamp 1698431365
transform 1 0 32928 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_346
timestamp 1698431365
transform 1 0 40096 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_53_352
timestamp 1698431365
transform 1 0 40768 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_416
timestamp 1698431365
transform 1 0 47936 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_53_422
timestamp 1698431365
transform 1 0 48608 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_486
timestamp 1698431365
transform 1 0 55776 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_53_492
timestamp 1698431365
transform 1 0 56448 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_556
timestamp 1698431365
transform 1 0 63616 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_53_562
timestamp 1698431365
transform 1 0 64288 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_626
timestamp 1698431365
transform 1 0 71456 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_53_632
timestamp 1698431365
transform 1 0 72128 0 -1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_53_664
timestamp 1698431365
transform 1 0 75712 0 -1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_2
timestamp 1698431365
transform 1 0 1568 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_4
timestamp 1698431365
transform 1 0 1792 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_23
timestamp 1698431365
transform 1 0 3920 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_27
timestamp 1698431365
transform 1 0 4368 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_54_37
timestamp 1698431365
transform 1 0 5488 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_101
timestamp 1698431365
transform 1 0 12656 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_54_107
timestamp 1698431365
transform 1 0 13328 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_171
timestamp 1698431365
transform 1 0 20496 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_54_177
timestamp 1698431365
transform 1 0 21168 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_241
timestamp 1698431365
transform 1 0 28336 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_54_247
timestamp 1698431365
transform 1 0 29008 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_311
timestamp 1698431365
transform 1 0 36176 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_54_317
timestamp 1698431365
transform 1 0 36848 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_381
timestamp 1698431365
transform 1 0 44016 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_54_387
timestamp 1698431365
transform 1 0 44688 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_451
timestamp 1698431365
transform 1 0 51856 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_54_457
timestamp 1698431365
transform 1 0 52528 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_521
timestamp 1698431365
transform 1 0 59696 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_54_527
timestamp 1698431365
transform 1 0 60368 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_591
timestamp 1698431365
transform 1 0 67536 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_54_597
timestamp 1698431365
transform 1 0 68208 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_661
timestamp 1698431365
transform 1 0 75376 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_667
timestamp 1698431365
transform 1 0 76048 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_675
timestamp 1698431365
transform 1 0 76944 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_679
timestamp 1698431365
transform 1 0 77392 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_55_28
timestamp 1698431365
transform 1 0 4480 0 -1 47040
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_55_60
timestamp 1698431365
transform 1 0 8064 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_68
timestamp 1698431365
transform 1 0 8960 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_55_72
timestamp 1698431365
transform 1 0 9408 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_136
timestamp 1698431365
transform 1 0 16576 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_55_142
timestamp 1698431365
transform 1 0 17248 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_206
timestamp 1698431365
transform 1 0 24416 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_55_212
timestamp 1698431365
transform 1 0 25088 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_276
timestamp 1698431365
transform 1 0 32256 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_55_282
timestamp 1698431365
transform 1 0 32928 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_346
timestamp 1698431365
transform 1 0 40096 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_55_352
timestamp 1698431365
transform 1 0 40768 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_416
timestamp 1698431365
transform 1 0 47936 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_55_422
timestamp 1698431365
transform 1 0 48608 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_486
timestamp 1698431365
transform 1 0 55776 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_55_492
timestamp 1698431365
transform 1 0 56448 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_556
timestamp 1698431365
transform 1 0 63616 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_55_562
timestamp 1698431365
transform 1 0 64288 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_626
timestamp 1698431365
transform 1 0 71456 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_55_632
timestamp 1698431365
transform 1 0 72128 0 -1 47040
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_55_664
timestamp 1698431365
transform 1 0 75712 0 -1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_55_680
timestamp 1698431365
transform 1 0 77504 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_28
timestamp 1698431365
transform 1 0 4480 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_32
timestamp 1698431365
transform 1 0 4928 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_34
timestamp 1698431365
transform 1 0 5152 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_56_37
timestamp 1698431365
transform 1 0 5488 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_101
timestamp 1698431365
transform 1 0 12656 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_56_107
timestamp 1698431365
transform 1 0 13328 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_171
timestamp 1698431365
transform 1 0 20496 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_56_177
timestamp 1698431365
transform 1 0 21168 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_241
timestamp 1698431365
transform 1 0 28336 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_56_247
timestamp 1698431365
transform 1 0 29008 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_311
timestamp 1698431365
transform 1 0 36176 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_56_317
timestamp 1698431365
transform 1 0 36848 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_381
timestamp 1698431365
transform 1 0 44016 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_56_387
timestamp 1698431365
transform 1 0 44688 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_451
timestamp 1698431365
transform 1 0 51856 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_56_457
timestamp 1698431365
transform 1 0 52528 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_521
timestamp 1698431365
transform 1 0 59696 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_56_527
timestamp 1698431365
transform 1 0 60368 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_591
timestamp 1698431365
transform 1 0 67536 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_56_597
timestamp 1698431365
transform 1 0 68208 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_661
timestamp 1698431365
transform 1 0 75376 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_56_667
timestamp 1698431365
transform 1 0 76048 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_675
timestamp 1698431365
transform 1 0 76944 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_679
timestamp 1698431365
transform 1 0 77392 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_2
timestamp 1698431365
transform 1 0 1568 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_4
timestamp 1698431365
transform 1 0 1792 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_57_23
timestamp 1698431365
transform 1 0 3920 0 -1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_57_55
timestamp 1698431365
transform 1 0 7504 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_63
timestamp 1698431365
transform 1 0 8400 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_67
timestamp 1698431365
transform 1 0 8848 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_69
timestamp 1698431365
transform 1 0 9072 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_57_72
timestamp 1698431365
transform 1 0 9408 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_136
timestamp 1698431365
transform 1 0 16576 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_57_142
timestamp 1698431365
transform 1 0 17248 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_206
timestamp 1698431365
transform 1 0 24416 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_57_212
timestamp 1698431365
transform 1 0 25088 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_276
timestamp 1698431365
transform 1 0 32256 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_57_282
timestamp 1698431365
transform 1 0 32928 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_346
timestamp 1698431365
transform 1 0 40096 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_57_352
timestamp 1698431365
transform 1 0 40768 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_416
timestamp 1698431365
transform 1 0 47936 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_57_422
timestamp 1698431365
transform 1 0 48608 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_486
timestamp 1698431365
transform 1 0 55776 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_57_492
timestamp 1698431365
transform 1 0 56448 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_556
timestamp 1698431365
transform 1 0 63616 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_57_562
timestamp 1698431365
transform 1 0 64288 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_626
timestamp 1698431365
transform 1 0 71456 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_57_632
timestamp 1698431365
transform 1 0 72128 0 -1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_57_664
timestamp 1698431365
transform 1 0 75712 0 -1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_28
timestamp 1698431365
transform 1 0 4480 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_32
timestamp 1698431365
transform 1 0 4928 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_34
timestamp 1698431365
transform 1 0 5152 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_58_37
timestamp 1698431365
transform 1 0 5488 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_101
timestamp 1698431365
transform 1 0 12656 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_58_107
timestamp 1698431365
transform 1 0 13328 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_171
timestamp 1698431365
transform 1 0 20496 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_58_177
timestamp 1698431365
transform 1 0 21168 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_241
timestamp 1698431365
transform 1 0 28336 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_58_247
timestamp 1698431365
transform 1 0 29008 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_311
timestamp 1698431365
transform 1 0 36176 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_58_317
timestamp 1698431365
transform 1 0 36848 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_381
timestamp 1698431365
transform 1 0 44016 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_58_387
timestamp 1698431365
transform 1 0 44688 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_451
timestamp 1698431365
transform 1 0 51856 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_58_457
timestamp 1698431365
transform 1 0 52528 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_521
timestamp 1698431365
transform 1 0 59696 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_58_527
timestamp 1698431365
transform 1 0 60368 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_591
timestamp 1698431365
transform 1 0 67536 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_58_597
timestamp 1698431365
transform 1 0 68208 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_661
timestamp 1698431365
transform 1 0 75376 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_58_667
timestamp 1698431365
transform 1 0 76048 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_675
timestamp 1698431365
transform 1 0 76944 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_679
timestamp 1698431365
transform 1 0 77392 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_59_28
timestamp 1698431365
transform 1 0 4480 0 -1 50176
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_59_60
timestamp 1698431365
transform 1 0 8064 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_68
timestamp 1698431365
transform 1 0 8960 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_59_72
timestamp 1698431365
transform 1 0 9408 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_136
timestamp 1698431365
transform 1 0 16576 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_59_142
timestamp 1698431365
transform 1 0 17248 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_206
timestamp 1698431365
transform 1 0 24416 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_59_212
timestamp 1698431365
transform 1 0 25088 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_276
timestamp 1698431365
transform 1 0 32256 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_59_282
timestamp 1698431365
transform 1 0 32928 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_346
timestamp 1698431365
transform 1 0 40096 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_59_352
timestamp 1698431365
transform 1 0 40768 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_416
timestamp 1698431365
transform 1 0 47936 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_59_422
timestamp 1698431365
transform 1 0 48608 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_486
timestamp 1698431365
transform 1 0 55776 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_59_492
timestamp 1698431365
transform 1 0 56448 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_556
timestamp 1698431365
transform 1 0 63616 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_59_562
timestamp 1698431365
transform 1 0 64288 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_626
timestamp 1698431365
transform 1 0 71456 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_59_632
timestamp 1698431365
transform 1 0 72128 0 -1 50176
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_59_664
timestamp 1698431365
transform 1 0 75712 0 -1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_59_680
timestamp 1698431365
transform 1 0 77504 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_28
timestamp 1698431365
transform 1 0 4480 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_32
timestamp 1698431365
transform 1 0 4928 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_34
timestamp 1698431365
transform 1 0 5152 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_60_37
timestamp 1698431365
transform 1 0 5488 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_101
timestamp 1698431365
transform 1 0 12656 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_60_107
timestamp 1698431365
transform 1 0 13328 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_171
timestamp 1698431365
transform 1 0 20496 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_60_177
timestamp 1698431365
transform 1 0 21168 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_241
timestamp 1698431365
transform 1 0 28336 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_60_247
timestamp 1698431365
transform 1 0 29008 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_311
timestamp 1698431365
transform 1 0 36176 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_60_317
timestamp 1698431365
transform 1 0 36848 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_381
timestamp 1698431365
transform 1 0 44016 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_60_387
timestamp 1698431365
transform 1 0 44688 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_451
timestamp 1698431365
transform 1 0 51856 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_60_457
timestamp 1698431365
transform 1 0 52528 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_521
timestamp 1698431365
transform 1 0 59696 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_60_527
timestamp 1698431365
transform 1 0 60368 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_591
timestamp 1698431365
transform 1 0 67536 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_60_597
timestamp 1698431365
transform 1 0 68208 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_661
timestamp 1698431365
transform 1 0 75376 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_60_667
timestamp 1698431365
transform 1 0 76048 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_675
timestamp 1698431365
transform 1 0 76944 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_679
timestamp 1698431365
transform 1 0 77392 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_2
timestamp 1698431365
transform 1 0 1568 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_61_24
timestamp 1698431365
transform 1 0 4032 0 -1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_61_56
timestamp 1698431365
transform 1 0 7616 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_64
timestamp 1698431365
transform 1 0 8512 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_68
timestamp 1698431365
transform 1 0 8960 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_61_72
timestamp 1698431365
transform 1 0 9408 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_136
timestamp 1698431365
transform 1 0 16576 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_61_142
timestamp 1698431365
transform 1 0 17248 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_206
timestamp 1698431365
transform 1 0 24416 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_61_212
timestamp 1698431365
transform 1 0 25088 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_276
timestamp 1698431365
transform 1 0 32256 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_61_282
timestamp 1698431365
transform 1 0 32928 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_346
timestamp 1698431365
transform 1 0 40096 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_61_352
timestamp 1698431365
transform 1 0 40768 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_416
timestamp 1698431365
transform 1 0 47936 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_61_422
timestamp 1698431365
transform 1 0 48608 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_486
timestamp 1698431365
transform 1 0 55776 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_61_492
timestamp 1698431365
transform 1 0 56448 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_556
timestamp 1698431365
transform 1 0 63616 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_61_562
timestamp 1698431365
transform 1 0 64288 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_626
timestamp 1698431365
transform 1 0 71456 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_61_632
timestamp 1698431365
transform 1 0 72128 0 -1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_61_664
timestamp 1698431365
transform 1 0 75712 0 -1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_28
timestamp 1698431365
transform 1 0 4480 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_32
timestamp 1698431365
transform 1 0 4928 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_34
timestamp 1698431365
transform 1 0 5152 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_62_37
timestamp 1698431365
transform 1 0 5488 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_101
timestamp 1698431365
transform 1 0 12656 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_62_107
timestamp 1698431365
transform 1 0 13328 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_171
timestamp 1698431365
transform 1 0 20496 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_62_177
timestamp 1698431365
transform 1 0 21168 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_241
timestamp 1698431365
transform 1 0 28336 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_62_247
timestamp 1698431365
transform 1 0 29008 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_311
timestamp 1698431365
transform 1 0 36176 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_62_317
timestamp 1698431365
transform 1 0 36848 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_381
timestamp 1698431365
transform 1 0 44016 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_62_387
timestamp 1698431365
transform 1 0 44688 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_451
timestamp 1698431365
transform 1 0 51856 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_62_457
timestamp 1698431365
transform 1 0 52528 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_521
timestamp 1698431365
transform 1 0 59696 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_62_527
timestamp 1698431365
transform 1 0 60368 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_591
timestamp 1698431365
transform 1 0 67536 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_62_597
timestamp 1698431365
transform 1 0 68208 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_661
timestamp 1698431365
transform 1 0 75376 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_62_667
timestamp 1698431365
transform 1 0 76048 0 1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_683
timestamp 1698431365
transform 1 0 77840 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_687
timestamp 1698431365
transform 1 0 78288 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_63_28
timestamp 1698431365
transform 1 0 4480 0 -1 53312
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_63_60
timestamp 1698431365
transform 1 0 8064 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_68
timestamp 1698431365
transform 1 0 8960 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_63_72
timestamp 1698431365
transform 1 0 9408 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_136
timestamp 1698431365
transform 1 0 16576 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_63_142
timestamp 1698431365
transform 1 0 17248 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_206
timestamp 1698431365
transform 1 0 24416 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_63_212
timestamp 1698431365
transform 1 0 25088 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_276
timestamp 1698431365
transform 1 0 32256 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_63_282
timestamp 1698431365
transform 1 0 32928 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_346
timestamp 1698431365
transform 1 0 40096 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_63_352
timestamp 1698431365
transform 1 0 40768 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_416
timestamp 1698431365
transform 1 0 47936 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_63_422
timestamp 1698431365
transform 1 0 48608 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_486
timestamp 1698431365
transform 1 0 55776 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_63_492
timestamp 1698431365
transform 1 0 56448 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_556
timestamp 1698431365
transform 1 0 63616 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_63_562
timestamp 1698431365
transform 1 0 64288 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_626
timestamp 1698431365
transform 1 0 71456 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_63_632
timestamp 1698431365
transform 1 0 72128 0 -1 53312
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_63_664
timestamp 1698431365
transform 1 0 75712 0 -1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_2
timestamp 1698431365
transform 1 0 1568 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_64_24
timestamp 1698431365
transform 1 0 4032 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_32
timestamp 1698431365
transform 1 0 4928 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_34
timestamp 1698431365
transform 1 0 5152 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_64_37
timestamp 1698431365
transform 1 0 5488 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_101
timestamp 1698431365
transform 1 0 12656 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_64_107
timestamp 1698431365
transform 1 0 13328 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_171
timestamp 1698431365
transform 1 0 20496 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_64_177
timestamp 1698431365
transform 1 0 21168 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_241
timestamp 1698431365
transform 1 0 28336 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_64_247
timestamp 1698431365
transform 1 0 29008 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_311
timestamp 1698431365
transform 1 0 36176 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_64_317
timestamp 1698431365
transform 1 0 36848 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_381
timestamp 1698431365
transform 1 0 44016 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_64_387
timestamp 1698431365
transform 1 0 44688 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_451
timestamp 1698431365
transform 1 0 51856 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_64_457
timestamp 1698431365
transform 1 0 52528 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_521
timestamp 1698431365
transform 1 0 59696 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_64_527
timestamp 1698431365
transform 1 0 60368 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_591
timestamp 1698431365
transform 1 0 67536 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_64_597
timestamp 1698431365
transform 1 0 68208 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_661
timestamp 1698431365
transform 1 0 75376 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_64_667
timestamp 1698431365
transform 1 0 76048 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_675
timestamp 1698431365
transform 1 0 76944 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_679
timestamp 1698431365
transform 1 0 77392 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_65_28
timestamp 1698431365
transform 1 0 4480 0 -1 54880
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_65_60
timestamp 1698431365
transform 1 0 8064 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_68
timestamp 1698431365
transform 1 0 8960 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_65_72
timestamp 1698431365
transform 1 0 9408 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_136
timestamp 1698431365
transform 1 0 16576 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_65_142
timestamp 1698431365
transform 1 0 17248 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_206
timestamp 1698431365
transform 1 0 24416 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_65_212
timestamp 1698431365
transform 1 0 25088 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_276
timestamp 1698431365
transform 1 0 32256 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_65_282
timestamp 1698431365
transform 1 0 32928 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_346
timestamp 1698431365
transform 1 0 40096 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_65_352
timestamp 1698431365
transform 1 0 40768 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_416
timestamp 1698431365
transform 1 0 47936 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_65_422
timestamp 1698431365
transform 1 0 48608 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_486
timestamp 1698431365
transform 1 0 55776 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_65_492
timestamp 1698431365
transform 1 0 56448 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_556
timestamp 1698431365
transform 1 0 63616 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_65_562
timestamp 1698431365
transform 1 0 64288 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_626
timestamp 1698431365
transform 1 0 71456 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_65_632
timestamp 1698431365
transform 1 0 72128 0 -1 54880
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_65_664
timestamp 1698431365
transform 1 0 75712 0 -1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_65_680
timestamp 1698431365
transform 1 0 77504 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_28
timestamp 1698431365
transform 1 0 4480 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_32
timestamp 1698431365
transform 1 0 4928 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_34
timestamp 1698431365
transform 1 0 5152 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_66_37
timestamp 1698431365
transform 1 0 5488 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_101
timestamp 1698431365
transform 1 0 12656 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_66_107
timestamp 1698431365
transform 1 0 13328 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_171
timestamp 1698431365
transform 1 0 20496 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_66_177
timestamp 1698431365
transform 1 0 21168 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_241
timestamp 1698431365
transform 1 0 28336 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_66_247
timestamp 1698431365
transform 1 0 29008 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_311
timestamp 1698431365
transform 1 0 36176 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_66_317
timestamp 1698431365
transform 1 0 36848 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_381
timestamp 1698431365
transform 1 0 44016 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_66_387
timestamp 1698431365
transform 1 0 44688 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_451
timestamp 1698431365
transform 1 0 51856 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_66_457
timestamp 1698431365
transform 1 0 52528 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_521
timestamp 1698431365
transform 1 0 59696 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_66_527
timestamp 1698431365
transform 1 0 60368 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_591
timestamp 1698431365
transform 1 0 67536 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_66_597
timestamp 1698431365
transform 1 0 68208 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_661
timestamp 1698431365
transform 1 0 75376 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_66_667
timestamp 1698431365
transform 1 0 76048 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_675
timestamp 1698431365
transform 1 0 76944 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_679
timestamp 1698431365
transform 1 0 77392 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_2
timestamp 1698431365
transform 1 0 1568 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_4
timestamp 1698431365
transform 1 0 1792 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_67_23
timestamp 1698431365
transform 1 0 3920 0 -1 56448
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_55
timestamp 1698431365
transform 1 0 7504 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_63
timestamp 1698431365
transform 1 0 8400 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_67
timestamp 1698431365
transform 1 0 8848 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_69
timestamp 1698431365
transform 1 0 9072 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_67_72
timestamp 1698431365
transform 1 0 9408 0 -1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_136
timestamp 1698431365
transform 1 0 16576 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_67_142
timestamp 1698431365
transform 1 0 17248 0 -1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_206
timestamp 1698431365
transform 1 0 24416 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_67_212
timestamp 1698431365
transform 1 0 25088 0 -1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_276
timestamp 1698431365
transform 1 0 32256 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_67_282
timestamp 1698431365
transform 1 0 32928 0 -1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_346
timestamp 1698431365
transform 1 0 40096 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_67_352
timestamp 1698431365
transform 1 0 40768 0 -1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_416
timestamp 1698431365
transform 1 0 47936 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_67_422
timestamp 1698431365
transform 1 0 48608 0 -1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_486
timestamp 1698431365
transform 1 0 55776 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_67_492
timestamp 1698431365
transform 1 0 56448 0 -1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_556
timestamp 1698431365
transform 1 0 63616 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_67_562
timestamp 1698431365
transform 1 0 64288 0 -1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_626
timestamp 1698431365
transform 1 0 71456 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_67_632
timestamp 1698431365
transform 1 0 72128 0 -1 56448
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_67_664
timestamp 1698431365
transform 1 0 75712 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_68_34
timestamp 1698431365
transform 1 0 5152 0 1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_68_37
timestamp 1698431365
transform 1 0 5488 0 1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_68_101
timestamp 1698431365
transform 1 0 12656 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_68_107
timestamp 1698431365
transform 1 0 13328 0 1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_68_171
timestamp 1698431365
transform 1 0 20496 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_68_177
timestamp 1698431365
transform 1 0 21168 0 1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_68_241
timestamp 1698431365
transform 1 0 28336 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_68_247
timestamp 1698431365
transform 1 0 29008 0 1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_68_311
timestamp 1698431365
transform 1 0 36176 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_68_317
timestamp 1698431365
transform 1 0 36848 0 1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_68_381
timestamp 1698431365
transform 1 0 44016 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_68_387
timestamp 1698431365
transform 1 0 44688 0 1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_68_451
timestamp 1698431365
transform 1 0 51856 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_68_457
timestamp 1698431365
transform 1 0 52528 0 1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_68_521
timestamp 1698431365
transform 1 0 59696 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_68_527
timestamp 1698431365
transform 1 0 60368 0 1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_68_591
timestamp 1698431365
transform 1 0 67536 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_68_597
timestamp 1698431365
transform 1 0 68208 0 1 56448
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_68_661
timestamp 1698431365
transform 1 0 75376 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_68_667
timestamp 1698431365
transform 1 0 76048 0 1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_68_675
timestamp 1698431365
transform 1 0 76944 0 1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_68_679
timestamp 1698431365
transform 1 0 77392 0 1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_69_28
timestamp 1698431365
transform 1 0 4480 0 -1 58016
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_69_60
timestamp 1698431365
transform 1 0 8064 0 -1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_69_68
timestamp 1698431365
transform 1 0 8960 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_69_72
timestamp 1698431365
transform 1 0 9408 0 -1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_69_136
timestamp 1698431365
transform 1 0 16576 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_69_142
timestamp 1698431365
transform 1 0 17248 0 -1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_69_206
timestamp 1698431365
transform 1 0 24416 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_69_212
timestamp 1698431365
transform 1 0 25088 0 -1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_69_276
timestamp 1698431365
transform 1 0 32256 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_69_282
timestamp 1698431365
transform 1 0 32928 0 -1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_69_346
timestamp 1698431365
transform 1 0 40096 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_69_352
timestamp 1698431365
transform 1 0 40768 0 -1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_69_416
timestamp 1698431365
transform 1 0 47936 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_69_422
timestamp 1698431365
transform 1 0 48608 0 -1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_69_486
timestamp 1698431365
transform 1 0 55776 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_69_492
timestamp 1698431365
transform 1 0 56448 0 -1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_69_556
timestamp 1698431365
transform 1 0 63616 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_69_562
timestamp 1698431365
transform 1 0 64288 0 -1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_69_626
timestamp 1698431365
transform 1 0 71456 0 -1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_69_632
timestamp 1698431365
transform 1 0 72128 0 -1 58016
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_69_664
timestamp 1698431365
transform 1 0 75712 0 -1 58016
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_69_680
timestamp 1698431365
transform 1 0 77504 0 -1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_70_28
timestamp 1698431365
transform 1 0 4480 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_70_32
timestamp 1698431365
transform 1 0 4928 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_70_34
timestamp 1698431365
transform 1 0 5152 0 1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_70_37
timestamp 1698431365
transform 1 0 5488 0 1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_70_101
timestamp 1698431365
transform 1 0 12656 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_70_107
timestamp 1698431365
transform 1 0 13328 0 1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_70_171
timestamp 1698431365
transform 1 0 20496 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_70_177
timestamp 1698431365
transform 1 0 21168 0 1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_70_241
timestamp 1698431365
transform 1 0 28336 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_70_247
timestamp 1698431365
transform 1 0 29008 0 1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_70_311
timestamp 1698431365
transform 1 0 36176 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_70_317
timestamp 1698431365
transform 1 0 36848 0 1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_70_381
timestamp 1698431365
transform 1 0 44016 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_70_387
timestamp 1698431365
transform 1 0 44688 0 1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_70_451
timestamp 1698431365
transform 1 0 51856 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_70_457
timestamp 1698431365
transform 1 0 52528 0 1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_70_521
timestamp 1698431365
transform 1 0 59696 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_70_527
timestamp 1698431365
transform 1 0 60368 0 1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_70_591
timestamp 1698431365
transform 1 0 67536 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_70_597
timestamp 1698431365
transform 1 0 68208 0 1 58016
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_70_661
timestamp 1698431365
transform 1 0 75376 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_70_667
timestamp 1698431365
transform 1 0 76048 0 1 58016
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_70_675
timestamp 1698431365
transform 1 0 76944 0 1 58016
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_70_679
timestamp 1698431365
transform 1 0 77392 0 1 58016
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_2
timestamp 1698431365
transform 1 0 1568 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_71_4
timestamp 1698431365
transform 1 0 1792 0 -1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_17
timestamp 1698431365
transform 1 0 3248 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_71_21
timestamp 1698431365
transform 1 0 3696 0 -1 59584
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_71_53
timestamp 1698431365
transform 1 0 7280 0 -1 59584
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_71_69
timestamp 1698431365
transform 1 0 9072 0 -1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_71_72
timestamp 1698431365
transform 1 0 9408 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_71_136
timestamp 1698431365
transform 1 0 16576 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_71_142
timestamp 1698431365
transform 1 0 17248 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_71_206
timestamp 1698431365
transform 1 0 24416 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_71_212
timestamp 1698431365
transform 1 0 25088 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_71_276
timestamp 1698431365
transform 1 0 32256 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_71_282
timestamp 1698431365
transform 1 0 32928 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_71_346
timestamp 1698431365
transform 1 0 40096 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_71_352
timestamp 1698431365
transform 1 0 40768 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_71_416
timestamp 1698431365
transform 1 0 47936 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_71_422
timestamp 1698431365
transform 1 0 48608 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_71_486
timestamp 1698431365
transform 1 0 55776 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_71_492
timestamp 1698431365
transform 1 0 56448 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_71_556
timestamp 1698431365
transform 1 0 63616 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_71_562
timestamp 1698431365
transform 1 0 64288 0 -1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_71_626
timestamp 1698431365
transform 1 0 71456 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_71_632
timestamp 1698431365
transform 1 0 72128 0 -1 59584
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_71_664
timestamp 1698431365
transform 1 0 75712 0 -1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_71_672
timestamp 1698431365
transform 1 0 76608 0 -1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_71_676
timestamp 1698431365
transform 1 0 77056 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_72_28
timestamp 1698431365
transform 1 0 4480 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_72_32
timestamp 1698431365
transform 1 0 4928 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_72_34
timestamp 1698431365
transform 1 0 5152 0 1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_72_37
timestamp 1698431365
transform 1 0 5488 0 1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_72_101
timestamp 1698431365
transform 1 0 12656 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_72_107
timestamp 1698431365
transform 1 0 13328 0 1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_72_171
timestamp 1698431365
transform 1 0 20496 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_72_177
timestamp 1698431365
transform 1 0 21168 0 1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_72_241
timestamp 1698431365
transform 1 0 28336 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_72_247
timestamp 1698431365
transform 1 0 29008 0 1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_72_311
timestamp 1698431365
transform 1 0 36176 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_72_317
timestamp 1698431365
transform 1 0 36848 0 1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_72_381
timestamp 1698431365
transform 1 0 44016 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_72_387
timestamp 1698431365
transform 1 0 44688 0 1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_72_451
timestamp 1698431365
transform 1 0 51856 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_72_457
timestamp 1698431365
transform 1 0 52528 0 1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_72_521
timestamp 1698431365
transform 1 0 59696 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_72_527
timestamp 1698431365
transform 1 0 60368 0 1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_72_591
timestamp 1698431365
transform 1 0 67536 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_72_597
timestamp 1698431365
transform 1 0 68208 0 1 59584
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_72_661
timestamp 1698431365
transform 1 0 75376 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_72_667
timestamp 1698431365
transform 1 0 76048 0 1 59584
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_72_683
timestamp 1698431365
transform 1 0 77840 0 1 59584
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_72_687
timestamp 1698431365
transform 1 0 78288 0 1 59584
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_73_28
timestamp 1698431365
transform 1 0 4480 0 -1 61152
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_73_60
timestamp 1698431365
transform 1 0 8064 0 -1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_73_68
timestamp 1698431365
transform 1 0 8960 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_73_72
timestamp 1698431365
transform 1 0 9408 0 -1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_73_136
timestamp 1698431365
transform 1 0 16576 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_73_142
timestamp 1698431365
transform 1 0 17248 0 -1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_73_206
timestamp 1698431365
transform 1 0 24416 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_73_212
timestamp 1698431365
transform 1 0 25088 0 -1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_73_276
timestamp 1698431365
transform 1 0 32256 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_73_282
timestamp 1698431365
transform 1 0 32928 0 -1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_73_346
timestamp 1698431365
transform 1 0 40096 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_73_352
timestamp 1698431365
transform 1 0 40768 0 -1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_73_416
timestamp 1698431365
transform 1 0 47936 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_73_422
timestamp 1698431365
transform 1 0 48608 0 -1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_73_486
timestamp 1698431365
transform 1 0 55776 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_73_492
timestamp 1698431365
transform 1 0 56448 0 -1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_73_556
timestamp 1698431365
transform 1 0 63616 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_73_562
timestamp 1698431365
transform 1 0 64288 0 -1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_73_626
timestamp 1698431365
transform 1 0 71456 0 -1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_73_632
timestamp 1698431365
transform 1 0 72128 0 -1 61152
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_73_664
timestamp 1698431365
transform 1 0 75712 0 -1 61152
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_74_2
timestamp 1698431365
transform 1 0 1568 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_74_4
timestamp 1698431365
transform 1 0 1792 0 1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_74_23
timestamp 1698431365
transform 1 0 3920 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_74_27
timestamp 1698431365
transform 1 0 4368 0 1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_74_37
timestamp 1698431365
transform 1 0 5488 0 1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_74_101
timestamp 1698431365
transform 1 0 12656 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_74_107
timestamp 1698431365
transform 1 0 13328 0 1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_74_171
timestamp 1698431365
transform 1 0 20496 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_74_177
timestamp 1698431365
transform 1 0 21168 0 1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_74_241
timestamp 1698431365
transform 1 0 28336 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_74_247
timestamp 1698431365
transform 1 0 29008 0 1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_74_311
timestamp 1698431365
transform 1 0 36176 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_74_317
timestamp 1698431365
transform 1 0 36848 0 1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_74_381
timestamp 1698431365
transform 1 0 44016 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_74_387
timestamp 1698431365
transform 1 0 44688 0 1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_74_451
timestamp 1698431365
transform 1 0 51856 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_74_457
timestamp 1698431365
transform 1 0 52528 0 1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_74_521
timestamp 1698431365
transform 1 0 59696 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_74_527
timestamp 1698431365
transform 1 0 60368 0 1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_74_591
timestamp 1698431365
transform 1 0 67536 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_74_597
timestamp 1698431365
transform 1 0 68208 0 1 61152
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_74_661
timestamp 1698431365
transform 1 0 75376 0 1 61152
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_74_667
timestamp 1698431365
transform 1 0 76048 0 1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_74_675
timestamp 1698431365
transform 1 0 76944 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_74_677
timestamp 1698431365
transform 1 0 77168 0 1 61152
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_75_28
timestamp 1698431365
transform 1 0 4480 0 -1 62720
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_75_60
timestamp 1698431365
transform 1 0 8064 0 -1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_75_68
timestamp 1698431365
transform 1 0 8960 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_75_72
timestamp 1698431365
transform 1 0 9408 0 -1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_75_136
timestamp 1698431365
transform 1 0 16576 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_75_142
timestamp 1698431365
transform 1 0 17248 0 -1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_75_206
timestamp 1698431365
transform 1 0 24416 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_75_212
timestamp 1698431365
transform 1 0 25088 0 -1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_75_276
timestamp 1698431365
transform 1 0 32256 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_75_282
timestamp 1698431365
transform 1 0 32928 0 -1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_75_346
timestamp 1698431365
transform 1 0 40096 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_75_352
timestamp 1698431365
transform 1 0 40768 0 -1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_75_416
timestamp 1698431365
transform 1 0 47936 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_75_422
timestamp 1698431365
transform 1 0 48608 0 -1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_75_486
timestamp 1698431365
transform 1 0 55776 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_75_492
timestamp 1698431365
transform 1 0 56448 0 -1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_75_556
timestamp 1698431365
transform 1 0 63616 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_75_562
timestamp 1698431365
transform 1 0 64288 0 -1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_75_626
timestamp 1698431365
transform 1 0 71456 0 -1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_75_632
timestamp 1698431365
transform 1 0 72128 0 -1 62720
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_75_664
timestamp 1698431365
transform 1 0 75712 0 -1 62720
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_75_680
timestamp 1698431365
transform 1 0 77504 0 -1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_76_28
timestamp 1698431365
transform 1 0 4480 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_76_32
timestamp 1698431365
transform 1 0 4928 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_76_34
timestamp 1698431365
transform 1 0 5152 0 1 62720
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_76_37
timestamp 1698431365
transform 1 0 5488 0 1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_76_101
timestamp 1698431365
transform 1 0 12656 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_76_107
timestamp 1698431365
transform 1 0 13328 0 1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_76_171
timestamp 1698431365
transform 1 0 20496 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_76_177
timestamp 1698431365
transform 1 0 21168 0 1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_76_241
timestamp 1698431365
transform 1 0 28336 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_76_247
timestamp 1698431365
transform 1 0 29008 0 1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_76_311
timestamp 1698431365
transform 1 0 36176 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_76_317
timestamp 1698431365
transform 1 0 36848 0 1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_76_381
timestamp 1698431365
transform 1 0 44016 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_76_387
timestamp 1698431365
transform 1 0 44688 0 1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_76_451
timestamp 1698431365
transform 1 0 51856 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_76_457
timestamp 1698431365
transform 1 0 52528 0 1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_76_521
timestamp 1698431365
transform 1 0 59696 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_76_527
timestamp 1698431365
transform 1 0 60368 0 1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_76_591
timestamp 1698431365
transform 1 0 67536 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_76_597
timestamp 1698431365
transform 1 0 68208 0 1 62720
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_76_661
timestamp 1698431365
transform 1 0 75376 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_76_667
timestamp 1698431365
transform 1 0 76048 0 1 62720
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_76_675
timestamp 1698431365
transform 1 0 76944 0 1 62720
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_76_679
timestamp 1698431365
transform 1 0 77392 0 1 62720
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_77_2
timestamp 1698431365
transform 1 0 1568 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_77_24
timestamp 1698431365
transform 1 0 4032 0 -1 64288
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_77_56
timestamp 1698431365
transform 1 0 7616 0 -1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_77_64
timestamp 1698431365
transform 1 0 8512 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_77_68
timestamp 1698431365
transform 1 0 8960 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_77_72
timestamp 1698431365
transform 1 0 9408 0 -1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_77_136
timestamp 1698431365
transform 1 0 16576 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_77_142
timestamp 1698431365
transform 1 0 17248 0 -1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_77_206
timestamp 1698431365
transform 1 0 24416 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_77_212
timestamp 1698431365
transform 1 0 25088 0 -1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_77_276
timestamp 1698431365
transform 1 0 32256 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_77_282
timestamp 1698431365
transform 1 0 32928 0 -1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_77_346
timestamp 1698431365
transform 1 0 40096 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_77_352
timestamp 1698431365
transform 1 0 40768 0 -1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_77_416
timestamp 1698431365
transform 1 0 47936 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_77_422
timestamp 1698431365
transform 1 0 48608 0 -1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_77_486
timestamp 1698431365
transform 1 0 55776 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_77_492
timestamp 1698431365
transform 1 0 56448 0 -1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_77_556
timestamp 1698431365
transform 1 0 63616 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_77_562
timestamp 1698431365
transform 1 0 64288 0 -1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_77_626
timestamp 1698431365
transform 1 0 71456 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_77_632
timestamp 1698431365
transform 1 0 72128 0 -1 64288
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_77_664
timestamp 1698431365
transform 1 0 75712 0 -1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_77_672
timestamp 1698431365
transform 1 0 76608 0 -1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_77_676
timestamp 1698431365
transform 1 0 77056 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_78_34
timestamp 1698431365
transform 1 0 5152 0 1 64288
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_78_37
timestamp 1698431365
transform 1 0 5488 0 1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_78_101
timestamp 1698431365
transform 1 0 12656 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_78_107
timestamp 1698431365
transform 1 0 13328 0 1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_78_171
timestamp 1698431365
transform 1 0 20496 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_78_177
timestamp 1698431365
transform 1 0 21168 0 1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_78_241
timestamp 1698431365
transform 1 0 28336 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_78_247
timestamp 1698431365
transform 1 0 29008 0 1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_78_311
timestamp 1698431365
transform 1 0 36176 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_78_317
timestamp 1698431365
transform 1 0 36848 0 1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_78_381
timestamp 1698431365
transform 1 0 44016 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_78_387
timestamp 1698431365
transform 1 0 44688 0 1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_78_451
timestamp 1698431365
transform 1 0 51856 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_78_457
timestamp 1698431365
transform 1 0 52528 0 1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_78_521
timestamp 1698431365
transform 1 0 59696 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_78_527
timestamp 1698431365
transform 1 0 60368 0 1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_78_591
timestamp 1698431365
transform 1 0 67536 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_78_597
timestamp 1698431365
transform 1 0 68208 0 1 64288
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_78_661
timestamp 1698431365
transform 1 0 75376 0 1 64288
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_78_667
timestamp 1698431365
transform 1 0 76048 0 1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_78_675
timestamp 1698431365
transform 1 0 76944 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_78_677
timestamp 1698431365
transform 1 0 77168 0 1 64288
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_79_28
timestamp 1698431365
transform 1 0 4480 0 -1 65856
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_79_60
timestamp 1698431365
transform 1 0 8064 0 -1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_79_68
timestamp 1698431365
transform 1 0 8960 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_79_72
timestamp 1698431365
transform 1 0 9408 0 -1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_79_136
timestamp 1698431365
transform 1 0 16576 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_79_142
timestamp 1698431365
transform 1 0 17248 0 -1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_79_206
timestamp 1698431365
transform 1 0 24416 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_79_212
timestamp 1698431365
transform 1 0 25088 0 -1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_79_276
timestamp 1698431365
transform 1 0 32256 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_79_282
timestamp 1698431365
transform 1 0 32928 0 -1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_79_346
timestamp 1698431365
transform 1 0 40096 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_79_352
timestamp 1698431365
transform 1 0 40768 0 -1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_79_416
timestamp 1698431365
transform 1 0 47936 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_79_422
timestamp 1698431365
transform 1 0 48608 0 -1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_79_486
timestamp 1698431365
transform 1 0 55776 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_79_492
timestamp 1698431365
transform 1 0 56448 0 -1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_79_556
timestamp 1698431365
transform 1 0 63616 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_79_562
timestamp 1698431365
transform 1 0 64288 0 -1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_79_626
timestamp 1698431365
transform 1 0 71456 0 -1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_79_632
timestamp 1698431365
transform 1 0 72128 0 -1 65856
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_79_664
timestamp 1698431365
transform 1 0 75712 0 -1 65856
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_79_680
timestamp 1698431365
transform 1 0 77504 0 -1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_80_28
timestamp 1698431365
transform 1 0 4480 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_80_32
timestamp 1698431365
transform 1 0 4928 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_80_34
timestamp 1698431365
transform 1 0 5152 0 1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_80_37
timestamp 1698431365
transform 1 0 5488 0 1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_80_101
timestamp 1698431365
transform 1 0 12656 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_80_107
timestamp 1698431365
transform 1 0 13328 0 1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_80_171
timestamp 1698431365
transform 1 0 20496 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_80_177
timestamp 1698431365
transform 1 0 21168 0 1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_80_241
timestamp 1698431365
transform 1 0 28336 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_80_247
timestamp 1698431365
transform 1 0 29008 0 1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_80_311
timestamp 1698431365
transform 1 0 36176 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_80_317
timestamp 1698431365
transform 1 0 36848 0 1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_80_381
timestamp 1698431365
transform 1 0 44016 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_80_387
timestamp 1698431365
transform 1 0 44688 0 1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_80_451
timestamp 1698431365
transform 1 0 51856 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_80_457
timestamp 1698431365
transform 1 0 52528 0 1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_80_521
timestamp 1698431365
transform 1 0 59696 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_80_527
timestamp 1698431365
transform 1 0 60368 0 1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_80_591
timestamp 1698431365
transform 1 0 67536 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_80_597
timestamp 1698431365
transform 1 0 68208 0 1 65856
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_80_661
timestamp 1698431365
transform 1 0 75376 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_80_667
timestamp 1698431365
transform 1 0 76048 0 1 65856
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_80_675
timestamp 1698431365
transform 1 0 76944 0 1 65856
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_80_679
timestamp 1698431365
transform 1 0 77392 0 1 65856
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_81_2
timestamp 1698431365
transform 1 0 1568 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_81_4
timestamp 1698431365
transform 1 0 1792 0 -1 67424
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_81_23
timestamp 1698431365
transform 1 0 3920 0 -1 67424
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_81_55
timestamp 1698431365
transform 1 0 7504 0 -1 67424
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_81_63
timestamp 1698431365
transform 1 0 8400 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_81_67
timestamp 1698431365
transform 1 0 8848 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_81_69
timestamp 1698431365
transform 1 0 9072 0 -1 67424
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_81_72
timestamp 1698431365
transform 1 0 9408 0 -1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_81_136
timestamp 1698431365
transform 1 0 16576 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_81_142
timestamp 1698431365
transform 1 0 17248 0 -1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_81_206
timestamp 1698431365
transform 1 0 24416 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_81_212
timestamp 1698431365
transform 1 0 25088 0 -1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_81_276
timestamp 1698431365
transform 1 0 32256 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_81_282
timestamp 1698431365
transform 1 0 32928 0 -1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_81_346
timestamp 1698431365
transform 1 0 40096 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_81_352
timestamp 1698431365
transform 1 0 40768 0 -1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_81_416
timestamp 1698431365
transform 1 0 47936 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_81_422
timestamp 1698431365
transform 1 0 48608 0 -1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_81_486
timestamp 1698431365
transform 1 0 55776 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_81_492
timestamp 1698431365
transform 1 0 56448 0 -1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_81_556
timestamp 1698431365
transform 1 0 63616 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_81_562
timestamp 1698431365
transform 1 0 64288 0 -1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_81_626
timestamp 1698431365
transform 1 0 71456 0 -1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_81_632
timestamp 1698431365
transform 1 0 72128 0 -1 67424
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_81_664
timestamp 1698431365
transform 1 0 75712 0 -1 67424
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_82_28
timestamp 1698431365
transform 1 0 4480 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_82_32
timestamp 1698431365
transform 1 0 4928 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_82_34
timestamp 1698431365
transform 1 0 5152 0 1 67424
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_82_37
timestamp 1698431365
transform 1 0 5488 0 1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_82_101
timestamp 1698431365
transform 1 0 12656 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_82_107
timestamp 1698431365
transform 1 0 13328 0 1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_82_171
timestamp 1698431365
transform 1 0 20496 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_82_177
timestamp 1698431365
transform 1 0 21168 0 1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_82_241
timestamp 1698431365
transform 1 0 28336 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_82_247
timestamp 1698431365
transform 1 0 29008 0 1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_82_311
timestamp 1698431365
transform 1 0 36176 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_82_317
timestamp 1698431365
transform 1 0 36848 0 1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_82_381
timestamp 1698431365
transform 1 0 44016 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_82_387
timestamp 1698431365
transform 1 0 44688 0 1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_82_451
timestamp 1698431365
transform 1 0 51856 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_82_457
timestamp 1698431365
transform 1 0 52528 0 1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_82_521
timestamp 1698431365
transform 1 0 59696 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_82_527
timestamp 1698431365
transform 1 0 60368 0 1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_82_591
timestamp 1698431365
transform 1 0 67536 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_82_597
timestamp 1698431365
transform 1 0 68208 0 1 67424
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_82_661
timestamp 1698431365
transform 1 0 75376 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_82_667
timestamp 1698431365
transform 1 0 76048 0 1 67424
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_82_683
timestamp 1698431365
transform 1 0 77840 0 1 67424
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_82_687
timestamp 1698431365
transform 1 0 78288 0 1 67424
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_83_28
timestamp 1698431365
transform 1 0 4480 0 -1 68992
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_83_60
timestamp 1698431365
transform 1 0 8064 0 -1 68992
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_83_68
timestamp 1698431365
transform 1 0 8960 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_83_72
timestamp 1698431365
transform 1 0 9408 0 -1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_83_136
timestamp 1698431365
transform 1 0 16576 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_83_142
timestamp 1698431365
transform 1 0 17248 0 -1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_83_206
timestamp 1698431365
transform 1 0 24416 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_83_212
timestamp 1698431365
transform 1 0 25088 0 -1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_83_276
timestamp 1698431365
transform 1 0 32256 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_83_282
timestamp 1698431365
transform 1 0 32928 0 -1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_83_346
timestamp 1698431365
transform 1 0 40096 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_83_352
timestamp 1698431365
transform 1 0 40768 0 -1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_83_416
timestamp 1698431365
transform 1 0 47936 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_83_422
timestamp 1698431365
transform 1 0 48608 0 -1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_83_486
timestamp 1698431365
transform 1 0 55776 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_83_492
timestamp 1698431365
transform 1 0 56448 0 -1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_83_556
timestamp 1698431365
transform 1 0 63616 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_83_562
timestamp 1698431365
transform 1 0 64288 0 -1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_83_626
timestamp 1698431365
transform 1 0 71456 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_83_632
timestamp 1698431365
transform 1 0 72128 0 -1 68992
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_83_664
timestamp 1698431365
transform 1 0 75712 0 -1 68992
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_83_672
timestamp 1698431365
transform 1 0 76608 0 -1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_83_676
timestamp 1698431365
transform 1 0 77056 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_84_2
timestamp 1698431365
transform 1 0 1568 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_84_4
timestamp 1698431365
transform 1 0 1792 0 1 68992
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_84_17
timestamp 1698431365
transform 1 0 3248 0 1 68992
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_84_33
timestamp 1698431365
transform 1 0 5040 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_84_37
timestamp 1698431365
transform 1 0 5488 0 1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_84_101
timestamp 1698431365
transform 1 0 12656 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_84_107
timestamp 1698431365
transform 1 0 13328 0 1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_84_171
timestamp 1698431365
transform 1 0 20496 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_84_177
timestamp 1698431365
transform 1 0 21168 0 1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_84_241
timestamp 1698431365
transform 1 0 28336 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_84_247
timestamp 1698431365
transform 1 0 29008 0 1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_84_311
timestamp 1698431365
transform 1 0 36176 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_84_317
timestamp 1698431365
transform 1 0 36848 0 1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_84_381
timestamp 1698431365
transform 1 0 44016 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_84_387
timestamp 1698431365
transform 1 0 44688 0 1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_84_451
timestamp 1698431365
transform 1 0 51856 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_84_457
timestamp 1698431365
transform 1 0 52528 0 1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_84_521
timestamp 1698431365
transform 1 0 59696 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_84_527
timestamp 1698431365
transform 1 0 60368 0 1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_84_591
timestamp 1698431365
transform 1 0 67536 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_84_597
timestamp 1698431365
transform 1 0 68208 0 1 68992
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_84_661
timestamp 1698431365
transform 1 0 75376 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_84_667
timestamp 1698431365
transform 1 0 76048 0 1 68992
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_84_675
timestamp 1698431365
transform 1 0 76944 0 1 68992
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_84_679
timestamp 1698431365
transform 1 0 77392 0 1 68992
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_85_28
timestamp 1698431365
transform 1 0 4480 0 -1 70560
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_85_60
timestamp 1698431365
transform 1 0 8064 0 -1 70560
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_85_68
timestamp 1698431365
transform 1 0 8960 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_85_72
timestamp 1698431365
transform 1 0 9408 0 -1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_85_136
timestamp 1698431365
transform 1 0 16576 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_85_142
timestamp 1698431365
transform 1 0 17248 0 -1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_85_206
timestamp 1698431365
transform 1 0 24416 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_85_212
timestamp 1698431365
transform 1 0 25088 0 -1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_85_276
timestamp 1698431365
transform 1 0 32256 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_85_282
timestamp 1698431365
transform 1 0 32928 0 -1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_85_346
timestamp 1698431365
transform 1 0 40096 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_85_352
timestamp 1698431365
transform 1 0 40768 0 -1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_85_416
timestamp 1698431365
transform 1 0 47936 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_85_422
timestamp 1698431365
transform 1 0 48608 0 -1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_85_486
timestamp 1698431365
transform 1 0 55776 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_85_492
timestamp 1698431365
transform 1 0 56448 0 -1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_85_556
timestamp 1698431365
transform 1 0 63616 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_85_562
timestamp 1698431365
transform 1 0 64288 0 -1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_85_626
timestamp 1698431365
transform 1 0 71456 0 -1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_85_632
timestamp 1698431365
transform 1 0 72128 0 -1 70560
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_85_664
timestamp 1698431365
transform 1 0 75712 0 -1 70560
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_85_680
timestamp 1698431365
transform 1 0 77504 0 -1 70560
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_86_28
timestamp 1698431365
transform 1 0 4480 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_86_32
timestamp 1698431365
transform 1 0 4928 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_86_34
timestamp 1698431365
transform 1 0 5152 0 1 70560
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_86_37
timestamp 1698431365
transform 1 0 5488 0 1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_86_101
timestamp 1698431365
transform 1 0 12656 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_86_107
timestamp 1698431365
transform 1 0 13328 0 1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_86_171
timestamp 1698431365
transform 1 0 20496 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_86_177
timestamp 1698431365
transform 1 0 21168 0 1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_86_241
timestamp 1698431365
transform 1 0 28336 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_86_247
timestamp 1698431365
transform 1 0 29008 0 1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_86_311
timestamp 1698431365
transform 1 0 36176 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_86_317
timestamp 1698431365
transform 1 0 36848 0 1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_86_381
timestamp 1698431365
transform 1 0 44016 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_86_387
timestamp 1698431365
transform 1 0 44688 0 1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_86_451
timestamp 1698431365
transform 1 0 51856 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_86_457
timestamp 1698431365
transform 1 0 52528 0 1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_86_521
timestamp 1698431365
transform 1 0 59696 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_86_527
timestamp 1698431365
transform 1 0 60368 0 1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_86_591
timestamp 1698431365
transform 1 0 67536 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_86_597
timestamp 1698431365
transform 1 0 68208 0 1 70560
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_86_661
timestamp 1698431365
transform 1 0 75376 0 1 70560
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_86_667
timestamp 1698431365
transform 1 0 76048 0 1 70560
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_86_675
timestamp 1698431365
transform 1 0 76944 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_86_677
timestamp 1698431365
transform 1 0 77168 0 1 70560
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_87_2
timestamp 1698431365
transform 1 0 1568 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_87_30
timestamp 1698431365
transform 1 0 4704 0 -1 72128
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_87_62
timestamp 1698431365
transform 1 0 8288 0 -1 72128
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_87_72
timestamp 1698431365
transform 1 0 9408 0 -1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_87_136
timestamp 1698431365
transform 1 0 16576 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_87_142
timestamp 1698431365
transform 1 0 17248 0 -1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_87_206
timestamp 1698431365
transform 1 0 24416 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_87_212
timestamp 1698431365
transform 1 0 25088 0 -1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_87_276
timestamp 1698431365
transform 1 0 32256 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_87_282
timestamp 1698431365
transform 1 0 32928 0 -1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_87_346
timestamp 1698431365
transform 1 0 40096 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_87_352
timestamp 1698431365
transform 1 0 40768 0 -1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_87_416
timestamp 1698431365
transform 1 0 47936 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_87_422
timestamp 1698431365
transform 1 0 48608 0 -1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_87_486
timestamp 1698431365
transform 1 0 55776 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_87_492
timestamp 1698431365
transform 1 0 56448 0 -1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_87_556
timestamp 1698431365
transform 1 0 63616 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_87_562
timestamp 1698431365
transform 1 0 64288 0 -1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_87_626
timestamp 1698431365
transform 1 0 71456 0 -1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_87_632
timestamp 1698431365
transform 1 0 72128 0 -1 72128
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_87_664
timestamp 1698431365
transform 1 0 75712 0 -1 72128
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_88_28
timestamp 1698431365
transform 1 0 4480 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_88_32
timestamp 1698431365
transform 1 0 4928 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_88_34
timestamp 1698431365
transform 1 0 5152 0 1 72128
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_88_37
timestamp 1698431365
transform 1 0 5488 0 1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_88_101
timestamp 1698431365
transform 1 0 12656 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_88_107
timestamp 1698431365
transform 1 0 13328 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_88_111
timestamp 1698431365
transform 1 0 13776 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_88_113
timestamp 1698431365
transform 1 0 14000 0 1 72128
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_88_116
timestamp 1698431365
transform 1 0 14336 0 1 72128
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_88_148
timestamp 1698431365
transform 1 0 17920 0 1 72128
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_88_164
timestamp 1698431365
transform 1 0 19712 0 1 72128
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_88_172
timestamp 1698431365
transform 1 0 20608 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_88_174
timestamp 1698431365
transform 1 0 20832 0 1 72128
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_88_177
timestamp 1698431365
transform 1 0 21168 0 1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_88_241
timestamp 1698431365
transform 1 0 28336 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_88_247
timestamp 1698431365
transform 1 0 29008 0 1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_88_311
timestamp 1698431365
transform 1 0 36176 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_88_317
timestamp 1698431365
transform 1 0 36848 0 1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_88_381
timestamp 1698431365
transform 1 0 44016 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_88_387
timestamp 1698431365
transform 1 0 44688 0 1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_88_451
timestamp 1698431365
transform 1 0 51856 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_88_457
timestamp 1698431365
transform 1 0 52528 0 1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_88_521
timestamp 1698431365
transform 1 0 59696 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_88_527
timestamp 1698431365
transform 1 0 60368 0 1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_88_591
timestamp 1698431365
transform 1 0 67536 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_88_597
timestamp 1698431365
transform 1 0 68208 0 1 72128
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_88_661
timestamp 1698431365
transform 1 0 75376 0 1 72128
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_88_667
timestamp 1698431365
transform 1 0 76048 0 1 72128
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_88_675
timestamp 1698431365
transform 1 0 76944 0 1 72128
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_88_678
timestamp 1698431365
transform 1 0 77280 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_89_34
timestamp 1698431365
transform 1 0 5152 0 -1 73696
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_89_66
timestamp 1698431365
transform 1 0 8736 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_89_72
timestamp 1698431365
transform 1 0 9408 0 -1 73696
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_89_142
timestamp 1698431365
transform 1 0 17248 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_89_146
timestamp 1698431365
transform 1 0 17696 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_89_148
timestamp 1698431365
transform 1 0 17920 0 -1 73696
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_89_151
timestamp 1698431365
transform 1 0 18256 0 -1 73696
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_89_183
timestamp 1698431365
transform 1 0 21840 0 -1 73696
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_89_199
timestamp 1698431365
transform 1 0 23632 0 -1 73696
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_89_207
timestamp 1698431365
transform 1 0 24528 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_89_209
timestamp 1698431365
transform 1 0 24752 0 -1 73696
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_89_212
timestamp 1698431365
transform 1 0 25088 0 -1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_89_276
timestamp 1698431365
transform 1 0 32256 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_89_282
timestamp 1698431365
transform 1 0 32928 0 -1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_89_346
timestamp 1698431365
transform 1 0 40096 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_89_352
timestamp 1698431365
transform 1 0 40768 0 -1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_89_416
timestamp 1698431365
transform 1 0 47936 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_89_422
timestamp 1698431365
transform 1 0 48608 0 -1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_89_486
timestamp 1698431365
transform 1 0 55776 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_89_492
timestamp 1698431365
transform 1 0 56448 0 -1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_89_556
timestamp 1698431365
transform 1 0 63616 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_89_562
timestamp 1698431365
transform 1 0 64288 0 -1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_89_626
timestamp 1698431365
transform 1 0 71456 0 -1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_89_632
timestamp 1698431365
transform 1 0 72128 0 -1 73696
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_89_664
timestamp 1698431365
transform 1 0 75712 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_89_666
timestamp 1698431365
transform 1 0 75936 0 -1 73696
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_89_669
timestamp 1698431365
transform 1 0 76272 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_89_673
timestamp 1698431365
transform 1 0 76720 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_89_675
timestamp 1698431365
transform 1 0 76944 0 -1 73696
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_89_678
timestamp 1698431365
transform 1 0 77280 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_90_34
timestamp 1698431365
transform 1 0 5152 0 1 73696
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_90_37
timestamp 1698431365
transform 1 0 5488 0 1 73696
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_90_69
timestamp 1698431365
transform 1 0 9072 0 1 73696
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_90_77
timestamp 1698431365
transform 1 0 9968 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_90_107
timestamp 1698431365
transform 1 0 13328 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_90_111
timestamp 1698431365
transform 1 0 13776 0 1 73696
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_90_114
timestamp 1698431365
transform 1 0 14112 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_90_118
timestamp 1698431365
transform 1 0 14560 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_90_122
timestamp 1698431365
transform 1 0 15008 0 1 73696
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_90_177
timestamp 1698431365
transform 1 0 21168 0 1 73696
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_90_195
timestamp 1698431365
transform 1 0 23184 0 1 73696
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_90_227
timestamp 1698431365
transform 1 0 26768 0 1 73696
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_90_243
timestamp 1698431365
transform 1 0 28560 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_90_247
timestamp 1698431365
transform 1 0 29008 0 1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_90_311
timestamp 1698431365
transform 1 0 36176 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_90_317
timestamp 1698431365
transform 1 0 36848 0 1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_90_381
timestamp 1698431365
transform 1 0 44016 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_90_387
timestamp 1698431365
transform 1 0 44688 0 1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_90_451
timestamp 1698431365
transform 1 0 51856 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_90_457
timestamp 1698431365
transform 1 0 52528 0 1 73696
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_90_489
timestamp 1698431365
transform 1 0 56112 0 1 73696
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_90_505
timestamp 1698431365
transform 1 0 57904 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_90_509
timestamp 1698431365
transform 1 0 58352 0 1 73696
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_90_512
timestamp 1698431365
transform 1 0 58688 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_90_514
timestamp 1698431365
transform 1 0 58912 0 1 73696
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_90_517
timestamp 1698431365
transform 1 0 59248 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_90_521
timestamp 1698431365
transform 1 0 59696 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_90_527
timestamp 1698431365
transform 1 0 60368 0 1 73696
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_90_591
timestamp 1698431365
transform 1 0 67536 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_90_597
timestamp 1698431365
transform 1 0 68208 0 1 73696
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_90_629
timestamp 1698431365
transform 1 0 71792 0 1 73696
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_90_645
timestamp 1698431365
transform 1 0 73584 0 1 73696
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_90_653
timestamp 1698431365
transform 1 0 74480 0 1 73696
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_90_657
timestamp 1698431365
transform 1 0 74928 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_90_661
timestamp 1698431365
transform 1 0 75376 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_90_667
timestamp 1698431365
transform 1 0 76048 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_90_671
timestamp 1698431365
transform 1 0 76496 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_90_673
timestamp 1698431365
transform 1 0 76720 0 1 73696
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_91_34
timestamp 1698431365
transform 1 0 5152 0 -1 75264
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_91_66
timestamp 1698431365
transform 1 0 8736 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_91_72
timestamp 1698431365
transform 1 0 9408 0 -1 75264
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_91_142
timestamp 1698431365
transform 1 0 17248 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_91_146
timestamp 1698431365
transform 1 0 17696 0 -1 75264
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_91_149
timestamp 1698431365
transform 1 0 18032 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_91_153
timestamp 1698431365
transform 1 0 18480 0 -1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_91_163
timestamp 1698431365
transform 1 0 19600 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_91_201
timestamp 1698431365
transform 1 0 23856 0 -1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_91_209
timestamp 1698431365
transform 1 0 24752 0 -1 75264
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_91_212
timestamp 1698431365
transform 1 0 25088 0 -1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_91_276
timestamp 1698431365
transform 1 0 32256 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_91_282
timestamp 1698431365
transform 1 0 32928 0 -1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_91_290
timestamp 1698431365
transform 1 0 33824 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_91_294
timestamp 1698431365
transform 1 0 34272 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_91_296
timestamp 1698431365
transform 1 0 34496 0 -1 75264
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_91_299
timestamp 1698431365
transform 1 0 34832 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_91_303
timestamp 1698431365
transform 1 0 35280 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_91_307
timestamp 1698431365
transform 1 0 35728 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_91_311
timestamp 1698431365
transform 1 0 36176 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_91_315
timestamp 1698431365
transform 1 0 36624 0 -1 75264
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_91_318
timestamp 1698431365
transform 1 0 36960 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_91_322
timestamp 1698431365
transform 1 0 37408 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_91_326
timestamp 1698431365
transform 1 0 37856 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_91_328
timestamp 1698431365
transform 1 0 38080 0 -1 75264
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_91_331
timestamp 1698431365
transform 1 0 38416 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_91_335
timestamp 1698431365
transform 1 0 38864 0 -1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_91_343
timestamp 1698431365
transform 1 0 39760 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_91_347
timestamp 1698431365
transform 1 0 40208 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_91_349
timestamp 1698431365
transform 1 0 40432 0 -1 75264
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_91_352
timestamp 1698431365
transform 1 0 40768 0 -1 75264
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_91_384
timestamp 1698431365
transform 1 0 44352 0 -1 75264
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_91_400
timestamp 1698431365
transform 1 0 46144 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_91_404
timestamp 1698431365
transform 1 0 46592 0 -1 75264
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_91_407
timestamp 1698431365
transform 1 0 46928 0 -1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_91_415
timestamp 1698431365
transform 1 0 47824 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_91_419
timestamp 1698431365
transform 1 0 48272 0 -1 75264
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_91_422
timestamp 1698431365
transform 1 0 48608 0 -1 75264
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_91_454
timestamp 1698431365
transform 1 0 52192 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_91_460
timestamp 1698431365
transform 1 0 52864 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_91_464
timestamp 1698431365
transform 1 0 53312 0 -1 75264
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_91_467
timestamp 1698431365
transform 1 0 53648 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_91_471
timestamp 1698431365
transform 1 0 54096 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_91_475
timestamp 1698431365
transform 1 0 54544 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_91_479
timestamp 1698431365
transform 1 0 54992 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_91_483
timestamp 1698431365
transform 1 0 55440 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_91_487
timestamp 1698431365
transform 1 0 55888 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_91_489
timestamp 1698431365
transform 1 0 56112 0 -1 75264
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_91_492
timestamp 1698431365
transform 1 0 56448 0 -1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_91_500
timestamp 1698431365
transform 1 0 57344 0 -1 75264
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_91_529
timestamp 1698431365
transform 1 0 60592 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_91_533
timestamp 1698431365
transform 1 0 61040 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_91_537
timestamp 1698431365
transform 1 0 61488 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_91_541
timestamp 1698431365
transform 1 0 61936 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_91_545
timestamp 1698431365
transform 1 0 62384 0 -1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_91_553
timestamp 1698431365
transform 1 0 63280 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_91_557
timestamp 1698431365
transform 1 0 63728 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_91_559
timestamp 1698431365
transform 1 0 63952 0 -1 75264
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_91_562
timestamp 1698431365
transform 1 0 64288 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_91_566
timestamp 1698431365
transform 1 0 64736 0 -1 75264
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_91_632
timestamp 1698431365
transform 1 0 72128 0 -1 75264
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_91_650
timestamp 1698431365
transform 1 0 74144 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_91_654
timestamp 1698431365
transform 1 0 74592 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_91_658
timestamp 1698431365
transform 1 0 75040 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_91_684
timestamp 1698431365
transform 1 0 77952 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_92_34
timestamp 1698431365
transform 1 0 5152 0 1 75264
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_92_37
timestamp 1698431365
transform 1 0 5488 0 1 75264
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_92_69
timestamp 1698431365
transform 1 0 9072 0 1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_77
timestamp 1698431365
transform 1 0 9968 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_107
timestamp 1698431365
transform 1 0 13328 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_111
timestamp 1698431365
transform 1 0 13776 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_92_113
timestamp 1698431365
transform 1 0 14000 0 1 75264
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_116
timestamp 1698431365
transform 1 0 14336 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_120
timestamp 1698431365
transform 1 0 14784 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_92_122
timestamp 1698431365
transform 1 0 15008 0 1 75264
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_207
timestamp 1698431365
transform 1 0 24528 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_211
timestamp 1698431365
transform 1 0 24976 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_92_215
timestamp 1698431365
transform 1 0 25424 0 1 75264
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_92_231
timestamp 1698431365
transform 1 0 27216 0 1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_92_239
timestamp 1698431365
transform 1 0 28112 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_243
timestamp 1698431365
transform 1 0 28560 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_92_247
timestamp 1698431365
transform 1 0 29008 0 1 75264
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_313
timestamp 1698431365
transform 1 0 36400 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_317
timestamp 1698431365
transform 1 0 36848 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_337
timestamp 1698431365
transform 1 0 39088 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_92_339
timestamp 1698431365
transform 1 0 39312 0 1 75264
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_92_342
timestamp 1698431365
transform 1 0 39648 0 1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_350
timestamp 1698431365
transform 1 0 40544 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_92_352
timestamp 1698431365
transform 1 0 40768 0 1 75264
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_355
timestamp 1698431365
transform 1 0 41104 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_365
timestamp 1698431365
transform 1 0 42224 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_92_369
timestamp 1698431365
transform 1 0 42672 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_92_373
timestamp 1698431365
transform 1 0 43120 0 1 75264
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_376
timestamp 1698431365
transform 1 0 43456 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_92_378
timestamp 1698431365
transform 1 0 43680 0 1 75264
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_381
timestamp 1698431365
transform 1 0 44016 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_387
timestamp 1698431365
transform 1 0 44688 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_397
timestamp 1698431365
transform 1 0 45808 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_401
timestamp 1698431365
transform 1 0 46256 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_405
timestamp 1698431365
transform 1 0 46704 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_415
timestamp 1698431365
transform 1 0 47824 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_419
timestamp 1698431365
transform 1 0 48272 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_423
timestamp 1698431365
transform 1 0 48720 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_427
timestamp 1698431365
transform 1 0 49168 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_439
timestamp 1698431365
transform 1 0 50512 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_443
timestamp 1698431365
transform 1 0 50960 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_447
timestamp 1698431365
transform 1 0 51408 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_451
timestamp 1698431365
transform 1 0 51856 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_465
timestamp 1698431365
transform 1 0 53424 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_523
timestamp 1698431365
transform 1 0 59920 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_547
timestamp 1698431365
transform 1 0 62608 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_551
timestamp 1698431365
transform 1 0 63056 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_555
timestamp 1698431365
transform 1 0 63504 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_559
timestamp 1698431365
transform 1 0 63952 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_92_563
timestamp 1698431365
transform 1 0 64400 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_575
timestamp 1698431365
transform 1 0 65744 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_579
timestamp 1698431365
transform 1 0 66192 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_583
timestamp 1698431365
transform 1 0 66640 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_587
timestamp 1698431365
transform 1 0 67088 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_92_589
timestamp 1698431365
transform 1 0 67312 0 1 75264
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_592
timestamp 1698431365
transform 1 0 67648 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_92_594
timestamp 1698431365
transform 1 0 67872 0 1 75264
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_597
timestamp 1698431365
transform 1 0 68208 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_601
timestamp 1698431365
transform 1 0 68656 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_92_603
timestamp 1698431365
transform 1 0 68880 0 1 75264
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_92_606
timestamp 1698431365
transform 1 0 69216 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_610
timestamp 1698431365
transform 1 0 69664 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_92_614
timestamp 1698431365
transform 1 0 70112 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_92_620
timestamp 1698431365
transform 1 0 70784 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_626
timestamp 1698431365
transform 1 0 71456 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_92_628
timestamp 1698431365
transform 1 0 71680 0 1 75264
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_631
timestamp 1698431365
transform 1 0 72016 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_641
timestamp 1698431365
transform 1 0 73136 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_645
timestamp 1698431365
transform 1 0 73584 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_649
timestamp 1698431365
transform 1 0 74032 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_92_651
timestamp 1698431365
transform 1 0 74256 0 1 75264
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_92_654
timestamp 1698431365
transform 1 0 74592 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_92_656
timestamp 1698431365
transform 1 0 74816 0 1 75264
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_92_679
timestamp 1698431365
transform 1 0 77392 0 1 75264
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_93_42
timestamp 1698431365
transform 1 0 6048 0 -1 76832
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_93_58
timestamp 1698431365
transform 1 0 7840 0 -1 76832
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_93_66
timestamp 1698431365
transform 1 0 8736 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_93_70
timestamp 1698431365
transform 1 0 9184 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_93_74
timestamp 1698431365
transform 1 0 9632 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_93_104
timestamp 1698431365
transform 1 0 12992 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_93_108
timestamp 1698431365
transform 1 0 13440 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_93_138
timestamp 1698431365
transform 1 0 16800 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_93_142
timestamp 1698431365
transform 1 0 17248 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_93_172
timestamp 1698431365
transform 1 0 20608 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_93_206
timestamp 1698431365
transform 1 0 24416 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_93_208
timestamp 1698431365
transform 1 0 24640 0 -1 76832
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_93_213
timestamp 1698431365
transform 1 0 25200 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_93_219
timestamp 1698431365
transform 1 0 25872 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_93_225
timestamp 1698431365
transform 1 0 26544 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_93_231
timestamp 1698431365
transform 1 0 27216 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_93_237
timestamp 1698431365
transform 1 0 27888 0 -1 76832
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_93_244
timestamp 1698431365
transform 1 0 28672 0 -1 76832
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_93_249
timestamp 1698431365
transform 1 0 29232 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_93_255
timestamp 1698431365
transform 1 0 29904 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_93_261
timestamp 1698431365
transform 1 0 30576 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_93_267
timestamp 1698431365
transform 1 0 31248 0 -1 76832
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_93_274
timestamp 1698431365
transform 1 0 32032 0 -1 76832
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_93_279
timestamp 1698431365
transform 1 0 32592 0 -1 76832
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_93_308
timestamp 1698431365
transform 1 0 35840 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_93_342
timestamp 1698431365
transform 1 0 39648 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_93_344
timestamp 1698431365
transform 1 0 39872 0 -1 76832
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_93_361
timestamp 1698431365
transform 1 0 41776 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_93_373
timestamp 1698431365
transform 1 0 43120 0 -1 76832
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_93_478
timestamp 1698431365
transform 1 0 54880 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_93_482
timestamp 1698431365
transform 1 0 55328 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_93_576
timestamp 1698431365
transform 1 0 65856 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_93_644
timestamp 1698431365
transform 1 0 73472 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input1
timestamp 1698431365
transform 1 0 25200 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input2
timestamp 1698431365
transform 1 0 33600 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input3
timestamp 1698431365
transform 1 0 31136 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input4
timestamp 1698431365
transform 1 0 27328 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input5
timestamp 1698431365
transform 1 0 28448 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input6
timestamp 1698431365
transform 1 0 35280 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input7
timestamp 1698431365
transform 1 0 29120 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input8
timestamp 1698431365
transform 1 0 29792 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input9
timestamp 1698431365
transform 1 0 35952 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input10
timestamp 1698431365
transform 1 0 30464 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input11
timestamp 1698431365
transform 1 0 36960 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input12
timestamp 1698431365
transform 1 0 23520 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input13
timestamp 1698431365
transform 1 0 37632 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input14
timestamp 1698431365
transform -1 0 49504 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input15
timestamp 1698431365
transform 1 0 31136 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input16
timestamp 1698431365
transform -1 0 48832 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input17
timestamp 1698431365
transform -1 0 49280 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input18
timestamp 1698431365
transform -1 0 42112 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input19
timestamp 1698431365
transform -1 0 50176 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input20
timestamp 1698431365
transform -1 0 50848 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input21
timestamp 1698431365
transform -1 0 46592 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input22
timestamp 1698431365
transform -1 0 48272 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input23
timestamp 1698431365
transform 1 0 22176 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input24
timestamp 1698431365
transform -1 0 49504 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input25
timestamp 1698431365
transform -1 0 50176 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input26
timestamp 1698431365
transform 1 0 24640 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input27
timestamp 1698431365
transform 1 0 29792 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input28
timestamp 1698431365
transform 1 0 24192 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input29
timestamp 1698431365
transform 1 0 23520 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input30
timestamp 1698431365
transform 1 0 25984 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input31
timestamp 1698431365
transform 1 0 28112 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input32
timestamp 1698431365
transform 1 0 26656 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input33
timestamp 1698431365
transform -1 0 49504 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input34
timestamp 1698431365
transform 1 0 3808 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input35
timestamp 1698431365
transform 1 0 10192 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input36
timestamp 1698431365
transform 1 0 8288 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input37
timestamp 1698431365
transform 1 0 13440 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input38
timestamp 1698431365
transform 1 0 9520 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input39
timestamp 1698431365
transform 1 0 9408 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input40
timestamp 1698431365
transform 1 0 10080 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input41
timestamp 1698431365
transform 1 0 14336 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input42
timestamp 1698431365
transform 1 0 12096 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input43
timestamp 1698431365
transform 1 0 13888 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input44
timestamp 1698431365
transform 1 0 14560 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input45
timestamp 1698431365
transform 1 0 5712 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input46
timestamp 1698431365
transform 1 0 15232 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input47
timestamp 1698431365
transform 1 0 18144 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input48
timestamp 1698431365
transform 1 0 17024 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input49
timestamp 1698431365
transform 1 0 18816 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input50
timestamp 1698431365
transform 1 0 17696 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input51
timestamp 1698431365
transform 1 0 19488 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input52
timestamp 1698431365
transform 1 0 18368 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input53
timestamp 1698431365
transform 1 0 19040 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input54
timestamp 1698431365
transform 1 0 19712 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input55
timestamp 1698431365
transform 1 0 22176 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input56
timestamp 1698431365
transform 1 0 4480 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input57
timestamp 1698431365
transform 1 0 20832 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input58
timestamp 1698431365
transform 1 0 21504 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input59
timestamp 1698431365
transform 1 0 6272 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input60
timestamp 1698431365
transform 1 0 6496 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input61
timestamp 1698431365
transform 1 0 5600 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input62
timestamp 1698431365
transform 1 0 6272 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input63
timestamp 1698431365
transform 1 0 6944 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input64
timestamp 1698431365
transform 1 0 8512 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input65
timestamp 1698431365
transform 1 0 7616 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input66
timestamp 1698431365
transform -1 0 51968 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input67
timestamp 1698431365
transform -1 0 52640 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input68
timestamp 1698431365
transform -1 0 53312 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input69
timestamp 1698431365
transform -1 0 53984 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input70
timestamp 1698431365
transform 1 0 2240 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input71
timestamp 1698431365
transform 1 0 1568 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input72
timestamp 1698431365
transform 1 0 1568 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input73
timestamp 1698431365
transform 1 0 1568 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input74
timestamp 1698431365
transform 1 0 1568 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input75
timestamp 1698431365
transform 1 0 1568 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input76
timestamp 1698431365
transform 1 0 1568 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input77
timestamp 1698431365
transform 1 0 1568 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input78
timestamp 1698431365
transform 1 0 1568 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input79
timestamp 1698431365
transform 1 0 1568 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input80
timestamp 1698431365
transform 1 0 1568 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input81
timestamp 1698431365
transform 1 0 1568 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input82
timestamp 1698431365
transform 1 0 1568 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input83
timestamp 1698431365
transform 1 0 1568 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input84
timestamp 1698431365
transform 1 0 1568 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input85
timestamp 1698431365
transform 1 0 1568 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input86
timestamp 1698431365
transform 1 0 1568 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input87
timestamp 1698431365
transform 1 0 1568 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input88
timestamp 1698431365
transform 1 0 1568 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input89
timestamp 1698431365
transform 1 0 1568 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input90
timestamp 1698431365
transform 1 0 1568 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input91
timestamp 1698431365
transform 1 0 1568 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input92
timestamp 1698431365
transform 1 0 1568 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input93
timestamp 1698431365
transform 1 0 1568 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input94
timestamp 1698431365
transform 1 0 1568 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input95
timestamp 1698431365
transform 1 0 1568 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input96
timestamp 1698431365
transform 1 0 1568 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input97
timestamp 1698431365
transform 1 0 1568 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input98
timestamp 1698431365
transform 1 0 1568 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input99
timestamp 1698431365
transform 1 0 1568 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input100
timestamp 1698431365
transform 1 0 1568 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input101
timestamp 1698431365
transform 1 0 1568 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input102
timestamp 1698431365
transform 1 0 76048 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input103
timestamp 1698431365
transform -1 0 78400 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input104
timestamp 1698431365
transform -1 0 78400 0 1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input105
timestamp 1698431365
transform -1 0 78400 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input106
timestamp 1698431365
transform -1 0 78400 0 1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input107
timestamp 1698431365
transform -1 0 78400 0 1 58016
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input108
timestamp 1698431365
transform -1 0 78400 0 -1 59584
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input109
timestamp 1698431365
transform -1 0 78400 0 -1 61152
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input110
timestamp 1698431365
transform -1 0 78400 0 1 61152
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input111
timestamp 1698431365
transform -1 0 78400 0 1 62720
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input112
timestamp 1698431365
transform -1 0 78400 0 -1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input113
timestamp 1698431365
transform -1 0 78400 0 1 64288
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input114
timestamp 1698431365
transform -1 0 78400 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input115
timestamp 1698431365
transform -1 0 78400 0 1 65856
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input116
timestamp 1698431365
transform -1 0 78400 0 -1 67424
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input117
timestamp 1698431365
transform -1 0 78400 0 -1 68992
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input118
timestamp 1698431365
transform -1 0 78400 0 1 68992
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input119
timestamp 1698431365
transform -1 0 78400 0 1 70560
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input120
timestamp 1698431365
transform -1 0 78400 0 -1 72128
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input121
timestamp 1698431365
transform -1 0 78400 0 1 72128
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input122
timestamp 1698431365
transform -1 0 78400 0 1 73696
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input123
timestamp 1698431365
transform -1 0 78400 0 -1 73696
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input124
timestamp 1698431365
transform -1 0 78400 0 1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input125
timestamp 1698431365
transform -1 0 78400 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input126
timestamp 1698431365
transform -1 0 77056 0 -1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input127
timestamp 1698431365
transform -1 0 77728 0 1 73696
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input128
timestamp 1698431365
transform -1 0 78400 0 1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input129
timestamp 1698431365
transform -1 0 78400 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input130
timestamp 1698431365
transform -1 0 78400 0 1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input131
timestamp 1698431365
transform -1 0 78400 0 1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input132
timestamp 1698431365
transform -1 0 78400 0 -1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input133
timestamp 1698431365
transform -1 0 78400 0 -1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input134
timestamp 1698431365
transform -1 0 78400 0 1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input135
timestamp 1698431365
transform -1 0 77504 0 -1 76832
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input136
timestamp 1698431365
transform -1 0 77728 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input137
timestamp 1698431365
transform -1 0 78400 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input138
timestamp 1698431365
transform -1 0 78400 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input139
timestamp 1698431365
transform 1 0 77056 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input140
timestamp 1698431365
transform -1 0 78400 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input141
timestamp 1698431365
transform 1 0 74704 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input142
timestamp 1698431365
transform -1 0 78400 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input143
timestamp 1698431365
transform -1 0 78400 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input144
timestamp 1698431365
transform 1 0 74480 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input145
timestamp 1698431365
transform -1 0 78400 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input146
timestamp 1698431365
transform -1 0 76944 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input147
timestamp 1698431365
transform -1 0 78400 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input148
timestamp 1698431365
transform -1 0 77728 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input149
timestamp 1698431365
transform -1 0 78400 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input150
timestamp 1698431365
transform -1 0 78400 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input151
timestamp 1698431365
transform -1 0 78400 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input152
timestamp 1698431365
transform -1 0 78400 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input153
timestamp 1698431365
transform 1 0 74144 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input154
timestamp 1698431365
transform 1 0 74816 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input155
timestamp 1698431365
transform 1 0 75488 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input156
timestamp 1698431365
transform 1 0 74480 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input157
timestamp 1698431365
transform 1 0 77728 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input158
timestamp 1698431365
transform -1 0 77728 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input159
timestamp 1698431365
transform -1 0 78400 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input160
timestamp 1698431365
transform 1 0 74816 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input161
timestamp 1698431365
transform -1 0 78400 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input162
timestamp 1698431365
transform -1 0 78400 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input163
timestamp 1698431365
transform -1 0 77728 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input164
timestamp 1698431365
transform -1 0 78400 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input165
timestamp 1698431365
transform -1 0 78400 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input166
timestamp 1698431365
transform -1 0 78400 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input167
timestamp 1698431365
transform -1 0 78400 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input168
timestamp 1698431365
transform 1 0 33712 0 1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input169
timestamp 1698431365
transform 1 0 40880 0 -1 76832
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input170
timestamp 1698431365
transform 1 0 41552 0 1 75264
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input171
timestamp 1698431365
transform 1 0 42224 0 -1 76832
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input172
timestamp 1698431365
transform 1 0 43456 0 -1 76832
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input173
timestamp 1698431365
transform 1 0 44352 0 -1 76832
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input174
timestamp 1698431365
transform -1 0 46144 0 -1 76832
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input175
timestamp 1698431365
transform 1 0 44912 0 1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input176
timestamp 1698431365
transform -1 0 47040 0 -1 76832
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input177
timestamp 1698431365
transform -1 0 48160 0 -1 76832
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input178
timestamp 1698431365
transform 1 0 46928 0 1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input179
timestamp 1698431365
transform 1 0 34608 0 1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input180
timestamp 1698431365
transform 1 0 48160 0 -1 76832
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input181
timestamp 1698431365
transform 1 0 49056 0 -1 76832
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input182
timestamp 1698431365
transform 1 0 49952 0 -1 76832
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input183
timestamp 1698431365
transform 1 0 49616 0 1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input184
timestamp 1698431365
transform 1 0 51072 0 -1 76832
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input185
timestamp 1698431365
transform 1 0 51968 0 -1 76832
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input186
timestamp 1698431365
transform 1 0 52864 0 -1 76832
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input187
timestamp 1698431365
transform 1 0 52528 0 1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input188
timestamp 1698431365
transform 1 0 53760 0 -1 76832
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input189
timestamp 1698431365
transform 1 0 53648 0 1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input190
timestamp 1698431365
transform 1 0 35504 0 1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input191
timestamp 1698431365
transform 1 0 54544 0 1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input192
timestamp 1698431365
transform 1 0 55440 0 1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input193
timestamp 1698431365
transform -1 0 36736 0 -1 76832
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input194
timestamp 1698431365
transform 1 0 36736 0 -1 76832
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input195
timestamp 1698431365
transform 1 0 37296 0 1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input196
timestamp 1698431365
transform 1 0 38192 0 1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input197
timestamp 1698431365
transform -1 0 38528 0 -1 76832
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input198
timestamp 1698431365
transform -1 0 39424 0 -1 76832
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input199
timestamp 1698431365
transform 1 0 39984 0 -1 76832
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input200
timestamp 1698431365
transform 1 0 32816 0 1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input201
timestamp 1698431365
transform 1 0 59248 0 1 75264
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input202
timestamp 1698431365
transform 1 0 65072 0 1 75264
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input203
timestamp 1698431365
transform 1 0 66304 0 -1 76832
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input204
timestamp 1698431365
transform 1 0 66976 0 -1 76832
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input205
timestamp 1698431365
transform 1 0 67648 0 -1 76832
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input206
timestamp 1698431365
transform 1 0 68320 0 -1 76832
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input207
timestamp 1698431365
transform 1 0 69216 0 -1 76832
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input208
timestamp 1698431365
transform 1 0 70112 0 -1 76832
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input209
timestamp 1698431365
transform 1 0 70784 0 -1 76832
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input210
timestamp 1698431365
transform 1 0 71456 0 -1 76832
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input211
timestamp 1698431365
transform 1 0 72128 0 -1 76832
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input212
timestamp 1698431365
transform 1 0 60368 0 1 75264
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input213
timestamp 1698431365
transform -1 0 73472 0 -1 76832
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input214
timestamp 1698431365
transform 1 0 72464 0 1 75264
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input215
timestamp 1698431365
transform -1 0 74592 0 -1 76832
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input216
timestamp 1698431365
transform -1 0 75264 0 -1 76832
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input217
timestamp 1698431365
transform -1 0 75936 0 -1 76832
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input218
timestamp 1698431365
transform -1 0 76608 0 -1 76832
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input219
timestamp 1698431365
transform 1 0 76048 0 1 75264
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input220
timestamp 1698431365
transform 1 0 76720 0 1 75264
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input221
timestamp 1698431365
transform 1 0 77728 0 -1 76832
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input222
timestamp 1698431365
transform 1 0 77056 0 -1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input223
timestamp 1698431365
transform -1 0 62272 0 -1 76832
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input224
timestamp 1698431365
transform 1 0 75152 0 1 75264
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input225
timestamp 1698431365
transform -1 0 76160 0 -1 75264
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input226
timestamp 1698431365
transform 1 0 61040 0 1 75264
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input227
timestamp 1698431365
transform 1 0 61936 0 1 75264
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input228
timestamp 1698431365
transform -1 0 63168 0 -1 76832
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input229
timestamp 1698431365
transform 1 0 63168 0 -1 76832
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input230
timestamp 1698431365
transform 1 0 63840 0 -1 76832
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input231
timestamp 1698431365
transform 1 0 64512 0 -1 76832
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input232
timestamp 1698431365
transform 1 0 65184 0 -1 76832
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output233 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 13104 0 1 73696
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output234
timestamp 1698431365
transform 1 0 18032 0 1 73696
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output235
timestamp 1698431365
transform -1 0 20944 0 1 75264
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output236
timestamp 1698431365
transform 1 0 17472 0 -1 76832
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output237
timestamp 1698431365
transform -1 0 22960 0 -1 75264
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output238
timestamp 1698431365
transform -1 0 24080 0 1 75264
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output239
timestamp 1698431365
transform -1 0 24192 0 -1 76832
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output240
timestamp 1698431365
transform -1 0 14112 0 -1 73696
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output241
timestamp 1698431365
transform -1 0 13104 0 1 75264
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output242
timestamp 1698431365
transform -1 0 14112 0 -1 75264
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output243
timestamp 1698431365
transform -1 0 12768 0 -1 76832
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output244
timestamp 1698431365
transform -1 0 17024 0 -1 73696
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output245
timestamp 1698431365
transform -1 0 17024 0 -1 75264
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output246
timestamp 1698431365
transform -1 0 18032 0 1 73696
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output247
timestamp 1698431365
transform -1 0 16576 0 -1 76832
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output248
timestamp 1698431365
transform -1 0 18032 0 1 75264
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output249
timestamp 1698431365
transform 1 0 52752 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output250
timestamp 1698431365
transform 1 0 59696 0 -1 6272
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output251
timestamp 1698431365
transform 1 0 60368 0 1 6272
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output252
timestamp 1698431365
transform 1 0 63280 0 1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output253
timestamp 1698431365
transform 1 0 64288 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output254
timestamp 1698431365
transform 1 0 66304 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output255
timestamp 1698431365
transform 1 0 63280 0 1 6272
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output256
timestamp 1698431365
transform 1 0 64288 0 -1 6272
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output257
timestamp 1698431365
transform 1 0 67200 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output258
timestamp 1698431365
transform 1 0 70112 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output259
timestamp 1698431365
transform 1 0 67200 0 -1 6272
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output260
timestamp 1698431365
transform 1 0 54880 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output261
timestamp 1698431365
transform 1 0 68208 0 1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output262
timestamp 1698431365
transform 1 0 66864 0 -1 7840
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output263
timestamp 1698431365
transform 1 0 68208 0 1 6272
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output264
timestamp 1698431365
transform 1 0 71120 0 1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output265
timestamp 1698431365
transform 1 0 72128 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output266
timestamp 1698431365
transform 1 0 73920 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output267
timestamp 1698431365
transform 1 0 71120 0 1 6272
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output268
timestamp 1698431365
transform 1 0 72128 0 -1 6272
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output269
timestamp 1698431365
transform 1 0 75040 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output270
timestamp 1698431365
transform 1 0 72240 0 -1 7840
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output271
timestamp 1698431365
transform 1 0 54096 0 1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output272
timestamp 1698431365
transform 1 0 75040 0 -1 6272
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output273
timestamp 1698431365
transform 1 0 75152 0 -1 7840
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output274
timestamp 1698431365
transform 1 0 56448 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output275
timestamp 1698431365
transform -1 0 61600 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output276
timestamp 1698431365
transform 1 0 57008 0 1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output277
timestamp 1698431365
transform 1 0 56784 0 -1 6272
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output278
timestamp 1698431365
transform -1 0 62272 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output279
timestamp 1698431365
transform 1 0 62496 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output280
timestamp 1698431365
transform 1 0 60368 0 1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output281
timestamp 1698431365
transform 1 0 49392 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output282
timestamp 1698431365
transform 1 0 1568 0 -1 39200
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output283
timestamp 1698431365
transform -1 0 4480 0 1 39200
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output284
timestamp 1698431365
transform -1 0 4480 0 1 40768
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output285
timestamp 1698431365
transform -1 0 4480 0 -1 42336
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output286
timestamp 1698431365
transform -1 0 4480 0 1 42336
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output287
timestamp 1698431365
transform -1 0 4480 0 -1 54880
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output288
timestamp 1698431365
transform 1 0 1568 0 1 54880
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output289
timestamp 1698431365
transform -1 0 4480 0 1 56448
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output290
timestamp 1698431365
transform -1 0 4480 0 -1 58016
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output291
timestamp 1698431365
transform 1 0 1568 0 1 58016
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output292
timestamp 1698431365
transform -1 0 4480 0 1 59584
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output293
timestamp 1698431365
transform 1 0 1568 0 -1 61152
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output294
timestamp 1698431365
transform -1 0 4480 0 -1 62720
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output295
timestamp 1698431365
transform -1 0 4480 0 1 62720
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output296
timestamp 1698431365
transform -1 0 4480 0 1 64288
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output297
timestamp 1698431365
transform 1 0 1568 0 1 43904
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output298
timestamp 1698431365
transform -1 0 4480 0 -1 65856
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output299
timestamp 1698431365
transform 1 0 1568 0 1 65856
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output300
timestamp 1698431365
transform -1 0 4480 0 1 67424
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output301
timestamp 1698431365
transform 1 0 1568 0 -1 68992
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output302
timestamp 1698431365
transform -1 0 4480 0 -1 70560
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output303
timestamp 1698431365
transform -1 0 4480 0 1 70560
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output304
timestamp 1698431365
transform -1 0 4480 0 1 72128
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output305
timestamp 1698431365
transform -1 0 4480 0 -1 73696
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output306
timestamp 1698431365
transform -1 0 4480 0 1 73696
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output307
timestamp 1698431365
transform -1 0 4480 0 1 75264
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output308
timestamp 1698431365
transform 1 0 1568 0 -1 45472
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output309
timestamp 1698431365
transform -1 0 4480 0 -1 76832
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output310
timestamp 1698431365
transform -1 0 4480 0 -1 75264
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output311
timestamp 1698431365
transform -1 0 4480 0 -1 47040
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output312
timestamp 1698431365
transform 1 0 1568 0 1 47040
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output313
timestamp 1698431365
transform -1 0 4480 0 1 48608
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output314
timestamp 1698431365
transform -1 0 4480 0 -1 50176
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output315
timestamp 1698431365
transform -1 0 4480 0 1 50176
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output316
timestamp 1698431365
transform -1 0 4480 0 1 51744
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output317
timestamp 1698431365
transform -1 0 4480 0 -1 53312
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output318
timestamp 1698431365
transform 1 0 75488 0 -1 42336
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output319
timestamp 1698431365
transform -1 0 78400 0 -1 40768
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output320
timestamp 1698431365
transform -1 0 75824 0 1 7840
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output321
timestamp 1698431365
transform -1 0 78400 0 -1 10976
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output322
timestamp 1698431365
transform -1 0 75488 0 -1 9408
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output323
timestamp 1698431365
transform -1 0 78400 0 -1 9408
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output324
timestamp 1698431365
transform -1 0 35616 0 -1 76832
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output325
timestamp 1698431365
transform -1 0 58464 0 -1 76832
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output326
timestamp 1698431365
transform -1 0 59248 0 1 75264
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output327
timestamp 1698431365
transform 1 0 58688 0 -1 76832
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output328
timestamp 1698431365
transform -1 0 60592 0 -1 75264
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_94 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698431365
transform -1 0 78624 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_95
timestamp 1698431365
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698431365
transform -1 0 78624 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_96
timestamp 1698431365
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698431365
transform -1 0 78624 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_97
timestamp 1698431365
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698431365
transform -1 0 78624 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_98
timestamp 1698431365
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698431365
transform -1 0 78624 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_99
timestamp 1698431365
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698431365
transform -1 0 78624 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_100
timestamp 1698431365
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698431365
transform -1 0 78624 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_101
timestamp 1698431365
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698431365
transform -1 0 78624 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_102
timestamp 1698431365
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698431365
transform -1 0 78624 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_103
timestamp 1698431365
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698431365
transform -1 0 78624 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_104
timestamp 1698431365
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698431365
transform -1 0 78624 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_105
timestamp 1698431365
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698431365
transform -1 0 78624 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_106
timestamp 1698431365
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698431365
transform -1 0 78624 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_107
timestamp 1698431365
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698431365
transform -1 0 78624 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_108
timestamp 1698431365
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698431365
transform -1 0 78624 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_109
timestamp 1698431365
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698431365
transform -1 0 78624 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_110
timestamp 1698431365
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698431365
transform -1 0 78624 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_111
timestamp 1698431365
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698431365
transform -1 0 78624 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_112
timestamp 1698431365
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698431365
transform -1 0 78624 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_113
timestamp 1698431365
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698431365
transform -1 0 78624 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_114
timestamp 1698431365
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698431365
transform -1 0 78624 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_115
timestamp 1698431365
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698431365
transform -1 0 78624 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_116
timestamp 1698431365
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1698431365
transform -1 0 78624 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_117
timestamp 1698431365
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1698431365
transform -1 0 78624 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_118
timestamp 1698431365
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1698431365
transform -1 0 78624 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_119
timestamp 1698431365
transform 1 0 1344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1698431365
transform -1 0 78624 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_120
timestamp 1698431365
transform 1 0 1344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1698431365
transform -1 0 78624 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_121
timestamp 1698431365
transform 1 0 1344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1698431365
transform -1 0 78624 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_122
timestamp 1698431365
transform 1 0 1344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1698431365
transform -1 0 78624 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_123
timestamp 1698431365
transform 1 0 1344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1698431365
transform -1 0 78624 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Left_124
timestamp 1698431365
transform 1 0 1344 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1698431365
transform -1 0 78624 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Left_125
timestamp 1698431365
transform 1 0 1344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1698431365
transform -1 0 78624 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Left_126
timestamp 1698431365
transform 1 0 1344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1698431365
transform -1 0 78624 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Left_127
timestamp 1698431365
transform 1 0 1344 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1698431365
transform -1 0 78624 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Left_128
timestamp 1698431365
transform 1 0 1344 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1698431365
transform -1 0 78624 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Left_129
timestamp 1698431365
transform 1 0 1344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Right_35
timestamp 1698431365
transform -1 0 78624 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Left_130
timestamp 1698431365
transform 1 0 1344 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Right_36
timestamp 1698431365
transform -1 0 78624 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Left_131
timestamp 1698431365
transform 1 0 1344 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Right_37
timestamp 1698431365
transform -1 0 78624 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Left_132
timestamp 1698431365
transform 1 0 1344 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Right_38
timestamp 1698431365
transform -1 0 78624 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Left_133
timestamp 1698431365
transform 1 0 1344 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Right_39
timestamp 1698431365
transform -1 0 78624 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Left_134
timestamp 1698431365
transform 1 0 1344 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Right_40
timestamp 1698431365
transform -1 0 78624 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Left_135
timestamp 1698431365
transform 1 0 1344 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Right_41
timestamp 1698431365
transform -1 0 78624 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Left_136
timestamp 1698431365
transform 1 0 1344 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Right_42
timestamp 1698431365
transform -1 0 78624 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Left_137
timestamp 1698431365
transform 1 0 1344 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Right_43
timestamp 1698431365
transform -1 0 78624 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Left_138
timestamp 1698431365
transform 1 0 1344 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Right_44
timestamp 1698431365
transform -1 0 78624 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_45_Left_139
timestamp 1698431365
transform 1 0 1344 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_45_Right_45
timestamp 1698431365
transform -1 0 78624 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_46_Left_140
timestamp 1698431365
transform 1 0 1344 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_46_Right_46
timestamp 1698431365
transform -1 0 78624 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_47_Left_141
timestamp 1698431365
transform 1 0 1344 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_47_Right_47
timestamp 1698431365
transform -1 0 78624 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_48_Left_142
timestamp 1698431365
transform 1 0 1344 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_48_Right_48
timestamp 1698431365
transform -1 0 78624 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_49_Left_143
timestamp 1698431365
transform 1 0 1344 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_49_Right_49
timestamp 1698431365
transform -1 0 78624 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_50_Left_144
timestamp 1698431365
transform 1 0 1344 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_50_Right_50
timestamp 1698431365
transform -1 0 78624 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_51_Left_145
timestamp 1698431365
transform 1 0 1344 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_51_Right_51
timestamp 1698431365
transform -1 0 78624 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_52_Left_146
timestamp 1698431365
transform 1 0 1344 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_52_Right_52
timestamp 1698431365
transform -1 0 78624 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_53_Left_147
timestamp 1698431365
transform 1 0 1344 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_53_Right_53
timestamp 1698431365
transform -1 0 78624 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_54_Left_148
timestamp 1698431365
transform 1 0 1344 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_54_Right_54
timestamp 1698431365
transform -1 0 78624 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_55_Left_149
timestamp 1698431365
transform 1 0 1344 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_55_Right_55
timestamp 1698431365
transform -1 0 78624 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_56_Left_150
timestamp 1698431365
transform 1 0 1344 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_56_Right_56
timestamp 1698431365
transform -1 0 78624 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_57_Left_151
timestamp 1698431365
transform 1 0 1344 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_57_Right_57
timestamp 1698431365
transform -1 0 78624 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_58_Left_152
timestamp 1698431365
transform 1 0 1344 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_58_Right_58
timestamp 1698431365
transform -1 0 78624 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_59_Left_153
timestamp 1698431365
transform 1 0 1344 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_59_Right_59
timestamp 1698431365
transform -1 0 78624 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_60_Left_154
timestamp 1698431365
transform 1 0 1344 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_60_Right_60
timestamp 1698431365
transform -1 0 78624 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_61_Left_155
timestamp 1698431365
transform 1 0 1344 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_61_Right_61
timestamp 1698431365
transform -1 0 78624 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_62_Left_156
timestamp 1698431365
transform 1 0 1344 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_62_Right_62
timestamp 1698431365
transform -1 0 78624 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_63_Left_157
timestamp 1698431365
transform 1 0 1344 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_63_Right_63
timestamp 1698431365
transform -1 0 78624 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_64_Left_158
timestamp 1698431365
transform 1 0 1344 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_64_Right_64
timestamp 1698431365
transform -1 0 78624 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_65_Left_159
timestamp 1698431365
transform 1 0 1344 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_65_Right_65
timestamp 1698431365
transform -1 0 78624 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_66_Left_160
timestamp 1698431365
transform 1 0 1344 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_66_Right_66
timestamp 1698431365
transform -1 0 78624 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_67_Left_161
timestamp 1698431365
transform 1 0 1344 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_67_Right_67
timestamp 1698431365
transform -1 0 78624 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_68_Left_162
timestamp 1698431365
transform 1 0 1344 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_68_Right_68
timestamp 1698431365
transform -1 0 78624 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_69_Left_163
timestamp 1698431365
transform 1 0 1344 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_69_Right_69
timestamp 1698431365
transform -1 0 78624 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_70_Left_164
timestamp 1698431365
transform 1 0 1344 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_70_Right_70
timestamp 1698431365
transform -1 0 78624 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_71_Left_165
timestamp 1698431365
transform 1 0 1344 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_71_Right_71
timestamp 1698431365
transform -1 0 78624 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_72_Left_166
timestamp 1698431365
transform 1 0 1344 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_72_Right_72
timestamp 1698431365
transform -1 0 78624 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_73_Left_167
timestamp 1698431365
transform 1 0 1344 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_73_Right_73
timestamp 1698431365
transform -1 0 78624 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_74_Left_168
timestamp 1698431365
transform 1 0 1344 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_74_Right_74
timestamp 1698431365
transform -1 0 78624 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_75_Left_169
timestamp 1698431365
transform 1 0 1344 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_75_Right_75
timestamp 1698431365
transform -1 0 78624 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_76_Left_170
timestamp 1698431365
transform 1 0 1344 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_76_Right_76
timestamp 1698431365
transform -1 0 78624 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_77_Left_171
timestamp 1698431365
transform 1 0 1344 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_77_Right_77
timestamp 1698431365
transform -1 0 78624 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_78_Left_172
timestamp 1698431365
transform 1 0 1344 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_78_Right_78
timestamp 1698431365
transform -1 0 78624 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_79_Left_173
timestamp 1698431365
transform 1 0 1344 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_79_Right_79
timestamp 1698431365
transform -1 0 78624 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_80_Left_174
timestamp 1698431365
transform 1 0 1344 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_80_Right_80
timestamp 1698431365
transform -1 0 78624 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_81_Left_175
timestamp 1698431365
transform 1 0 1344 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_81_Right_81
timestamp 1698431365
transform -1 0 78624 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_82_Left_176
timestamp 1698431365
transform 1 0 1344 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_82_Right_82
timestamp 1698431365
transform -1 0 78624 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_83_Left_177
timestamp 1698431365
transform 1 0 1344 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_83_Right_83
timestamp 1698431365
transform -1 0 78624 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_84_Left_178
timestamp 1698431365
transform 1 0 1344 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_84_Right_84
timestamp 1698431365
transform -1 0 78624 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_85_Left_179
timestamp 1698431365
transform 1 0 1344 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_85_Right_85
timestamp 1698431365
transform -1 0 78624 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_86_Left_180
timestamp 1698431365
transform 1 0 1344 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_86_Right_86
timestamp 1698431365
transform -1 0 78624 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_87_Left_181
timestamp 1698431365
transform 1 0 1344 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_87_Right_87
timestamp 1698431365
transform -1 0 78624 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_88_Left_182
timestamp 1698431365
transform 1 0 1344 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_88_Right_88
timestamp 1698431365
transform -1 0 78624 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_89_Left_183
timestamp 1698431365
transform 1 0 1344 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_89_Right_89
timestamp 1698431365
transform -1 0 78624 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_90_Left_184
timestamp 1698431365
transform 1 0 1344 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_90_Right_90
timestamp 1698431365
transform -1 0 78624 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_91_Left_185
timestamp 1698431365
transform 1 0 1344 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_91_Right_91
timestamp 1698431365
transform -1 0 78624 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_92_Left_186
timestamp 1698431365
transform 1 0 1344 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_92_Right_92
timestamp 1698431365
transform -1 0 78624 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_93_Left_187
timestamp 1698431365
transform 1 0 1344 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_93_Right_93
timestamp 1698431365
transform -1 0 78624 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  simple_interconnect_343 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 20832 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  simple_interconnect_344
timestamp 1698431365
transform -1 0 23408 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  simple_interconnect_345
timestamp 1698431365
transform -1 0 23856 0 -1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  simple_interconnect_346
timestamp 1698431365
transform -1 0 24528 0 1 75264
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  simple_interconnect_347
timestamp 1698431365
transform -1 0 25200 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  simple_interconnect_348
timestamp 1698431365
transform -1 0 25872 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  simple_interconnect_349
timestamp 1698431365
transform -1 0 26544 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  simple_interconnect_350
timestamp 1698431365
transform -1 0 27216 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  simple_interconnect_351
timestamp 1698431365
transform -1 0 27888 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  simple_interconnect_352
timestamp 1698431365
transform -1 0 28672 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  simple_interconnect_353
timestamp 1698431365
transform -1 0 29232 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  simple_interconnect_354
timestamp 1698431365
transform -1 0 29904 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  simple_interconnect_355
timestamp 1698431365
transform -1 0 30576 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  simple_interconnect_356
timestamp 1698431365
transform -1 0 31248 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  simple_interconnect_357
timestamp 1698431365
transform -1 0 31808 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  simple_interconnect_358
timestamp 1698431365
transform -1 0 32592 0 -1 76832
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_188 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5152 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_189
timestamp 1698431365
transform 1 0 8960 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_190
timestamp 1698431365
transform 1 0 12768 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_191
timestamp 1698431365
transform 1 0 16576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_192
timestamp 1698431365
transform 1 0 20384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_193
timestamp 1698431365
transform 1 0 24192 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_194
timestamp 1698431365
transform 1 0 28000 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_195
timestamp 1698431365
transform 1 0 31808 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_196
timestamp 1698431365
transform 1 0 35616 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_197
timestamp 1698431365
transform 1 0 39424 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_198
timestamp 1698431365
transform 1 0 43232 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_199
timestamp 1698431365
transform 1 0 47040 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_200
timestamp 1698431365
transform 1 0 50848 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_201
timestamp 1698431365
transform 1 0 54656 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_202
timestamp 1698431365
transform 1 0 58464 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_203
timestamp 1698431365
transform 1 0 62272 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_204
timestamp 1698431365
transform 1 0 66080 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_205
timestamp 1698431365
transform 1 0 69888 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_206
timestamp 1698431365
transform 1 0 73696 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_207
timestamp 1698431365
transform 1 0 77504 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_208
timestamp 1698431365
transform 1 0 9184 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_209
timestamp 1698431365
transform 1 0 17024 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_210
timestamp 1698431365
transform 1 0 24864 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_211
timestamp 1698431365
transform 1 0 32704 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_212
timestamp 1698431365
transform 1 0 40544 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_213
timestamp 1698431365
transform 1 0 48384 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_214
timestamp 1698431365
transform 1 0 56224 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_215
timestamp 1698431365
transform 1 0 64064 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_216
timestamp 1698431365
transform 1 0 71904 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_217
timestamp 1698431365
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_218
timestamp 1698431365
transform 1 0 13104 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_219
timestamp 1698431365
transform 1 0 20944 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_220
timestamp 1698431365
transform 1 0 28784 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_221
timestamp 1698431365
transform 1 0 36624 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_222
timestamp 1698431365
transform 1 0 44464 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_223
timestamp 1698431365
transform 1 0 52304 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_224
timestamp 1698431365
transform 1 0 60144 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_225
timestamp 1698431365
transform 1 0 67984 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_226
timestamp 1698431365
transform 1 0 75824 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_227
timestamp 1698431365
transform 1 0 9184 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_228
timestamp 1698431365
transform 1 0 17024 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_229
timestamp 1698431365
transform 1 0 24864 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_230
timestamp 1698431365
transform 1 0 32704 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_231
timestamp 1698431365
transform 1 0 40544 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_232
timestamp 1698431365
transform 1 0 48384 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_233
timestamp 1698431365
transform 1 0 56224 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_234
timestamp 1698431365
transform 1 0 64064 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_235
timestamp 1698431365
transform 1 0 71904 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_236
timestamp 1698431365
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_237
timestamp 1698431365
transform 1 0 13104 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_238
timestamp 1698431365
transform 1 0 20944 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_239
timestamp 1698431365
transform 1 0 28784 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_240
timestamp 1698431365
transform 1 0 36624 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_241
timestamp 1698431365
transform 1 0 44464 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_242
timestamp 1698431365
transform 1 0 52304 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_243
timestamp 1698431365
transform 1 0 60144 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_244
timestamp 1698431365
transform 1 0 67984 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_245
timestamp 1698431365
transform 1 0 75824 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_246
timestamp 1698431365
transform 1 0 9184 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_247
timestamp 1698431365
transform 1 0 17024 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_248
timestamp 1698431365
transform 1 0 24864 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_249
timestamp 1698431365
transform 1 0 32704 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_250
timestamp 1698431365
transform 1 0 40544 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_251
timestamp 1698431365
transform 1 0 48384 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_252
timestamp 1698431365
transform 1 0 56224 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_253
timestamp 1698431365
transform 1 0 64064 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_254
timestamp 1698431365
transform 1 0 71904 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_255
timestamp 1698431365
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_256
timestamp 1698431365
transform 1 0 13104 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_257
timestamp 1698431365
transform 1 0 20944 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_258
timestamp 1698431365
transform 1 0 28784 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_259
timestamp 1698431365
transform 1 0 36624 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_260
timestamp 1698431365
transform 1 0 44464 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_261
timestamp 1698431365
transform 1 0 52304 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_262
timestamp 1698431365
transform 1 0 60144 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_263
timestamp 1698431365
transform 1 0 67984 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_264
timestamp 1698431365
transform 1 0 75824 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_265
timestamp 1698431365
transform 1 0 9184 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_266
timestamp 1698431365
transform 1 0 17024 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_267
timestamp 1698431365
transform 1 0 24864 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_268
timestamp 1698431365
transform 1 0 32704 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_269
timestamp 1698431365
transform 1 0 40544 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_270
timestamp 1698431365
transform 1 0 48384 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_271
timestamp 1698431365
transform 1 0 56224 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_272
timestamp 1698431365
transform 1 0 64064 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_273
timestamp 1698431365
transform 1 0 71904 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_274
timestamp 1698431365
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_275
timestamp 1698431365
transform 1 0 13104 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_276
timestamp 1698431365
transform 1 0 20944 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_277
timestamp 1698431365
transform 1 0 28784 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_278
timestamp 1698431365
transform 1 0 36624 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_279
timestamp 1698431365
transform 1 0 44464 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_280
timestamp 1698431365
transform 1 0 52304 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_281
timestamp 1698431365
transform 1 0 60144 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_282
timestamp 1698431365
transform 1 0 67984 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_283
timestamp 1698431365
transform 1 0 75824 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_284
timestamp 1698431365
transform 1 0 9184 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_285
timestamp 1698431365
transform 1 0 17024 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_286
timestamp 1698431365
transform 1 0 24864 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_287
timestamp 1698431365
transform 1 0 32704 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_288
timestamp 1698431365
transform 1 0 40544 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_289
timestamp 1698431365
transform 1 0 48384 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_290
timestamp 1698431365
transform 1 0 56224 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_291
timestamp 1698431365
transform 1 0 64064 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_292
timestamp 1698431365
transform 1 0 71904 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_293
timestamp 1698431365
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_294
timestamp 1698431365
transform 1 0 13104 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_295
timestamp 1698431365
transform 1 0 20944 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_296
timestamp 1698431365
transform 1 0 28784 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_297
timestamp 1698431365
transform 1 0 36624 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_298
timestamp 1698431365
transform 1 0 44464 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_299
timestamp 1698431365
transform 1 0 52304 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_300
timestamp 1698431365
transform 1 0 60144 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_301
timestamp 1698431365
transform 1 0 67984 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_302
timestamp 1698431365
transform 1 0 75824 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_303
timestamp 1698431365
transform 1 0 9184 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_304
timestamp 1698431365
transform 1 0 17024 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_305
timestamp 1698431365
transform 1 0 24864 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_306
timestamp 1698431365
transform 1 0 32704 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_307
timestamp 1698431365
transform 1 0 40544 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_308
timestamp 1698431365
transform 1 0 48384 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_309
timestamp 1698431365
transform 1 0 56224 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_310
timestamp 1698431365
transform 1 0 64064 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_311
timestamp 1698431365
transform 1 0 71904 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_312
timestamp 1698431365
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_313
timestamp 1698431365
transform 1 0 13104 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_314
timestamp 1698431365
transform 1 0 20944 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_315
timestamp 1698431365
transform 1 0 28784 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_316
timestamp 1698431365
transform 1 0 36624 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_317
timestamp 1698431365
transform 1 0 44464 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_318
timestamp 1698431365
transform 1 0 52304 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_319
timestamp 1698431365
transform 1 0 60144 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_320
timestamp 1698431365
transform 1 0 67984 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_321
timestamp 1698431365
transform 1 0 75824 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_322
timestamp 1698431365
transform 1 0 9184 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_323
timestamp 1698431365
transform 1 0 17024 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_324
timestamp 1698431365
transform 1 0 24864 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_325
timestamp 1698431365
transform 1 0 32704 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_326
timestamp 1698431365
transform 1 0 40544 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_327
timestamp 1698431365
transform 1 0 48384 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_328
timestamp 1698431365
transform 1 0 56224 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_329
timestamp 1698431365
transform 1 0 64064 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_330
timestamp 1698431365
transform 1 0 71904 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_331
timestamp 1698431365
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_332
timestamp 1698431365
transform 1 0 13104 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_333
timestamp 1698431365
transform 1 0 20944 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_334
timestamp 1698431365
transform 1 0 28784 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_335
timestamp 1698431365
transform 1 0 36624 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_336
timestamp 1698431365
transform 1 0 44464 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_337
timestamp 1698431365
transform 1 0 52304 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_338
timestamp 1698431365
transform 1 0 60144 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_339
timestamp 1698431365
transform 1 0 67984 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_340
timestamp 1698431365
transform 1 0 75824 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_341
timestamp 1698431365
transform 1 0 9184 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_342
timestamp 1698431365
transform 1 0 17024 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_343
timestamp 1698431365
transform 1 0 24864 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_344
timestamp 1698431365
transform 1 0 32704 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_345
timestamp 1698431365
transform 1 0 40544 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_346
timestamp 1698431365
transform 1 0 48384 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_347
timestamp 1698431365
transform 1 0 56224 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_348
timestamp 1698431365
transform 1 0 64064 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_349
timestamp 1698431365
transform 1 0 71904 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_350
timestamp 1698431365
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_351
timestamp 1698431365
transform 1 0 13104 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_352
timestamp 1698431365
transform 1 0 20944 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_353
timestamp 1698431365
transform 1 0 28784 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_354
timestamp 1698431365
transform 1 0 36624 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_355
timestamp 1698431365
transform 1 0 44464 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_356
timestamp 1698431365
transform 1 0 52304 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_357
timestamp 1698431365
transform 1 0 60144 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_358
timestamp 1698431365
transform 1 0 67984 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_359
timestamp 1698431365
transform 1 0 75824 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_360
timestamp 1698431365
transform 1 0 9184 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_361
timestamp 1698431365
transform 1 0 17024 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_362
timestamp 1698431365
transform 1 0 24864 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_363
timestamp 1698431365
transform 1 0 32704 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_364
timestamp 1698431365
transform 1 0 40544 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_365
timestamp 1698431365
transform 1 0 48384 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_366
timestamp 1698431365
transform 1 0 56224 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_367
timestamp 1698431365
transform 1 0 64064 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_368
timestamp 1698431365
transform 1 0 71904 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_369
timestamp 1698431365
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_370
timestamp 1698431365
transform 1 0 13104 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_371
timestamp 1698431365
transform 1 0 20944 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_372
timestamp 1698431365
transform 1 0 28784 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_373
timestamp 1698431365
transform 1 0 36624 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_374
timestamp 1698431365
transform 1 0 44464 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_375
timestamp 1698431365
transform 1 0 52304 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_376
timestamp 1698431365
transform 1 0 60144 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_377
timestamp 1698431365
transform 1 0 67984 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_378
timestamp 1698431365
transform 1 0 75824 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_379
timestamp 1698431365
transform 1 0 9184 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_380
timestamp 1698431365
transform 1 0 17024 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_381
timestamp 1698431365
transform 1 0 24864 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_382
timestamp 1698431365
transform 1 0 32704 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_383
timestamp 1698431365
transform 1 0 40544 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_384
timestamp 1698431365
transform 1 0 48384 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_385
timestamp 1698431365
transform 1 0 56224 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_386
timestamp 1698431365
transform 1 0 64064 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_387
timestamp 1698431365
transform 1 0 71904 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_388
timestamp 1698431365
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_389
timestamp 1698431365
transform 1 0 13104 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_390
timestamp 1698431365
transform 1 0 20944 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_391
timestamp 1698431365
transform 1 0 28784 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_392
timestamp 1698431365
transform 1 0 36624 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_393
timestamp 1698431365
transform 1 0 44464 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_394
timestamp 1698431365
transform 1 0 52304 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_395
timestamp 1698431365
transform 1 0 60144 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_396
timestamp 1698431365
transform 1 0 67984 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_397
timestamp 1698431365
transform 1 0 75824 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_398
timestamp 1698431365
transform 1 0 9184 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_399
timestamp 1698431365
transform 1 0 17024 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_400
timestamp 1698431365
transform 1 0 24864 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_401
timestamp 1698431365
transform 1 0 32704 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_402
timestamp 1698431365
transform 1 0 40544 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_403
timestamp 1698431365
transform 1 0 48384 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_404
timestamp 1698431365
transform 1 0 56224 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_405
timestamp 1698431365
transform 1 0 64064 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_406
timestamp 1698431365
transform 1 0 71904 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_407
timestamp 1698431365
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_408
timestamp 1698431365
transform 1 0 13104 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_409
timestamp 1698431365
transform 1 0 20944 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_410
timestamp 1698431365
transform 1 0 28784 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_411
timestamp 1698431365
transform 1 0 36624 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_412
timestamp 1698431365
transform 1 0 44464 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_413
timestamp 1698431365
transform 1 0 52304 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_414
timestamp 1698431365
transform 1 0 60144 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_415
timestamp 1698431365
transform 1 0 67984 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_416
timestamp 1698431365
transform 1 0 75824 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_417
timestamp 1698431365
transform 1 0 9184 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_418
timestamp 1698431365
transform 1 0 17024 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_419
timestamp 1698431365
transform 1 0 24864 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_420
timestamp 1698431365
transform 1 0 32704 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_421
timestamp 1698431365
transform 1 0 40544 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_422
timestamp 1698431365
transform 1 0 48384 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_423
timestamp 1698431365
transform 1 0 56224 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_424
timestamp 1698431365
transform 1 0 64064 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_425
timestamp 1698431365
transform 1 0 71904 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_426
timestamp 1698431365
transform 1 0 5264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_427
timestamp 1698431365
transform 1 0 13104 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_428
timestamp 1698431365
transform 1 0 20944 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_429
timestamp 1698431365
transform 1 0 28784 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_430
timestamp 1698431365
transform 1 0 36624 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_431
timestamp 1698431365
transform 1 0 44464 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_432
timestamp 1698431365
transform 1 0 52304 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_433
timestamp 1698431365
transform 1 0 60144 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_434
timestamp 1698431365
transform 1 0 67984 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_435
timestamp 1698431365
transform 1 0 75824 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_436
timestamp 1698431365
transform 1 0 9184 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_437
timestamp 1698431365
transform 1 0 17024 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_438
timestamp 1698431365
transform 1 0 24864 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_439
timestamp 1698431365
transform 1 0 32704 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_440
timestamp 1698431365
transform 1 0 40544 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_441
timestamp 1698431365
transform 1 0 48384 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_442
timestamp 1698431365
transform 1 0 56224 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_443
timestamp 1698431365
transform 1 0 64064 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_444
timestamp 1698431365
transform 1 0 71904 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_445
timestamp 1698431365
transform 1 0 5264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_446
timestamp 1698431365
transform 1 0 13104 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_447
timestamp 1698431365
transform 1 0 20944 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_448
timestamp 1698431365
transform 1 0 28784 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_449
timestamp 1698431365
transform 1 0 36624 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_450
timestamp 1698431365
transform 1 0 44464 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_451
timestamp 1698431365
transform 1 0 52304 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_452
timestamp 1698431365
transform 1 0 60144 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_453
timestamp 1698431365
transform 1 0 67984 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_454
timestamp 1698431365
transform 1 0 75824 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_455
timestamp 1698431365
transform 1 0 9184 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_456
timestamp 1698431365
transform 1 0 17024 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_457
timestamp 1698431365
transform 1 0 24864 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_458
timestamp 1698431365
transform 1 0 32704 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_459
timestamp 1698431365
transform 1 0 40544 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_460
timestamp 1698431365
transform 1 0 48384 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_461
timestamp 1698431365
transform 1 0 56224 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_462
timestamp 1698431365
transform 1 0 64064 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_463
timestamp 1698431365
transform 1 0 71904 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_464
timestamp 1698431365
transform 1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_465
timestamp 1698431365
transform 1 0 13104 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_466
timestamp 1698431365
transform 1 0 20944 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_467
timestamp 1698431365
transform 1 0 28784 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_468
timestamp 1698431365
transform 1 0 36624 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_469
timestamp 1698431365
transform 1 0 44464 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_470
timestamp 1698431365
transform 1 0 52304 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_471
timestamp 1698431365
transform 1 0 60144 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_472
timestamp 1698431365
transform 1 0 67984 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_473
timestamp 1698431365
transform 1 0 75824 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_474
timestamp 1698431365
transform 1 0 9184 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_475
timestamp 1698431365
transform 1 0 17024 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_476
timestamp 1698431365
transform 1 0 24864 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_477
timestamp 1698431365
transform 1 0 32704 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_478
timestamp 1698431365
transform 1 0 40544 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_479
timestamp 1698431365
transform 1 0 48384 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_480
timestamp 1698431365
transform 1 0 56224 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_481
timestamp 1698431365
transform 1 0 64064 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_482
timestamp 1698431365
transform 1 0 71904 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_483
timestamp 1698431365
transform 1 0 5264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_484
timestamp 1698431365
transform 1 0 13104 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_485
timestamp 1698431365
transform 1 0 20944 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_486
timestamp 1698431365
transform 1 0 28784 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_487
timestamp 1698431365
transform 1 0 36624 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_488
timestamp 1698431365
transform 1 0 44464 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_489
timestamp 1698431365
transform 1 0 52304 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_490
timestamp 1698431365
transform 1 0 60144 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_491
timestamp 1698431365
transform 1 0 67984 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_492
timestamp 1698431365
transform 1 0 75824 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_493
timestamp 1698431365
transform 1 0 9184 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_494
timestamp 1698431365
transform 1 0 17024 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_495
timestamp 1698431365
transform 1 0 24864 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_496
timestamp 1698431365
transform 1 0 32704 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_497
timestamp 1698431365
transform 1 0 40544 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_498
timestamp 1698431365
transform 1 0 48384 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_499
timestamp 1698431365
transform 1 0 56224 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_500
timestamp 1698431365
transform 1 0 64064 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_501
timestamp 1698431365
transform 1 0 71904 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_502
timestamp 1698431365
transform 1 0 5264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_503
timestamp 1698431365
transform 1 0 13104 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_504
timestamp 1698431365
transform 1 0 20944 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_505
timestamp 1698431365
transform 1 0 28784 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_506
timestamp 1698431365
transform 1 0 36624 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_507
timestamp 1698431365
transform 1 0 44464 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_508
timestamp 1698431365
transform 1 0 52304 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_509
timestamp 1698431365
transform 1 0 60144 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_510
timestamp 1698431365
transform 1 0 67984 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_511
timestamp 1698431365
transform 1 0 75824 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_512
timestamp 1698431365
transform 1 0 9184 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_513
timestamp 1698431365
transform 1 0 17024 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_514
timestamp 1698431365
transform 1 0 24864 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_515
timestamp 1698431365
transform 1 0 32704 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_516
timestamp 1698431365
transform 1 0 40544 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_517
timestamp 1698431365
transform 1 0 48384 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_518
timestamp 1698431365
transform 1 0 56224 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_519
timestamp 1698431365
transform 1 0 64064 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_520
timestamp 1698431365
transform 1 0 71904 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_521
timestamp 1698431365
transform 1 0 5264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_522
timestamp 1698431365
transform 1 0 13104 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_523
timestamp 1698431365
transform 1 0 20944 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_524
timestamp 1698431365
transform 1 0 28784 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_525
timestamp 1698431365
transform 1 0 36624 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_526
timestamp 1698431365
transform 1 0 44464 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_527
timestamp 1698431365
transform 1 0 52304 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_528
timestamp 1698431365
transform 1 0 60144 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_529
timestamp 1698431365
transform 1 0 67984 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_530
timestamp 1698431365
transform 1 0 75824 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_531
timestamp 1698431365
transform 1 0 9184 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_532
timestamp 1698431365
transform 1 0 17024 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_533
timestamp 1698431365
transform 1 0 24864 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_534
timestamp 1698431365
transform 1 0 32704 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_535
timestamp 1698431365
transform 1 0 40544 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_536
timestamp 1698431365
transform 1 0 48384 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_537
timestamp 1698431365
transform 1 0 56224 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_538
timestamp 1698431365
transform 1 0 64064 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_539
timestamp 1698431365
transform 1 0 71904 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_540
timestamp 1698431365
transform 1 0 5264 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_541
timestamp 1698431365
transform 1 0 13104 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_542
timestamp 1698431365
transform 1 0 20944 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_543
timestamp 1698431365
transform 1 0 28784 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_544
timestamp 1698431365
transform 1 0 36624 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_545
timestamp 1698431365
transform 1 0 44464 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_546
timestamp 1698431365
transform 1 0 52304 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_547
timestamp 1698431365
transform 1 0 60144 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_548
timestamp 1698431365
transform 1 0 67984 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_549
timestamp 1698431365
transform 1 0 75824 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_550
timestamp 1698431365
transform 1 0 9184 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_551
timestamp 1698431365
transform 1 0 17024 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_552
timestamp 1698431365
transform 1 0 24864 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_553
timestamp 1698431365
transform 1 0 32704 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_554
timestamp 1698431365
transform 1 0 40544 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_555
timestamp 1698431365
transform 1 0 48384 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_556
timestamp 1698431365
transform 1 0 56224 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_557
timestamp 1698431365
transform 1 0 64064 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_558
timestamp 1698431365
transform 1 0 71904 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_559
timestamp 1698431365
transform 1 0 5264 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_560
timestamp 1698431365
transform 1 0 13104 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_561
timestamp 1698431365
transform 1 0 20944 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_562
timestamp 1698431365
transform 1 0 28784 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_563
timestamp 1698431365
transform 1 0 36624 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_564
timestamp 1698431365
transform 1 0 44464 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_565
timestamp 1698431365
transform 1 0 52304 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_566
timestamp 1698431365
transform 1 0 60144 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_567
timestamp 1698431365
transform 1 0 67984 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_568
timestamp 1698431365
transform 1 0 75824 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_569
timestamp 1698431365
transform 1 0 9184 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_570
timestamp 1698431365
transform 1 0 17024 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_571
timestamp 1698431365
transform 1 0 24864 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_572
timestamp 1698431365
transform 1 0 32704 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_573
timestamp 1698431365
transform 1 0 40544 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_574
timestamp 1698431365
transform 1 0 48384 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_575
timestamp 1698431365
transform 1 0 56224 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_576
timestamp 1698431365
transform 1 0 64064 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_577
timestamp 1698431365
transform 1 0 71904 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_578
timestamp 1698431365
transform 1 0 5264 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_579
timestamp 1698431365
transform 1 0 13104 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_580
timestamp 1698431365
transform 1 0 20944 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_581
timestamp 1698431365
transform 1 0 28784 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_582
timestamp 1698431365
transform 1 0 36624 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_583
timestamp 1698431365
transform 1 0 44464 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_584
timestamp 1698431365
transform 1 0 52304 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_585
timestamp 1698431365
transform 1 0 60144 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_586
timestamp 1698431365
transform 1 0 67984 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_587
timestamp 1698431365
transform 1 0 75824 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_588
timestamp 1698431365
transform 1 0 9184 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_589
timestamp 1698431365
transform 1 0 17024 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_590
timestamp 1698431365
transform 1 0 24864 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_591
timestamp 1698431365
transform 1 0 32704 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_592
timestamp 1698431365
transform 1 0 40544 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_593
timestamp 1698431365
transform 1 0 48384 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_594
timestamp 1698431365
transform 1 0 56224 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_595
timestamp 1698431365
transform 1 0 64064 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_596
timestamp 1698431365
transform 1 0 71904 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_597
timestamp 1698431365
transform 1 0 5264 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_598
timestamp 1698431365
transform 1 0 13104 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_599
timestamp 1698431365
transform 1 0 20944 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_600
timestamp 1698431365
transform 1 0 28784 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_601
timestamp 1698431365
transform 1 0 36624 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_602
timestamp 1698431365
transform 1 0 44464 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_603
timestamp 1698431365
transform 1 0 52304 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_604
timestamp 1698431365
transform 1 0 60144 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_605
timestamp 1698431365
transform 1 0 67984 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_606
timestamp 1698431365
transform 1 0 75824 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_607
timestamp 1698431365
transform 1 0 9184 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_608
timestamp 1698431365
transform 1 0 17024 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_609
timestamp 1698431365
transform 1 0 24864 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_610
timestamp 1698431365
transform 1 0 32704 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_611
timestamp 1698431365
transform 1 0 40544 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_612
timestamp 1698431365
transform 1 0 48384 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_613
timestamp 1698431365
transform 1 0 56224 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_614
timestamp 1698431365
transform 1 0 64064 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_615
timestamp 1698431365
transform 1 0 71904 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_616
timestamp 1698431365
transform 1 0 5264 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_617
timestamp 1698431365
transform 1 0 13104 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_618
timestamp 1698431365
transform 1 0 20944 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_619
timestamp 1698431365
transform 1 0 28784 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_620
timestamp 1698431365
transform 1 0 36624 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_621
timestamp 1698431365
transform 1 0 44464 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_622
timestamp 1698431365
transform 1 0 52304 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_623
timestamp 1698431365
transform 1 0 60144 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_624
timestamp 1698431365
transform 1 0 67984 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_625
timestamp 1698431365
transform 1 0 75824 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_626
timestamp 1698431365
transform 1 0 9184 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_627
timestamp 1698431365
transform 1 0 17024 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_628
timestamp 1698431365
transform 1 0 24864 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_629
timestamp 1698431365
transform 1 0 32704 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_630
timestamp 1698431365
transform 1 0 40544 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_631
timestamp 1698431365
transform 1 0 48384 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_632
timestamp 1698431365
transform 1 0 56224 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_633
timestamp 1698431365
transform 1 0 64064 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_634
timestamp 1698431365
transform 1 0 71904 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_635
timestamp 1698431365
transform 1 0 5264 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_636
timestamp 1698431365
transform 1 0 13104 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_637
timestamp 1698431365
transform 1 0 20944 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_638
timestamp 1698431365
transform 1 0 28784 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_639
timestamp 1698431365
transform 1 0 36624 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_640
timestamp 1698431365
transform 1 0 44464 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_641
timestamp 1698431365
transform 1 0 52304 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_642
timestamp 1698431365
transform 1 0 60144 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_643
timestamp 1698431365
transform 1 0 67984 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_644
timestamp 1698431365
transform 1 0 75824 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_645
timestamp 1698431365
transform 1 0 9184 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_646
timestamp 1698431365
transform 1 0 17024 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_647
timestamp 1698431365
transform 1 0 24864 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_648
timestamp 1698431365
transform 1 0 32704 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_649
timestamp 1698431365
transform 1 0 40544 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_650
timestamp 1698431365
transform 1 0 48384 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_651
timestamp 1698431365
transform 1 0 56224 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_652
timestamp 1698431365
transform 1 0 64064 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_653
timestamp 1698431365
transform 1 0 71904 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_654
timestamp 1698431365
transform 1 0 5264 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_655
timestamp 1698431365
transform 1 0 13104 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_656
timestamp 1698431365
transform 1 0 20944 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_657
timestamp 1698431365
transform 1 0 28784 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_658
timestamp 1698431365
transform 1 0 36624 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_659
timestamp 1698431365
transform 1 0 44464 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_660
timestamp 1698431365
transform 1 0 52304 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_661
timestamp 1698431365
transform 1 0 60144 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_662
timestamp 1698431365
transform 1 0 67984 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_663
timestamp 1698431365
transform 1 0 75824 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_664
timestamp 1698431365
transform 1 0 9184 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_665
timestamp 1698431365
transform 1 0 17024 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_666
timestamp 1698431365
transform 1 0 24864 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_667
timestamp 1698431365
transform 1 0 32704 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_668
timestamp 1698431365
transform 1 0 40544 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_669
timestamp 1698431365
transform 1 0 48384 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_670
timestamp 1698431365
transform 1 0 56224 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_671
timestamp 1698431365
transform 1 0 64064 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_672
timestamp 1698431365
transform 1 0 71904 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_673
timestamp 1698431365
transform 1 0 5264 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_674
timestamp 1698431365
transform 1 0 13104 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_675
timestamp 1698431365
transform 1 0 20944 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_676
timestamp 1698431365
transform 1 0 28784 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_677
timestamp 1698431365
transform 1 0 36624 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_678
timestamp 1698431365
transform 1 0 44464 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_679
timestamp 1698431365
transform 1 0 52304 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_680
timestamp 1698431365
transform 1 0 60144 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_681
timestamp 1698431365
transform 1 0 67984 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_682
timestamp 1698431365
transform 1 0 75824 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_683
timestamp 1698431365
transform 1 0 9184 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_684
timestamp 1698431365
transform 1 0 17024 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_685
timestamp 1698431365
transform 1 0 24864 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_686
timestamp 1698431365
transform 1 0 32704 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_687
timestamp 1698431365
transform 1 0 40544 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_688
timestamp 1698431365
transform 1 0 48384 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_689
timestamp 1698431365
transform 1 0 56224 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_690
timestamp 1698431365
transform 1 0 64064 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_691
timestamp 1698431365
transform 1 0 71904 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_692
timestamp 1698431365
transform 1 0 5264 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_693
timestamp 1698431365
transform 1 0 13104 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_694
timestamp 1698431365
transform 1 0 20944 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_695
timestamp 1698431365
transform 1 0 28784 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_696
timestamp 1698431365
transform 1 0 36624 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_697
timestamp 1698431365
transform 1 0 44464 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_698
timestamp 1698431365
transform 1 0 52304 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_699
timestamp 1698431365
transform 1 0 60144 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_700
timestamp 1698431365
transform 1 0 67984 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_701
timestamp 1698431365
transform 1 0 75824 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_702
timestamp 1698431365
transform 1 0 9184 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_703
timestamp 1698431365
transform 1 0 17024 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_704
timestamp 1698431365
transform 1 0 24864 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_705
timestamp 1698431365
transform 1 0 32704 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_706
timestamp 1698431365
transform 1 0 40544 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_707
timestamp 1698431365
transform 1 0 48384 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_708
timestamp 1698431365
transform 1 0 56224 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_709
timestamp 1698431365
transform 1 0 64064 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_710
timestamp 1698431365
transform 1 0 71904 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_711
timestamp 1698431365
transform 1 0 5264 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_712
timestamp 1698431365
transform 1 0 13104 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_713
timestamp 1698431365
transform 1 0 20944 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_714
timestamp 1698431365
transform 1 0 28784 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_715
timestamp 1698431365
transform 1 0 36624 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_716
timestamp 1698431365
transform 1 0 44464 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_717
timestamp 1698431365
transform 1 0 52304 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_718
timestamp 1698431365
transform 1 0 60144 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_719
timestamp 1698431365
transform 1 0 67984 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_720
timestamp 1698431365
transform 1 0 75824 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_721
timestamp 1698431365
transform 1 0 9184 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_722
timestamp 1698431365
transform 1 0 17024 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_723
timestamp 1698431365
transform 1 0 24864 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_724
timestamp 1698431365
transform 1 0 32704 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_725
timestamp 1698431365
transform 1 0 40544 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_726
timestamp 1698431365
transform 1 0 48384 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_727
timestamp 1698431365
transform 1 0 56224 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_728
timestamp 1698431365
transform 1 0 64064 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_729
timestamp 1698431365
transform 1 0 71904 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_730
timestamp 1698431365
transform 1 0 5264 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_731
timestamp 1698431365
transform 1 0 13104 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_732
timestamp 1698431365
transform 1 0 20944 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_733
timestamp 1698431365
transform 1 0 28784 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_734
timestamp 1698431365
transform 1 0 36624 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_735
timestamp 1698431365
transform 1 0 44464 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_736
timestamp 1698431365
transform 1 0 52304 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_737
timestamp 1698431365
transform 1 0 60144 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_738
timestamp 1698431365
transform 1 0 67984 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_739
timestamp 1698431365
transform 1 0 75824 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_740
timestamp 1698431365
transform 1 0 9184 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_741
timestamp 1698431365
transform 1 0 17024 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_742
timestamp 1698431365
transform 1 0 24864 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_743
timestamp 1698431365
transform 1 0 32704 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_744
timestamp 1698431365
transform 1 0 40544 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_745
timestamp 1698431365
transform 1 0 48384 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_746
timestamp 1698431365
transform 1 0 56224 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_747
timestamp 1698431365
transform 1 0 64064 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_748
timestamp 1698431365
transform 1 0 71904 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_749
timestamp 1698431365
transform 1 0 5264 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_750
timestamp 1698431365
transform 1 0 13104 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_751
timestamp 1698431365
transform 1 0 20944 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_752
timestamp 1698431365
transform 1 0 28784 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_753
timestamp 1698431365
transform 1 0 36624 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_754
timestamp 1698431365
transform 1 0 44464 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_755
timestamp 1698431365
transform 1 0 52304 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_756
timestamp 1698431365
transform 1 0 60144 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_757
timestamp 1698431365
transform 1 0 67984 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_758
timestamp 1698431365
transform 1 0 75824 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_759
timestamp 1698431365
transform 1 0 9184 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_760
timestamp 1698431365
transform 1 0 17024 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_761
timestamp 1698431365
transform 1 0 24864 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_762
timestamp 1698431365
transform 1 0 32704 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_763
timestamp 1698431365
transform 1 0 40544 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_764
timestamp 1698431365
transform 1 0 48384 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_765
timestamp 1698431365
transform 1 0 56224 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_766
timestamp 1698431365
transform 1 0 64064 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_767
timestamp 1698431365
transform 1 0 71904 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_768
timestamp 1698431365
transform 1 0 5264 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_769
timestamp 1698431365
transform 1 0 13104 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_770
timestamp 1698431365
transform 1 0 20944 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_771
timestamp 1698431365
transform 1 0 28784 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_772
timestamp 1698431365
transform 1 0 36624 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_773
timestamp 1698431365
transform 1 0 44464 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_774
timestamp 1698431365
transform 1 0 52304 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_775
timestamp 1698431365
transform 1 0 60144 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_776
timestamp 1698431365
transform 1 0 67984 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_777
timestamp 1698431365
transform 1 0 75824 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_778
timestamp 1698431365
transform 1 0 9184 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_779
timestamp 1698431365
transform 1 0 17024 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_780
timestamp 1698431365
transform 1 0 24864 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_781
timestamp 1698431365
transform 1 0 32704 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_782
timestamp 1698431365
transform 1 0 40544 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_783
timestamp 1698431365
transform 1 0 48384 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_784
timestamp 1698431365
transform 1 0 56224 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_785
timestamp 1698431365
transform 1 0 64064 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_786
timestamp 1698431365
transform 1 0 71904 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_787
timestamp 1698431365
transform 1 0 5264 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_788
timestamp 1698431365
transform 1 0 13104 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_789
timestamp 1698431365
transform 1 0 20944 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_790
timestamp 1698431365
transform 1 0 28784 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_791
timestamp 1698431365
transform 1 0 36624 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_792
timestamp 1698431365
transform 1 0 44464 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_793
timestamp 1698431365
transform 1 0 52304 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_794
timestamp 1698431365
transform 1 0 60144 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_795
timestamp 1698431365
transform 1 0 67984 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_796
timestamp 1698431365
transform 1 0 75824 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_797
timestamp 1698431365
transform 1 0 9184 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_798
timestamp 1698431365
transform 1 0 17024 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_799
timestamp 1698431365
transform 1 0 24864 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_800
timestamp 1698431365
transform 1 0 32704 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_801
timestamp 1698431365
transform 1 0 40544 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_802
timestamp 1698431365
transform 1 0 48384 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_803
timestamp 1698431365
transform 1 0 56224 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_804
timestamp 1698431365
transform 1 0 64064 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_805
timestamp 1698431365
transform 1 0 71904 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_806
timestamp 1698431365
transform 1 0 5264 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_807
timestamp 1698431365
transform 1 0 13104 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_808
timestamp 1698431365
transform 1 0 20944 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_809
timestamp 1698431365
transform 1 0 28784 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_810
timestamp 1698431365
transform 1 0 36624 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_811
timestamp 1698431365
transform 1 0 44464 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_812
timestamp 1698431365
transform 1 0 52304 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_813
timestamp 1698431365
transform 1 0 60144 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_814
timestamp 1698431365
transform 1 0 67984 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_815
timestamp 1698431365
transform 1 0 75824 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_816
timestamp 1698431365
transform 1 0 9184 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_817
timestamp 1698431365
transform 1 0 17024 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_818
timestamp 1698431365
transform 1 0 24864 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_819
timestamp 1698431365
transform 1 0 32704 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_820
timestamp 1698431365
transform 1 0 40544 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_821
timestamp 1698431365
transform 1 0 48384 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_822
timestamp 1698431365
transform 1 0 56224 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_823
timestamp 1698431365
transform 1 0 64064 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_824
timestamp 1698431365
transform 1 0 71904 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_825
timestamp 1698431365
transform 1 0 5264 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_826
timestamp 1698431365
transform 1 0 13104 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_827
timestamp 1698431365
transform 1 0 20944 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_828
timestamp 1698431365
transform 1 0 28784 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_829
timestamp 1698431365
transform 1 0 36624 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_830
timestamp 1698431365
transform 1 0 44464 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_831
timestamp 1698431365
transform 1 0 52304 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_832
timestamp 1698431365
transform 1 0 60144 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_833
timestamp 1698431365
transform 1 0 67984 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_834
timestamp 1698431365
transform 1 0 75824 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_835
timestamp 1698431365
transform 1 0 9184 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_836
timestamp 1698431365
transform 1 0 17024 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_837
timestamp 1698431365
transform 1 0 24864 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_838
timestamp 1698431365
transform 1 0 32704 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_839
timestamp 1698431365
transform 1 0 40544 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_840
timestamp 1698431365
transform 1 0 48384 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_841
timestamp 1698431365
transform 1 0 56224 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_842
timestamp 1698431365
transform 1 0 64064 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_843
timestamp 1698431365
transform 1 0 71904 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_68_844
timestamp 1698431365
transform 1 0 5264 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_68_845
timestamp 1698431365
transform 1 0 13104 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_68_846
timestamp 1698431365
transform 1 0 20944 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_68_847
timestamp 1698431365
transform 1 0 28784 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_68_848
timestamp 1698431365
transform 1 0 36624 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_68_849
timestamp 1698431365
transform 1 0 44464 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_68_850
timestamp 1698431365
transform 1 0 52304 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_68_851
timestamp 1698431365
transform 1 0 60144 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_68_852
timestamp 1698431365
transform 1 0 67984 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_68_853
timestamp 1698431365
transform 1 0 75824 0 1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_69_854
timestamp 1698431365
transform 1 0 9184 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_69_855
timestamp 1698431365
transform 1 0 17024 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_69_856
timestamp 1698431365
transform 1 0 24864 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_69_857
timestamp 1698431365
transform 1 0 32704 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_69_858
timestamp 1698431365
transform 1 0 40544 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_69_859
timestamp 1698431365
transform 1 0 48384 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_69_860
timestamp 1698431365
transform 1 0 56224 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_69_861
timestamp 1698431365
transform 1 0 64064 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_69_862
timestamp 1698431365
transform 1 0 71904 0 -1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_863
timestamp 1698431365
transform 1 0 5264 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_864
timestamp 1698431365
transform 1 0 13104 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_865
timestamp 1698431365
transform 1 0 20944 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_866
timestamp 1698431365
transform 1 0 28784 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_867
timestamp 1698431365
transform 1 0 36624 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_868
timestamp 1698431365
transform 1 0 44464 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_869
timestamp 1698431365
transform 1 0 52304 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_870
timestamp 1698431365
transform 1 0 60144 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_871
timestamp 1698431365
transform 1 0 67984 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_70_872
timestamp 1698431365
transform 1 0 75824 0 1 58016
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_71_873
timestamp 1698431365
transform 1 0 9184 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_71_874
timestamp 1698431365
transform 1 0 17024 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_71_875
timestamp 1698431365
transform 1 0 24864 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_71_876
timestamp 1698431365
transform 1 0 32704 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_71_877
timestamp 1698431365
transform 1 0 40544 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_71_878
timestamp 1698431365
transform 1 0 48384 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_71_879
timestamp 1698431365
transform 1 0 56224 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_71_880
timestamp 1698431365
transform 1 0 64064 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_71_881
timestamp 1698431365
transform 1 0 71904 0 -1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_72_882
timestamp 1698431365
transform 1 0 5264 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_72_883
timestamp 1698431365
transform 1 0 13104 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_72_884
timestamp 1698431365
transform 1 0 20944 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_72_885
timestamp 1698431365
transform 1 0 28784 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_72_886
timestamp 1698431365
transform 1 0 36624 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_72_887
timestamp 1698431365
transform 1 0 44464 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_72_888
timestamp 1698431365
transform 1 0 52304 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_72_889
timestamp 1698431365
transform 1 0 60144 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_72_890
timestamp 1698431365
transform 1 0 67984 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_72_891
timestamp 1698431365
transform 1 0 75824 0 1 59584
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_73_892
timestamp 1698431365
transform 1 0 9184 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_73_893
timestamp 1698431365
transform 1 0 17024 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_73_894
timestamp 1698431365
transform 1 0 24864 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_73_895
timestamp 1698431365
transform 1 0 32704 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_73_896
timestamp 1698431365
transform 1 0 40544 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_73_897
timestamp 1698431365
transform 1 0 48384 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_73_898
timestamp 1698431365
transform 1 0 56224 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_73_899
timestamp 1698431365
transform 1 0 64064 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_73_900
timestamp 1698431365
transform 1 0 71904 0 -1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_74_901
timestamp 1698431365
transform 1 0 5264 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_74_902
timestamp 1698431365
transform 1 0 13104 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_74_903
timestamp 1698431365
transform 1 0 20944 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_74_904
timestamp 1698431365
transform 1 0 28784 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_74_905
timestamp 1698431365
transform 1 0 36624 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_74_906
timestamp 1698431365
transform 1 0 44464 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_74_907
timestamp 1698431365
transform 1 0 52304 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_74_908
timestamp 1698431365
transform 1 0 60144 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_74_909
timestamp 1698431365
transform 1 0 67984 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_74_910
timestamp 1698431365
transform 1 0 75824 0 1 61152
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_75_911
timestamp 1698431365
transform 1 0 9184 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_75_912
timestamp 1698431365
transform 1 0 17024 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_75_913
timestamp 1698431365
transform 1 0 24864 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_75_914
timestamp 1698431365
transform 1 0 32704 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_75_915
timestamp 1698431365
transform 1 0 40544 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_75_916
timestamp 1698431365
transform 1 0 48384 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_75_917
timestamp 1698431365
transform 1 0 56224 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_75_918
timestamp 1698431365
transform 1 0 64064 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_75_919
timestamp 1698431365
transform 1 0 71904 0 -1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_76_920
timestamp 1698431365
transform 1 0 5264 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_76_921
timestamp 1698431365
transform 1 0 13104 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_76_922
timestamp 1698431365
transform 1 0 20944 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_76_923
timestamp 1698431365
transform 1 0 28784 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_76_924
timestamp 1698431365
transform 1 0 36624 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_76_925
timestamp 1698431365
transform 1 0 44464 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_76_926
timestamp 1698431365
transform 1 0 52304 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_76_927
timestamp 1698431365
transform 1 0 60144 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_76_928
timestamp 1698431365
transform 1 0 67984 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_76_929
timestamp 1698431365
transform 1 0 75824 0 1 62720
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_77_930
timestamp 1698431365
transform 1 0 9184 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_77_931
timestamp 1698431365
transform 1 0 17024 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_77_932
timestamp 1698431365
transform 1 0 24864 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_77_933
timestamp 1698431365
transform 1 0 32704 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_77_934
timestamp 1698431365
transform 1 0 40544 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_77_935
timestamp 1698431365
transform 1 0 48384 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_77_936
timestamp 1698431365
transform 1 0 56224 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_77_937
timestamp 1698431365
transform 1 0 64064 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_77_938
timestamp 1698431365
transform 1 0 71904 0 -1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_78_939
timestamp 1698431365
transform 1 0 5264 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_78_940
timestamp 1698431365
transform 1 0 13104 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_78_941
timestamp 1698431365
transform 1 0 20944 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_78_942
timestamp 1698431365
transform 1 0 28784 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_78_943
timestamp 1698431365
transform 1 0 36624 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_78_944
timestamp 1698431365
transform 1 0 44464 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_78_945
timestamp 1698431365
transform 1 0 52304 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_78_946
timestamp 1698431365
transform 1 0 60144 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_78_947
timestamp 1698431365
transform 1 0 67984 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_78_948
timestamp 1698431365
transform 1 0 75824 0 1 64288
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_79_949
timestamp 1698431365
transform 1 0 9184 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_79_950
timestamp 1698431365
transform 1 0 17024 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_79_951
timestamp 1698431365
transform 1 0 24864 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_79_952
timestamp 1698431365
transform 1 0 32704 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_79_953
timestamp 1698431365
transform 1 0 40544 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_79_954
timestamp 1698431365
transform 1 0 48384 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_79_955
timestamp 1698431365
transform 1 0 56224 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_79_956
timestamp 1698431365
transform 1 0 64064 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_79_957
timestamp 1698431365
transform 1 0 71904 0 -1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_80_958
timestamp 1698431365
transform 1 0 5264 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_80_959
timestamp 1698431365
transform 1 0 13104 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_80_960
timestamp 1698431365
transform 1 0 20944 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_80_961
timestamp 1698431365
transform 1 0 28784 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_80_962
timestamp 1698431365
transform 1 0 36624 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_80_963
timestamp 1698431365
transform 1 0 44464 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_80_964
timestamp 1698431365
transform 1 0 52304 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_80_965
timestamp 1698431365
transform 1 0 60144 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_80_966
timestamp 1698431365
transform 1 0 67984 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_80_967
timestamp 1698431365
transform 1 0 75824 0 1 65856
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_81_968
timestamp 1698431365
transform 1 0 9184 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_81_969
timestamp 1698431365
transform 1 0 17024 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_81_970
timestamp 1698431365
transform 1 0 24864 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_81_971
timestamp 1698431365
transform 1 0 32704 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_81_972
timestamp 1698431365
transform 1 0 40544 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_81_973
timestamp 1698431365
transform 1 0 48384 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_81_974
timestamp 1698431365
transform 1 0 56224 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_81_975
timestamp 1698431365
transform 1 0 64064 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_81_976
timestamp 1698431365
transform 1 0 71904 0 -1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_82_977
timestamp 1698431365
transform 1 0 5264 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_82_978
timestamp 1698431365
transform 1 0 13104 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_82_979
timestamp 1698431365
transform 1 0 20944 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_82_980
timestamp 1698431365
transform 1 0 28784 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_82_981
timestamp 1698431365
transform 1 0 36624 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_82_982
timestamp 1698431365
transform 1 0 44464 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_82_983
timestamp 1698431365
transform 1 0 52304 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_82_984
timestamp 1698431365
transform 1 0 60144 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_82_985
timestamp 1698431365
transform 1 0 67984 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_82_986
timestamp 1698431365
transform 1 0 75824 0 1 67424
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_83_987
timestamp 1698431365
transform 1 0 9184 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_83_988
timestamp 1698431365
transform 1 0 17024 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_83_989
timestamp 1698431365
transform 1 0 24864 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_83_990
timestamp 1698431365
transform 1 0 32704 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_83_991
timestamp 1698431365
transform 1 0 40544 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_83_992
timestamp 1698431365
transform 1 0 48384 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_83_993
timestamp 1698431365
transform 1 0 56224 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_83_994
timestamp 1698431365
transform 1 0 64064 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_83_995
timestamp 1698431365
transform 1 0 71904 0 -1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_84_996
timestamp 1698431365
transform 1 0 5264 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_84_997
timestamp 1698431365
transform 1 0 13104 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_84_998
timestamp 1698431365
transform 1 0 20944 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_84_999
timestamp 1698431365
transform 1 0 28784 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_84_1000
timestamp 1698431365
transform 1 0 36624 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_84_1001
timestamp 1698431365
transform 1 0 44464 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_84_1002
timestamp 1698431365
transform 1 0 52304 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_84_1003
timestamp 1698431365
transform 1 0 60144 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_84_1004
timestamp 1698431365
transform 1 0 67984 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_84_1005
timestamp 1698431365
transform 1 0 75824 0 1 68992
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_85_1006
timestamp 1698431365
transform 1 0 9184 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_85_1007
timestamp 1698431365
transform 1 0 17024 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_85_1008
timestamp 1698431365
transform 1 0 24864 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_85_1009
timestamp 1698431365
transform 1 0 32704 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_85_1010
timestamp 1698431365
transform 1 0 40544 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_85_1011
timestamp 1698431365
transform 1 0 48384 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_85_1012
timestamp 1698431365
transform 1 0 56224 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_85_1013
timestamp 1698431365
transform 1 0 64064 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_85_1014
timestamp 1698431365
transform 1 0 71904 0 -1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_86_1015
timestamp 1698431365
transform 1 0 5264 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_86_1016
timestamp 1698431365
transform 1 0 13104 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_86_1017
timestamp 1698431365
transform 1 0 20944 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_86_1018
timestamp 1698431365
transform 1 0 28784 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_86_1019
timestamp 1698431365
transform 1 0 36624 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_86_1020
timestamp 1698431365
transform 1 0 44464 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_86_1021
timestamp 1698431365
transform 1 0 52304 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_86_1022
timestamp 1698431365
transform 1 0 60144 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_86_1023
timestamp 1698431365
transform 1 0 67984 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_86_1024
timestamp 1698431365
transform 1 0 75824 0 1 70560
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_87_1025
timestamp 1698431365
transform 1 0 9184 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_87_1026
timestamp 1698431365
transform 1 0 17024 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_87_1027
timestamp 1698431365
transform 1 0 24864 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_87_1028
timestamp 1698431365
transform 1 0 32704 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_87_1029
timestamp 1698431365
transform 1 0 40544 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_87_1030
timestamp 1698431365
transform 1 0 48384 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_87_1031
timestamp 1698431365
transform 1 0 56224 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_87_1032
timestamp 1698431365
transform 1 0 64064 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_87_1033
timestamp 1698431365
transform 1 0 71904 0 -1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_88_1034
timestamp 1698431365
transform 1 0 5264 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_88_1035
timestamp 1698431365
transform 1 0 13104 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_88_1036
timestamp 1698431365
transform 1 0 20944 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_88_1037
timestamp 1698431365
transform 1 0 28784 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_88_1038
timestamp 1698431365
transform 1 0 36624 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_88_1039
timestamp 1698431365
transform 1 0 44464 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_88_1040
timestamp 1698431365
transform 1 0 52304 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_88_1041
timestamp 1698431365
transform 1 0 60144 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_88_1042
timestamp 1698431365
transform 1 0 67984 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_88_1043
timestamp 1698431365
transform 1 0 75824 0 1 72128
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_89_1044
timestamp 1698431365
transform 1 0 9184 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_89_1045
timestamp 1698431365
transform 1 0 17024 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_89_1046
timestamp 1698431365
transform 1 0 24864 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_89_1047
timestamp 1698431365
transform 1 0 32704 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_89_1048
timestamp 1698431365
transform 1 0 40544 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_89_1049
timestamp 1698431365
transform 1 0 48384 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_89_1050
timestamp 1698431365
transform 1 0 56224 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_89_1051
timestamp 1698431365
transform 1 0 64064 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_89_1052
timestamp 1698431365
transform 1 0 71904 0 -1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_90_1053
timestamp 1698431365
transform 1 0 5264 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_90_1054
timestamp 1698431365
transform 1 0 13104 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_90_1055
timestamp 1698431365
transform 1 0 20944 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_90_1056
timestamp 1698431365
transform 1 0 28784 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_90_1057
timestamp 1698431365
transform 1 0 36624 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_90_1058
timestamp 1698431365
transform 1 0 44464 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_90_1059
timestamp 1698431365
transform 1 0 52304 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_90_1060
timestamp 1698431365
transform 1 0 60144 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_90_1061
timestamp 1698431365
transform 1 0 67984 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_90_1062
timestamp 1698431365
transform 1 0 75824 0 1 73696
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_91_1063
timestamp 1698431365
transform 1 0 9184 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_91_1064
timestamp 1698431365
transform 1 0 17024 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_91_1065
timestamp 1698431365
transform 1 0 24864 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_91_1066
timestamp 1698431365
transform 1 0 32704 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_91_1067
timestamp 1698431365
transform 1 0 40544 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_91_1068
timestamp 1698431365
transform 1 0 48384 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_91_1069
timestamp 1698431365
transform 1 0 56224 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_91_1070
timestamp 1698431365
transform 1 0 64064 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_91_1071
timestamp 1698431365
transform 1 0 71904 0 -1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_92_1072
timestamp 1698431365
transform 1 0 5264 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_92_1073
timestamp 1698431365
transform 1 0 13104 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_92_1074
timestamp 1698431365
transform 1 0 20944 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_92_1075
timestamp 1698431365
transform 1 0 28784 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_92_1076
timestamp 1698431365
transform 1 0 36624 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_92_1077
timestamp 1698431365
transform 1 0 44464 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_92_1078
timestamp 1698431365
transform 1 0 52304 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_92_1079
timestamp 1698431365
transform 1 0 60144 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_92_1080
timestamp 1698431365
transform 1 0 67984 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_92_1081
timestamp 1698431365
transform 1 0 75824 0 1 75264
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_93_1082
timestamp 1698431365
transform 1 0 5152 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_93_1083
timestamp 1698431365
transform 1 0 8960 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_93_1084
timestamp 1698431365
transform 1 0 12768 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_93_1085
timestamp 1698431365
transform 1 0 16576 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_93_1086
timestamp 1698431365
transform 1 0 20384 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_93_1087
timestamp 1698431365
transform 1 0 24192 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_93_1088
timestamp 1698431365
transform 1 0 28000 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_93_1089
timestamp 1698431365
transform 1 0 31808 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_93_1090
timestamp 1698431365
transform 1 0 35616 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_93_1091
timestamp 1698431365
transform 1 0 39424 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_93_1092
timestamp 1698431365
transform 1 0 43232 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_93_1093
timestamp 1698431365
transform 1 0 47040 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_93_1094
timestamp 1698431365
transform 1 0 50848 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_93_1095
timestamp 1698431365
transform 1 0 54656 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_93_1096
timestamp 1698431365
transform 1 0 58464 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_93_1097
timestamp 1698431365
transform 1 0 62272 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_93_1098
timestamp 1698431365
transform 1 0 66080 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_93_1099
timestamp 1698431365
transform 1 0 69888 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_93_1100
timestamp 1698431365
transform 1 0 73696 0 -1 76832
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_93_1101
timestamp 1698431365
transform 1 0 77504 0 -1 76832
box -86 -86 310 870
<< labels >>
flabel metal2 s 74144 0 74256 800 0 FreeSans 448 90 0 0 clk
port 0 nsew signal input
flabel metal2 s 448 79200 560 80000 0 FreeSans 448 90 0 0 gpio_in[0]
port 1 nsew signal input
flabel metal2 s 7168 79200 7280 80000 0 FreeSans 448 90 0 0 gpio_in[10]
port 2 nsew signal input
flabel metal2 s 7840 79200 7952 80000 0 FreeSans 448 90 0 0 gpio_in[11]
port 3 nsew signal input
flabel metal2 s 8512 79200 8624 80000 0 FreeSans 448 90 0 0 gpio_in[12]
port 4 nsew signal input
flabel metal2 s 9184 79200 9296 80000 0 FreeSans 448 90 0 0 gpio_in[13]
port 5 nsew signal input
flabel metal2 s 9856 79200 9968 80000 0 FreeSans 448 90 0 0 gpio_in[14]
port 6 nsew signal input
flabel metal2 s 10528 79200 10640 80000 0 FreeSans 448 90 0 0 gpio_in[15]
port 7 nsew signal input
flabel metal2 s 1120 79200 1232 80000 0 FreeSans 448 90 0 0 gpio_in[1]
port 8 nsew signal input
flabel metal2 s 1792 79200 1904 80000 0 FreeSans 448 90 0 0 gpio_in[2]
port 9 nsew signal input
flabel metal2 s 2464 79200 2576 80000 0 FreeSans 448 90 0 0 gpio_in[3]
port 10 nsew signal input
flabel metal2 s 3136 79200 3248 80000 0 FreeSans 448 90 0 0 gpio_in[4]
port 11 nsew signal input
flabel metal2 s 3808 79200 3920 80000 0 FreeSans 448 90 0 0 gpio_in[5]
port 12 nsew signal input
flabel metal2 s 4480 79200 4592 80000 0 FreeSans 448 90 0 0 gpio_in[6]
port 13 nsew signal input
flabel metal2 s 5152 79200 5264 80000 0 FreeSans 448 90 0 0 gpio_in[7]
port 14 nsew signal input
flabel metal2 s 5824 79200 5936 80000 0 FreeSans 448 90 0 0 gpio_in[8]
port 15 nsew signal input
flabel metal2 s 6496 79200 6608 80000 0 FreeSans 448 90 0 0 gpio_in[9]
port 16 nsew signal input
flabel metal2 s 21952 79200 22064 80000 0 FreeSans 448 90 0 0 gpio_oeb[0]
port 17 nsew signal tristate
flabel metal2 s 28672 79200 28784 80000 0 FreeSans 448 90 0 0 gpio_oeb[10]
port 18 nsew signal tristate
flabel metal2 s 29344 79200 29456 80000 0 FreeSans 448 90 0 0 gpio_oeb[11]
port 19 nsew signal tristate
flabel metal2 s 30016 79200 30128 80000 0 FreeSans 448 90 0 0 gpio_oeb[12]
port 20 nsew signal tristate
flabel metal2 s 30688 79200 30800 80000 0 FreeSans 448 90 0 0 gpio_oeb[13]
port 21 nsew signal tristate
flabel metal2 s 31360 79200 31472 80000 0 FreeSans 448 90 0 0 gpio_oeb[14]
port 22 nsew signal tristate
flabel metal2 s 32032 79200 32144 80000 0 FreeSans 448 90 0 0 gpio_oeb[15]
port 23 nsew signal tristate
flabel metal2 s 22624 79200 22736 80000 0 FreeSans 448 90 0 0 gpio_oeb[1]
port 24 nsew signal tristate
flabel metal2 s 23296 79200 23408 80000 0 FreeSans 448 90 0 0 gpio_oeb[2]
port 25 nsew signal tristate
flabel metal2 s 23968 79200 24080 80000 0 FreeSans 448 90 0 0 gpio_oeb[3]
port 26 nsew signal tristate
flabel metal2 s 24640 79200 24752 80000 0 FreeSans 448 90 0 0 gpio_oeb[4]
port 27 nsew signal tristate
flabel metal2 s 25312 79200 25424 80000 0 FreeSans 448 90 0 0 gpio_oeb[5]
port 28 nsew signal tristate
flabel metal2 s 25984 79200 26096 80000 0 FreeSans 448 90 0 0 gpio_oeb[6]
port 29 nsew signal tristate
flabel metal2 s 26656 79200 26768 80000 0 FreeSans 448 90 0 0 gpio_oeb[7]
port 30 nsew signal tristate
flabel metal2 s 27328 79200 27440 80000 0 FreeSans 448 90 0 0 gpio_oeb[8]
port 31 nsew signal tristate
flabel metal2 s 28000 79200 28112 80000 0 FreeSans 448 90 0 0 gpio_oeb[9]
port 32 nsew signal tristate
flabel metal2 s 11200 79200 11312 80000 0 FreeSans 448 90 0 0 gpio_out[0]
port 33 nsew signal tristate
flabel metal2 s 17920 79200 18032 80000 0 FreeSans 448 90 0 0 gpio_out[10]
port 34 nsew signal tristate
flabel metal2 s 18592 79200 18704 80000 0 FreeSans 448 90 0 0 gpio_out[11]
port 35 nsew signal tristate
flabel metal2 s 19264 79200 19376 80000 0 FreeSans 448 90 0 0 gpio_out[12]
port 36 nsew signal tristate
flabel metal2 s 19936 79200 20048 80000 0 FreeSans 448 90 0 0 gpio_out[13]
port 37 nsew signal tristate
flabel metal2 s 20608 79200 20720 80000 0 FreeSans 448 90 0 0 gpio_out[14]
port 38 nsew signal tristate
flabel metal2 s 21280 79200 21392 80000 0 FreeSans 448 90 0 0 gpio_out[15]
port 39 nsew signal tristate
flabel metal2 s 11872 79200 11984 80000 0 FreeSans 448 90 0 0 gpio_out[1]
port 40 nsew signal tristate
flabel metal2 s 12544 79200 12656 80000 0 FreeSans 448 90 0 0 gpio_out[2]
port 41 nsew signal tristate
flabel metal2 s 13216 79200 13328 80000 0 FreeSans 448 90 0 0 gpio_out[3]
port 42 nsew signal tristate
flabel metal2 s 13888 79200 14000 80000 0 FreeSans 448 90 0 0 gpio_out[4]
port 43 nsew signal tristate
flabel metal2 s 14560 79200 14672 80000 0 FreeSans 448 90 0 0 gpio_out[5]
port 44 nsew signal tristate
flabel metal2 s 15232 79200 15344 80000 0 FreeSans 448 90 0 0 gpio_out[6]
port 45 nsew signal tristate
flabel metal2 s 15904 79200 16016 80000 0 FreeSans 448 90 0 0 gpio_out[7]
port 46 nsew signal tristate
flabel metal2 s 16576 79200 16688 80000 0 FreeSans 448 90 0 0 gpio_out[8]
port 47 nsew signal tristate
flabel metal2 s 17248 79200 17360 80000 0 FreeSans 448 90 0 0 gpio_out[9]
port 48 nsew signal tristate
flabel metal2 s 26432 0 26544 800 0 FreeSans 448 90 0 0 mem_addr[0]
port 49 nsew signal input
flabel metal2 s 33152 0 33264 800 0 FreeSans 448 90 0 0 mem_addr[10]
port 50 nsew signal input
flabel metal2 s 33824 0 33936 800 0 FreeSans 448 90 0 0 mem_addr[11]
port 51 nsew signal input
flabel metal2 s 34496 0 34608 800 0 FreeSans 448 90 0 0 mem_addr[12]
port 52 nsew signal input
flabel metal2 s 35168 0 35280 800 0 FreeSans 448 90 0 0 mem_addr[13]
port 53 nsew signal input
flabel metal2 s 35840 0 35952 800 0 FreeSans 448 90 0 0 mem_addr[14]
port 54 nsew signal input
flabel metal2 s 36512 0 36624 800 0 FreeSans 448 90 0 0 mem_addr[15]
port 55 nsew signal input
flabel metal2 s 37184 0 37296 800 0 FreeSans 448 90 0 0 mem_addr[16]
port 56 nsew signal input
flabel metal2 s 37856 0 37968 800 0 FreeSans 448 90 0 0 mem_addr[17]
port 57 nsew signal input
flabel metal2 s 38528 0 38640 800 0 FreeSans 448 90 0 0 mem_addr[18]
port 58 nsew signal input
flabel metal2 s 39200 0 39312 800 0 FreeSans 448 90 0 0 mem_addr[19]
port 59 nsew signal input
flabel metal2 s 27104 0 27216 800 0 FreeSans 448 90 0 0 mem_addr[1]
port 60 nsew signal input
flabel metal2 s 39872 0 39984 800 0 FreeSans 448 90 0 0 mem_addr[20]
port 61 nsew signal input
flabel metal2 s 40544 0 40656 800 0 FreeSans 448 90 0 0 mem_addr[21]
port 62 nsew signal input
flabel metal2 s 41216 0 41328 800 0 FreeSans 448 90 0 0 mem_addr[22]
port 63 nsew signal input
flabel metal2 s 41888 0 42000 800 0 FreeSans 448 90 0 0 mem_addr[23]
port 64 nsew signal input
flabel metal2 s 42560 0 42672 800 0 FreeSans 448 90 0 0 mem_addr[24]
port 65 nsew signal input
flabel metal2 s 43232 0 43344 800 0 FreeSans 448 90 0 0 mem_addr[25]
port 66 nsew signal input
flabel metal2 s 43904 0 44016 800 0 FreeSans 448 90 0 0 mem_addr[26]
port 67 nsew signal input
flabel metal2 s 44576 0 44688 800 0 FreeSans 448 90 0 0 mem_addr[27]
port 68 nsew signal input
flabel metal2 s 45248 0 45360 800 0 FreeSans 448 90 0 0 mem_addr[28]
port 69 nsew signal input
flabel metal2 s 45920 0 46032 800 0 FreeSans 448 90 0 0 mem_addr[29]
port 70 nsew signal input
flabel metal2 s 27776 0 27888 800 0 FreeSans 448 90 0 0 mem_addr[2]
port 71 nsew signal input
flabel metal2 s 46592 0 46704 800 0 FreeSans 448 90 0 0 mem_addr[30]
port 72 nsew signal input
flabel metal2 s 47264 0 47376 800 0 FreeSans 448 90 0 0 mem_addr[31]
port 73 nsew signal input
flabel metal2 s 28448 0 28560 800 0 FreeSans 448 90 0 0 mem_addr[3]
port 74 nsew signal input
flabel metal2 s 29120 0 29232 800 0 FreeSans 448 90 0 0 mem_addr[4]
port 75 nsew signal input
flabel metal2 s 29792 0 29904 800 0 FreeSans 448 90 0 0 mem_addr[5]
port 76 nsew signal input
flabel metal2 s 30464 0 30576 800 0 FreeSans 448 90 0 0 mem_addr[6]
port 77 nsew signal input
flabel metal2 s 31136 0 31248 800 0 FreeSans 448 90 0 0 mem_addr[7]
port 78 nsew signal input
flabel metal2 s 31808 0 31920 800 0 FreeSans 448 90 0 0 mem_addr[8]
port 79 nsew signal input
flabel metal2 s 32480 0 32592 800 0 FreeSans 448 90 0 0 mem_addr[9]
port 80 nsew signal input
flabel metal2 s 48608 0 48720 800 0 FreeSans 448 90 0 0 mem_instr
port 81 nsew signal input
flabel metal2 s 52640 0 52752 800 0 FreeSans 448 90 0 0 mem_rdata[0]
port 82 nsew signal tristate
flabel metal2 s 59360 0 59472 800 0 FreeSans 448 90 0 0 mem_rdata[10]
port 83 nsew signal tristate
flabel metal2 s 60032 0 60144 800 0 FreeSans 448 90 0 0 mem_rdata[11]
port 84 nsew signal tristate
flabel metal2 s 60704 0 60816 800 0 FreeSans 448 90 0 0 mem_rdata[12]
port 85 nsew signal tristate
flabel metal2 s 61376 0 61488 800 0 FreeSans 448 90 0 0 mem_rdata[13]
port 86 nsew signal tristate
flabel metal2 s 62048 0 62160 800 0 FreeSans 448 90 0 0 mem_rdata[14]
port 87 nsew signal tristate
flabel metal2 s 62720 0 62832 800 0 FreeSans 448 90 0 0 mem_rdata[15]
port 88 nsew signal tristate
flabel metal2 s 63392 0 63504 800 0 FreeSans 448 90 0 0 mem_rdata[16]
port 89 nsew signal tristate
flabel metal2 s 64064 0 64176 800 0 FreeSans 448 90 0 0 mem_rdata[17]
port 90 nsew signal tristate
flabel metal2 s 64736 0 64848 800 0 FreeSans 448 90 0 0 mem_rdata[18]
port 91 nsew signal tristate
flabel metal2 s 65408 0 65520 800 0 FreeSans 448 90 0 0 mem_rdata[19]
port 92 nsew signal tristate
flabel metal2 s 53312 0 53424 800 0 FreeSans 448 90 0 0 mem_rdata[1]
port 93 nsew signal tristate
flabel metal2 s 66080 0 66192 800 0 FreeSans 448 90 0 0 mem_rdata[20]
port 94 nsew signal tristate
flabel metal2 s 66752 0 66864 800 0 FreeSans 448 90 0 0 mem_rdata[21]
port 95 nsew signal tristate
flabel metal2 s 67424 0 67536 800 0 FreeSans 448 90 0 0 mem_rdata[22]
port 96 nsew signal tristate
flabel metal2 s 68096 0 68208 800 0 FreeSans 448 90 0 0 mem_rdata[23]
port 97 nsew signal tristate
flabel metal2 s 68768 0 68880 800 0 FreeSans 448 90 0 0 mem_rdata[24]
port 98 nsew signal tristate
flabel metal2 s 69440 0 69552 800 0 FreeSans 448 90 0 0 mem_rdata[25]
port 99 nsew signal tristate
flabel metal2 s 70112 0 70224 800 0 FreeSans 448 90 0 0 mem_rdata[26]
port 100 nsew signal tristate
flabel metal2 s 70784 0 70896 800 0 FreeSans 448 90 0 0 mem_rdata[27]
port 101 nsew signal tristate
flabel metal2 s 71456 0 71568 800 0 FreeSans 448 90 0 0 mem_rdata[28]
port 102 nsew signal tristate
flabel metal2 s 72128 0 72240 800 0 FreeSans 448 90 0 0 mem_rdata[29]
port 103 nsew signal tristate
flabel metal2 s 53984 0 54096 800 0 FreeSans 448 90 0 0 mem_rdata[2]
port 104 nsew signal tristate
flabel metal2 s 72800 0 72912 800 0 FreeSans 448 90 0 0 mem_rdata[30]
port 105 nsew signal tristate
flabel metal2 s 73472 0 73584 800 0 FreeSans 448 90 0 0 mem_rdata[31]
port 106 nsew signal tristate
flabel metal2 s 54656 0 54768 800 0 FreeSans 448 90 0 0 mem_rdata[3]
port 107 nsew signal tristate
flabel metal2 s 55328 0 55440 800 0 FreeSans 448 90 0 0 mem_rdata[4]
port 108 nsew signal tristate
flabel metal2 s 56000 0 56112 800 0 FreeSans 448 90 0 0 mem_rdata[5]
port 109 nsew signal tristate
flabel metal2 s 56672 0 56784 800 0 FreeSans 448 90 0 0 mem_rdata[6]
port 110 nsew signal tristate
flabel metal2 s 57344 0 57456 800 0 FreeSans 448 90 0 0 mem_rdata[7]
port 111 nsew signal tristate
flabel metal2 s 58016 0 58128 800 0 FreeSans 448 90 0 0 mem_rdata[8]
port 112 nsew signal tristate
flabel metal2 s 58688 0 58800 800 0 FreeSans 448 90 0 0 mem_rdata[9]
port 113 nsew signal tristate
flabel metal2 s 49280 0 49392 800 0 FreeSans 448 90 0 0 mem_ready
port 114 nsew signal tristate
flabel metal2 s 47936 0 48048 800 0 FreeSans 448 90 0 0 mem_valid
port 115 nsew signal input
flabel metal2 s 4928 0 5040 800 0 FreeSans 448 90 0 0 mem_wdata[0]
port 116 nsew signal input
flabel metal2 s 11648 0 11760 800 0 FreeSans 448 90 0 0 mem_wdata[10]
port 117 nsew signal input
flabel metal2 s 12320 0 12432 800 0 FreeSans 448 90 0 0 mem_wdata[11]
port 118 nsew signal input
flabel metal2 s 12992 0 13104 800 0 FreeSans 448 90 0 0 mem_wdata[12]
port 119 nsew signal input
flabel metal2 s 13664 0 13776 800 0 FreeSans 448 90 0 0 mem_wdata[13]
port 120 nsew signal input
flabel metal2 s 14336 0 14448 800 0 FreeSans 448 90 0 0 mem_wdata[14]
port 121 nsew signal input
flabel metal2 s 15008 0 15120 800 0 FreeSans 448 90 0 0 mem_wdata[15]
port 122 nsew signal input
flabel metal2 s 15680 0 15792 800 0 FreeSans 448 90 0 0 mem_wdata[16]
port 123 nsew signal input
flabel metal2 s 16352 0 16464 800 0 FreeSans 448 90 0 0 mem_wdata[17]
port 124 nsew signal input
flabel metal2 s 17024 0 17136 800 0 FreeSans 448 90 0 0 mem_wdata[18]
port 125 nsew signal input
flabel metal2 s 17696 0 17808 800 0 FreeSans 448 90 0 0 mem_wdata[19]
port 126 nsew signal input
flabel metal2 s 5600 0 5712 800 0 FreeSans 448 90 0 0 mem_wdata[1]
port 127 nsew signal input
flabel metal2 s 18368 0 18480 800 0 FreeSans 448 90 0 0 mem_wdata[20]
port 128 nsew signal input
flabel metal2 s 19040 0 19152 800 0 FreeSans 448 90 0 0 mem_wdata[21]
port 129 nsew signal input
flabel metal2 s 19712 0 19824 800 0 FreeSans 448 90 0 0 mem_wdata[22]
port 130 nsew signal input
flabel metal2 s 20384 0 20496 800 0 FreeSans 448 90 0 0 mem_wdata[23]
port 131 nsew signal input
flabel metal2 s 21056 0 21168 800 0 FreeSans 448 90 0 0 mem_wdata[24]
port 132 nsew signal input
flabel metal2 s 21728 0 21840 800 0 FreeSans 448 90 0 0 mem_wdata[25]
port 133 nsew signal input
flabel metal2 s 22400 0 22512 800 0 FreeSans 448 90 0 0 mem_wdata[26]
port 134 nsew signal input
flabel metal2 s 23072 0 23184 800 0 FreeSans 448 90 0 0 mem_wdata[27]
port 135 nsew signal input
flabel metal2 s 23744 0 23856 800 0 FreeSans 448 90 0 0 mem_wdata[28]
port 136 nsew signal input
flabel metal2 s 24416 0 24528 800 0 FreeSans 448 90 0 0 mem_wdata[29]
port 137 nsew signal input
flabel metal2 s 6272 0 6384 800 0 FreeSans 448 90 0 0 mem_wdata[2]
port 138 nsew signal input
flabel metal2 s 25088 0 25200 800 0 FreeSans 448 90 0 0 mem_wdata[30]
port 139 nsew signal input
flabel metal2 s 25760 0 25872 800 0 FreeSans 448 90 0 0 mem_wdata[31]
port 140 nsew signal input
flabel metal2 s 6944 0 7056 800 0 FreeSans 448 90 0 0 mem_wdata[3]
port 141 nsew signal input
flabel metal2 s 7616 0 7728 800 0 FreeSans 448 90 0 0 mem_wdata[4]
port 142 nsew signal input
flabel metal2 s 8288 0 8400 800 0 FreeSans 448 90 0 0 mem_wdata[5]
port 143 nsew signal input
flabel metal2 s 8960 0 9072 800 0 FreeSans 448 90 0 0 mem_wdata[6]
port 144 nsew signal input
flabel metal2 s 9632 0 9744 800 0 FreeSans 448 90 0 0 mem_wdata[7]
port 145 nsew signal input
flabel metal2 s 10304 0 10416 800 0 FreeSans 448 90 0 0 mem_wdata[8]
port 146 nsew signal input
flabel metal2 s 10976 0 11088 800 0 FreeSans 448 90 0 0 mem_wdata[9]
port 147 nsew signal input
flabel metal2 s 49952 0 50064 800 0 FreeSans 448 90 0 0 mem_wstrb[0]
port 148 nsew signal input
flabel metal2 s 50624 0 50736 800 0 FreeSans 448 90 0 0 mem_wstrb[1]
port 149 nsew signal input
flabel metal2 s 51296 0 51408 800 0 FreeSans 448 90 0 0 mem_wstrb[2]
port 150 nsew signal input
flabel metal2 s 51968 0 52080 800 0 FreeSans 448 90 0 0 mem_wstrb[3]
port 151 nsew signal input
flabel metal3 s 0 38080 800 38192 0 FreeSans 448 0 0 0 ram_gwenb[0]
port 152 nsew signal tristate
flabel metal3 s 0 39200 800 39312 0 FreeSans 448 0 0 0 ram_gwenb[1]
port 153 nsew signal tristate
flabel metal3 s 0 40320 800 40432 0 FreeSans 448 0 0 0 ram_gwenb[2]
port 154 nsew signal tristate
flabel metal3 s 0 41440 800 41552 0 FreeSans 448 0 0 0 ram_gwenb[3]
port 155 nsew signal tristate
flabel metal3 s 0 2240 800 2352 0 FreeSans 448 0 0 0 ram_rdata[0]
port 156 nsew signal input
flabel metal3 s 0 13440 800 13552 0 FreeSans 448 0 0 0 ram_rdata[10]
port 157 nsew signal input
flabel metal3 s 0 14560 800 14672 0 FreeSans 448 0 0 0 ram_rdata[11]
port 158 nsew signal input
flabel metal3 s 0 15680 800 15792 0 FreeSans 448 0 0 0 ram_rdata[12]
port 159 nsew signal input
flabel metal3 s 0 16800 800 16912 0 FreeSans 448 0 0 0 ram_rdata[13]
port 160 nsew signal input
flabel metal3 s 0 17920 800 18032 0 FreeSans 448 0 0 0 ram_rdata[14]
port 161 nsew signal input
flabel metal3 s 0 19040 800 19152 0 FreeSans 448 0 0 0 ram_rdata[15]
port 162 nsew signal input
flabel metal3 s 0 20160 800 20272 0 FreeSans 448 0 0 0 ram_rdata[16]
port 163 nsew signal input
flabel metal3 s 0 21280 800 21392 0 FreeSans 448 0 0 0 ram_rdata[17]
port 164 nsew signal input
flabel metal3 s 0 22400 800 22512 0 FreeSans 448 0 0 0 ram_rdata[18]
port 165 nsew signal input
flabel metal3 s 0 23520 800 23632 0 FreeSans 448 0 0 0 ram_rdata[19]
port 166 nsew signal input
flabel metal3 s 0 3360 800 3472 0 FreeSans 448 0 0 0 ram_rdata[1]
port 167 nsew signal input
flabel metal3 s 0 24640 800 24752 0 FreeSans 448 0 0 0 ram_rdata[20]
port 168 nsew signal input
flabel metal3 s 0 25760 800 25872 0 FreeSans 448 0 0 0 ram_rdata[21]
port 169 nsew signal input
flabel metal3 s 0 26880 800 26992 0 FreeSans 448 0 0 0 ram_rdata[22]
port 170 nsew signal input
flabel metal3 s 0 28000 800 28112 0 FreeSans 448 0 0 0 ram_rdata[23]
port 171 nsew signal input
flabel metal3 s 0 29120 800 29232 0 FreeSans 448 0 0 0 ram_rdata[24]
port 172 nsew signal input
flabel metal3 s 0 30240 800 30352 0 FreeSans 448 0 0 0 ram_rdata[25]
port 173 nsew signal input
flabel metal3 s 0 31360 800 31472 0 FreeSans 448 0 0 0 ram_rdata[26]
port 174 nsew signal input
flabel metal3 s 0 32480 800 32592 0 FreeSans 448 0 0 0 ram_rdata[27]
port 175 nsew signal input
flabel metal3 s 0 33600 800 33712 0 FreeSans 448 0 0 0 ram_rdata[28]
port 176 nsew signal input
flabel metal3 s 0 34720 800 34832 0 FreeSans 448 0 0 0 ram_rdata[29]
port 177 nsew signal input
flabel metal3 s 0 4480 800 4592 0 FreeSans 448 0 0 0 ram_rdata[2]
port 178 nsew signal input
flabel metal3 s 0 35840 800 35952 0 FreeSans 448 0 0 0 ram_rdata[30]
port 179 nsew signal input
flabel metal3 s 0 36960 800 37072 0 FreeSans 448 0 0 0 ram_rdata[31]
port 180 nsew signal input
flabel metal3 s 0 5600 800 5712 0 FreeSans 448 0 0 0 ram_rdata[3]
port 181 nsew signal input
flabel metal3 s 0 6720 800 6832 0 FreeSans 448 0 0 0 ram_rdata[4]
port 182 nsew signal input
flabel metal3 s 0 7840 800 7952 0 FreeSans 448 0 0 0 ram_rdata[5]
port 183 nsew signal input
flabel metal3 s 0 8960 800 9072 0 FreeSans 448 0 0 0 ram_rdata[6]
port 184 nsew signal input
flabel metal3 s 0 10080 800 10192 0 FreeSans 448 0 0 0 ram_rdata[7]
port 185 nsew signal input
flabel metal3 s 0 11200 800 11312 0 FreeSans 448 0 0 0 ram_rdata[8]
port 186 nsew signal input
flabel metal3 s 0 12320 800 12432 0 FreeSans 448 0 0 0 ram_rdata[9]
port 187 nsew signal input
flabel metal3 s 0 42560 800 42672 0 FreeSans 448 0 0 0 ram_wenb[0]
port 188 nsew signal tristate
flabel metal3 s 0 53760 800 53872 0 FreeSans 448 0 0 0 ram_wenb[10]
port 189 nsew signal tristate
flabel metal3 s 0 54880 800 54992 0 FreeSans 448 0 0 0 ram_wenb[11]
port 190 nsew signal tristate
flabel metal3 s 0 56000 800 56112 0 FreeSans 448 0 0 0 ram_wenb[12]
port 191 nsew signal tristate
flabel metal3 s 0 57120 800 57232 0 FreeSans 448 0 0 0 ram_wenb[13]
port 192 nsew signal tristate
flabel metal3 s 0 58240 800 58352 0 FreeSans 448 0 0 0 ram_wenb[14]
port 193 nsew signal tristate
flabel metal3 s 0 59360 800 59472 0 FreeSans 448 0 0 0 ram_wenb[15]
port 194 nsew signal tristate
flabel metal3 s 0 60480 800 60592 0 FreeSans 448 0 0 0 ram_wenb[16]
port 195 nsew signal tristate
flabel metal3 s 0 61600 800 61712 0 FreeSans 448 0 0 0 ram_wenb[17]
port 196 nsew signal tristate
flabel metal3 s 0 62720 800 62832 0 FreeSans 448 0 0 0 ram_wenb[18]
port 197 nsew signal tristate
flabel metal3 s 0 63840 800 63952 0 FreeSans 448 0 0 0 ram_wenb[19]
port 198 nsew signal tristate
flabel metal3 s 0 43680 800 43792 0 FreeSans 448 0 0 0 ram_wenb[1]
port 199 nsew signal tristate
flabel metal3 s 0 64960 800 65072 0 FreeSans 448 0 0 0 ram_wenb[20]
port 200 nsew signal tristate
flabel metal3 s 0 66080 800 66192 0 FreeSans 448 0 0 0 ram_wenb[21]
port 201 nsew signal tristate
flabel metal3 s 0 67200 800 67312 0 FreeSans 448 0 0 0 ram_wenb[22]
port 202 nsew signal tristate
flabel metal3 s 0 68320 800 68432 0 FreeSans 448 0 0 0 ram_wenb[23]
port 203 nsew signal tristate
flabel metal3 s 0 69440 800 69552 0 FreeSans 448 0 0 0 ram_wenb[24]
port 204 nsew signal tristate
flabel metal3 s 0 70560 800 70672 0 FreeSans 448 0 0 0 ram_wenb[25]
port 205 nsew signal tristate
flabel metal3 s 0 71680 800 71792 0 FreeSans 448 0 0 0 ram_wenb[26]
port 206 nsew signal tristate
flabel metal3 s 0 72800 800 72912 0 FreeSans 448 0 0 0 ram_wenb[27]
port 207 nsew signal tristate
flabel metal3 s 0 73920 800 74032 0 FreeSans 448 0 0 0 ram_wenb[28]
port 208 nsew signal tristate
flabel metal3 s 0 75040 800 75152 0 FreeSans 448 0 0 0 ram_wenb[29]
port 209 nsew signal tristate
flabel metal3 s 0 44800 800 44912 0 FreeSans 448 0 0 0 ram_wenb[2]
port 210 nsew signal tristate
flabel metal3 s 0 76160 800 76272 0 FreeSans 448 0 0 0 ram_wenb[30]
port 211 nsew signal tristate
flabel metal3 s 0 77280 800 77392 0 FreeSans 448 0 0 0 ram_wenb[31]
port 212 nsew signal tristate
flabel metal3 s 0 45920 800 46032 0 FreeSans 448 0 0 0 ram_wenb[3]
port 213 nsew signal tristate
flabel metal3 s 0 47040 800 47152 0 FreeSans 448 0 0 0 ram_wenb[4]
port 214 nsew signal tristate
flabel metal3 s 0 48160 800 48272 0 FreeSans 448 0 0 0 ram_wenb[5]
port 215 nsew signal tristate
flabel metal3 s 0 49280 800 49392 0 FreeSans 448 0 0 0 ram_wenb[6]
port 216 nsew signal tristate
flabel metal3 s 0 50400 800 50512 0 FreeSans 448 0 0 0 ram_wenb[7]
port 217 nsew signal tristate
flabel metal3 s 0 51520 800 51632 0 FreeSans 448 0 0 0 ram_wenb[8]
port 218 nsew signal tristate
flabel metal3 s 0 52640 800 52752 0 FreeSans 448 0 0 0 ram_wenb[9]
port 219 nsew signal tristate
flabel metal2 s 74816 0 74928 800 0 FreeSans 448 90 0 0 resetn
port 220 nsew signal input
flabel metal3 s 79200 42112 80000 42224 0 FreeSans 448 0 0 0 simpleuart_dat_re
port 221 nsew signal tristate
flabel metal3 s 79200 40992 80000 41104 0 FreeSans 448 0 0 0 simpleuart_dat_we
port 222 nsew signal tristate
flabel metal3 s 79200 672 80000 784 0 FreeSans 448 0 0 0 simpleuart_div_we[0]
port 223 nsew signal tristate
flabel metal3 s 79200 1792 80000 1904 0 FreeSans 448 0 0 0 simpleuart_div_we[1]
port 224 nsew signal tristate
flabel metal3 s 79200 2912 80000 3024 0 FreeSans 448 0 0 0 simpleuart_div_we[2]
port 225 nsew signal tristate
flabel metal3 s 79200 4032 80000 4144 0 FreeSans 448 0 0 0 simpleuart_div_we[3]
port 226 nsew signal tristate
flabel metal3 s 79200 43232 80000 43344 0 FreeSans 448 0 0 0 simpleuart_reg_dat_do[0]
port 227 nsew signal input
flabel metal3 s 79200 54432 80000 54544 0 FreeSans 448 0 0 0 simpleuart_reg_dat_do[10]
port 228 nsew signal input
flabel metal3 s 79200 55552 80000 55664 0 FreeSans 448 0 0 0 simpleuart_reg_dat_do[11]
port 229 nsew signal input
flabel metal3 s 79200 56672 80000 56784 0 FreeSans 448 0 0 0 simpleuart_reg_dat_do[12]
port 230 nsew signal input
flabel metal3 s 79200 57792 80000 57904 0 FreeSans 448 0 0 0 simpleuart_reg_dat_do[13]
port 231 nsew signal input
flabel metal3 s 79200 58912 80000 59024 0 FreeSans 448 0 0 0 simpleuart_reg_dat_do[14]
port 232 nsew signal input
flabel metal3 s 79200 60032 80000 60144 0 FreeSans 448 0 0 0 simpleuart_reg_dat_do[15]
port 233 nsew signal input
flabel metal3 s 79200 61152 80000 61264 0 FreeSans 448 0 0 0 simpleuart_reg_dat_do[16]
port 234 nsew signal input
flabel metal3 s 79200 62272 80000 62384 0 FreeSans 448 0 0 0 simpleuart_reg_dat_do[17]
port 235 nsew signal input
flabel metal3 s 79200 63392 80000 63504 0 FreeSans 448 0 0 0 simpleuart_reg_dat_do[18]
port 236 nsew signal input
flabel metal3 s 79200 64512 80000 64624 0 FreeSans 448 0 0 0 simpleuart_reg_dat_do[19]
port 237 nsew signal input
flabel metal3 s 79200 44352 80000 44464 0 FreeSans 448 0 0 0 simpleuart_reg_dat_do[1]
port 238 nsew signal input
flabel metal3 s 79200 65632 80000 65744 0 FreeSans 448 0 0 0 simpleuart_reg_dat_do[20]
port 239 nsew signal input
flabel metal3 s 79200 66752 80000 66864 0 FreeSans 448 0 0 0 simpleuart_reg_dat_do[21]
port 240 nsew signal input
flabel metal3 s 79200 67872 80000 67984 0 FreeSans 448 0 0 0 simpleuart_reg_dat_do[22]
port 241 nsew signal input
flabel metal3 s 79200 68992 80000 69104 0 FreeSans 448 0 0 0 simpleuart_reg_dat_do[23]
port 242 nsew signal input
flabel metal3 s 79200 70112 80000 70224 0 FreeSans 448 0 0 0 simpleuart_reg_dat_do[24]
port 243 nsew signal input
flabel metal3 s 79200 71232 80000 71344 0 FreeSans 448 0 0 0 simpleuart_reg_dat_do[25]
port 244 nsew signal input
flabel metal3 s 79200 72352 80000 72464 0 FreeSans 448 0 0 0 simpleuart_reg_dat_do[26]
port 245 nsew signal input
flabel metal3 s 79200 73472 80000 73584 0 FreeSans 448 0 0 0 simpleuart_reg_dat_do[27]
port 246 nsew signal input
flabel metal3 s 79200 74592 80000 74704 0 FreeSans 448 0 0 0 simpleuart_reg_dat_do[28]
port 247 nsew signal input
flabel metal3 s 79200 75712 80000 75824 0 FreeSans 448 0 0 0 simpleuart_reg_dat_do[29]
port 248 nsew signal input
flabel metal3 s 79200 45472 80000 45584 0 FreeSans 448 0 0 0 simpleuart_reg_dat_do[2]
port 249 nsew signal input
flabel metal3 s 79200 76832 80000 76944 0 FreeSans 448 0 0 0 simpleuart_reg_dat_do[30]
port 250 nsew signal input
flabel metal3 s 79200 77952 80000 78064 0 FreeSans 448 0 0 0 simpleuart_reg_dat_do[31]
port 251 nsew signal input
flabel metal3 s 79200 46592 80000 46704 0 FreeSans 448 0 0 0 simpleuart_reg_dat_do[3]
port 252 nsew signal input
flabel metal3 s 79200 47712 80000 47824 0 FreeSans 448 0 0 0 simpleuart_reg_dat_do[4]
port 253 nsew signal input
flabel metal3 s 79200 48832 80000 48944 0 FreeSans 448 0 0 0 simpleuart_reg_dat_do[5]
port 254 nsew signal input
flabel metal3 s 79200 49952 80000 50064 0 FreeSans 448 0 0 0 simpleuart_reg_dat_do[6]
port 255 nsew signal input
flabel metal3 s 79200 51072 80000 51184 0 FreeSans 448 0 0 0 simpleuart_reg_dat_do[7]
port 256 nsew signal input
flabel metal3 s 79200 52192 80000 52304 0 FreeSans 448 0 0 0 simpleuart_reg_dat_do[8]
port 257 nsew signal input
flabel metal3 s 79200 53312 80000 53424 0 FreeSans 448 0 0 0 simpleuart_reg_dat_do[9]
port 258 nsew signal input
flabel metal3 s 79200 79072 80000 79184 0 FreeSans 448 0 0 0 simpleuart_reg_dat_wait
port 259 nsew signal input
flabel metal3 s 79200 5152 80000 5264 0 FreeSans 448 0 0 0 simpleuart_reg_div_do[0]
port 260 nsew signal input
flabel metal3 s 79200 16352 80000 16464 0 FreeSans 448 0 0 0 simpleuart_reg_div_do[10]
port 261 nsew signal input
flabel metal3 s 79200 17472 80000 17584 0 FreeSans 448 0 0 0 simpleuart_reg_div_do[11]
port 262 nsew signal input
flabel metal3 s 79200 18592 80000 18704 0 FreeSans 448 0 0 0 simpleuart_reg_div_do[12]
port 263 nsew signal input
flabel metal3 s 79200 19712 80000 19824 0 FreeSans 448 0 0 0 simpleuart_reg_div_do[13]
port 264 nsew signal input
flabel metal3 s 79200 20832 80000 20944 0 FreeSans 448 0 0 0 simpleuart_reg_div_do[14]
port 265 nsew signal input
flabel metal3 s 79200 21952 80000 22064 0 FreeSans 448 0 0 0 simpleuart_reg_div_do[15]
port 266 nsew signal input
flabel metal3 s 79200 23072 80000 23184 0 FreeSans 448 0 0 0 simpleuart_reg_div_do[16]
port 267 nsew signal input
flabel metal3 s 79200 24192 80000 24304 0 FreeSans 448 0 0 0 simpleuart_reg_div_do[17]
port 268 nsew signal input
flabel metal3 s 79200 25312 80000 25424 0 FreeSans 448 0 0 0 simpleuart_reg_div_do[18]
port 269 nsew signal input
flabel metal3 s 79200 26432 80000 26544 0 FreeSans 448 0 0 0 simpleuart_reg_div_do[19]
port 270 nsew signal input
flabel metal3 s 79200 6272 80000 6384 0 FreeSans 448 0 0 0 simpleuart_reg_div_do[1]
port 271 nsew signal input
flabel metal3 s 79200 27552 80000 27664 0 FreeSans 448 0 0 0 simpleuart_reg_div_do[20]
port 272 nsew signal input
flabel metal3 s 79200 28672 80000 28784 0 FreeSans 448 0 0 0 simpleuart_reg_div_do[21]
port 273 nsew signal input
flabel metal3 s 79200 29792 80000 29904 0 FreeSans 448 0 0 0 simpleuart_reg_div_do[22]
port 274 nsew signal input
flabel metal3 s 79200 30912 80000 31024 0 FreeSans 448 0 0 0 simpleuart_reg_div_do[23]
port 275 nsew signal input
flabel metal3 s 79200 32032 80000 32144 0 FreeSans 448 0 0 0 simpleuart_reg_div_do[24]
port 276 nsew signal input
flabel metal3 s 79200 33152 80000 33264 0 FreeSans 448 0 0 0 simpleuart_reg_div_do[25]
port 277 nsew signal input
flabel metal3 s 79200 34272 80000 34384 0 FreeSans 448 0 0 0 simpleuart_reg_div_do[26]
port 278 nsew signal input
flabel metal3 s 79200 35392 80000 35504 0 FreeSans 448 0 0 0 simpleuart_reg_div_do[27]
port 279 nsew signal input
flabel metal3 s 79200 36512 80000 36624 0 FreeSans 448 0 0 0 simpleuart_reg_div_do[28]
port 280 nsew signal input
flabel metal3 s 79200 37632 80000 37744 0 FreeSans 448 0 0 0 simpleuart_reg_div_do[29]
port 281 nsew signal input
flabel metal3 s 79200 7392 80000 7504 0 FreeSans 448 0 0 0 simpleuart_reg_div_do[2]
port 282 nsew signal input
flabel metal3 s 79200 38752 80000 38864 0 FreeSans 448 0 0 0 simpleuart_reg_div_do[30]
port 283 nsew signal input
flabel metal3 s 79200 39872 80000 39984 0 FreeSans 448 0 0 0 simpleuart_reg_div_do[31]
port 284 nsew signal input
flabel metal3 s 79200 8512 80000 8624 0 FreeSans 448 0 0 0 simpleuart_reg_div_do[3]
port 285 nsew signal input
flabel metal3 s 79200 9632 80000 9744 0 FreeSans 448 0 0 0 simpleuart_reg_div_do[4]
port 286 nsew signal input
flabel metal3 s 79200 10752 80000 10864 0 FreeSans 448 0 0 0 simpleuart_reg_div_do[5]
port 287 nsew signal input
flabel metal3 s 79200 11872 80000 11984 0 FreeSans 448 0 0 0 simpleuart_reg_div_do[6]
port 288 nsew signal input
flabel metal3 s 79200 12992 80000 13104 0 FreeSans 448 0 0 0 simpleuart_reg_div_do[7]
port 289 nsew signal input
flabel metal3 s 79200 14112 80000 14224 0 FreeSans 448 0 0 0 simpleuart_reg_div_do[8]
port 290 nsew signal input
flabel metal3 s 79200 15232 80000 15344 0 FreeSans 448 0 0 0 simpleuart_reg_div_do[9]
port 291 nsew signal input
flabel metal2 s 34048 79200 34160 80000 0 FreeSans 448 90 0 0 spimem_rdata[0]
port 292 nsew signal input
flabel metal2 s 40768 79200 40880 80000 0 FreeSans 448 90 0 0 spimem_rdata[10]
port 293 nsew signal input
flabel metal2 s 41440 79200 41552 80000 0 FreeSans 448 90 0 0 spimem_rdata[11]
port 294 nsew signal input
flabel metal2 s 42112 79200 42224 80000 0 FreeSans 448 90 0 0 spimem_rdata[12]
port 295 nsew signal input
flabel metal2 s 42784 79200 42896 80000 0 FreeSans 448 90 0 0 spimem_rdata[13]
port 296 nsew signal input
flabel metal2 s 43456 79200 43568 80000 0 FreeSans 448 90 0 0 spimem_rdata[14]
port 297 nsew signal input
flabel metal2 s 44128 79200 44240 80000 0 FreeSans 448 90 0 0 spimem_rdata[15]
port 298 nsew signal input
flabel metal2 s 44800 79200 44912 80000 0 FreeSans 448 90 0 0 spimem_rdata[16]
port 299 nsew signal input
flabel metal2 s 45472 79200 45584 80000 0 FreeSans 448 90 0 0 spimem_rdata[17]
port 300 nsew signal input
flabel metal2 s 46144 79200 46256 80000 0 FreeSans 448 90 0 0 spimem_rdata[18]
port 301 nsew signal input
flabel metal2 s 46816 79200 46928 80000 0 FreeSans 448 90 0 0 spimem_rdata[19]
port 302 nsew signal input
flabel metal2 s 34720 79200 34832 80000 0 FreeSans 448 90 0 0 spimem_rdata[1]
port 303 nsew signal input
flabel metal2 s 47488 79200 47600 80000 0 FreeSans 448 90 0 0 spimem_rdata[20]
port 304 nsew signal input
flabel metal2 s 48160 79200 48272 80000 0 FreeSans 448 90 0 0 spimem_rdata[21]
port 305 nsew signal input
flabel metal2 s 48832 79200 48944 80000 0 FreeSans 448 90 0 0 spimem_rdata[22]
port 306 nsew signal input
flabel metal2 s 49504 79200 49616 80000 0 FreeSans 448 90 0 0 spimem_rdata[23]
port 307 nsew signal input
flabel metal2 s 50176 79200 50288 80000 0 FreeSans 448 90 0 0 spimem_rdata[24]
port 308 nsew signal input
flabel metal2 s 50848 79200 50960 80000 0 FreeSans 448 90 0 0 spimem_rdata[25]
port 309 nsew signal input
flabel metal2 s 51520 79200 51632 80000 0 FreeSans 448 90 0 0 spimem_rdata[26]
port 310 nsew signal input
flabel metal2 s 52192 79200 52304 80000 0 FreeSans 448 90 0 0 spimem_rdata[27]
port 311 nsew signal input
flabel metal2 s 52864 79200 52976 80000 0 FreeSans 448 90 0 0 spimem_rdata[28]
port 312 nsew signal input
flabel metal2 s 53536 79200 53648 80000 0 FreeSans 448 90 0 0 spimem_rdata[29]
port 313 nsew signal input
flabel metal2 s 35392 79200 35504 80000 0 FreeSans 448 90 0 0 spimem_rdata[2]
port 314 nsew signal input
flabel metal2 s 54208 79200 54320 80000 0 FreeSans 448 90 0 0 spimem_rdata[30]
port 315 nsew signal input
flabel metal2 s 54880 79200 54992 80000 0 FreeSans 448 90 0 0 spimem_rdata[31]
port 316 nsew signal input
flabel metal2 s 36064 79200 36176 80000 0 FreeSans 448 90 0 0 spimem_rdata[3]
port 317 nsew signal input
flabel metal2 s 36736 79200 36848 80000 0 FreeSans 448 90 0 0 spimem_rdata[4]
port 318 nsew signal input
flabel metal2 s 37408 79200 37520 80000 0 FreeSans 448 90 0 0 spimem_rdata[5]
port 319 nsew signal input
flabel metal2 s 38080 79200 38192 80000 0 FreeSans 448 90 0 0 spimem_rdata[6]
port 320 nsew signal input
flabel metal2 s 38752 79200 38864 80000 0 FreeSans 448 90 0 0 spimem_rdata[7]
port 321 nsew signal input
flabel metal2 s 39424 79200 39536 80000 0 FreeSans 448 90 0 0 spimem_rdata[8]
port 322 nsew signal input
flabel metal2 s 40096 79200 40208 80000 0 FreeSans 448 90 0 0 spimem_rdata[9]
port 323 nsew signal input
flabel metal2 s 32704 79200 32816 80000 0 FreeSans 448 90 0 0 spimem_ready
port 324 nsew signal input
flabel metal2 s 33376 79200 33488 80000 0 FreeSans 448 90 0 0 spimem_valid
port 325 nsew signal tristate
flabel metal2 s 58240 79200 58352 80000 0 FreeSans 448 90 0 0 spimemio_cfgreg_do[0]
port 326 nsew signal input
flabel metal2 s 64960 79200 65072 80000 0 FreeSans 448 90 0 0 spimemio_cfgreg_do[10]
port 327 nsew signal input
flabel metal2 s 65632 79200 65744 80000 0 FreeSans 448 90 0 0 spimemio_cfgreg_do[11]
port 328 nsew signal input
flabel metal2 s 66304 79200 66416 80000 0 FreeSans 448 90 0 0 spimemio_cfgreg_do[12]
port 329 nsew signal input
flabel metal2 s 66976 79200 67088 80000 0 FreeSans 448 90 0 0 spimemio_cfgreg_do[13]
port 330 nsew signal input
flabel metal2 s 67648 79200 67760 80000 0 FreeSans 448 90 0 0 spimemio_cfgreg_do[14]
port 331 nsew signal input
flabel metal2 s 68320 79200 68432 80000 0 FreeSans 448 90 0 0 spimemio_cfgreg_do[15]
port 332 nsew signal input
flabel metal2 s 68992 79200 69104 80000 0 FreeSans 448 90 0 0 spimemio_cfgreg_do[16]
port 333 nsew signal input
flabel metal2 s 69664 79200 69776 80000 0 FreeSans 448 90 0 0 spimemio_cfgreg_do[17]
port 334 nsew signal input
flabel metal2 s 70336 79200 70448 80000 0 FreeSans 448 90 0 0 spimemio_cfgreg_do[18]
port 335 nsew signal input
flabel metal2 s 71008 79200 71120 80000 0 FreeSans 448 90 0 0 spimemio_cfgreg_do[19]
port 336 nsew signal input
flabel metal2 s 58912 79200 59024 80000 0 FreeSans 448 90 0 0 spimemio_cfgreg_do[1]
port 337 nsew signal input
flabel metal2 s 71680 79200 71792 80000 0 FreeSans 448 90 0 0 spimemio_cfgreg_do[20]
port 338 nsew signal input
flabel metal2 s 72352 79200 72464 80000 0 FreeSans 448 90 0 0 spimemio_cfgreg_do[21]
port 339 nsew signal input
flabel metal2 s 73024 79200 73136 80000 0 FreeSans 448 90 0 0 spimemio_cfgreg_do[22]
port 340 nsew signal input
flabel metal2 s 73696 79200 73808 80000 0 FreeSans 448 90 0 0 spimemio_cfgreg_do[23]
port 341 nsew signal input
flabel metal2 s 74368 79200 74480 80000 0 FreeSans 448 90 0 0 spimemio_cfgreg_do[24]
port 342 nsew signal input
flabel metal2 s 75040 79200 75152 80000 0 FreeSans 448 90 0 0 spimemio_cfgreg_do[25]
port 343 nsew signal input
flabel metal2 s 75712 79200 75824 80000 0 FreeSans 448 90 0 0 spimemio_cfgreg_do[26]
port 344 nsew signal input
flabel metal2 s 76384 79200 76496 80000 0 FreeSans 448 90 0 0 spimemio_cfgreg_do[27]
port 345 nsew signal input
flabel metal2 s 77056 79200 77168 80000 0 FreeSans 448 90 0 0 spimemio_cfgreg_do[28]
port 346 nsew signal input
flabel metal2 s 77728 79200 77840 80000 0 FreeSans 448 90 0 0 spimemio_cfgreg_do[29]
port 347 nsew signal input
flabel metal2 s 59584 79200 59696 80000 0 FreeSans 448 90 0 0 spimemio_cfgreg_do[2]
port 348 nsew signal input
flabel metal2 s 78400 79200 78512 80000 0 FreeSans 448 90 0 0 spimemio_cfgreg_do[30]
port 349 nsew signal input
flabel metal2 s 79072 79200 79184 80000 0 FreeSans 448 90 0 0 spimemio_cfgreg_do[31]
port 350 nsew signal input
flabel metal2 s 60256 79200 60368 80000 0 FreeSans 448 90 0 0 spimemio_cfgreg_do[3]
port 351 nsew signal input
flabel metal2 s 60928 79200 61040 80000 0 FreeSans 448 90 0 0 spimemio_cfgreg_do[4]
port 352 nsew signal input
flabel metal2 s 61600 79200 61712 80000 0 FreeSans 448 90 0 0 spimemio_cfgreg_do[5]
port 353 nsew signal input
flabel metal2 s 62272 79200 62384 80000 0 FreeSans 448 90 0 0 spimemio_cfgreg_do[6]
port 354 nsew signal input
flabel metal2 s 62944 79200 63056 80000 0 FreeSans 448 90 0 0 spimemio_cfgreg_do[7]
port 355 nsew signal input
flabel metal2 s 63616 79200 63728 80000 0 FreeSans 448 90 0 0 spimemio_cfgreg_do[8]
port 356 nsew signal input
flabel metal2 s 64288 79200 64400 80000 0 FreeSans 448 90 0 0 spimemio_cfgreg_do[9]
port 357 nsew signal input
flabel metal2 s 55552 79200 55664 80000 0 FreeSans 448 90 0 0 spimemio_cfgreg_we[0]
port 358 nsew signal tristate
flabel metal2 s 56224 79200 56336 80000 0 FreeSans 448 90 0 0 spimemio_cfgreg_we[1]
port 359 nsew signal tristate
flabel metal2 s 56896 79200 57008 80000 0 FreeSans 448 90 0 0 spimemio_cfgreg_we[2]
port 360 nsew signal tristate
flabel metal2 s 57568 79200 57680 80000 0 FreeSans 448 90 0 0 spimemio_cfgreg_we[3]
port 361 nsew signal tristate
flabel metal4 s 4448 3076 4768 76892 0 FreeSans 1280 90 0 0 vdd
port 362 nsew power bidirectional
flabel metal4 s 35168 3076 35488 76892 0 FreeSans 1280 90 0 0 vdd
port 362 nsew power bidirectional
flabel metal4 s 65888 3076 66208 76892 0 FreeSans 1280 90 0 0 vdd
port 362 nsew power bidirectional
flabel metal4 s 19808 3076 20128 76892 0 FreeSans 1280 90 0 0 vss
port 363 nsew ground bidirectional
flabel metal4 s 50528 3076 50848 76892 0 FreeSans 1280 90 0 0 vss
port 363 nsew ground bidirectional
rlabel metal1 39984 76048 39984 76048 0 vdd
rlabel metal1 39984 76832 39984 76832 0 vss
rlabel metal2 41664 24808 41664 24808 0 _0000_
rlabel metal3 16912 9240 16912 9240 0 _0001_
rlabel metal2 14560 9128 14560 9128 0 _0002_
rlabel metal2 15736 7896 15736 7896 0 _0003_
rlabel metal2 17416 5880 17416 5880 0 _0004_
rlabel metal2 17696 12040 17696 12040 0 _0005_
rlabel metal2 20440 13384 20440 13384 0 _0006_
rlabel metal2 19376 10696 19376 10696 0 _0007_
rlabel metal2 19600 7336 19600 7336 0 _0008_
rlabel metal3 24640 4200 24640 4200 0 _0009_
rlabel metal2 24024 5488 24024 5488 0 _0010_
rlabel metal3 23352 6664 23352 6664 0 _0011_
rlabel metal2 27496 8624 27496 8624 0 _0012_
rlabel metal2 22904 9408 22904 9408 0 _0013_
rlabel metal2 26488 11760 26488 11760 0 _0014_
rlabel metal2 22568 11760 22568 11760 0 _0015_
rlabel metal2 23296 11480 23296 11480 0 _0016_
rlabel metal2 30184 8624 30184 8624 0 _0017_
rlabel metal2 34216 10584 34216 10584 0 _0018_
rlabel metal2 30184 11760 30184 11760 0 _0019_
rlabel metal2 29176 10248 29176 10248 0 _0020_
rlabel metal2 35000 9520 35000 9520 0 _0021_
rlabel metal2 34104 4816 34104 4816 0 _0022_
rlabel metal2 31472 5656 31472 5656 0 _0023_
rlabel metal2 34552 6328 34552 6328 0 _0024_
rlabel metal3 28112 23016 28112 23016 0 _0025_
rlabel metal2 25032 24304 25032 24304 0 _0026_
rlabel metal2 28000 24024 28000 24024 0 _0027_
rlabel metal2 25144 22568 25144 22568 0 _0028_
rlabel metal2 17640 24304 17640 24304 0 _0029_
rlabel metal2 21784 24304 21784 24304 0 _0030_
rlabel metal2 17752 21784 17752 21784 0 _0031_
rlabel metal2 21784 22736 21784 22736 0 _0032_
rlabel metal2 20272 19320 20272 19320 0 _0033_
rlabel metal2 20664 18032 20664 18032 0 _0034_
rlabel metal2 22512 17752 22512 17752 0 _0035_
rlabel metal2 22848 19320 22848 19320 0 _0036_
rlabel metal2 27160 18592 27160 18592 0 _0037_
rlabel metal3 30856 17528 30856 17528 0 _0038_
rlabel metal2 28504 20328 28504 20328 0 _0039_
rlabel metal2 31528 20440 31528 20440 0 _0040_
rlabel metal2 35896 14896 35896 14896 0 _0041_
rlabel metal2 35224 12600 35224 12600 0 _0042_
rlabel metal2 33544 14168 33544 14168 0 _0043_
rlabel metal2 33544 15736 33544 15736 0 _0044_
rlabel metal2 26712 16464 26712 16464 0 _0045_
rlabel metal2 28168 16520 28168 16520 0 _0046_
rlabel metal2 25704 15232 25704 15232 0 _0047_
rlabel metal2 29792 15960 29792 15960 0 _0048_
rlabel metal2 40264 13328 40264 13328 0 _0049_
rlabel metal2 43176 13328 43176 13328 0 _0050_
rlabel metal2 42952 15148 42952 15148 0 _0051_
rlabel metal2 40040 15148 40040 15148 0 _0052_
rlabel metal2 39480 11032 39480 11032 0 _0053_
rlabel metal2 43512 9856 43512 9856 0 _0054_
rlabel metal2 38808 9352 38808 9352 0 _0055_
rlabel metal2 44072 9464 44072 9464 0 _0056_
rlabel metal2 37968 6664 37968 6664 0 _0057_
rlabel metal2 9352 8624 9352 8624 0 _0058_
rlabel metal2 9464 10192 9464 10192 0 _0059_
rlabel metal2 9800 11760 9800 11760 0 _0060_
rlabel metal2 13272 11424 13272 11424 0 _0061_
rlabel metal2 11144 7056 11144 7056 0 _0062_
rlabel metal2 10808 5488 10808 5488 0 _0063_
rlabel metal2 11816 4648 11816 4648 0 _0064_
rlabel metal2 15176 5264 15176 5264 0 _0065_
rlabel metal2 32088 6048 32088 6048 0 _0066_
rlabel metal2 29624 5096 29624 5096 0 _0067_
rlabel metal2 34776 6216 34776 6216 0 _0068_
rlabel metal3 25480 19096 25480 19096 0 _0069_
rlabel metal2 22568 20384 22568 20384 0 _0070_
rlabel metal2 25816 24024 25816 24024 0 _0071_
rlabel metal2 19992 22232 19992 22232 0 _0072_
rlabel metal2 23688 24024 23688 24024 0 _0073_
rlabel metal2 24192 23352 24192 23352 0 _0074_
rlabel metal2 25368 24976 25368 24976 0 _0075_
rlabel metal3 25760 23912 25760 23912 0 _0076_
rlabel metal2 24248 22456 24248 22456 0 _0077_
rlabel metal3 17584 21560 17584 21560 0 _0078_
rlabel metal2 19544 23520 19544 23520 0 _0079_
rlabel metal2 18200 23968 18200 23968 0 _0080_
rlabel metal3 21000 23912 21000 23912 0 _0081_
rlabel metal2 17528 22344 17528 22344 0 _0082_
rlabel metal3 20552 22344 20552 22344 0 _0083_
rlabel metal2 22008 19152 22008 19152 0 _0084_
rlabel metal2 19208 18368 19208 18368 0 _0085_
rlabel metal2 19768 19712 19768 19712 0 _0086_
rlabel metal3 19824 17640 19824 17640 0 _0087_
rlabel metal2 22008 17920 22008 17920 0 _0088_
rlabel metal3 21336 18984 21336 18984 0 _0089_
rlabel metal2 31640 18816 31640 18816 0 _0090_
rlabel metal2 25704 20720 25704 20720 0 _0091_
rlabel metal2 26880 19208 26880 19208 0 _0092_
rlabel metal2 26600 19040 26600 19040 0 _0093_
rlabel metal2 29064 20720 29064 20720 0 _0094_
rlabel metal2 30968 20048 30968 20048 0 _0095_
rlabel metal3 38724 13832 38724 13832 0 _0096_
rlabel metal3 34496 13944 34496 13944 0 _0097_
rlabel metal2 37128 12040 37128 12040 0 _0098_
rlabel metal3 31472 13720 31472 13720 0 _0099_
rlabel metal2 30968 14112 30968 14112 0 _0100_
rlabel metal2 34664 12264 34664 12264 0 _0101_
rlabel metal3 32480 13720 32480 13720 0 _0102_
rlabel metal2 32984 15204 32984 15204 0 _0103_
rlabel metal2 26824 15792 26824 15792 0 _0104_
rlabel metal3 29512 13832 29512 13832 0 _0105_
rlabel metal2 26376 15484 26376 15484 0 _0106_
rlabel metal2 28728 15596 28728 15596 0 _0107_
rlabel metal2 27272 14896 27272 14896 0 _0108_
rlabel metal2 28840 14224 28840 14224 0 _0109_
rlabel metal2 42952 14224 42952 14224 0 _0110_
rlabel metal2 39704 13608 39704 13608 0 _0111_
rlabel metal3 39424 13720 39424 13720 0 _0112_
rlabel metal3 41944 12376 41944 12376 0 _0113_
rlabel metal2 38584 14112 38584 14112 0 _0114_
rlabel metal2 39424 15288 39424 15288 0 _0115_
rlabel metal2 39592 11144 39592 11144 0 _0116_
rlabel metal3 36792 9800 36792 9800 0 _0117_
rlabel metal2 37464 10304 37464 10304 0 _0118_
rlabel metal3 39928 9632 39928 9632 0 _0119_
rlabel metal2 39368 9800 39368 9800 0 _0120_
rlabel metal3 44408 9800 44408 9800 0 _0121_
rlabel metal2 38248 7952 38248 7952 0 _0122_
rlabel metal3 20104 2408 20104 2408 0 _0123_
rlabel metal3 8792 6776 8792 6776 0 _0124_
rlabel metal2 9408 6888 9408 6888 0 _0125_
rlabel metal2 13384 9688 13384 9688 0 _0126_
rlabel metal2 11816 9968 11816 9968 0 _0127_
rlabel metal2 12376 10976 12376 10976 0 _0128_
rlabel metal3 10696 8120 10696 8120 0 _0129_
rlabel metal2 8344 8176 8344 8176 0 _0130_
rlabel metal3 10752 9688 10752 9688 0 _0131_
rlabel metal2 9016 9464 9016 9464 0 _0132_
rlabel metal3 10864 12040 10864 12040 0 _0133_
rlabel metal2 8792 7112 8792 7112 0 _0134_
rlabel metal2 13496 10696 13496 10696 0 _0135_
rlabel metal3 9576 4984 9576 4984 0 _0136_
rlabel metal2 7448 4536 7448 4536 0 _0137_
rlabel metal2 14168 6104 14168 6104 0 _0138_
rlabel metal3 13608 5096 13608 5096 0 _0139_
rlabel metal3 12712 6888 12712 6888 0 _0140_
rlabel metal2 8232 4872 8232 4872 0 _0141_
rlabel metal3 12264 5208 12264 5208 0 _0142_
rlabel metal3 10192 5096 10192 5096 0 _0143_
rlabel metal3 12208 5096 12208 5096 0 _0144_
rlabel metal2 13384 3864 13384 3864 0 _0145_
rlabel metal2 13776 3752 13776 3752 0 _0146_
rlabel metal2 47320 4984 47320 4984 0 _0147_
rlabel metal2 46648 5432 46648 5432 0 _0148_
rlabel metal3 43400 5992 43400 5992 0 _0149_
rlabel metal2 41384 3584 41384 3584 0 _0150_
rlabel metal2 43064 3472 43064 3472 0 _0151_
rlabel metal2 42504 3472 42504 3472 0 _0152_
rlabel metal2 44296 4032 44296 4032 0 _0153_
rlabel metal2 43736 3864 43736 3864 0 _0154_
rlabel metal2 33992 4200 33992 4200 0 _0155_
rlabel metal2 33656 3808 33656 3808 0 _0156_
rlabel metal2 42280 3864 42280 3864 0 _0157_
rlabel metal2 39256 4312 39256 4312 0 _0158_
rlabel metal2 36568 8344 36568 8344 0 _0159_
rlabel metal3 40880 3752 40880 3752 0 _0160_
rlabel metal2 43960 16352 43960 16352 0 _0161_
rlabel metal3 44464 15848 44464 15848 0 _0162_
rlabel metal2 41048 9072 41048 9072 0 _0163_
rlabel metal2 38920 5488 38920 5488 0 _0164_
rlabel metal2 40040 4928 40040 4928 0 _0165_
rlabel metal2 43736 20524 43736 20524 0 _0166_
rlabel metal2 42840 5096 42840 5096 0 _0167_
rlabel metal2 46424 16912 46424 16912 0 _0168_
rlabel metal2 44184 7280 44184 7280 0 _0169_
rlabel metal2 43120 8232 43120 8232 0 _0170_
rlabel metal2 43624 8512 43624 8512 0 _0171_
rlabel metal3 45304 17024 45304 17024 0 _0172_
rlabel metal2 43960 17752 43960 17752 0 _0173_
rlabel metal3 41720 7336 41720 7336 0 _0174_
rlabel metal2 44408 5152 44408 5152 0 _0175_
rlabel metal2 43064 7280 43064 7280 0 _0176_
rlabel metal2 42448 22344 42448 22344 0 _0177_
rlabel metal2 70840 18928 70840 18928 0 _0178_
rlabel metal2 74984 39536 74984 39536 0 _0179_
rlabel metal2 74088 41216 74088 41216 0 _0180_
rlabel metal2 51184 6664 51184 6664 0 _0181_
rlabel metal2 50792 6496 50792 6496 0 _0182_
rlabel metal3 48888 23184 48888 23184 0 _0183_
rlabel metal2 72128 41272 72128 41272 0 _0184_
rlabel metal2 74648 41440 74648 41440 0 _0185_
rlabel metal2 42056 9016 42056 9016 0 _0186_
rlabel metal2 74648 13048 74648 13048 0 _0187_
rlabel metal2 68376 40824 68376 40824 0 _0188_
rlabel metal2 61096 39984 61096 39984 0 _0189_
rlabel metal3 58072 41720 58072 41720 0 _0190_
rlabel metal2 55048 42336 55048 42336 0 _0191_
rlabel metal2 55832 41552 55832 41552 0 _0192_
rlabel metal2 57176 42448 57176 42448 0 _0193_
rlabel metal2 58072 42448 58072 42448 0 _0194_
rlabel metal2 72464 38920 72464 38920 0 _0195_
rlabel metal2 72856 39312 72856 39312 0 _0196_
rlabel metal3 73528 34720 73528 34720 0 _0197_
rlabel metal2 77224 4816 77224 4816 0 _0198_
rlabel metal2 77784 12432 77784 12432 0 _0199_
rlabel metal3 76608 3528 76608 3528 0 _0200_
rlabel metal2 77784 5768 77784 5768 0 _0201_
rlabel metal2 77000 4200 77000 4200 0 _0202_
rlabel metal3 33152 22344 33152 22344 0 _0203_
rlabel metal3 41440 20440 41440 20440 0 _0204_
rlabel metal2 39816 22736 39816 22736 0 _0205_
rlabel metal2 37352 21952 37352 21952 0 _0206_
rlabel metal2 74200 26600 74200 26600 0 _0207_
rlabel metal3 75768 23800 75768 23800 0 _0208_
rlabel metal2 76272 24136 76272 24136 0 _0209_
rlabel metal2 75432 25144 75432 25144 0 _0210_
rlabel metal3 44632 22624 44632 22624 0 _0211_
rlabel metal3 65800 38808 65800 38808 0 _0212_
rlabel metal2 63224 40040 63224 40040 0 _0213_
rlabel metal2 73304 26096 73304 26096 0 _0214_
rlabel metal3 68264 26152 68264 26152 0 _0215_
rlabel metal2 37352 18928 37352 18928 0 _0216_
rlabel metal3 36288 20664 36288 20664 0 _0217_
rlabel metal2 33992 20496 33992 20496 0 _0218_
rlabel metal2 45640 24584 45640 24584 0 _0219_
rlabel metal2 39032 20720 39032 20720 0 _0220_
rlabel metal3 36176 21560 36176 21560 0 _0221_
rlabel metal2 34440 22008 34440 22008 0 _0222_
rlabel metal2 34328 22736 34328 22736 0 _0223_
rlabel metal2 41832 24472 41832 24472 0 _0224_
rlabel metal3 35336 26936 35336 26936 0 _0225_
rlabel metal2 41888 25256 41888 25256 0 _0226_
rlabel metal3 35168 27048 35168 27048 0 _0227_
rlabel metal2 33544 23352 33544 23352 0 _0228_
rlabel metal2 28504 24024 28504 24024 0 _0229_
rlabel metal2 74816 27496 74816 27496 0 _0230_
rlabel metal3 75880 25480 75880 25480 0 _0231_
rlabel metal2 74200 25592 74200 25592 0 _0232_
rlabel metal2 35336 25312 35336 25312 0 _0233_
rlabel metal2 34888 20272 34888 20272 0 _0234_
rlabel metal2 36232 22344 36232 22344 0 _0235_
rlabel metal2 35112 24304 35112 24304 0 _0236_
rlabel metal2 35616 26600 35616 26600 0 _0237_
rlabel metal3 34216 24696 34216 24696 0 _0238_
rlabel metal2 72184 34160 72184 34160 0 _0239_
rlabel metal3 73192 34664 73192 34664 0 _0240_
rlabel metal3 74536 23912 74536 23912 0 _0241_
rlabel metal2 72296 23800 72296 23800 0 _0242_
rlabel metal2 36624 28392 36624 28392 0 _0243_
rlabel metal3 34608 20216 34608 20216 0 _0244_
rlabel metal2 35448 22176 35448 22176 0 _0245_
rlabel metal2 36008 24416 36008 24416 0 _0246_
rlabel metal2 35784 25480 35784 25480 0 _0247_
rlabel metal3 25592 23016 25592 23016 0 _0248_
rlabel metal2 71736 33376 71736 33376 0 _0249_
rlabel metal2 73080 25648 73080 25648 0 _0250_
rlabel metal2 76552 24416 76552 24416 0 _0251_
rlabel metal2 63336 41552 63336 41552 0 _0252_
rlabel metal3 67760 24920 67760 24920 0 _0253_
rlabel metal2 34944 27272 34944 27272 0 _0254_
rlabel metal2 33544 20384 33544 20384 0 _0255_
rlabel metal2 35224 20888 35224 20888 0 _0256_
rlabel metal2 35112 22680 35112 22680 0 _0257_
rlabel metal2 36344 21728 36344 21728 0 _0258_
rlabel metal2 19768 24136 19768 24136 0 _0259_
rlabel metal2 40488 24584 40488 24584 0 _0260_
rlabel metal2 64008 25032 64008 25032 0 _0261_
rlabel metal2 77168 23800 77168 23800 0 _0262_
rlabel metal2 63448 24136 63448 24136 0 _0263_
rlabel metal2 64344 40376 64344 40376 0 _0264_
rlabel metal2 62776 29988 62776 29988 0 _0265_
rlabel metal2 63336 24360 63336 24360 0 _0266_
rlabel metal2 35616 17640 35616 17640 0 _0267_
rlabel metal2 35112 17696 35112 17696 0 _0268_
rlabel metal2 35840 17640 35840 17640 0 _0269_
rlabel metal2 35336 17808 35336 17808 0 _0270_
rlabel metal2 38192 23688 38192 23688 0 _0271_
rlabel metal2 38808 25984 38808 25984 0 _0272_
rlabel metal2 37912 28224 37912 28224 0 _0273_
rlabel metal2 38080 25480 38080 25480 0 _0274_
rlabel metal2 40376 23800 40376 23800 0 _0275_
rlabel metal3 67256 34104 67256 34104 0 _0276_
rlabel metal2 63560 24248 63560 24248 0 _0277_
rlabel metal2 62888 26992 62888 26992 0 _0278_
rlabel metal2 43736 25424 43736 25424 0 _0279_
rlabel metal2 33936 17864 33936 17864 0 _0280_
rlabel metal2 39592 22568 39592 22568 0 _0281_
rlabel metal2 39480 24192 39480 24192 0 _0282_
rlabel metal2 38248 24864 38248 24864 0 _0283_
rlabel metal2 39256 21504 39256 21504 0 _0284_
rlabel metal2 71792 29512 71792 29512 0 _0285_
rlabel metal2 70952 32144 70952 32144 0 _0286_
rlabel metal3 72800 25480 72800 25480 0 _0287_
rlabel metal2 73864 24416 73864 24416 0 _0288_
rlabel metal3 67760 26264 67760 26264 0 _0289_
rlabel metal2 38920 25256 38920 25256 0 _0290_
rlabel metal3 35672 17528 35672 17528 0 _0291_
rlabel metal2 37240 19600 37240 19600 0 _0292_
rlabel metal2 37520 23688 37520 23688 0 _0293_
rlabel metal2 37464 22288 37464 22288 0 _0294_
rlabel metal2 39032 22176 39032 22176 0 _0295_
rlabel metal2 73304 30912 73304 30912 0 _0296_
rlabel metal2 71848 26180 71848 26180 0 _0297_
rlabel metal2 72184 25312 72184 25312 0 _0298_
rlabel metal2 65856 40376 65856 40376 0 _0299_
rlabel metal2 70504 25704 70504 25704 0 _0300_
rlabel metal3 43848 25200 43848 25200 0 _0301_
rlabel metal2 35784 15624 35784 15624 0 _0302_
rlabel metal2 41608 21336 41608 21336 0 _0303_
rlabel metal2 41384 22624 41384 22624 0 _0304_
rlabel metal3 39816 22232 39816 22232 0 _0305_
rlabel metal2 40768 16184 40768 16184 0 _0306_
rlabel metal3 42504 20776 42504 20776 0 _0307_
rlabel metal2 72072 26152 72072 26152 0 _0308_
rlabel metal3 75880 19992 75880 19992 0 _0309_
rlabel metal2 72184 20048 72184 20048 0 _0310_
rlabel metal2 66808 40768 66808 40768 0 _0311_
rlabel metal2 70952 21784 70952 21784 0 _0312_
rlabel metal3 49560 17136 49560 17136 0 _0313_
rlabel metal3 40320 17528 40320 17528 0 _0314_
rlabel metal2 39256 17528 39256 17528 0 _0315_
rlabel metal2 39816 18312 39816 18312 0 _0316_
rlabel metal2 40264 17360 40264 17360 0 _0317_
rlabel metal2 40656 17640 40656 17640 0 _0318_
rlabel metal3 41160 26936 41160 26936 0 _0319_
rlabel metal2 39928 26208 39928 26208 0 _0320_
rlabel metal2 41832 23464 41832 23464 0 _0321_
rlabel metal2 43400 19320 43400 19320 0 _0322_
rlabel metal4 71400 27272 71400 27272 0 _0323_
rlabel metal2 71624 21504 71624 21504 0 _0324_
rlabel metal3 67872 21784 67872 21784 0 _0325_
rlabel metal2 44968 17640 44968 17640 0 _0326_
rlabel metal2 39256 16352 39256 16352 0 _0327_
rlabel metal2 39592 16352 39592 16352 0 _0328_
rlabel metal2 42280 18144 42280 18144 0 _0329_
rlabel metal2 39816 25424 39816 25424 0 _0330_
rlabel metal2 43176 17808 43176 17808 0 _0331_
rlabel metal4 72744 29288 72744 29288 0 _0332_
rlabel metal2 72576 26712 72576 26712 0 _0333_
rlabel metal2 73080 20440 73080 20440 0 _0334_
rlabel metal3 69888 21560 69888 21560 0 _0335_
rlabel metal2 45080 17416 45080 17416 0 _0336_
rlabel metal2 38472 17304 38472 17304 0 _0337_
rlabel metal2 41384 17192 41384 17192 0 _0338_
rlabel metal2 41720 17360 41720 17360 0 _0339_
rlabel metal2 41496 21840 41496 21840 0 _0340_
rlabel metal2 41048 16968 41048 16968 0 _0341_
rlabel metal3 75320 26936 75320 26936 0 _0342_
rlabel metal2 73528 27440 73528 27440 0 _0343_
rlabel metal2 73192 23800 73192 23800 0 _0344_
rlabel metal2 73864 20496 73864 20496 0 _0345_
rlabel metal3 68152 37464 68152 37464 0 _0346_
rlabel metal2 69496 38920 69496 38920 0 _0347_
rlabel metal3 69720 20776 69720 20776 0 _0348_
rlabel metal2 40600 18928 40600 18928 0 _0349_
rlabel metal2 38584 16184 38584 16184 0 _0350_
rlabel metal2 39480 17360 39480 17360 0 _0351_
rlabel metal2 40824 19432 40824 19432 0 _0352_
rlabel metal2 41160 23744 41160 23744 0 _0353_
rlabel metal2 46648 19432 46648 19432 0 _0354_
rlabel metal2 46200 21616 46200 21616 0 _0355_
rlabel metal2 73304 22960 73304 22960 0 _0356_
rlabel metal2 77224 21896 77224 21896 0 _0357_
rlabel metal2 73640 22176 73640 22176 0 _0358_
rlabel metal2 68600 39200 68600 39200 0 _0359_
rlabel metal3 69944 22456 69944 22456 0 _0360_
rlabel metal2 41720 18984 41720 18984 0 _0361_
rlabel via2 39256 19320 39256 19320 0 _0362_
rlabel metal2 38808 18480 38808 18480 0 _0363_
rlabel metal2 39928 19600 39928 19600 0 _0364_
rlabel metal2 41608 18760 41608 18760 0 _0365_
rlabel metal2 44744 19208 44744 19208 0 _0366_
rlabel metal2 44968 25088 44968 25088 0 _0367_
rlabel metal2 44184 25088 44184 25088 0 _0368_
rlabel metal2 43512 22680 43512 22680 0 _0369_
rlabel metal2 47096 19544 47096 19544 0 _0370_
rlabel metal2 72912 23128 72912 23128 0 _0371_
rlabel metal2 73528 22624 73528 22624 0 _0372_
rlabel metal3 70616 23352 70616 23352 0 _0373_
rlabel metal2 45864 16240 45864 16240 0 _0374_
rlabel metal2 39032 19152 39032 19152 0 _0375_
rlabel metal2 39704 20188 39704 20188 0 _0376_
rlabel metal2 45416 18424 45416 18424 0 _0377_
rlabel metal2 44464 25144 44464 25144 0 _0378_
rlabel metal2 44184 22848 44184 22848 0 _0379_
rlabel metal2 75880 28224 75880 28224 0 _0380_
rlabel metal2 74984 22960 74984 22960 0 _0381_
rlabel metal3 76048 20552 76048 20552 0 _0382_
rlabel metal2 71736 22792 71736 22792 0 _0383_
rlabel metal2 47880 24248 47880 24248 0 _0384_
rlabel metal2 38024 18480 38024 18480 0 _0385_
rlabel metal2 43624 24024 43624 24024 0 _0386_
rlabel metal2 44016 23688 44016 23688 0 _0387_
rlabel metal2 46536 23352 46536 23352 0 _0388_
rlabel metal3 39480 21448 39480 21448 0 _0389_
rlabel metal2 76664 29008 76664 29008 0 _0390_
rlabel metal2 75992 24080 75992 24080 0 _0391_
rlabel metal2 76216 22624 76216 22624 0 _0392_
rlabel metal3 69944 39592 69944 39592 0 _0393_
rlabel metal2 68992 39704 68992 39704 0 _0394_
rlabel metal2 49392 23688 49392 23688 0 _0395_
rlabel metal3 36736 20104 36736 20104 0 _0396_
rlabel metal3 44856 23744 44856 23744 0 _0397_
rlabel metal2 45024 21560 45024 21560 0 _0398_
rlabel metal2 44072 22008 44072 22008 0 _0399_
rlabel metal2 48776 16800 48776 16800 0 _0400_
rlabel metal3 46872 15512 46872 15512 0 _0401_
rlabel metal2 49448 15680 49448 15680 0 _0402_
rlabel metal2 71232 27048 71232 27048 0 _0403_
rlabel metal3 78344 26824 78344 26824 0 _0404_
rlabel metal3 76104 26712 76104 26712 0 _0405_
rlabel metal2 71288 26600 71288 26600 0 _0406_
rlabel metal2 74200 38752 74200 38752 0 _0407_
rlabel metal2 71400 39200 71400 39200 0 _0408_
rlabel metal2 70616 28392 70616 28392 0 _0409_
rlabel metal2 47768 24248 47768 24248 0 _0410_
rlabel metal2 45864 26152 45864 26152 0 _0411_
rlabel metal2 46592 23912 46592 23912 0 _0412_
rlabel metal2 48048 20216 48048 20216 0 _0413_
rlabel metal2 46312 25256 46312 25256 0 _0414_
rlabel metal2 46760 23968 46760 23968 0 _0415_
rlabel metal2 47768 22176 47768 22176 0 _0416_
rlabel metal2 47488 21112 47488 21112 0 _0417_
rlabel metal2 49112 21840 49112 21840 0 _0418_
rlabel metal2 47544 17752 47544 17752 0 _0419_
rlabel metal2 47544 22960 47544 22960 0 _0420_
rlabel metal3 45752 20776 45752 20776 0 _0421_
rlabel metal2 46984 18088 46984 18088 0 _0422_
rlabel metal2 48776 13664 48776 13664 0 _0423_
rlabel metal3 73360 28056 73360 28056 0 _0424_
rlabel metal3 70952 27776 70952 27776 0 _0425_
rlabel metal2 70616 38668 70616 38668 0 _0426_
rlabel metal2 48104 22456 48104 22456 0 _0427_
rlabel metal3 46032 22232 46032 22232 0 _0428_
rlabel metal2 47992 22176 47992 22176 0 _0429_
rlabel metal2 47768 14840 47768 14840 0 _0430_
rlabel metal2 46312 14952 46312 14952 0 _0431_
rlabel metal3 50652 14280 50652 14280 0 _0432_
rlabel metal2 76216 31136 76216 31136 0 _0433_
rlabel metal2 71176 26096 71176 26096 0 _0434_
rlabel metal2 71400 25816 71400 25816 0 _0435_
rlabel metal2 69104 30744 69104 30744 0 _0436_
rlabel metal2 48048 23240 48048 23240 0 _0437_
rlabel metal2 46088 22624 46088 22624 0 _0438_
rlabel metal2 46424 22624 46424 22624 0 _0439_
rlabel metal3 49112 20328 49112 20328 0 _0440_
rlabel metal3 48272 15400 48272 15400 0 _0441_
rlabel metal2 49000 15848 49000 15848 0 _0442_
rlabel metal3 75936 30968 75936 30968 0 _0443_
rlabel metal3 75600 30184 75600 30184 0 _0444_
rlabel metal3 75936 27272 75936 27272 0 _0445_
rlabel metal2 71736 37744 71736 37744 0 _0446_
rlabel metal2 71848 33600 71848 33600 0 _0447_
rlabel metal3 49784 23688 49784 23688 0 _0448_
rlabel metal2 46088 23800 46088 23800 0 _0449_
rlabel metal2 47096 23744 47096 23744 0 _0450_
rlabel metal2 47824 21000 47824 21000 0 _0451_
rlabel metal2 47096 20524 47096 20524 0 _0452_
rlabel metal2 26600 16240 26600 16240 0 _0453_
rlabel metal2 51128 19544 51128 19544 0 _0454_
rlabel metal2 72688 29624 72688 29624 0 _0455_
rlabel metal3 76496 29176 76496 29176 0 _0456_
rlabel metal2 72856 28784 72856 28784 0 _0457_
rlabel metal2 73416 36736 73416 36736 0 _0458_
rlabel metal2 72408 29960 72408 29960 0 _0459_
rlabel metal2 49448 26432 49448 26432 0 _0460_
rlabel metal3 47208 26376 47208 26376 0 _0461_
rlabel metal2 47096 25984 47096 25984 0 _0462_
rlabel metal2 46872 25816 46872 25816 0 _0463_
rlabel metal2 49336 26432 49336 26432 0 _0464_
rlabel metal2 49504 26040 49504 26040 0 _0465_
rlabel metal2 48664 21168 48664 21168 0 _0466_
rlabel metal3 49616 20776 49616 20776 0 _0467_
rlabel metal2 49224 20356 49224 20356 0 _0468_
rlabel metal2 50008 17528 50008 17528 0 _0469_
rlabel metal2 73528 29792 73528 29792 0 _0470_
rlabel metal3 73752 29344 73752 29344 0 _0471_
rlabel metal2 73360 29624 73360 29624 0 _0472_
rlabel metal3 49504 26376 49504 26376 0 _0473_
rlabel metal3 45696 26264 45696 26264 0 _0474_
rlabel metal3 47656 26264 47656 26264 0 _0475_
rlabel metal2 48944 26040 48944 26040 0 _0476_
rlabel metal2 48888 20972 48888 20972 0 _0477_
rlabel metal2 47432 16688 47432 16688 0 _0478_
rlabel metal2 76776 32200 76776 32200 0 _0479_
rlabel metal3 75600 31528 75600 31528 0 _0480_
rlabel metal2 77336 29512 77336 29512 0 _0481_
rlabel metal2 73640 35784 73640 35784 0 _0482_
rlabel metal2 49280 26824 49280 26824 0 _0483_
rlabel metal2 47096 26992 47096 26992 0 _0484_
rlabel metal3 48216 27048 48216 27048 0 _0485_
rlabel metal2 49728 23912 49728 23912 0 _0486_
rlabel metal2 49336 19432 49336 19432 0 _0487_
rlabel metal3 43680 19712 43680 19712 0 _0488_
rlabel metal2 77112 33488 77112 33488 0 _0489_
rlabel metal2 74200 32928 74200 32928 0 _0490_
rlabel metal2 77448 30016 77448 30016 0 _0491_
rlabel metal2 74704 38808 74704 38808 0 _0492_
rlabel metal2 73696 32536 73696 32536 0 _0493_
rlabel metal3 50092 26936 50092 26936 0 _0494_
rlabel metal2 46200 27328 46200 27328 0 _0495_
rlabel metal2 49672 27104 49672 27104 0 _0496_
rlabel metal2 50008 25172 50008 25172 0 _0497_
rlabel metal2 50904 20776 50904 20776 0 _0498_
rlabel metal2 41272 14280 41272 14280 0 _0499_
rlabel metal3 53368 14728 53368 14728 0 _0500_
rlabel metal3 76328 33320 76328 33320 0 _0501_
rlabel metal2 73976 33992 73976 33992 0 _0502_
rlabel metal3 74368 33432 74368 33432 0 _0503_
rlabel metal2 75432 38976 75432 38976 0 _0504_
rlabel metal2 74480 35672 74480 35672 0 _0505_
rlabel metal3 55328 30184 55328 30184 0 _0506_
rlabel metal3 46872 31080 46872 31080 0 _0507_
rlabel metal2 45192 29848 45192 29848 0 _0508_
rlabel metal2 46648 31360 46648 31360 0 _0509_
rlabel metal3 48440 30184 48440 30184 0 _0510_
rlabel metal2 51520 19432 51520 19432 0 _0511_
rlabel metal2 51352 20384 51352 20384 0 _0512_
rlabel metal2 53256 19152 53256 19152 0 _0513_
rlabel metal2 52696 16744 52696 16744 0 _0514_
rlabel metal2 45416 14448 45416 14448 0 _0515_
rlabel metal2 75544 33264 75544 33264 0 _0516_
rlabel metal2 77672 30352 77672 30352 0 _0517_
rlabel metal3 75040 38248 75040 38248 0 _0518_
rlabel metal2 52360 31752 52360 31752 0 _0519_
rlabel metal2 44968 30352 44968 30352 0 _0520_
rlabel metal2 50568 30912 50568 30912 0 _0521_
rlabel metal2 51184 14616 51184 14616 0 _0522_
rlabel metal2 52808 16464 52808 16464 0 _0523_
rlabel metal3 44128 14504 44128 14504 0 _0524_
rlabel metal2 76552 37128 76552 37128 0 _0525_
rlabel metal2 76888 35056 76888 35056 0 _0526_
rlabel metal2 77672 32368 77672 32368 0 _0527_
rlabel metal2 75208 37072 75208 37072 0 _0528_
rlabel metal2 52864 31192 52864 31192 0 _0529_
rlabel metal3 45360 30968 45360 30968 0 _0530_
rlabel metal3 48664 30968 48664 30968 0 _0531_
rlabel metal2 51128 20552 51128 20552 0 _0532_
rlabel metal2 52360 19208 52360 19208 0 _0533_
rlabel metal3 40880 15288 40880 15288 0 _0534_
rlabel metal2 76216 38808 76216 38808 0 _0535_
rlabel metal2 76832 38248 76832 38248 0 _0536_
rlabel metal2 77896 32984 77896 32984 0 _0537_
rlabel metal2 76776 41272 76776 41272 0 _0538_
rlabel metal2 76608 36456 76608 36456 0 _0539_
rlabel metal2 52808 34272 52808 34272 0 _0540_
rlabel metal2 45976 31696 45976 31696 0 _0541_
rlabel metal3 48664 31752 48664 31752 0 _0542_
rlabel metal3 54544 13944 54544 13944 0 _0543_
rlabel metal3 53760 13832 53760 13832 0 _0544_
rlabel metal2 40264 11256 40264 11256 0 _0545_
rlabel metal2 53424 18536 53424 18536 0 _0546_
rlabel metal2 77336 36568 77336 36568 0 _0547_
rlabel metal2 77840 39480 77840 39480 0 _0548_
rlabel metal2 75544 36848 75544 36848 0 _0549_
rlabel metal2 77672 39928 77672 39928 0 _0550_
rlabel metal2 77224 40040 77224 40040 0 _0551_
rlabel metal2 54152 34776 54152 34776 0 _0552_
rlabel metal2 46200 35280 46200 35280 0 _0553_
rlabel metal2 45304 33824 45304 33824 0 _0554_
rlabel metal3 46816 34104 46816 34104 0 _0555_
rlabel metal2 46088 33656 46088 33656 0 _0556_
rlabel metal2 52360 22568 52360 22568 0 _0557_
rlabel metal3 55776 20664 55776 20664 0 _0558_
rlabel metal2 54152 20832 54152 20832 0 _0559_
rlabel metal2 53536 17528 53536 17528 0 _0560_
rlabel metal3 53284 11144 53284 11144 0 _0561_
rlabel metal3 77000 37464 77000 37464 0 _0562_
rlabel metal2 78008 37016 78008 37016 0 _0563_
rlabel metal2 77336 38668 77336 38668 0 _0564_
rlabel metal3 57960 35000 57960 35000 0 _0565_
rlabel metal2 46648 34832 46648 34832 0 _0566_
rlabel metal3 50400 34888 50400 34888 0 _0567_
rlabel metal2 53928 23044 53928 23044 0 _0568_
rlabel metal2 54152 19824 54152 19824 0 _0569_
rlabel metal2 41608 13608 41608 13608 0 _0570_
rlabel metal2 75320 39480 75320 39480 0 _0571_
rlabel metal3 76608 38920 76608 38920 0 _0572_
rlabel metal2 77112 41888 77112 41888 0 _0573_
rlabel metal3 76216 39368 76216 39368 0 _0574_
rlabel metal2 45752 35000 45752 35000 0 _0575_
rlabel metal2 46088 34944 46088 34944 0 _0576_
rlabel metal2 56840 17360 56840 17360 0 _0577_
rlabel metal2 55048 20664 55048 20664 0 _0578_
rlabel metal2 52920 10192 52920 10192 0 _0579_
rlabel metal2 73192 40040 73192 40040 0 _0580_
rlabel metal2 78008 39984 78008 39984 0 _0581_
rlabel metal2 73640 40488 73640 40488 0 _0582_
rlabel metal3 63616 40152 63616 40152 0 _0583_
rlabel metal3 45472 35672 45472 35672 0 _0584_
rlabel metal3 50008 35672 50008 35672 0 _0585_
rlabel metal3 56168 18424 56168 18424 0 _0586_
rlabel metal2 55720 19544 55720 19544 0 _0587_
rlabel metal2 75544 41552 75544 41552 0 _0588_
rlabel metal2 42280 7112 42280 7112 0 _0589_
rlabel metal2 29568 5992 29568 5992 0 _0590_
rlabel metal2 16240 4424 16240 4424 0 _0591_
rlabel metal3 13720 3304 13720 3304 0 _0592_
rlabel metal2 15624 7560 15624 7560 0 _0593_
rlabel metal2 30072 6160 30072 6160 0 _0594_
rlabel metal2 20104 6552 20104 6552 0 _0595_
rlabel metal2 18200 7056 18200 7056 0 _0596_
rlabel metal2 26544 7672 26544 7672 0 _0597_
rlabel metal3 18648 9240 18648 9240 0 _0598_
rlabel metal2 17808 9128 17808 9128 0 _0599_
rlabel metal2 11144 4816 11144 4816 0 _0600_
rlabel metal2 18536 9464 18536 9464 0 _0601_
rlabel metal3 15316 7448 15316 7448 0 _0602_
rlabel metal2 15848 7784 15848 7784 0 _0603_
rlabel metal2 15400 4760 15400 4760 0 _0604_
rlabel metal2 17808 5880 17808 5880 0 _0605_
rlabel metal2 16856 3752 16856 3752 0 _0606_
rlabel metal2 17976 6328 17976 6328 0 _0607_
rlabel metal2 19880 14336 19880 14336 0 _0608_
rlabel metal2 20552 8176 20552 8176 0 _0609_
rlabel metal2 18088 12936 18088 12936 0 _0610_
rlabel metal2 18648 6608 18648 6608 0 _0611_
rlabel metal2 20104 13552 20104 13552 0 _0612_
rlabel metal2 16744 6496 16744 6496 0 _0613_
rlabel metal2 19656 11368 19656 11368 0 _0614_
rlabel metal2 17864 4704 17864 4704 0 _0615_
rlabel metal2 19992 7504 19992 7504 0 _0616_
rlabel metal2 22456 6888 22456 6888 0 _0617_
rlabel metal3 23072 4984 23072 4984 0 _0618_
rlabel metal2 20328 3920 20328 3920 0 _0619_
rlabel metal2 27272 8120 27272 8120 0 _0620_
rlabel metal2 26040 7448 26040 7448 0 _0621_
rlabel metal2 26824 6384 26824 6384 0 _0622_
rlabel metal2 23352 4760 23352 4760 0 _0623_
rlabel metal2 21672 4704 21672 4704 0 _0624_
rlabel metal2 24136 6440 24136 6440 0 _0625_
rlabel metal2 23240 6664 23240 6664 0 _0626_
rlabel metal2 23576 6552 23576 6552 0 _0627_
rlabel metal2 21112 4424 21112 4424 0 _0628_
rlabel metal3 27160 8344 27160 8344 0 _0629_
rlabel metal2 22232 6216 22232 6216 0 _0630_
rlabel metal2 22680 8344 22680 8344 0 _0631_
rlabel metal2 26712 10136 26712 10136 0 _0632_
rlabel metal2 24696 9576 24696 9576 0 _0633_
rlabel metal2 25648 10696 25648 10696 0 _0634_
rlabel metal3 24192 10472 24192 10472 0 _0635_
rlabel metal2 21336 6832 21336 6832 0 _0636_
rlabel metal2 26600 10976 26600 10976 0 _0637_
rlabel metal2 21784 6888 21784 6888 0 _0638_
rlabel metal3 23800 11256 23800 11256 0 _0639_
rlabel metal2 22120 7056 22120 7056 0 _0640_
rlabel metal2 23408 11256 23408 11256 0 _0641_
rlabel metal2 29288 6160 29288 6160 0 _0642_
rlabel metal3 24752 5656 24752 5656 0 _0643_
rlabel metal2 25928 7280 25928 7280 0 _0644_
rlabel metal2 32200 7280 32200 7280 0 _0645_
rlabel metal2 32144 9576 32144 9576 0 _0646_
rlabel metal2 32648 11424 32648 11424 0 _0647_
rlabel metal2 30296 8400 30296 8400 0 _0648_
rlabel metal2 27608 6944 27608 6944 0 _0649_
rlabel metal3 33544 10024 33544 10024 0 _0650_
rlabel metal2 27160 8176 27160 8176 0 _0651_
rlabel metal3 31136 11256 31136 11256 0 _0652_
rlabel metal2 23128 4256 23128 4256 0 _0653_
rlabel metal3 31360 9688 31360 9688 0 _0654_
rlabel metal3 31696 7560 31696 7560 0 _0655_
rlabel metal2 32480 7336 32480 7336 0 _0656_
rlabel metal2 33432 7840 33432 7840 0 _0657_
rlabel metal2 35056 6552 35056 6552 0 _0658_
rlabel metal2 34664 9016 34664 9016 0 _0659_
rlabel metal2 30744 5040 30744 5040 0 _0660_
rlabel metal2 30968 5880 30968 5880 0 _0661_
rlabel metal3 31080 5768 31080 5768 0 _0662_
rlabel metal2 74200 2478 74200 2478 0 clk
rlabel metal2 24696 19936 24696 19936 0 clknet_0_clk
rlabel metal2 15400 10640 15400 10640 0 clknet_3_0__leaf_clk
rlabel metal3 19096 9016 19096 9016 0 clknet_3_1__leaf_clk
rlabel metal2 18648 18480 18648 18480 0 clknet_3_2__leaf_clk
rlabel metal2 25256 16856 25256 16856 0 clknet_3_3__leaf_clk
rlabel metal2 34552 7616 34552 7616 0 clknet_3_4__leaf_clk
rlabel metal2 42112 15288 42112 15288 0 clknet_3_5__leaf_clk
rlabel metal2 27888 23128 27888 23128 0 clknet_3_6__leaf_clk
rlabel metal2 40376 22848 40376 22848 0 clknet_3_7__leaf_clk
rlabel metal3 26740 5880 26740 5880 0 gpio\[16\]
rlabel metal2 26264 7000 26264 7000 0 gpio\[17\]
rlabel metal2 25816 9240 25816 9240 0 gpio\[18\]
rlabel metal2 26824 8624 26824 8624 0 gpio\[19\]
rlabel metal2 25984 12488 25984 12488 0 gpio\[20\]
rlabel metal2 26376 10808 26376 10808 0 gpio\[21\]
rlabel metal2 24696 12824 24696 12824 0 gpio\[22\]
rlabel metal2 25480 13272 25480 13272 0 gpio\[23\]
rlabel metal2 32424 10416 32424 10416 0 gpio\[24\]
rlabel metal2 41048 11928 41048 11928 0 gpio\[25\]
rlabel metal2 38360 13720 38360 13720 0 gpio\[26\]
rlabel metal2 39704 12152 39704 12152 0 gpio\[27\]
rlabel metal2 37128 8848 37128 8848 0 gpio\[28\]
rlabel metal3 33992 6608 33992 6608 0 gpio\[29\]
rlabel metal3 39704 9464 39704 9464 0 gpio\[30\]
rlabel metal2 37464 7280 37464 7280 0 gpio\[31\]
rlabel metal2 11256 76706 11256 76706 0 gpio_out[0]
rlabel metal2 19208 74928 19208 74928 0 gpio_out[10]
rlabel metal2 18648 77490 18648 77490 0 gpio_out[11]
rlabel metal2 19320 77882 19320 77882 0 gpio_out[12]
rlabel metal2 20216 75040 20216 75040 0 gpio_out[13]
rlabel metal3 21336 75880 21336 75880 0 gpio_out[14]
rlabel metal2 21336 77770 21336 77770 0 gpio_out[15]
rlabel metal2 11928 77714 11928 77714 0 gpio_out[1]
rlabel metal2 12600 77546 12600 77546 0 gpio_out[2]
rlabel metal2 12936 75600 12936 75600 0 gpio_out[3]
rlabel metal2 11592 75880 11592 75880 0 gpio_out[4]
rlabel metal2 14616 76202 14616 76202 0 gpio_out[5]
rlabel metal2 15288 77098 15288 77098 0 gpio_out[6]
rlabel metal2 15960 76762 15960 76762 0 gpio_out[7]
rlabel metal3 16016 76664 16016 76664 0 gpio_out[8]
rlabel metal2 17304 77546 17304 77546 0 gpio_out[9]
rlabel metal2 30856 22680 30856 22680 0 iomem_rdata\[0\]
rlabel metal3 25032 18312 25032 18312 0 iomem_rdata\[10\]
rlabel metal2 25256 20496 25256 20496 0 iomem_rdata\[11\]
rlabel metal2 29232 18312 29232 18312 0 iomem_rdata\[12\]
rlabel metal3 33040 18312 33040 18312 0 iomem_rdata\[13\]
rlabel metal2 30632 20272 30632 20272 0 iomem_rdata\[14\]
rlabel metal2 33656 21168 33656 21168 0 iomem_rdata\[15\]
rlabel metal3 38472 15176 38472 15176 0 iomem_rdata\[16\]
rlabel metal3 37128 13048 37128 13048 0 iomem_rdata\[17\]
rlabel metal2 34664 14224 34664 14224 0 iomem_rdata\[18\]
rlabel metal2 35504 16184 35504 16184 0 iomem_rdata\[19\]
rlabel metal2 27160 24696 27160 24696 0 iomem_rdata\[1\]
rlabel metal2 28336 16744 28336 16744 0 iomem_rdata\[20\]
rlabel metal2 31808 16744 31808 16744 0 iomem_rdata\[21\]
rlabel metal2 27832 14168 27832 14168 0 iomem_rdata\[22\]
rlabel metal2 32032 15400 32032 15400 0 iomem_rdata\[23\]
rlabel metal2 42392 13720 42392 13720 0 iomem_rdata\[24\]
rlabel metal2 44968 13664 44968 13664 0 iomem_rdata\[25\]
rlabel metal2 45080 15232 45080 15232 0 iomem_rdata\[26\]
rlabel metal2 41944 15288 41944 15288 0 iomem_rdata\[27\]
rlabel metal2 40376 11368 40376 11368 0 iomem_rdata\[28\]
rlabel metal2 44296 10864 44296 10864 0 iomem_rdata\[29\]
rlabel metal2 30072 24640 30072 24640 0 iomem_rdata\[2\]
rlabel metal2 40432 8904 40432 8904 0 iomem_rdata\[30\]
rlabel metal2 44632 9912 44632 9912 0 iomem_rdata\[31\]
rlabel metal2 27608 22400 27608 22400 0 iomem_rdata\[3\]
rlabel metal2 20104 24304 20104 24304 0 iomem_rdata\[4\]
rlabel metal2 23744 24584 23744 24584 0 iomem_rdata\[5\]
rlabel metal3 19936 22456 19936 22456 0 iomem_rdata\[6\]
rlabel metal2 23184 22456 23184 22456 0 iomem_rdata\[7\]
rlabel metal2 21784 21168 21784 21168 0 iomem_rdata\[8\]
rlabel metal2 21448 18704 21448 18704 0 iomem_rdata\[9\]
rlabel metal2 44296 7000 44296 7000 0 iomem_ready
rlabel metal2 26488 1246 26488 1246 0 mem_addr[0]
rlabel metal2 33208 2058 33208 2058 0 mem_addr[10]
rlabel metal2 26712 5320 26712 5320 0 mem_addr[11]
rlabel metal2 21560 5376 21560 5376 0 mem_addr[12]
rlabel metal2 21560 2940 21560 2940 0 mem_addr[13]
rlabel metal2 35896 2058 35896 2058 0 mem_addr[14]
rlabel metal2 25088 6440 25088 6440 0 mem_addr[15]
rlabel metal2 21056 4872 21056 4872 0 mem_addr[16]
rlabel metal2 37912 2058 37912 2058 0 mem_addr[17]
rlabel metal2 30800 3528 30800 3528 0 mem_addr[18]
rlabel metal2 39368 3304 39368 3304 0 mem_addr[19]
rlabel metal2 23688 4928 23688 4928 0 mem_addr[1]
rlabel metal2 40936 8736 40936 8736 0 mem_addr[20]
rlabel metal3 49728 3304 49728 3304 0 mem_addr[21]
rlabel metal2 41160 3864 41160 3864 0 mem_addr[22]
rlabel metal2 48552 3696 48552 3696 0 mem_addr[23]
rlabel metal2 42616 2058 42616 2058 0 mem_addr[24]
rlabel metal3 42616 4312 42616 4312 0 mem_addr[25]
rlabel metal2 51800 4480 51800 4480 0 mem_addr[26]
rlabel metal2 50568 3640 50568 3640 0 mem_addr[27]
rlabel metal2 45304 2058 45304 2058 0 mem_addr[28]
rlabel metal2 47992 5712 47992 5712 0 mem_addr[29]
rlabel metal2 22344 3864 22344 3864 0 mem_addr[2]
rlabel metal2 50904 5376 50904 5376 0 mem_addr[30]
rlabel metal2 47432 3304 47432 3304 0 mem_addr[31]
rlabel metal2 24808 4424 24808 4424 0 mem_addr[3]
rlabel metal2 29960 6216 29960 6216 0 mem_addr[4]
rlabel metal2 24360 5768 24360 5768 0 mem_addr[5]
rlabel metal3 23968 3304 23968 3304 0 mem_addr[6]
rlabel metal2 26152 4032 26152 4032 0 mem_addr[7]
rlabel metal2 23576 6216 23576 6216 0 mem_addr[8]
rlabel metal3 24360 3192 24360 3192 0 mem_addr[9]
rlabel metal2 52696 2422 52696 2422 0 mem_rdata[0]
rlabel metal2 59416 3206 59416 3206 0 mem_rdata[10]
rlabel metal2 60088 3598 60088 3598 0 mem_rdata[11]
rlabel metal2 60760 2982 60760 2982 0 mem_rdata[12]
rlabel metal2 61432 2254 61432 2254 0 mem_rdata[13]
rlabel metal2 62104 2310 62104 2310 0 mem_rdata[14]
rlabel metal2 62776 3598 62776 3598 0 mem_rdata[15]
rlabel metal2 63448 854 63448 854 0 mem_rdata[16]
rlabel metal2 64120 2422 64120 2422 0 mem_rdata[17]
rlabel metal3 71288 3528 71288 3528 0 mem_rdata[18]
rlabel metal2 68936 4648 68936 4648 0 mem_rdata[19]
rlabel metal2 53368 2198 53368 2198 0 mem_rdata[1]
rlabel metal2 66136 1694 66136 1694 0 mem_rdata[20]
rlabel metal2 68600 6216 68600 6216 0 mem_rdata[21]
rlabel metal2 67480 1974 67480 1974 0 mem_rdata[22]
rlabel metal2 68152 2814 68152 2814 0 mem_rdata[23]
rlabel metal2 68824 2422 68824 2422 0 mem_rdata[24]
rlabel metal2 69496 2254 69496 2254 0 mem_rdata[25]
rlabel metal2 70168 854 70168 854 0 mem_rdata[26]
rlabel metal2 70840 3206 70840 3206 0 mem_rdata[27]
rlabel metal2 71512 2086 71512 2086 0 mem_rdata[28]
rlabel metal2 72184 2926 72184 2926 0 mem_rdata[29]
rlabel metal2 54040 2534 54040 2534 0 mem_rdata[2]
rlabel metal2 72856 2982 72856 2982 0 mem_rdata[30]
rlabel metal2 73528 3038 73528 3038 0 mem_rdata[31]
rlabel metal2 54712 2422 54712 2422 0 mem_rdata[3]
rlabel metal2 55384 2142 55384 2142 0 mem_rdata[4]
rlabel metal2 56056 1526 56056 1526 0 mem_rdata[5]
rlabel metal2 56728 3206 56728 3206 0 mem_rdata[6]
rlabel metal2 57400 2086 57400 2086 0 mem_rdata[7]
rlabel metal2 58072 1190 58072 1190 0 mem_rdata[8]
rlabel metal2 58744 2814 58744 2814 0 mem_rdata[9]
rlabel metal2 49336 2422 49336 2422 0 mem_ready
rlabel metal2 48048 3080 48048 3080 0 mem_valid
rlabel metal2 4424 728 4424 728 0 mem_wdata[0]
rlabel metal2 10360 4648 10360 4648 0 mem_wdata[10]
rlabel metal2 8456 3864 8456 3864 0 mem_wdata[11]
rlabel metal2 13048 2058 13048 2058 0 mem_wdata[12]
rlabel metal2 13608 3080 13608 3080 0 mem_wdata[13]
rlabel metal2 14336 2072 14336 2072 0 mem_wdata[14]
rlabel metal2 15008 3192 15008 3192 0 mem_wdata[15]
rlabel metal2 15736 1246 15736 1246 0 mem_wdata[16]
rlabel metal2 10472 6776 10472 6776 0 mem_wdata[17]
rlabel metal4 15176 4144 15176 4144 0 mem_wdata[18]
rlabel metal2 17752 2086 17752 2086 0 mem_wdata[19]
rlabel metal2 5768 2856 5768 2856 0 mem_wdata[1]
rlabel metal2 15400 3920 15400 3920 0 mem_wdata[20]
rlabel metal2 18312 4592 18312 4592 0 mem_wdata[21]
rlabel metal2 19768 854 19768 854 0 mem_wdata[22]
rlabel metal2 19096 4424 19096 4424 0 mem_wdata[23]
rlabel metal2 17864 3920 17864 3920 0 mem_wdata[24]
rlabel metal2 21784 2058 21784 2058 0 mem_wdata[25]
rlabel metal2 18648 3808 18648 3808 0 mem_wdata[26]
rlabel metal2 23128 854 23128 854 0 mem_wdata[27]
rlabel metal2 23800 1246 23800 1246 0 mem_wdata[28]
rlabel metal2 22456 4424 22456 4424 0 mem_wdata[29]
rlabel metal2 4760 3472 4760 3472 0 mem_wdata[2]
rlabel metal2 21000 3584 21000 3584 0 mem_wdata[30]
rlabel metal2 21784 3584 21784 3584 0 mem_wdata[31]
rlabel metal2 6832 3192 6832 3192 0 mem_wdata[3]
rlabel metal2 6776 4088 6776 4088 0 mem_wdata[4]
rlabel metal2 5768 3584 5768 3584 0 mem_wdata[5]
rlabel metal2 6440 4200 6440 4200 0 mem_wdata[6]
rlabel metal2 7224 3248 7224 3248 0 mem_wdata[7]
rlabel metal2 8792 4368 8792 4368 0 mem_wdata[8]
rlabel metal2 7896 3696 7896 3696 0 mem_wdata[9]
rlabel metal2 50064 2968 50064 2968 0 mem_wstrb[0]
rlabel metal2 52360 3472 52360 3472 0 mem_wstrb[1]
rlabel metal2 53032 3584 53032 3584 0 mem_wstrb[2]
rlabel metal3 52864 3528 52864 3528 0 mem_wstrb[3]
rlabel metal2 25648 6552 25648 6552 0 net1
rlabel metal2 30968 3752 30968 3752 0 net10
rlabel metal3 2072 10976 2072 10976 0 net100
rlabel metal2 2128 12824 2128 12824 0 net101
rlabel metal2 76664 5936 76664 5936 0 net102
rlabel metal3 76664 43624 76664 43624 0 net103
rlabel metal2 77896 54544 77896 54544 0 net104
rlabel metal2 65296 40712 65296 40712 0 net105
rlabel metal3 75768 46872 75768 46872 0 net106
rlabel metal2 73808 28728 73808 28728 0 net107
rlabel metal3 76328 59080 76328 59080 0 net108
rlabel metal3 77112 60872 77112 60872 0 net109
rlabel metal2 37520 8008 37520 8008 0 net11
rlabel metal3 76552 61544 76552 61544 0 net110
rlabel metal3 77056 62216 77056 62216 0 net111
rlabel metal3 77056 64008 77056 64008 0 net112
rlabel metal3 77392 64680 77392 64680 0 net113
rlabel metal3 75992 45192 75992 45192 0 net114
rlabel metal3 77280 66024 77280 66024 0 net115
rlabel metal2 78288 61544 78288 61544 0 net116
rlabel metal3 77280 68488 77280 68488 0 net117
rlabel metal3 77336 69160 77336 69160 0 net118
rlabel metal3 78232 70952 78232 70952 0 net119
rlabel metal2 24080 4424 24080 4424 0 net12
rlabel metal3 73248 71848 73248 71848 0 net120
rlabel metal3 77000 72408 77000 72408 0 net121
rlabel metal2 76552 39144 76552 39144 0 net122
rlabel metal3 71624 73416 71624 73416 0 net123
rlabel metal2 78736 40264 78736 40264 0 net124
rlabel metal2 77784 45136 77784 45136 0 net125
rlabel metal2 76720 72632 76720 72632 0 net126
rlabel metal3 75936 72296 75936 72296 0 net127
rlabel metal3 78344 47208 78344 47208 0 net128
rlabel metal3 78232 48328 78232 48328 0 net129
rlabel metal2 38136 6552 38136 6552 0 net13
rlabel metal2 77560 47376 77560 47376 0 net130
rlabel metal2 77336 47824 77336 47824 0 net131
rlabel metal4 72072 41216 72072 41216 0 net132
rlabel metal3 76440 46984 76440 46984 0 net133
rlabel metal2 77896 53704 77896 53704 0 net134
rlabel metal2 46144 22120 46144 22120 0 net135
rlabel metal2 77224 7224 77224 7224 0 net136
rlabel metal2 77840 17080 77840 17080 0 net137
rlabel metal2 77896 17976 77896 17976 0 net138
rlabel metal2 77616 18648 77616 18648 0 net139
rlabel metal2 43624 4648 43624 4648 0 net14
rlabel metal2 77896 19096 77896 19096 0 net140
rlabel metal2 76776 21224 76776 21224 0 net141
rlabel metal2 77896 20440 77896 20440 0 net142
rlabel metal2 77896 22064 77896 22064 0 net143
rlabel metal2 75152 24920 75152 24920 0 net144
rlabel metal2 77840 23800 77840 23800 0 net145
rlabel metal2 76384 26824 76384 26824 0 net146
rlabel metal2 77896 6776 77896 6776 0 net147
rlabel metal2 77224 26768 77224 26768 0 net148
rlabel metal2 77896 26600 77896 26600 0 net149
rlabel metal2 40488 3332 40488 3332 0 net15
rlabel metal2 77840 28056 77840 28056 0 net150
rlabel metal2 77896 28728 77896 28728 0 net151
rlabel metal2 73752 32928 73752 32928 0 net152
rlabel metal2 77896 30856 77896 30856 0 net153
rlabel metal2 77952 31752 77952 31752 0 net154
rlabel metal2 75992 33488 75992 33488 0 net155
rlabel metal2 75152 36456 75152 36456 0 net156
rlabel metal2 78176 34776 78176 34776 0 net157
rlabel metal2 77224 8260 77224 8260 0 net158
rlabel metal2 77784 36344 77784 36344 0 net159
rlabel metal2 42000 5096 42000 5096 0 net16
rlabel metal2 78120 39704 78120 39704 0 net160
rlabel metal3 77168 9352 77168 9352 0 net161
rlabel metal3 78288 9576 78288 9576 0 net162
rlabel metal2 77168 15176 77168 15176 0 net163
rlabel metal2 78008 11256 78008 11256 0 net164
rlabel metal2 76944 24808 76944 24808 0 net165
rlabel metal3 77392 14392 77392 14392 0 net166
rlabel metal3 76664 15960 76664 15960 0 net167
rlabel metal2 34776 27552 34776 27552 0 net168
rlabel metal3 42224 26488 42224 26488 0 net169
rlabel metal2 25928 2464 25928 2464 0 net17
rlabel metal2 42280 43680 42280 43680 0 net170
rlabel metal2 42504 25872 42504 25872 0 net171
rlabel metal3 44184 26488 44184 26488 0 net172
rlabel metal2 44856 26096 44856 26096 0 net173
rlabel metal3 47376 24920 47376 24920 0 net174
rlabel metal2 45696 24248 45696 24248 0 net175
rlabel metal2 45696 25256 45696 25256 0 net176
rlabel metal4 47376 55440 47376 55440 0 net177
rlabel metal3 47880 20776 47880 20776 0 net178
rlabel metal3 34440 27832 34440 27832 0 net179
rlabel metal2 44296 7840 44296 7840 0 net18
rlabel metal2 50232 22960 50232 22960 0 net180
rlabel metal2 49448 21840 49448 21840 0 net181
rlabel metal2 48664 50624 48664 50624 0 net182
rlabel metal2 51800 22960 51800 22960 0 net183
rlabel metal2 50288 26824 50288 26824 0 net184
rlabel metal2 52528 55440 52528 55440 0 net185
rlabel metal2 53592 67200 53592 67200 0 net186
rlabel metal3 53760 22456 53760 22456 0 net187
rlabel metal3 55776 20104 55776 20104 0 net188
rlabel metal2 54488 71736 54488 71736 0 net189
rlabel metal2 47096 5040 47096 5040 0 net19
rlabel metal2 36288 31920 36288 31920 0 net190
rlabel metal3 54880 71512 54880 71512 0 net191
rlabel metal2 56224 67200 56224 67200 0 net192
rlabel metal3 36456 28056 36456 28056 0 net193
rlabel metal2 37576 28784 37576 28784 0 net194
rlabel metal2 39032 28504 39032 28504 0 net195
rlabel metal2 39088 75656 39088 75656 0 net196
rlabel metal2 37688 28280 37688 28280 0 net197
rlabel metal2 38864 74984 38864 74984 0 net198
rlabel metal2 40712 57484 40712 57484 0 net199
rlabel metal2 34104 7000 34104 7000 0 net2
rlabel metal2 46536 5824 46536 5824 0 net20
rlabel metal3 44296 22176 44296 22176 0 net200
rlabel metal3 60648 41272 60648 41272 0 net201
rlabel metal3 66248 75432 66248 75432 0 net202
rlabel metal3 67312 39368 67312 39368 0 net203
rlabel metal2 67480 71876 67480 71876 0 net204
rlabel metal2 69944 38528 69944 38528 0 net205
rlabel metal1 69608 77000 69608 77000 0 net206
rlabel metal2 69720 71876 69720 71876 0 net207
rlabel metal3 70896 67256 70896 67256 0 net208
rlabel metal2 71064 67480 71064 67480 0 net209
rlabel metal2 46088 7056 46088 7056 0 net21
rlabel metal2 71904 76552 71904 76552 0 net210
rlabel metal2 72688 76552 72688 76552 0 net211
rlabel metal3 61152 67256 61152 67256 0 net212
rlabel metal2 72912 67368 72912 67368 0 net213
rlabel metal2 73136 75432 73136 75432 0 net214
rlabel metal3 72688 36456 72688 36456 0 net215
rlabel metal2 74480 68040 74480 68040 0 net216
rlabel metal3 73696 68712 73696 68712 0 net217
rlabel metal2 75096 38864 75096 38864 0 net218
rlabel metal3 77000 37240 77000 37240 0 net219
rlabel metal2 46760 5880 46760 5880 0 net22
rlabel metal2 76440 41944 76440 41944 0 net220
rlabel metal2 77448 41272 77448 41272 0 net221
rlabel metal2 77896 49000 77896 49000 0 net222
rlabel metal2 61320 67480 61320 67480 0 net223
rlabel metal2 77112 42784 77112 42784 0 net224
rlabel metal3 74816 68824 74816 68824 0 net225
rlabel metal2 62552 41328 62552 41328 0 net226
rlabel metal2 62608 75432 62608 75432 0 net227
rlabel metal2 62496 76552 62496 76552 0 net228
rlabel metal3 64008 41944 64008 41944 0 net229
rlabel metal2 22680 2352 22680 2352 0 net23
rlabel metal2 64848 71624 64848 71624 0 net230
rlabel metal3 65072 67256 65072 67256 0 net231
rlabel metal2 65688 71876 65688 71876 0 net232
rlabel metal3 13552 73976 13552 73976 0 net233
rlabel metal2 17864 18648 17864 18648 0 net234
rlabel metal2 20328 75208 20328 75208 0 net235
rlabel metal3 18760 76440 18760 76440 0 net236
rlabel metal2 22792 74424 22792 74424 0 net237
rlabel metal2 23912 75488 23912 75488 0 net238
rlabel metal3 25592 75656 25592 75656 0 net239
rlabel metal3 47992 5880 47992 5880 0 net24
rlabel metal2 13944 72800 13944 72800 0 net240
rlabel metal2 12600 74200 12600 74200 0 net241
rlabel metal3 12600 74872 12600 74872 0 net242
rlabel metal3 13776 76328 13776 76328 0 net243
rlabel metal2 14056 73640 14056 73640 0 net244
rlabel metal3 15624 75656 15624 75656 0 net245
rlabel metal2 18256 43680 18256 43680 0 net246
rlabel metal2 20608 31920 20608 31920 0 net247
rlabel metal2 18312 74368 18312 74368 0 net248
rlabel metal2 52640 5768 52640 5768 0 net249
rlabel metal3 49168 6552 49168 6552 0 net25
rlabel metal2 59528 7448 59528 7448 0 net250
rlabel metal2 43120 20552 43120 20552 0 net251
rlabel metal2 46536 20776 46536 20776 0 net252
rlabel metal2 46872 18816 46872 18816 0 net253
rlabel metal2 45640 23352 45640 23352 0 net254
rlabel metal3 62384 6664 62384 6664 0 net255
rlabel metal2 64456 5992 64456 5992 0 net256
rlabel metal2 67424 4872 67424 4872 0 net257
rlabel metal2 69832 5656 69832 5656 0 net258
rlabel metal2 67368 5936 67368 5936 0 net259
rlabel metal2 25368 2800 25368 2800 0 net26
rlabel metal2 55384 8176 55384 8176 0 net260
rlabel metal2 67424 6440 67424 6440 0 net261
rlabel metal2 67032 7560 67032 7560 0 net262
rlabel metal2 68152 6664 68152 6664 0 net263
rlabel metal2 71064 4816 71064 4816 0 net264
rlabel metal2 72296 4256 72296 4256 0 net265
rlabel metal2 70504 4088 70504 4088 0 net266
rlabel metal2 71288 6272 71288 6272 0 net267
rlabel metal2 72296 5824 72296 5824 0 net268
rlabel metal2 70504 5656 70504 5656 0 net269
rlabel metal2 30352 7560 30352 7560 0 net27
rlabel metal2 72408 7504 72408 7504 0 net270
rlabel metal2 54152 5208 54152 5208 0 net271
rlabel metal3 74816 5880 74816 5880 0 net272
rlabel metal2 76328 7728 76328 7728 0 net273
rlabel metal3 42280 20216 42280 20216 0 net274
rlabel metal3 60256 3528 60256 3528 0 net275
rlabel metal2 39032 23688 39032 23688 0 net276
rlabel metal3 56504 5880 56504 5880 0 net277
rlabel metal2 40600 22288 40600 22288 0 net278
rlabel metal2 42840 20664 42840 20664 0 net279
rlabel metal3 28000 4424 28000 4424 0 net28
rlabel metal2 43960 19544 43960 19544 0 net280
rlabel metal2 43792 18200 43792 18200 0 net281
rlabel metal2 2856 45808 2856 45808 0 net282
rlabel metal3 4088 40376 4088 40376 0 net283
rlabel metal3 4872 40488 4872 40488 0 net284
rlabel metal3 3864 40600 3864 40600 0 net285
rlabel metal2 2744 43176 2744 43176 0 net286
rlabel metal2 3528 54040 3528 54040 0 net287
rlabel metal2 2072 55720 2072 55720 0 net288
rlabel metal2 3752 56560 3752 56560 0 net289
rlabel metal2 24024 3640 24024 3640 0 net29
rlabel metal2 4480 56728 4480 56728 0 net290
rlabel metal2 2072 58856 2072 58856 0 net291
rlabel metal2 2744 59696 2744 59696 0 net292
rlabel metal2 2072 61040 2072 61040 0 net293
rlabel metal2 3416 61880 3416 61880 0 net294
rlabel metal2 3192 63560 3192 63560 0 net295
rlabel metal2 3864 64400 3864 64400 0 net296
rlabel metal2 2072 44016 2072 44016 0 net297
rlabel metal2 4648 64736 4648 64736 0 net298
rlabel metal2 2072 66696 2072 66696 0 net299
rlabel metal2 38696 6552 38696 6552 0 net3
rlabel metal2 26488 3864 26488 3864 0 net30
rlabel metal2 3416 67536 3416 67536 0 net300
rlabel metal2 2072 68880 2072 68880 0 net301
rlabel metal2 2744 69720 2744 69720 0 net302
rlabel metal3 3584 71960 3584 71960 0 net303
rlabel metal2 3528 72240 3528 72240 0 net304
rlabel metal2 4312 73360 4312 73360 0 net305
rlabel metal2 4648 74032 4648 74032 0 net306
rlabel metal2 4592 75096 4592 75096 0 net307
rlabel metal2 2072 45360 2072 45360 0 net308
rlabel metal2 4648 75712 4648 75712 0 net309
rlabel metal2 28616 5208 28616 5208 0 net31
rlabel metal2 4200 75768 4200 75768 0 net310
rlabel metal2 3416 46200 3416 46200 0 net311
rlabel metal2 2072 47880 2072 47880 0 net312
rlabel metal2 2744 48720 2744 48720 0 net313
rlabel metal2 3416 49112 3416 49112 0 net314
rlabel metal2 2856 51016 2856 51016 0 net315
rlabel metal2 3528 51856 3528 51856 0 net316
rlabel metal3 3584 53592 3584 53592 0 net317
rlabel metal2 75320 42000 75320 42000 0 net318
rlabel metal2 78176 42504 78176 42504 0 net319
rlabel metal2 27160 3976 27160 3976 0 net32
rlabel metal3 76496 10024 76496 10024 0 net320
rlabel metal2 78344 3416 78344 3416 0 net321
rlabel metal2 77560 5656 77560 5656 0 net322
rlabel metal2 77336 5908 77336 5908 0 net323
rlabel metal2 42728 10080 42728 10080 0 net324
rlabel metal2 55832 44072 55832 44072 0 net325
rlabel metal2 56728 43232 56728 43232 0 net326
rlabel metal2 57624 75768 57624 75768 0 net327
rlabel metal3 59248 42840 59248 42840 0 net328
rlabel metal2 3640 64232 3640 64232 0 net329
rlabel metal2 40152 6048 40152 6048 0 net33
rlabel metal2 3080 67088 3080 67088 0 net330
rlabel metal2 2296 64064 2296 64064 0 net331
rlabel metal2 4424 41272 4424 41272 0 net332
rlabel metal2 2408 57680 2408 57680 0 net333
rlabel metal2 3864 53144 3864 53144 0 net334
rlabel metal2 2072 53480 2072 53480 0 net335
rlabel metal2 2688 48216 2688 48216 0 net336
rlabel metal2 3192 50456 3192 50456 0 net337
rlabel metal2 2632 45080 2632 45080 0 net338
rlabel metal2 4200 72072 4200 72072 0 net339
rlabel metal2 4312 4536 4312 4536 0 net34
rlabel metal2 5264 76552 5264 76552 0 net340
rlabel metal3 5152 71848 5152 71848 0 net341
rlabel metal2 1904 71624 1904 71624 0 net342
rlabel metal3 21560 76664 21560 76664 0 net343
rlabel metal2 23128 76160 23128 76160 0 net344
rlabel metal2 23464 75096 23464 75096 0 net345
rlabel metal2 24136 75544 24136 75544 0 net346
rlabel metal2 24808 76664 24808 76664 0 net347
rlabel metal2 25480 76664 25480 76664 0 net348
rlabel metal2 26152 76664 26152 76664 0 net349
rlabel metal2 11536 3528 11536 3528 0 net35
rlabel metal2 26712 77938 26712 77938 0 net350
rlabel metal2 27496 76664 27496 76664 0 net351
rlabel metal2 28392 77280 28392 77280 0 net352
rlabel metal2 28840 76664 28840 76664 0 net353
rlabel metal2 29512 76664 29512 76664 0 net354
rlabel metal2 30184 76664 30184 76664 0 net355
rlabel metal2 30856 76664 30856 76664 0 net356
rlabel metal2 31472 76664 31472 76664 0 net357
rlabel metal2 32200 76664 32200 76664 0 net358
rlabel metal2 8792 3248 8792 3248 0 net36
rlabel metal2 17864 5320 17864 5320 0 net37
rlabel metal2 18816 5096 18816 5096 0 net38
rlabel metal2 9912 3864 9912 3864 0 net39
rlabel metal2 27832 3080 27832 3080 0 net4
rlabel metal2 17528 3976 17528 3976 0 net40
rlabel metal2 20328 4368 20328 4368 0 net41
rlabel metal2 21784 4200 21784 4200 0 net42
rlabel metal2 14392 2800 14392 2800 0 net43
rlabel metal2 20888 4088 20888 4088 0 net44
rlabel metal2 6272 4536 6272 4536 0 net45
rlabel metal2 15904 3416 15904 3416 0 net46
rlabel metal2 18816 4536 18816 4536 0 net47
rlabel metal2 17472 3416 17472 3416 0 net48
rlabel metal2 19376 4536 19376 4536 0 net49
rlabel metal2 28952 3136 28952 3136 0 net5
rlabel metal2 18144 3416 18144 3416 0 net50
rlabel metal2 27496 3164 27496 3164 0 net51
rlabel metal2 18872 2296 18872 2296 0 net52
rlabel metal3 21280 3528 21280 3528 0 net53
rlabel metal2 20440 7280 20440 7280 0 net54
rlabel metal2 22680 4648 22680 4648 0 net55
rlabel metal2 4984 4368 4984 4368 0 net56
rlabel metal2 21336 2464 21336 2464 0 net57
rlabel metal2 22456 5040 22456 5040 0 net58
rlabel metal2 6776 5432 6776 5432 0 net59
rlabel metal2 35728 8008 35728 8008 0 net6
rlabel metal2 7336 4368 7336 4368 0 net60
rlabel metal2 6104 3864 6104 3864 0 net61
rlabel metal2 6832 3416 6832 3416 0 net62
rlabel metal2 7448 3752 7448 3752 0 net63
rlabel metal2 15288 5656 15288 5656 0 net64
rlabel metal2 10920 3472 10920 3472 0 net65
rlabel metal2 51240 3360 51240 3360 0 net66
rlabel metal2 51016 5544 51016 5544 0 net67
rlabel metal2 51576 6384 51576 6384 0 net68
rlabel metal2 53480 5712 53480 5712 0 net69
rlabel metal2 29624 4032 29624 4032 0 net7
rlabel metal2 2744 5096 2744 5096 0 net70
rlabel metal2 38360 16240 38360 16240 0 net71
rlabel metal3 20272 15400 20272 15400 0 net72
rlabel metal2 2072 16128 2072 16128 0 net73
rlabel metal2 2072 17248 2072 17248 0 net74
rlabel metal2 2072 18200 2072 18200 0 net75
rlabel metal2 2072 19712 2072 19712 0 net76
rlabel metal2 2128 20664 2128 20664 0 net77
rlabel metal2 2072 22176 2072 22176 0 net78
rlabel metal2 2072 23072 2072 23072 0 net79
rlabel metal2 38696 3976 38696 3976 0 net8
rlabel metal2 2072 23912 2072 23912 0 net80
rlabel metal2 2072 4088 2072 4088 0 net81
rlabel metal2 2128 25368 2128 25368 0 net82
rlabel metal2 44408 26600 44408 26600 0 net83
rlabel metal2 2072 27272 2072 27272 0 net84
rlabel metal2 2072 28560 2072 28560 0 net85
rlabel metal2 44968 29512 44968 29512 0 net86
rlabel metal2 26936 30576 26936 30576 0 net87
rlabel metal2 44296 31360 44296 31360 0 net88
rlabel metal2 28504 32368 28504 32368 0 net89
rlabel metal2 36568 5432 36568 5432 0 net9
rlabel metal2 2072 33768 2072 33768 0 net90
rlabel metal2 45192 34720 45192 34720 0 net91
rlabel metal2 2072 5376 2072 5376 0 net92
rlabel metal2 44744 36064 44744 36064 0 net93
rlabel metal2 26936 36848 26936 36848 0 net94
rlabel metal2 2016 6104 2016 6104 0 net95
rlabel metal2 34664 17192 34664 17192 0 net96
rlabel metal2 2072 8260 2072 8260 0 net97
rlabel metal2 2072 9856 2072 9856 0 net98
rlabel metal2 2128 10808 2128 10808 0 net99
rlabel metal3 2086 38136 2086 38136 0 ram_gwenb[0]
rlabel metal3 1358 39256 1358 39256 0 ram_gwenb[1]
rlabel metal3 1358 40376 1358 40376 0 ram_gwenb[2]
rlabel metal3 1358 41496 1358 41496 0 ram_gwenb[3]
rlabel metal2 2408 2856 2408 2856 0 ram_rdata[0]
rlabel metal2 1736 13608 1736 13608 0 ram_rdata[10]
rlabel metal2 1736 14952 1736 14952 0 ram_rdata[11]
rlabel metal2 1736 15848 1736 15848 0 ram_rdata[12]
rlabel metal2 1736 17192 1736 17192 0 ram_rdata[13]
rlabel metal2 1736 18200 1736 18200 0 ram_rdata[14]
rlabel metal3 1246 19096 1246 19096 0 ram_rdata[15]
rlabel metal2 1736 20384 1736 20384 0 ram_rdata[16]
rlabel metal2 1736 21448 1736 21448 0 ram_rdata[17]
rlabel metal2 1736 22792 1736 22792 0 ram_rdata[18]
rlabel metal2 1736 23688 1736 23688 0 ram_rdata[19]
rlabel metal3 1246 3416 1246 3416 0 ram_rdata[1]
rlabel metal2 1736 24976 1736 24976 0 ram_rdata[20]
rlabel metal2 1736 26040 1736 26040 0 ram_rdata[21]
rlabel metal3 1246 26936 1246 26936 0 ram_rdata[22]
rlabel metal2 1736 28336 1736 28336 0 ram_rdata[23]
rlabel metal2 1736 29288 1736 29288 0 ram_rdata[24]
rlabel metal2 1736 30632 1736 30632 0 ram_rdata[25]
rlabel metal2 1736 31528 1736 31528 0 ram_rdata[26]
rlabel metal2 1736 32816 1736 32816 0 ram_rdata[27]
rlabel metal2 1736 33880 1736 33880 0 ram_rdata[28]
rlabel metal3 1246 34776 1246 34776 0 ram_rdata[29]
rlabel metal2 1736 4816 1736 4816 0 ram_rdata[2]
rlabel metal2 1736 36120 1736 36120 0 ram_rdata[30]
rlabel metal2 1736 37128 1736 37128 0 ram_rdata[31]
rlabel metal2 1736 5768 1736 5768 0 ram_rdata[3]
rlabel metal2 1736 7112 1736 7112 0 ram_rdata[4]
rlabel metal2 1736 8008 1736 8008 0 ram_rdata[5]
rlabel metal2 1736 9352 1736 9352 0 ram_rdata[6]
rlabel metal2 1736 10360 1736 10360 0 ram_rdata[7]
rlabel metal3 1246 11256 1246 11256 0 ram_rdata[8]
rlabel metal2 1736 12600 1736 12600 0 ram_rdata[9]
rlabel metal2 43848 23464 43848 23464 0 ram_ready
rlabel metal3 1358 42616 1358 42616 0 ram_wenb[0]
rlabel metal3 1358 53816 1358 53816 0 ram_wenb[10]
rlabel metal3 1750 54936 1750 54936 0 ram_wenb[11]
rlabel metal3 1358 56056 1358 56056 0 ram_wenb[12]
rlabel metal3 1358 57176 1358 57176 0 ram_wenb[13]
rlabel metal3 1750 58296 1750 58296 0 ram_wenb[14]
rlabel metal3 1358 59416 1358 59416 0 ram_wenb[15]
rlabel metal3 1750 60536 1750 60536 0 ram_wenb[16]
rlabel metal3 1358 61656 1358 61656 0 ram_wenb[17]
rlabel metal3 1358 62776 1358 62776 0 ram_wenb[18]
rlabel metal3 1358 63896 1358 63896 0 ram_wenb[19]
rlabel metal3 854 43736 854 43736 0 ram_wenb[1]
rlabel metal3 1358 65016 1358 65016 0 ram_wenb[20]
rlabel metal3 1750 66136 1750 66136 0 ram_wenb[21]
rlabel metal3 1358 67256 1358 67256 0 ram_wenb[22]
rlabel metal3 1750 68376 1750 68376 0 ram_wenb[23]
rlabel metal3 1358 69496 1358 69496 0 ram_wenb[24]
rlabel metal3 1358 70616 1358 70616 0 ram_wenb[25]
rlabel metal3 1358 71736 1358 71736 0 ram_wenb[26]
rlabel metal3 1358 72856 1358 72856 0 ram_wenb[27]
rlabel metal3 1358 73976 1358 73976 0 ram_wenb[28]
rlabel metal3 1358 75096 1358 75096 0 ram_wenb[29]
rlabel metal3 1750 44856 1750 44856 0 ram_wenb[2]
rlabel metal3 1358 76216 1358 76216 0 ram_wenb[30]
rlabel metal3 1470 77336 1470 77336 0 ram_wenb[31]
rlabel metal3 1358 45976 1358 45976 0 ram_wenb[3]
rlabel metal3 1750 47096 1750 47096 0 ram_wenb[4]
rlabel metal3 1358 48216 1358 48216 0 ram_wenb[5]
rlabel metal3 1358 49336 1358 49336 0 ram_wenb[6]
rlabel metal3 1358 50456 1358 50456 0 ram_wenb[7]
rlabel metal3 1358 51576 1358 51576 0 ram_wenb[8]
rlabel metal3 1358 52696 1358 52696 0 ram_wenb[9]
rlabel metal3 75656 5096 75656 5096 0 resetn
rlabel metal2 78008 42000 78008 42000 0 simpleuart_dat_re
rlabel metal2 76552 40768 76552 40768 0 simpleuart_dat_we
rlabel metal3 76762 728 76762 728 0 simpleuart_div_we[0]
rlabel metal3 75992 7224 75992 7224 0 simpleuart_div_we[1]
rlabel metal3 73976 4984 73976 4984 0 simpleuart_div_we[2]
rlabel metal3 75208 7560 75208 7560 0 simpleuart_div_we[3]
rlabel metal2 78232 43400 78232 43400 0 simpleuart_reg_dat_do[0]
rlabel metal2 78232 54824 78232 54824 0 simpleuart_reg_dat_do[10]
rlabel metal2 78232 55832 78232 55832 0 simpleuart_reg_dat_do[11]
rlabel metal3 78722 56728 78722 56728 0 simpleuart_reg_dat_do[12]
rlabel metal2 78232 58016 78232 58016 0 simpleuart_reg_dat_do[13]
rlabel metal2 78232 59080 78232 59080 0 simpleuart_reg_dat_do[14]
rlabel metal2 78232 60424 78232 60424 0 simpleuart_reg_dat_do[15]
rlabel metal2 78232 61264 78232 61264 0 simpleuart_reg_dat_do[16]
rlabel metal2 78232 62664 78232 62664 0 simpleuart_reg_dat_do[17]
rlabel metal2 78232 63672 78232 63672 0 simpleuart_reg_dat_do[18]
rlabel metal3 78722 64568 78722 64568 0 simpleuart_reg_dat_do[19]
rlabel metal2 78232 44744 78232 44744 0 simpleuart_reg_dat_do[1]
rlabel metal2 78232 65856 78232 65856 0 simpleuart_reg_dat_do[20]
rlabel metal2 78232 66920 78232 66920 0 simpleuart_reg_dat_do[21]
rlabel metal2 78232 68264 78232 68264 0 simpleuart_reg_dat_do[22]
rlabel metal2 78232 69104 78232 69104 0 simpleuart_reg_dat_do[23]
rlabel metal2 78232 70448 78232 70448 0 simpleuart_reg_dat_do[24]
rlabel metal2 78232 71512 78232 71512 0 simpleuart_reg_dat_do[25]
rlabel metal3 78722 72408 78722 72408 0 simpleuart_reg_dat_do[26]
rlabel metal3 78834 73528 78834 73528 0 simpleuart_reg_dat_do[27]
rlabel metal2 78288 73528 78288 73528 0 simpleuart_reg_dat_do[28]
rlabel metal2 78176 75544 78176 75544 0 simpleuart_reg_dat_do[29]
rlabel metal2 78232 45640 78232 45640 0 simpleuart_reg_dat_do[2]
rlabel metal2 76944 75096 76944 75096 0 simpleuart_reg_dat_do[30]
rlabel metal3 78512 75096 78512 75096 0 simpleuart_reg_dat_do[31]
rlabel metal2 78232 46984 78232 46984 0 simpleuart_reg_dat_do[3]
rlabel metal2 78232 47992 78232 47992 0 simpleuart_reg_dat_do[4]
rlabel metal3 78722 48888 78722 48888 0 simpleuart_reg_dat_do[5]
rlabel metal2 78232 50232 78232 50232 0 simpleuart_reg_dat_do[6]
rlabel metal2 78232 51240 78232 51240 0 simpleuart_reg_dat_do[7]
rlabel metal2 78232 52584 78232 52584 0 simpleuart_reg_dat_do[8]
rlabel metal2 78232 53480 78232 53480 0 simpleuart_reg_dat_do[9]
rlabel metal2 77336 77896 77336 77896 0 simpleuart_reg_dat_wait
rlabel metal2 77616 6552 77616 6552 0 simpleuart_reg_div_do[0]
rlabel metal2 78232 16632 78232 16632 0 simpleuart_reg_div_do[10]
rlabel metal3 78722 17528 78722 17528 0 simpleuart_reg_div_do[11]
rlabel metal2 77336 18536 77336 18536 0 simpleuart_reg_div_do[12]
rlabel metal2 78232 19096 78232 19096 0 simpleuart_reg_div_do[13]
rlabel metal2 74872 21224 74872 21224 0 simpleuart_reg_div_do[14]
rlabel metal2 78120 21000 78120 21000 0 simpleuart_reg_div_do[15]
rlabel metal2 78232 22400 78232 22400 0 simpleuart_reg_div_do[16]
rlabel metal2 74648 24472 74648 24472 0 simpleuart_reg_div_do[17]
rlabel metal2 78232 23744 78232 23744 0 simpleuart_reg_div_do[18]
rlabel metal2 76776 25984 76776 25984 0 simpleuart_reg_div_do[19]
rlabel metal2 78344 6216 78344 6216 0 simpleuart_reg_div_do[1]
rlabel metal2 77672 26376 77672 26376 0 simpleuart_reg_div_do[20]
rlabel metal2 78232 26208 78232 26208 0 simpleuart_reg_div_do[21]
rlabel metal2 76496 22456 76496 22456 0 simpleuart_reg_div_do[22]
rlabel metal2 71288 28896 71288 28896 0 simpleuart_reg_div_do[23]
rlabel metal3 72436 31080 72436 31080 0 simpleuart_reg_div_do[24]
rlabel metal2 75264 31864 75264 31864 0 simpleuart_reg_div_do[25]
rlabel metal3 72436 33992 72436 33992 0 simpleuart_reg_div_do[26]
rlabel metal2 75768 34776 75768 34776 0 simpleuart_reg_div_do[27]
rlabel metal2 74760 36512 74760 36512 0 simpleuart_reg_div_do[28]
rlabel metal2 71176 33600 71176 33600 0 simpleuart_reg_div_do[29]
rlabel metal2 77560 7784 77560 7784 0 simpleuart_reg_div_do[2]
rlabel metal2 78176 38808 78176 38808 0 simpleuart_reg_div_do[30]
rlabel metal2 75992 39424 75992 39424 0 simpleuart_reg_div_do[31]
rlabel metal3 77504 8232 77504 8232 0 simpleuart_reg_div_do[3]
rlabel metal3 78722 9688 78722 9688 0 simpleuart_reg_div_do[4]
rlabel metal2 77560 11032 77560 11032 0 simpleuart_reg_div_do[5]
rlabel metal2 78232 11648 78232 11648 0 simpleuart_reg_div_do[6]
rlabel metal2 78232 13384 78232 13384 0 simpleuart_reg_div_do[7]
rlabel metal2 78232 14280 78232 14280 0 simpleuart_reg_div_do[8]
rlabel metal2 78232 15624 78232 15624 0 simpleuart_reg_div_do[9]
rlabel metal2 34048 75656 34048 75656 0 spimem_rdata[0]
rlabel metal2 40936 76664 40936 76664 0 spimem_rdata[10]
rlabel metal2 41496 77490 41496 77490 0 spimem_rdata[11]
rlabel metal2 42280 76664 42280 76664 0 spimem_rdata[12]
rlabel metal2 43624 76888 43624 76888 0 spimem_rdata[13]
rlabel metal2 44520 76832 44520 76832 0 spimem_rdata[14]
rlabel metal2 45976 76608 45976 76608 0 spimem_rdata[15]
rlabel metal2 45080 76216 45080 76216 0 spimem_rdata[16]
rlabel metal2 46760 76720 46760 76720 0 spimem_rdata[17]
rlabel metal2 47880 76552 47880 76552 0 spimem_rdata[18]
rlabel metal2 47096 76160 47096 76160 0 spimem_rdata[19]
rlabel metal2 34776 77434 34776 77434 0 spimem_rdata[1]
rlabel metal2 48328 76832 48328 76832 0 spimem_rdata[20]
rlabel metal3 48720 76664 48720 76664 0 spimem_rdata[21]
rlabel metal2 50120 76832 50120 76832 0 spimem_rdata[22]
rlabel metal2 49784 76216 49784 76216 0 spimem_rdata[23]
rlabel metal2 50232 77938 50232 77938 0 spimem_rdata[24]
rlabel metal2 52136 76888 52136 76888 0 spimem_rdata[25]
rlabel metal2 53032 76832 53032 76832 0 spimem_rdata[26]
rlabel metal2 52248 77490 52248 77490 0 spimem_rdata[27]
rlabel metal3 53424 76664 53424 76664 0 spimem_rdata[28]
rlabel metal2 53704 75656 53704 75656 0 spimem_rdata[29]
rlabel metal2 35672 76048 35672 76048 0 spimem_rdata[2]
rlabel metal2 54712 75880 54712 75880 0 spimem_rdata[30]
rlabel metal2 55720 76104 55720 76104 0 spimem_rdata[31]
rlabel metal2 36456 76608 36456 76608 0 spimem_rdata[3]
rlabel metal2 36904 76720 36904 76720 0 spimem_rdata[4]
rlabel metal2 37408 75656 37408 75656 0 spimem_rdata[5]
rlabel metal2 38248 75656 38248 75656 0 spimem_rdata[6]
rlabel metal2 38808 77938 38808 77938 0 spimem_rdata[7]
rlabel metal2 39368 76664 39368 76664 0 spimem_rdata[8]
rlabel metal2 40152 77938 40152 77938 0 spimem_rdata[9]
rlabel metal2 32760 77490 32760 77490 0 spimem_ready
rlabel metal2 33432 77770 33432 77770 0 spimem_valid
rlabel metal3 58800 75432 58800 75432 0 spimemio_cfgreg_do[0]
rlabel metal2 65072 75768 65072 75768 0 spimemio_cfgreg_do[10]
rlabel metal2 66472 76832 66472 76832 0 spimemio_cfgreg_do[11]
rlabel metal2 67144 76888 67144 76888 0 spimemio_cfgreg_do[12]
rlabel metal2 67816 76832 67816 76832 0 spimemio_cfgreg_do[13]
rlabel metal2 68488 76832 68488 76832 0 spimemio_cfgreg_do[14]
rlabel metal3 68880 76664 68880 76664 0 spimemio_cfgreg_do[15]
rlabel metal2 70280 76944 70280 76944 0 spimemio_cfgreg_do[16]
rlabel metal2 70952 76776 70952 76776 0 spimemio_cfgreg_do[17]
rlabel metal3 71008 76552 71008 76552 0 spimemio_cfgreg_do[18]
rlabel metal2 72296 76888 72296 76888 0 spimemio_cfgreg_do[19]
rlabel metal2 60536 75376 60536 75376 0 spimemio_cfgreg_do[1]
rlabel metal2 73192 76776 73192 76776 0 spimemio_cfgreg_do[20]
rlabel metal2 72408 77490 72408 77490 0 spimemio_cfgreg_do[21]
rlabel metal2 73080 78106 73080 78106 0 spimemio_cfgreg_do[22]
rlabel metal2 73752 78162 73752 78162 0 spimemio_cfgreg_do[23]
rlabel metal2 75768 76776 75768 76776 0 spimemio_cfgreg_do[24]
rlabel metal2 76440 76832 76440 76832 0 spimemio_cfgreg_do[25]
rlabel metal2 76216 76440 76216 76440 0 spimemio_cfgreg_do[26]
rlabel metal2 76888 76552 76888 76552 0 spimemio_cfgreg_do[27]
rlabel metal2 76272 73528 76272 73528 0 spimemio_cfgreg_do[28]
rlabel metal2 77224 72968 77224 72968 0 spimemio_cfgreg_do[29]
rlabel metal2 62888 75488 62888 75488 0 spimemio_cfgreg_do[2]
rlabel metal2 75432 75600 75432 75600 0 spimemio_cfgreg_do[30]
rlabel metal3 77560 74984 77560 74984 0 spimemio_cfgreg_do[31]
rlabel metal3 60760 75544 60760 75544 0 spimemio_cfgreg_do[3]
rlabel metal2 62104 75488 62104 75488 0 spimemio_cfgreg_do[4]
rlabel metal2 62888 76720 62888 76720 0 spimemio_cfgreg_do[5]
rlabel metal2 63336 76832 63336 76832 0 spimemio_cfgreg_do[6]
rlabel metal3 63504 76664 63504 76664 0 spimemio_cfgreg_do[7]
rlabel metal2 64680 76832 64680 76832 0 spimemio_cfgreg_do[8]
rlabel metal2 65352 76888 65352 76888 0 spimemio_cfgreg_do[9]
rlabel metal2 55608 78498 55608 78498 0 spimemio_cfgreg_we[0]
rlabel metal2 56728 76608 56728 76608 0 spimemio_cfgreg_we[1]
rlabel metal2 56952 77938 56952 77938 0 spimemio_cfgreg_we[2]
rlabel metal2 57624 78106 57624 78106 0 spimemio_cfgreg_we[3]
<< properties >>
string FIXED_BBOX 0 0 80000 80000
<< end >>

magic
tech gf180mcuD
magscale 1 10
timestamp 1702204438
<< metal1 >>
rect 1344 46282 48608 46316
rect 1344 46230 4478 46282
rect 4530 46230 4582 46282
rect 4634 46230 4686 46282
rect 4738 46230 35198 46282
rect 35250 46230 35302 46282
rect 35354 46230 35406 46282
rect 35458 46230 48608 46282
rect 1344 46196 48608 46230
rect 29374 46114 29426 46126
rect 29374 46050 29426 46062
rect 33182 46114 33234 46126
rect 33182 46050 33234 46062
rect 36990 46114 37042 46126
rect 36990 46050 37042 46062
rect 10670 46002 10722 46014
rect 10670 45938 10722 45950
rect 17726 46002 17778 46014
rect 26898 45950 26910 46002
rect 26962 45950 26974 46002
rect 17726 45938 17778 45950
rect 16270 45890 16322 45902
rect 13906 45838 13918 45890
rect 13970 45838 13982 45890
rect 15250 45838 15262 45890
rect 15314 45838 15326 45890
rect 16270 45826 16322 45838
rect 18398 45890 18450 45902
rect 18398 45826 18450 45838
rect 19630 45890 19682 45902
rect 20066 45838 20078 45890
rect 20130 45838 20142 45890
rect 23874 45838 23886 45890
rect 23938 45838 23950 45890
rect 25442 45838 25454 45890
rect 25506 45838 25518 45890
rect 28578 45838 28590 45890
rect 28642 45838 28654 45890
rect 31490 45838 31502 45890
rect 31554 45838 31566 45890
rect 32162 45838 32174 45890
rect 32226 45838 32238 45890
rect 35970 45838 35982 45890
rect 36034 45838 36046 45890
rect 39778 45838 39790 45890
rect 39842 45838 39854 45890
rect 42914 45838 42926 45890
rect 42978 45838 42990 45890
rect 44034 45838 44046 45890
rect 44098 45838 44110 45890
rect 19630 45826 19682 45838
rect 19406 45778 19458 45790
rect 19406 45714 19458 45726
rect 24558 45778 24610 45790
rect 24558 45714 24610 45726
rect 35422 45778 35474 45790
rect 35422 45714 35474 45726
rect 39230 45778 39282 45790
rect 39230 45714 39282 45726
rect 1710 45666 1762 45678
rect 1710 45602 1762 45614
rect 8094 45666 8146 45678
rect 8094 45602 8146 45614
rect 9550 45666 9602 45678
rect 9550 45602 9602 45614
rect 11118 45666 11170 45678
rect 11118 45602 11170 45614
rect 11678 45666 11730 45678
rect 11678 45602 11730 45614
rect 12126 45666 12178 45678
rect 12126 45602 12178 45614
rect 12574 45666 12626 45678
rect 12574 45602 12626 45614
rect 13470 45666 13522 45678
rect 14590 45666 14642 45678
rect 13682 45614 13694 45666
rect 13746 45614 13758 45666
rect 13470 45602 13522 45614
rect 14590 45602 14642 45614
rect 15038 45666 15090 45678
rect 15038 45602 15090 45614
rect 15822 45666 15874 45678
rect 15822 45602 15874 45614
rect 17166 45666 17218 45678
rect 17166 45602 17218 45614
rect 18174 45666 18226 45678
rect 18174 45602 18226 45614
rect 18734 45666 18786 45678
rect 18734 45602 18786 45614
rect 20974 45666 21026 45678
rect 20974 45602 21026 45614
rect 22990 45666 23042 45678
rect 22990 45602 23042 45614
rect 24894 45666 24946 45678
rect 24894 45602 24946 45614
rect 31278 45666 31330 45678
rect 31278 45602 31330 45614
rect 35086 45666 35138 45678
rect 35086 45602 35138 45614
rect 38894 45666 38946 45678
rect 38894 45602 38946 45614
rect 40798 45666 40850 45678
rect 40798 45602 40850 45614
rect 42702 45666 42754 45678
rect 42702 45602 42754 45614
rect 44606 45666 44658 45678
rect 44606 45602 44658 45614
rect 46846 45666 46898 45678
rect 46846 45602 46898 45614
rect 47742 45666 47794 45678
rect 47742 45602 47794 45614
rect 48190 45666 48242 45678
rect 48190 45602 48242 45614
rect 1344 45498 48608 45532
rect 1344 45446 19838 45498
rect 19890 45446 19942 45498
rect 19994 45446 20046 45498
rect 20098 45446 48608 45498
rect 1344 45412 48608 45446
rect 25342 45330 25394 45342
rect 25342 45266 25394 45278
rect 30158 45330 30210 45342
rect 30158 45266 30210 45278
rect 31278 45330 31330 45342
rect 31278 45266 31330 45278
rect 46062 45330 46114 45342
rect 46062 45266 46114 45278
rect 48190 45218 48242 45230
rect 26450 45166 26462 45218
rect 26514 45166 26526 45218
rect 29026 45166 29038 45218
rect 29090 45166 29102 45218
rect 31938 45166 31950 45218
rect 32002 45166 32014 45218
rect 32386 45166 32398 45218
rect 32450 45166 32462 45218
rect 34626 45166 34638 45218
rect 34690 45166 34702 45218
rect 37874 45166 37886 45218
rect 37938 45166 37950 45218
rect 42578 45166 42590 45218
rect 42642 45166 42654 45218
rect 48190 45154 48242 45166
rect 25678 45106 25730 45118
rect 13234 45054 13246 45106
rect 13298 45054 13310 45106
rect 13682 45054 13694 45106
rect 13746 45054 13758 45106
rect 17602 45054 17614 45106
rect 17666 45054 17678 45106
rect 20738 45054 20750 45106
rect 20802 45054 20814 45106
rect 24434 45054 24446 45106
rect 24498 45054 24510 45106
rect 26338 45054 26350 45106
rect 26402 45054 26414 45106
rect 29810 45054 29822 45106
rect 29874 45054 29886 45106
rect 30370 45054 30382 45106
rect 30434 45054 30446 45106
rect 33954 45054 33966 45106
rect 34018 45054 34030 45106
rect 37090 45054 37102 45106
rect 37154 45054 37166 45106
rect 41794 45054 41806 45106
rect 41858 45054 41870 45106
rect 45042 45054 45054 45106
rect 45106 45054 45118 45106
rect 25678 45042 25730 45054
rect 7422 44994 7474 45006
rect 7422 44930 7474 44942
rect 7982 44994 8034 45006
rect 7982 44930 8034 44942
rect 8430 44994 8482 45006
rect 8430 44930 8482 44942
rect 9102 44994 9154 45006
rect 9102 44930 9154 44942
rect 9662 44994 9714 45006
rect 9662 44930 9714 44942
rect 10110 44994 10162 45006
rect 16606 44994 16658 45006
rect 33294 44994 33346 45006
rect 41134 44994 41186 45006
rect 10434 44942 10446 44994
rect 10498 44942 10510 44994
rect 12562 44942 12574 44994
rect 12626 44942 12638 44994
rect 14466 44942 14478 44994
rect 14530 44942 14542 44994
rect 18274 44942 18286 44994
rect 18338 44942 18350 44994
rect 20402 44942 20414 44994
rect 20466 44942 20478 44994
rect 21522 44942 21534 44994
rect 21586 44942 21598 44994
rect 23650 44942 23662 44994
rect 23714 44942 23726 44994
rect 24098 44942 24110 44994
rect 24162 44942 24174 44994
rect 26898 44942 26910 44994
rect 26962 44942 26974 44994
rect 36754 44942 36766 44994
rect 36818 44942 36830 44994
rect 40002 44942 40014 44994
rect 40066 44942 40078 44994
rect 10110 44930 10162 44942
rect 16606 44930 16658 44942
rect 33294 44930 33346 44942
rect 41134 44930 41186 44942
rect 41582 44994 41634 45006
rect 44706 44942 44718 44994
rect 44770 44942 44782 44994
rect 41582 44930 41634 44942
rect 31614 44882 31666 44894
rect 7522 44830 7534 44882
rect 7586 44879 7598 44882
rect 8418 44879 8430 44882
rect 7586 44833 8430 44879
rect 7586 44830 7598 44833
rect 8418 44830 8430 44833
rect 8482 44830 8494 44882
rect 31614 44818 31666 44830
rect 1344 44714 48608 44748
rect 1344 44662 4478 44714
rect 4530 44662 4582 44714
rect 4634 44662 4686 44714
rect 4738 44662 35198 44714
rect 35250 44662 35302 44714
rect 35354 44662 35406 44714
rect 35458 44662 48608 44714
rect 1344 44628 48608 44662
rect 27358 44546 27410 44558
rect 27358 44482 27410 44494
rect 27694 44546 27746 44558
rect 27694 44482 27746 44494
rect 34526 44546 34578 44558
rect 34526 44482 34578 44494
rect 42030 44546 42082 44558
rect 42030 44482 42082 44494
rect 44942 44546 44994 44558
rect 44942 44482 44994 44494
rect 17390 44434 17442 44446
rect 37102 44434 37154 44446
rect 11666 44382 11678 44434
rect 11730 44382 11742 44434
rect 20626 44382 20638 44434
rect 20690 44382 20702 44434
rect 23090 44382 23102 44434
rect 23154 44382 23166 44434
rect 25218 44382 25230 44434
rect 25282 44382 25294 44434
rect 31042 44382 31054 44434
rect 31106 44382 31118 44434
rect 33170 44382 33182 44434
rect 33234 44382 33246 44434
rect 40674 44382 40686 44434
rect 40738 44382 40750 44434
rect 17390 44370 17442 44382
rect 37102 44370 37154 44382
rect 7422 44322 7474 44334
rect 7422 44258 7474 44270
rect 7870 44322 7922 44334
rect 7870 44258 7922 44270
rect 8094 44322 8146 44334
rect 21870 44322 21922 44334
rect 29934 44322 29986 44334
rect 45278 44322 45330 44334
rect 47182 44322 47234 44334
rect 8754 44270 8766 44322
rect 8818 44270 8830 44322
rect 17826 44270 17838 44322
rect 17890 44270 17902 44322
rect 25890 44270 25902 44322
rect 25954 44270 25966 44322
rect 28354 44270 28366 44322
rect 28418 44270 28430 44322
rect 30370 44270 30382 44322
rect 30434 44270 30446 44322
rect 33730 44270 33742 44322
rect 33794 44270 33806 44322
rect 37762 44270 37774 44322
rect 37826 44270 37838 44322
rect 41010 44270 41022 44322
rect 41074 44270 41086 44322
rect 44146 44270 44158 44322
rect 44210 44270 44222 44322
rect 45714 44270 45726 44322
rect 45778 44270 45790 44322
rect 8094 44258 8146 44270
rect 21870 44258 21922 44270
rect 29934 44258 29986 44270
rect 45278 44258 45330 44270
rect 47182 44258 47234 44270
rect 8430 44210 8482 44222
rect 12910 44210 12962 44222
rect 9538 44158 9550 44210
rect 9602 44158 9614 44210
rect 8430 44146 8482 44158
rect 12910 44146 12962 44158
rect 14702 44210 14754 44222
rect 14702 44146 14754 44158
rect 16382 44210 16434 44222
rect 16382 44146 16434 44158
rect 16494 44210 16546 44222
rect 18498 44158 18510 44210
rect 18562 44158 18574 44210
rect 22082 44158 22094 44210
rect 22146 44158 22158 44210
rect 22642 44158 22654 44210
rect 22706 44158 22718 44210
rect 28466 44158 28478 44210
rect 28530 44158 28542 44210
rect 38546 44158 38558 44210
rect 38610 44158 38622 44210
rect 45826 44158 45838 44210
rect 45890 44158 45902 44210
rect 47506 44158 47518 44210
rect 47570 44158 47582 44210
rect 47954 44158 47966 44210
rect 48018 44158 48030 44210
rect 16494 44146 16546 44158
rect 4846 44098 4898 44110
rect 4846 44034 4898 44046
rect 5854 44098 5906 44110
rect 5854 44034 5906 44046
rect 6414 44098 6466 44110
rect 6414 44034 6466 44046
rect 6862 44098 6914 44110
rect 6862 44034 6914 44046
rect 7198 44098 7250 44110
rect 7198 44034 7250 44046
rect 7310 44098 7362 44110
rect 7310 44034 7362 44046
rect 8318 44098 8370 44110
rect 8318 44034 8370 44046
rect 12014 44098 12066 44110
rect 12574 44098 12626 44110
rect 12338 44046 12350 44098
rect 12402 44046 12414 44098
rect 12014 44034 12066 44046
rect 12574 44034 12626 44046
rect 12798 44098 12850 44110
rect 12798 44034 12850 44046
rect 13694 44098 13746 44110
rect 13694 44034 13746 44046
rect 14142 44098 14194 44110
rect 14142 44034 14194 44046
rect 14366 44098 14418 44110
rect 14366 44034 14418 44046
rect 14590 44098 14642 44110
rect 14590 44034 14642 44046
rect 15486 44098 15538 44110
rect 15486 44034 15538 44046
rect 15822 44098 15874 44110
rect 15822 44034 15874 44046
rect 16158 44098 16210 44110
rect 16158 44034 16210 44046
rect 17054 44098 17106 44110
rect 17054 44034 17106 44046
rect 21534 44098 21586 44110
rect 21534 44034 21586 44046
rect 26462 44098 26514 44110
rect 26462 44034 26514 44046
rect 29374 44098 29426 44110
rect 29374 44034 29426 44046
rect 43934 44098 43986 44110
rect 43934 44034 43986 44046
rect 46846 44098 46898 44110
rect 46846 44034 46898 44046
rect 1344 43930 48608 43964
rect 1344 43878 19838 43930
rect 19890 43878 19942 43930
rect 19994 43878 20046 43930
rect 20098 43878 48608 43930
rect 1344 43844 48608 43878
rect 15598 43762 15650 43774
rect 15598 43698 15650 43710
rect 21422 43762 21474 43774
rect 21422 43698 21474 43710
rect 29150 43762 29202 43774
rect 29150 43698 29202 43710
rect 45278 43762 45330 43774
rect 45278 43698 45330 43710
rect 11454 43650 11506 43662
rect 6850 43598 6862 43650
rect 6914 43598 6926 43650
rect 11454 43586 11506 43598
rect 16494 43650 16546 43662
rect 18622 43650 18674 43662
rect 18274 43598 18286 43650
rect 18338 43598 18350 43650
rect 16494 43586 16546 43598
rect 18622 43586 18674 43598
rect 19070 43650 19122 43662
rect 25342 43650 25394 43662
rect 23650 43598 23662 43650
rect 23714 43598 23726 43650
rect 19070 43586 19122 43598
rect 25342 43586 25394 43598
rect 39006 43650 39058 43662
rect 40910 43650 40962 43662
rect 39554 43598 39566 43650
rect 39618 43598 39630 43650
rect 39890 43598 39902 43650
rect 39954 43598 39966 43650
rect 43922 43598 43934 43650
rect 43986 43598 43998 43650
rect 39006 43586 39058 43598
rect 40910 43586 40962 43598
rect 11342 43538 11394 43550
rect 6178 43486 6190 43538
rect 6242 43486 6254 43538
rect 9986 43486 9998 43538
rect 10050 43486 10062 43538
rect 10882 43486 10894 43538
rect 10946 43486 10958 43538
rect 11342 43474 11394 43486
rect 11566 43538 11618 43550
rect 15710 43538 15762 43550
rect 11890 43486 11902 43538
rect 11954 43486 11966 43538
rect 12450 43486 12462 43538
rect 12514 43486 12526 43538
rect 11566 43474 11618 43486
rect 15710 43474 15762 43486
rect 16270 43538 16322 43550
rect 16270 43474 16322 43486
rect 18958 43538 19010 43550
rect 18958 43474 19010 43486
rect 19294 43538 19346 43550
rect 39342 43538 39394 43550
rect 21634 43486 21646 43538
rect 21698 43486 21710 43538
rect 22530 43486 22542 43538
rect 22594 43486 22606 43538
rect 25890 43486 25902 43538
rect 25954 43486 25966 43538
rect 29698 43486 29710 43538
rect 29762 43486 29774 43538
rect 33282 43486 33294 43538
rect 33346 43486 33358 43538
rect 35970 43486 35982 43538
rect 36034 43486 36046 43538
rect 19294 43474 19346 43486
rect 39342 43474 39394 43486
rect 41246 43538 41298 43550
rect 44594 43486 44606 43538
rect 44658 43486 44670 43538
rect 45826 43486 45838 43538
rect 45890 43486 45902 43538
rect 41246 43474 41298 43486
rect 1822 43426 1874 43438
rect 1822 43362 1874 43374
rect 2270 43426 2322 43438
rect 2270 43362 2322 43374
rect 3950 43426 4002 43438
rect 3950 43362 4002 43374
rect 4398 43426 4450 43438
rect 4398 43362 4450 43374
rect 4846 43426 4898 43438
rect 4846 43362 4898 43374
rect 5406 43426 5458 43438
rect 5406 43362 5458 43374
rect 5854 43426 5906 43438
rect 9550 43426 9602 43438
rect 8978 43374 8990 43426
rect 9042 43374 9054 43426
rect 5854 43362 5906 43374
rect 9550 43362 9602 43374
rect 10446 43426 10498 43438
rect 17502 43426 17554 43438
rect 13122 43374 13134 43426
rect 13186 43374 13198 43426
rect 15250 43374 15262 43426
rect 15314 43374 15326 43426
rect 10446 43362 10498 43374
rect 17502 43362 17554 43374
rect 17950 43426 18002 43438
rect 17950 43362 18002 43374
rect 19742 43426 19794 43438
rect 19742 43362 19794 43374
rect 20638 43426 20690 43438
rect 20638 43362 20690 43374
rect 21086 43426 21138 43438
rect 34078 43426 34130 43438
rect 26562 43374 26574 43426
rect 26626 43374 26638 43426
rect 28690 43374 28702 43426
rect 28754 43374 28766 43426
rect 30370 43374 30382 43426
rect 30434 43374 30446 43426
rect 32498 43374 32510 43426
rect 32562 43374 32574 43426
rect 21086 43362 21138 43374
rect 34078 43362 34130 43374
rect 36990 43426 37042 43438
rect 41794 43374 41806 43426
rect 41858 43374 41870 43426
rect 36990 43362 37042 43374
rect 15934 43314 15986 43326
rect 3826 43262 3838 43314
rect 3890 43311 3902 43314
rect 4834 43311 4846 43314
rect 3890 43265 4846 43311
rect 3890 43262 3902 43265
rect 4834 43262 4846 43265
rect 4898 43262 4910 43314
rect 15934 43250 15986 43262
rect 47966 43314 48018 43326
rect 47966 43250 48018 43262
rect 1344 43146 48608 43180
rect 1344 43094 4478 43146
rect 4530 43094 4582 43146
rect 4634 43094 4686 43146
rect 4738 43094 35198 43146
rect 35250 43094 35302 43146
rect 35354 43094 35406 43146
rect 35458 43094 48608 43146
rect 1344 43060 48608 43094
rect 29598 42978 29650 42990
rect 29598 42914 29650 42926
rect 32174 42978 32226 42990
rect 32174 42914 32226 42926
rect 34526 42978 34578 42990
rect 34526 42914 34578 42926
rect 37214 42978 37266 42990
rect 37214 42914 37266 42926
rect 40126 42978 40178 42990
rect 40126 42914 40178 42926
rect 42926 42978 42978 42990
rect 42926 42914 42978 42926
rect 43262 42978 43314 42990
rect 43262 42914 43314 42926
rect 13694 42866 13746 42878
rect 19070 42866 19122 42878
rect 10098 42814 10110 42866
rect 10162 42814 10174 42866
rect 14578 42814 14590 42866
rect 14642 42814 14654 42866
rect 15698 42814 15710 42866
rect 15762 42814 15774 42866
rect 26114 42814 26126 42866
rect 26178 42814 26190 42866
rect 46946 42814 46958 42866
rect 47010 42814 47022 42866
rect 13694 42802 13746 42814
rect 19070 42802 19122 42814
rect 9102 42754 9154 42766
rect 13806 42754 13858 42766
rect 5618 42702 5630 42754
rect 5682 42702 5694 42754
rect 10994 42702 11006 42754
rect 11058 42702 11070 42754
rect 11330 42702 11342 42754
rect 11394 42702 11406 42754
rect 9102 42690 9154 42702
rect 13806 42690 13858 42702
rect 14254 42754 14306 42766
rect 20414 42754 20466 42766
rect 18610 42702 18622 42754
rect 18674 42702 18686 42754
rect 19954 42702 19966 42754
rect 20018 42702 20030 42754
rect 23314 42702 23326 42754
rect 23378 42702 23390 42754
rect 31154 42702 31166 42754
rect 31218 42702 31230 42754
rect 36194 42702 36206 42754
rect 36258 42702 36270 42754
rect 39330 42702 39342 42754
rect 39394 42702 39406 42754
rect 42018 42702 42030 42754
rect 42082 42702 42094 42754
rect 43698 42702 43710 42754
rect 43762 42702 43774 42754
rect 48178 42702 48190 42754
rect 48242 42702 48254 42754
rect 14254 42690 14306 42702
rect 20414 42690 20466 42702
rect 9214 42642 9266 42654
rect 19406 42642 19458 42654
rect 27022 42642 27074 42654
rect 6402 42590 6414 42642
rect 6466 42590 6478 42642
rect 10210 42590 10222 42642
rect 10274 42590 10286 42642
rect 11442 42590 11454 42642
rect 11506 42590 11518 42642
rect 17826 42590 17838 42642
rect 17890 42590 17902 42642
rect 23986 42590 23998 42642
rect 24050 42590 24062 42642
rect 9214 42578 9266 42590
rect 19406 42578 19458 42590
rect 27022 42578 27074 42590
rect 27358 42642 27410 42654
rect 27358 42578 27410 42590
rect 29262 42642 29314 42654
rect 45278 42642 45330 42654
rect 29922 42590 29934 42642
rect 29986 42590 29998 42642
rect 30258 42590 30270 42642
rect 30322 42590 30334 42642
rect 34738 42590 34750 42642
rect 34802 42590 34814 42642
rect 35074 42590 35086 42642
rect 35138 42590 35150 42642
rect 43810 42590 43822 42642
rect 43874 42590 43886 42642
rect 29262 42578 29314 42590
rect 45278 42578 45330 42590
rect 1822 42530 1874 42542
rect 1822 42466 1874 42478
rect 2494 42530 2546 42542
rect 2494 42466 2546 42478
rect 2942 42530 2994 42542
rect 2942 42466 2994 42478
rect 3390 42530 3442 42542
rect 3390 42466 3442 42478
rect 3950 42530 4002 42542
rect 3950 42466 4002 42478
rect 4398 42530 4450 42542
rect 4398 42466 4450 42478
rect 4846 42530 4898 42542
rect 9438 42530 9490 42542
rect 8642 42478 8654 42530
rect 8706 42478 8718 42530
rect 4846 42466 4898 42478
rect 9438 42466 9490 42478
rect 13582 42530 13634 42542
rect 13582 42466 13634 42478
rect 15038 42530 15090 42542
rect 15038 42466 15090 42478
rect 18958 42530 19010 42542
rect 18958 42466 19010 42478
rect 19182 42530 19234 42542
rect 19182 42466 19234 42478
rect 26574 42530 26626 42542
rect 26574 42466 26626 42478
rect 34190 42530 34242 42542
rect 34190 42466 34242 42478
rect 36430 42530 36482 42542
rect 36430 42466 36482 42478
rect 1344 42362 48608 42396
rect 1344 42310 19838 42362
rect 19890 42310 19942 42362
rect 19994 42310 20046 42362
rect 20098 42310 48608 42362
rect 1344 42276 48608 42310
rect 12462 42194 12514 42206
rect 7970 42142 7982 42194
rect 8034 42142 8046 42194
rect 12462 42130 12514 42142
rect 15262 42194 15314 42206
rect 24222 42194 24274 42206
rect 15586 42142 15598 42194
rect 15650 42142 15662 42194
rect 15262 42130 15314 42142
rect 24222 42130 24274 42142
rect 31278 42194 31330 42206
rect 31278 42130 31330 42142
rect 48190 42194 48242 42206
rect 48190 42130 48242 42142
rect 5854 42082 5906 42094
rect 16606 42082 16658 42094
rect 27694 42082 27746 42094
rect 4834 42030 4846 42082
rect 4898 42030 4910 42082
rect 8866 42030 8878 42082
rect 8930 42030 8942 42082
rect 11890 42030 11902 42082
rect 11954 42030 11966 42082
rect 18274 42030 18286 42082
rect 18338 42030 18350 42082
rect 18946 42030 18958 42082
rect 19010 42030 19022 42082
rect 26226 42030 26238 42082
rect 26290 42030 26302 42082
rect 5854 42018 5906 42030
rect 16606 42018 16658 42030
rect 27694 42018 27746 42030
rect 30382 42082 30434 42094
rect 30382 42018 30434 42030
rect 31614 42082 31666 42094
rect 31614 42018 31666 42030
rect 1710 41970 1762 41982
rect 1710 41906 1762 41918
rect 3838 41970 3890 41982
rect 3838 41906 3890 41918
rect 4286 41970 4338 41982
rect 10446 41970 10498 41982
rect 4610 41918 4622 41970
rect 4674 41918 4686 41970
rect 6962 41918 6974 41970
rect 7026 41918 7038 41970
rect 7410 41918 7422 41970
rect 7474 41918 7486 41970
rect 4286 41906 4338 41918
rect 10446 41906 10498 41918
rect 10670 41970 10722 41982
rect 10670 41906 10722 41918
rect 13358 41970 13410 41982
rect 13358 41906 13410 41918
rect 13582 41970 13634 41982
rect 13582 41906 13634 41918
rect 13806 41970 13858 41982
rect 13806 41906 13858 41918
rect 14030 41970 14082 41982
rect 14030 41906 14082 41918
rect 14366 41970 14418 41982
rect 14366 41906 14418 41918
rect 14926 41970 14978 41982
rect 14926 41906 14978 41918
rect 15934 41970 15986 41982
rect 24558 41970 24610 41982
rect 30718 41970 30770 41982
rect 18498 41918 18510 41970
rect 18562 41918 18574 41970
rect 20626 41918 20638 41970
rect 20690 41918 20702 41970
rect 23762 41918 23774 41970
rect 23826 41918 23838 41970
rect 26338 41918 26350 41970
rect 26402 41918 26414 41970
rect 27458 41918 27470 41970
rect 27522 41918 27534 41970
rect 15934 41906 15986 41918
rect 24558 41906 24610 41918
rect 30718 41906 30770 41918
rect 32510 41970 32562 41982
rect 39678 41970 39730 41982
rect 33170 41918 33182 41970
rect 33234 41918 33246 41970
rect 36306 41918 36318 41970
rect 36370 41918 36382 41970
rect 37090 41918 37102 41970
rect 37154 41918 37166 41970
rect 44482 41918 44494 41970
rect 44546 41918 44558 41970
rect 44818 41918 44830 41970
rect 44882 41918 44894 41970
rect 32510 41906 32562 41918
rect 39678 41906 39730 41918
rect 2270 41858 2322 41870
rect 2270 41794 2322 41806
rect 3166 41858 3218 41870
rect 3166 41794 3218 41806
rect 9774 41858 9826 41870
rect 25342 41858 25394 41870
rect 11554 41806 11566 41858
rect 11618 41806 11630 41858
rect 12898 41806 12910 41858
rect 12962 41806 12974 41858
rect 16146 41806 16158 41858
rect 16210 41806 16222 41858
rect 17490 41806 17502 41858
rect 17554 41806 17566 41858
rect 20962 41806 20974 41858
rect 21026 41806 21038 41858
rect 23090 41806 23102 41858
rect 23154 41806 23166 41858
rect 9774 41794 9826 41806
rect 25342 41794 25394 41806
rect 28814 41858 28866 41870
rect 28814 41794 28866 41806
rect 30046 41858 30098 41870
rect 40126 41858 40178 41870
rect 33842 41806 33854 41858
rect 33906 41806 33918 41858
rect 35970 41806 35982 41858
rect 36034 41806 36046 41858
rect 39218 41806 39230 41858
rect 39282 41806 39294 41858
rect 30046 41794 30098 41806
rect 40126 41794 40178 41806
rect 41022 41858 41074 41870
rect 41570 41806 41582 41858
rect 41634 41806 41646 41858
rect 43698 41806 43710 41858
rect 43762 41806 43774 41858
rect 45602 41806 45614 41858
rect 45666 41806 45678 41858
rect 47730 41806 47742 41858
rect 47794 41806 47806 41858
rect 41022 41794 41074 41806
rect 10334 41746 10386 41758
rect 10334 41682 10386 41694
rect 16718 41746 16770 41758
rect 16718 41682 16770 41694
rect 25678 41746 25730 41758
rect 25678 41682 25730 41694
rect 1344 41578 48608 41612
rect 1344 41526 4478 41578
rect 4530 41526 4582 41578
rect 4634 41526 4686 41578
rect 4738 41526 35198 41578
rect 35250 41526 35302 41578
rect 35354 41526 35406 41578
rect 35458 41526 48608 41578
rect 1344 41492 48608 41526
rect 34638 41410 34690 41422
rect 12674 41358 12686 41410
rect 12738 41358 12750 41410
rect 16258 41358 16270 41410
rect 16322 41358 16334 41410
rect 34638 41346 34690 41358
rect 37214 41410 37266 41422
rect 37214 41346 37266 41358
rect 37550 41410 37602 41422
rect 37550 41346 37602 41358
rect 17278 41298 17330 41310
rect 5058 41246 5070 41298
rect 5122 41246 5134 41298
rect 5842 41246 5854 41298
rect 5906 41246 5918 41298
rect 15026 41246 15038 41298
rect 15090 41246 15102 41298
rect 17278 41234 17330 41246
rect 18398 41298 18450 41310
rect 24110 41298 24162 41310
rect 21746 41246 21758 41298
rect 21810 41246 21822 41298
rect 18398 41234 18450 41246
rect 24110 41234 24162 41246
rect 24894 41298 24946 41310
rect 32734 41298 32786 41310
rect 25666 41246 25678 41298
rect 25730 41246 25742 41298
rect 27794 41246 27806 41298
rect 27858 41246 27870 41298
rect 30146 41246 30158 41298
rect 30210 41246 30222 41298
rect 32274 41246 32286 41298
rect 32338 41246 32350 41298
rect 24894 41234 24946 41246
rect 32734 41234 32786 41246
rect 43934 41298 43986 41310
rect 47842 41246 47854 41298
rect 47906 41246 47918 41298
rect 43934 41234 43986 41246
rect 9326 41186 9378 41198
rect 2146 41134 2158 41186
rect 2210 41134 2222 41186
rect 5618 41134 5630 41186
rect 5682 41134 5694 41186
rect 8754 41134 8766 41186
rect 8818 41134 8830 41186
rect 9326 41122 9378 41134
rect 11006 41186 11058 41198
rect 15710 41186 15762 41198
rect 17054 41186 17106 41198
rect 12898 41134 12910 41186
rect 12962 41134 12974 41186
rect 13794 41134 13806 41186
rect 13858 41134 13870 41186
rect 14914 41134 14926 41186
rect 14978 41134 14990 41186
rect 16370 41134 16382 41186
rect 16434 41134 16446 41186
rect 11006 41122 11058 41134
rect 15710 41122 15762 41134
rect 17054 41122 17106 41134
rect 17390 41186 17442 41198
rect 17390 41122 17442 41134
rect 18510 41186 18562 41198
rect 20414 41186 20466 41198
rect 19842 41134 19854 41186
rect 19906 41134 19918 41186
rect 18510 41122 18562 41134
rect 20414 41122 20466 41134
rect 21310 41186 21362 41198
rect 38894 41186 38946 41198
rect 28578 41134 28590 41186
rect 28642 41134 28654 41186
rect 29362 41134 29374 41186
rect 29426 41134 29438 41186
rect 33618 41134 33630 41186
rect 33682 41134 33694 41186
rect 35186 41134 35198 41186
rect 35250 41134 35262 41186
rect 36194 41134 36206 41186
rect 36258 41134 36270 41186
rect 21310 41122 21362 41134
rect 38894 41122 38946 41134
rect 39230 41186 39282 41198
rect 41470 41186 41522 41198
rect 39666 41134 39678 41186
rect 39730 41134 39742 41186
rect 40786 41134 40798 41186
rect 40850 41134 40862 41186
rect 39230 41122 39282 41134
rect 41470 41122 41522 41134
rect 41806 41186 41858 41198
rect 45602 41134 45614 41186
rect 45666 41134 45678 41186
rect 41806 41122 41858 41134
rect 9774 41074 9826 41086
rect 2930 41022 2942 41074
rect 2994 41022 3006 41074
rect 7074 41022 7086 41074
rect 7138 41022 7150 41074
rect 7970 41022 7982 41074
rect 8034 41022 8046 41074
rect 9774 41010 9826 41022
rect 12126 41074 12178 41086
rect 14254 41074 14306 41086
rect 16830 41074 16882 41086
rect 12338 41022 12350 41074
rect 12402 41022 12414 41074
rect 15922 41022 15934 41074
rect 15986 41022 15998 41074
rect 12126 41010 12178 41022
rect 14254 41010 14306 41022
rect 16830 41010 16882 41022
rect 18286 41074 18338 41086
rect 18286 41010 18338 41022
rect 18846 41074 18898 41086
rect 33854 41074 33906 41086
rect 19954 41022 19966 41074
rect 20018 41022 20030 41074
rect 20290 41022 20302 41074
rect 20354 41022 20366 41074
rect 22642 41022 22654 41074
rect 22706 41022 22718 41074
rect 18846 41010 18898 41022
rect 33854 41010 33906 41022
rect 34302 41074 34354 41086
rect 43150 41074 43202 41086
rect 35410 41022 35422 41074
rect 35474 41022 35486 41074
rect 37762 41022 37774 41074
rect 37826 41022 37838 41074
rect 38210 41022 38222 41074
rect 38274 41022 38286 41074
rect 39778 41022 39790 41074
rect 39842 41022 39854 41074
rect 42018 41022 42030 41074
rect 42082 41022 42094 41074
rect 42354 41022 42366 41074
rect 42418 41022 42430 41074
rect 34302 41010 34354 41022
rect 43150 41010 43202 41022
rect 44942 41074 44994 41086
rect 44942 41010 44994 41022
rect 45278 41074 45330 41086
rect 45278 41010 45330 41022
rect 1822 40962 1874 40974
rect 1822 40898 1874 40910
rect 9326 40962 9378 40974
rect 16494 40962 16546 40974
rect 12450 40910 12462 40962
rect 12514 40910 12526 40962
rect 13570 40910 13582 40962
rect 13634 40910 13646 40962
rect 9326 40898 9378 40910
rect 16494 40898 16546 40910
rect 17950 40962 18002 40974
rect 17950 40898 18002 40910
rect 19406 40962 19458 40974
rect 19406 40898 19458 40910
rect 22990 40962 23042 40974
rect 22990 40898 23042 40910
rect 36430 40962 36482 40974
rect 36430 40898 36482 40910
rect 41022 40962 41074 40974
rect 41022 40898 41074 40910
rect 43486 40962 43538 40974
rect 43486 40898 43538 40910
rect 1344 40794 48608 40828
rect 1344 40742 19838 40794
rect 19890 40742 19942 40794
rect 19994 40742 20046 40794
rect 20098 40742 48608 40794
rect 1344 40708 48608 40742
rect 6302 40626 6354 40638
rect 6302 40562 6354 40574
rect 7198 40626 7250 40638
rect 7198 40562 7250 40574
rect 15934 40626 15986 40638
rect 15934 40562 15986 40574
rect 18286 40626 18338 40638
rect 18286 40562 18338 40574
rect 19742 40626 19794 40638
rect 19742 40562 19794 40574
rect 28254 40626 28306 40638
rect 28254 40562 28306 40574
rect 30942 40626 30994 40638
rect 30942 40562 30994 40574
rect 36318 40626 36370 40638
rect 36318 40562 36370 40574
rect 43822 40626 43874 40638
rect 43822 40562 43874 40574
rect 44606 40626 44658 40638
rect 44606 40562 44658 40574
rect 10558 40514 10610 40526
rect 16830 40514 16882 40526
rect 20862 40514 20914 40526
rect 5282 40462 5294 40514
rect 5346 40462 5358 40514
rect 5954 40462 5966 40514
rect 6018 40462 6030 40514
rect 11890 40462 11902 40514
rect 11954 40462 11966 40514
rect 13010 40462 13022 40514
rect 13074 40462 13086 40514
rect 15474 40462 15486 40514
rect 15538 40462 15550 40514
rect 20402 40462 20414 40514
rect 20466 40462 20478 40514
rect 10558 40450 10610 40462
rect 16830 40450 16882 40462
rect 20862 40450 20914 40462
rect 22318 40514 22370 40526
rect 35646 40514 35698 40526
rect 45278 40514 45330 40526
rect 23202 40462 23214 40514
rect 23266 40462 23278 40514
rect 26450 40462 26462 40514
rect 26514 40462 26526 40514
rect 27010 40462 27022 40514
rect 27074 40462 27086 40514
rect 29250 40462 29262 40514
rect 29314 40462 29326 40514
rect 31490 40462 31502 40514
rect 31554 40462 31566 40514
rect 31938 40462 31950 40514
rect 32002 40462 32014 40514
rect 37426 40462 37438 40514
rect 37490 40462 37502 40514
rect 41682 40462 41694 40514
rect 41746 40462 41758 40514
rect 42018 40462 42030 40514
rect 42082 40462 42094 40514
rect 42914 40462 42926 40514
rect 42978 40462 42990 40514
rect 22318 40450 22370 40462
rect 35646 40450 35698 40462
rect 45278 40450 45330 40462
rect 8766 40402 8818 40414
rect 1810 40350 1822 40402
rect 1874 40350 1886 40402
rect 5058 40350 5070 40402
rect 5122 40350 5134 40402
rect 8766 40338 8818 40350
rect 11006 40402 11058 40414
rect 16718 40402 16770 40414
rect 11330 40350 11342 40402
rect 11394 40350 11406 40402
rect 13682 40350 13694 40402
rect 13746 40350 13758 40402
rect 14802 40350 14814 40402
rect 14866 40350 14878 40402
rect 11006 40338 11058 40350
rect 16718 40338 16770 40350
rect 18846 40402 18898 40414
rect 18846 40338 18898 40350
rect 19182 40402 19234 40414
rect 20638 40402 20690 40414
rect 20178 40350 20190 40402
rect 20242 40350 20254 40402
rect 19182 40338 19234 40350
rect 20638 40338 20690 40350
rect 20974 40402 21026 40414
rect 29934 40402 29986 40414
rect 33966 40402 34018 40414
rect 22754 40350 22766 40402
rect 22818 40350 22830 40402
rect 23426 40350 23438 40402
rect 23490 40350 23502 40402
rect 29138 40350 29150 40402
rect 29202 40350 29214 40402
rect 33170 40350 33182 40402
rect 33234 40350 33246 40402
rect 35186 40350 35198 40402
rect 35250 40350 35262 40402
rect 36642 40350 36654 40402
rect 36706 40350 36718 40402
rect 42690 40350 42702 40402
rect 42754 40350 42766 40402
rect 45042 40350 45054 40402
rect 45106 40350 45118 40402
rect 45602 40350 45614 40402
rect 45666 40350 45678 40402
rect 20974 40338 21026 40350
rect 29934 40338 29986 40350
rect 33966 40338 34018 40350
rect 6638 40290 6690 40302
rect 2482 40238 2494 40290
rect 2546 40238 2558 40290
rect 4610 40238 4622 40290
rect 4674 40238 4686 40290
rect 6638 40226 6690 40238
rect 8094 40290 8146 40302
rect 8094 40226 8146 40238
rect 9886 40290 9938 40302
rect 9886 40226 9938 40238
rect 10110 40290 10162 40302
rect 10110 40226 10162 40238
rect 10894 40290 10946 40302
rect 10894 40226 10946 40238
rect 16046 40290 16098 40302
rect 16046 40226 16098 40238
rect 17614 40290 17666 40302
rect 17614 40226 17666 40238
rect 17950 40290 18002 40302
rect 17950 40226 18002 40238
rect 19294 40290 19346 40302
rect 19294 40226 19346 40238
rect 26238 40290 26290 40302
rect 26238 40226 26290 40238
rect 31278 40290 31330 40302
rect 40014 40290 40066 40302
rect 33506 40238 33518 40290
rect 33570 40238 33582 40290
rect 34402 40238 34414 40290
rect 34466 40238 34478 40290
rect 39554 40238 39566 40290
rect 39618 40238 39630 40290
rect 31278 40226 31330 40238
rect 40014 40226 40066 40238
rect 7646 40178 7698 40190
rect 7646 40114 7698 40126
rect 8318 40178 8370 40190
rect 8318 40114 8370 40126
rect 8542 40178 8594 40190
rect 8542 40114 8594 40126
rect 9438 40178 9490 40190
rect 9438 40114 9490 40126
rect 10334 40178 10386 40190
rect 10334 40114 10386 40126
rect 16270 40178 16322 40190
rect 25902 40178 25954 40190
rect 19506 40126 19518 40178
rect 19570 40175 19582 40178
rect 19730 40175 19742 40178
rect 19570 40129 19742 40175
rect 19570 40126 19582 40129
rect 19730 40126 19742 40129
rect 19794 40126 19806 40178
rect 16270 40114 16322 40126
rect 25902 40114 25954 40126
rect 28590 40178 28642 40190
rect 28590 40114 28642 40126
rect 41022 40178 41074 40190
rect 41022 40114 41074 40126
rect 41358 40178 41410 40190
rect 41358 40114 41410 40126
rect 43486 40178 43538 40190
rect 43486 40114 43538 40126
rect 47966 40178 48018 40190
rect 47966 40114 48018 40126
rect 1344 40010 48608 40044
rect 1344 39958 4478 40010
rect 4530 39958 4582 40010
rect 4634 39958 4686 40010
rect 4738 39958 35198 40010
rect 35250 39958 35302 40010
rect 35354 39958 35406 40010
rect 35458 39958 48608 40010
rect 1344 39924 48608 39958
rect 6302 39842 6354 39854
rect 6302 39778 6354 39790
rect 7422 39842 7474 39854
rect 7422 39778 7474 39790
rect 7646 39842 7698 39854
rect 7646 39778 7698 39790
rect 7870 39842 7922 39854
rect 16830 39842 16882 39854
rect 13458 39790 13470 39842
rect 13522 39790 13534 39842
rect 16482 39790 16494 39842
rect 16546 39790 16558 39842
rect 7870 39778 7922 39790
rect 16830 39778 16882 39790
rect 17166 39842 17218 39854
rect 17166 39778 17218 39790
rect 38334 39842 38386 39854
rect 38334 39778 38386 39790
rect 38670 39842 38722 39854
rect 38670 39778 38722 39790
rect 43038 39842 43090 39854
rect 43038 39778 43090 39790
rect 43374 39842 43426 39854
rect 43374 39778 43426 39790
rect 2270 39730 2322 39742
rect 2270 39666 2322 39678
rect 3390 39730 3442 39742
rect 3390 39666 3442 39678
rect 7198 39730 7250 39742
rect 7198 39666 7250 39678
rect 18958 39730 19010 39742
rect 18958 39666 19010 39678
rect 22990 39730 23042 39742
rect 31614 39730 31666 39742
rect 36430 39730 36482 39742
rect 26786 39678 26798 39730
rect 26850 39678 26862 39730
rect 34850 39678 34862 39730
rect 34914 39678 34926 39730
rect 22990 39666 23042 39678
rect 31614 39666 31666 39678
rect 36430 39666 36482 39678
rect 37102 39730 37154 39742
rect 42018 39678 42030 39730
rect 42082 39678 42094 39730
rect 46050 39678 46062 39730
rect 46114 39678 46126 39730
rect 48178 39678 48190 39730
rect 48242 39678 48254 39730
rect 37102 39666 37154 39678
rect 1710 39618 1762 39630
rect 1710 39554 1762 39566
rect 2606 39618 2658 39630
rect 2606 39554 2658 39566
rect 3278 39618 3330 39630
rect 4062 39618 4114 39630
rect 15822 39618 15874 39630
rect 3826 39566 3838 39618
rect 3890 39566 3902 39618
rect 10322 39566 10334 39618
rect 10386 39566 10398 39618
rect 12338 39566 12350 39618
rect 12402 39566 12414 39618
rect 14242 39566 14254 39618
rect 14306 39566 14318 39618
rect 3278 39554 3330 39566
rect 4062 39554 4114 39566
rect 15822 39554 15874 39566
rect 16046 39618 16098 39630
rect 18622 39618 18674 39630
rect 20302 39618 20354 39630
rect 17154 39566 17166 39618
rect 17218 39566 17230 39618
rect 18386 39566 18398 39618
rect 18450 39566 18462 39618
rect 19842 39566 19854 39618
rect 19906 39566 19918 39618
rect 16046 39554 16098 39566
rect 18622 39554 18674 39566
rect 20302 39554 20354 39566
rect 22094 39618 22146 39630
rect 22094 39554 22146 39566
rect 22654 39618 22706 39630
rect 23426 39566 23438 39618
rect 23490 39566 23502 39618
rect 23986 39566 23998 39618
rect 24050 39566 24062 39618
rect 31938 39566 31950 39618
rect 32002 39566 32014 39618
rect 39106 39566 39118 39618
rect 39170 39566 39182 39618
rect 44146 39566 44158 39618
rect 44210 39566 44222 39618
rect 45378 39566 45390 39618
rect 45442 39566 45454 39618
rect 22654 39554 22706 39566
rect 2942 39506 2994 39518
rect 2942 39442 2994 39454
rect 4398 39506 4450 39518
rect 4398 39442 4450 39454
rect 5966 39506 6018 39518
rect 5966 39442 6018 39454
rect 6190 39506 6242 39518
rect 11230 39506 11282 39518
rect 8530 39454 8542 39506
rect 8594 39454 8606 39506
rect 6190 39442 6242 39454
rect 11230 39442 11282 39454
rect 13918 39506 13970 39518
rect 13918 39442 13970 39454
rect 14030 39506 14082 39518
rect 14030 39442 14082 39454
rect 14702 39506 14754 39518
rect 14702 39442 14754 39454
rect 15934 39506 15986 39518
rect 19070 39506 19122 39518
rect 18834 39454 18846 39506
rect 18898 39454 18910 39506
rect 15934 39442 15986 39454
rect 19070 39442 19122 39454
rect 19406 39506 19458 39518
rect 24658 39454 24670 39506
rect 24722 39454 24734 39506
rect 32722 39454 32734 39506
rect 32786 39454 32798 39506
rect 35186 39454 35198 39506
rect 35250 39454 35262 39506
rect 37762 39454 37774 39506
rect 37826 39454 37838 39506
rect 38098 39454 38110 39506
rect 38162 39454 38174 39506
rect 39890 39454 39902 39506
rect 39954 39454 39966 39506
rect 43922 39454 43934 39506
rect 43986 39454 43998 39506
rect 19406 39442 19458 39454
rect 3502 39394 3554 39406
rect 3502 39330 3554 39342
rect 4286 39394 4338 39406
rect 4286 39330 4338 39342
rect 4846 39394 4898 39406
rect 4846 39330 4898 39342
rect 6862 39394 6914 39406
rect 6862 39330 6914 39342
rect 8318 39394 8370 39406
rect 8318 39330 8370 39342
rect 9886 39394 9938 39406
rect 9886 39330 9938 39342
rect 13022 39394 13074 39406
rect 13022 39330 13074 39342
rect 14590 39394 14642 39406
rect 14590 39330 14642 39342
rect 15262 39394 15314 39406
rect 15262 39330 15314 39342
rect 18062 39394 18114 39406
rect 18062 39330 18114 39342
rect 21422 39394 21474 39406
rect 21422 39330 21474 39342
rect 27246 39394 27298 39406
rect 27246 39330 27298 39342
rect 29262 39394 29314 39406
rect 29262 39330 29314 39342
rect 35534 39394 35586 39406
rect 35534 39330 35586 39342
rect 42478 39394 42530 39406
rect 42478 39330 42530 39342
rect 45054 39394 45106 39406
rect 45054 39330 45106 39342
rect 1344 39226 48608 39260
rect 1344 39174 19838 39226
rect 19890 39174 19942 39226
rect 19994 39174 20046 39226
rect 20098 39174 48608 39226
rect 1344 39140 48608 39174
rect 6526 39058 6578 39070
rect 6526 38994 6578 39006
rect 6750 39058 6802 39070
rect 6750 38994 6802 39006
rect 8542 39058 8594 39070
rect 8542 38994 8594 39006
rect 9998 39058 10050 39070
rect 9998 38994 10050 39006
rect 10894 39058 10946 39070
rect 10894 38994 10946 39006
rect 16046 39058 16098 39070
rect 16046 38994 16098 39006
rect 20302 39058 20354 39070
rect 20302 38994 20354 39006
rect 21646 39058 21698 39070
rect 21646 38994 21698 39006
rect 21870 39058 21922 39070
rect 22990 39058 23042 39070
rect 22642 39006 22654 39058
rect 22706 39006 22718 39058
rect 21870 38994 21922 39006
rect 22990 38994 23042 39006
rect 23662 39058 23714 39070
rect 23662 38994 23714 39006
rect 25230 39058 25282 39070
rect 25230 38994 25282 39006
rect 31838 39058 31890 39070
rect 31838 38994 31890 39006
rect 33070 39058 33122 39070
rect 33070 38994 33122 39006
rect 40238 39058 40290 39070
rect 40238 38994 40290 39006
rect 40910 39058 40962 39070
rect 40910 38994 40962 39006
rect 41694 39058 41746 39070
rect 41694 38994 41746 39006
rect 5294 38946 5346 38958
rect 5294 38882 5346 38894
rect 7982 38946 8034 38958
rect 7982 38882 8034 38894
rect 11790 38946 11842 38958
rect 20526 38946 20578 38958
rect 12226 38894 12238 38946
rect 12290 38894 12302 38946
rect 18162 38894 18174 38946
rect 18226 38894 18238 38946
rect 19506 38894 19518 38946
rect 19570 38894 19582 38946
rect 11790 38882 11842 38894
rect 20526 38882 20578 38894
rect 21198 38946 21250 38958
rect 21198 38882 21250 38894
rect 21310 38946 21362 38958
rect 25566 38946 25618 38958
rect 31054 38946 31106 38958
rect 45950 38946 46002 38958
rect 23314 38894 23326 38946
rect 23378 38894 23390 38946
rect 30370 38894 30382 38946
rect 30434 38894 30446 38946
rect 35074 38894 35086 38946
rect 35138 38894 35150 38946
rect 39330 38894 39342 38946
rect 39394 38894 39406 38946
rect 39554 38894 39566 38946
rect 39618 38894 39630 38946
rect 43250 38894 43262 38946
rect 43314 38894 43326 38946
rect 47842 38894 47854 38946
rect 47906 38894 47918 38946
rect 21310 38882 21362 38894
rect 25566 38882 25618 38894
rect 31054 38882 31106 38894
rect 45950 38882 46002 38894
rect 5742 38834 5794 38846
rect 1810 38782 1822 38834
rect 1874 38782 1886 38834
rect 5742 38770 5794 38782
rect 5854 38834 5906 38846
rect 5854 38770 5906 38782
rect 6302 38834 6354 38846
rect 6302 38770 6354 38782
rect 7086 38834 7138 38846
rect 10446 38834 10498 38846
rect 7522 38782 7534 38834
rect 7586 38782 7598 38834
rect 7086 38770 7138 38782
rect 10446 38770 10498 38782
rect 13246 38834 13298 38846
rect 15486 38834 15538 38846
rect 13794 38782 13806 38834
rect 13858 38782 13870 38834
rect 14914 38782 14926 38834
rect 14978 38782 14990 38834
rect 13246 38770 13298 38782
rect 15486 38770 15538 38782
rect 21534 38834 21586 38846
rect 21534 38770 21586 38782
rect 21982 38834 22034 38846
rect 29822 38834 29874 38846
rect 33406 38834 33458 38846
rect 26114 38782 26126 38834
rect 26178 38782 26190 38834
rect 30482 38782 30494 38834
rect 30546 38782 30558 38834
rect 31266 38782 31278 38834
rect 31330 38782 31342 38834
rect 21982 38770 22034 38782
rect 29822 38770 29874 38782
rect 33406 38770 33458 38782
rect 34078 38834 34130 38846
rect 34078 38770 34130 38782
rect 34414 38834 34466 38846
rect 39902 38834 39954 38846
rect 46286 38834 46338 38846
rect 35186 38782 35198 38834
rect 35250 38782 35262 38834
rect 35858 38782 35870 38834
rect 35922 38782 35934 38834
rect 41122 38782 41134 38834
rect 41186 38782 41198 38834
rect 42466 38782 42478 38834
rect 42530 38782 42542 38834
rect 34414 38770 34466 38782
rect 39902 38770 39954 38782
rect 46286 38770 46338 38782
rect 46734 38834 46786 38846
rect 47506 38782 47518 38834
rect 47570 38782 47582 38834
rect 46734 38770 46786 38782
rect 5182 38722 5234 38734
rect 2482 38670 2494 38722
rect 2546 38670 2558 38722
rect 4722 38670 4734 38722
rect 4786 38670 4798 38722
rect 5182 38658 5234 38670
rect 6078 38722 6130 38734
rect 6078 38658 6130 38670
rect 8990 38722 9042 38734
rect 8990 38658 9042 38670
rect 11342 38722 11394 38734
rect 11342 38658 11394 38670
rect 15598 38722 15650 38734
rect 15598 38658 15650 38670
rect 16830 38722 16882 38734
rect 16830 38658 16882 38670
rect 17838 38722 17890 38734
rect 17838 38658 17890 38670
rect 19854 38722 19906 38734
rect 24110 38722 24162 38734
rect 29486 38722 29538 38734
rect 42142 38722 42194 38734
rect 20178 38670 20190 38722
rect 20242 38670 20254 38722
rect 26898 38670 26910 38722
rect 26962 38670 26974 38722
rect 29026 38670 29038 38722
rect 29090 38670 29102 38722
rect 36530 38670 36542 38722
rect 36594 38670 36606 38722
rect 38658 38670 38670 38722
rect 38722 38670 38734 38722
rect 47070 38722 47122 38734
rect 19854 38658 19906 38670
rect 24110 38658 24162 38670
rect 29486 38658 29538 38670
rect 42142 38658 42194 38670
rect 45378 38643 45390 38695
rect 45442 38643 45454 38695
rect 47070 38658 47122 38670
rect 6862 38610 6914 38622
rect 6862 38546 6914 38558
rect 11678 38610 11730 38622
rect 13806 38610 13858 38622
rect 12338 38558 12350 38610
rect 12402 38558 12414 38610
rect 11678 38546 11730 38558
rect 13806 38546 13858 38558
rect 1344 38442 48608 38476
rect 1344 38390 4478 38442
rect 4530 38390 4582 38442
rect 4634 38390 4686 38442
rect 4738 38390 35198 38442
rect 35250 38390 35302 38442
rect 35354 38390 35406 38442
rect 35458 38390 48608 38442
rect 1344 38356 48608 38390
rect 7758 38274 7810 38286
rect 7758 38210 7810 38222
rect 20078 38274 20130 38286
rect 37550 38274 37602 38286
rect 23650 38222 23662 38274
rect 23714 38271 23726 38274
rect 24098 38271 24110 38274
rect 23714 38225 24110 38271
rect 23714 38222 23726 38225
rect 24098 38222 24110 38225
rect 24162 38271 24174 38274
rect 24322 38271 24334 38274
rect 24162 38225 24334 38271
rect 24162 38222 24174 38225
rect 24322 38222 24334 38225
rect 24386 38222 24398 38274
rect 20078 38210 20130 38222
rect 37550 38210 37602 38222
rect 2270 38162 2322 38174
rect 2270 38098 2322 38110
rect 2718 38162 2770 38174
rect 4846 38162 4898 38174
rect 7646 38162 7698 38174
rect 3602 38110 3614 38162
rect 3666 38110 3678 38162
rect 6178 38110 6190 38162
rect 6242 38110 6254 38162
rect 2718 38098 2770 38110
rect 4846 38098 4898 38110
rect 7646 38098 7698 38110
rect 8318 38162 8370 38174
rect 8318 38098 8370 38110
rect 8654 38162 8706 38174
rect 13694 38162 13746 38174
rect 9874 38110 9886 38162
rect 9938 38110 9950 38162
rect 12786 38110 12798 38162
rect 12850 38110 12862 38162
rect 8654 38098 8706 38110
rect 13694 38098 13746 38110
rect 17390 38162 17442 38174
rect 17390 38098 17442 38110
rect 18622 38162 18674 38174
rect 18622 38098 18674 38110
rect 19406 38162 19458 38174
rect 19406 38098 19458 38110
rect 23662 38162 23714 38174
rect 23662 38098 23714 38110
rect 24110 38162 24162 38174
rect 32622 38162 32674 38174
rect 38894 38162 38946 38174
rect 42590 38162 42642 38174
rect 30034 38110 30046 38162
rect 30098 38110 30110 38162
rect 32162 38110 32174 38162
rect 32226 38110 32238 38162
rect 34514 38110 34526 38162
rect 34578 38110 34590 38162
rect 42130 38110 42142 38162
rect 42194 38110 42206 38162
rect 24110 38098 24162 38110
rect 32622 38098 32674 38110
rect 38894 38098 38946 38110
rect 42590 38098 42642 38110
rect 44942 38162 44994 38174
rect 48178 38110 48190 38162
rect 48242 38110 48254 38162
rect 44942 38098 44994 38110
rect 1710 38050 1762 38062
rect 1710 37986 1762 37998
rect 2830 38050 2882 38062
rect 2830 37986 2882 37998
rect 3278 38050 3330 38062
rect 8094 38050 8146 38062
rect 6514 37998 6526 38050
rect 6578 37998 6590 38050
rect 3278 37986 3330 37998
rect 8094 37986 8146 37998
rect 8542 38050 8594 38062
rect 11118 38050 11170 38062
rect 16494 38050 16546 38062
rect 9650 37998 9662 38050
rect 9714 37998 9726 38050
rect 11442 37998 11454 38050
rect 11506 37998 11518 38050
rect 12002 37998 12014 38050
rect 12066 37998 12078 38050
rect 12338 37998 12350 38050
rect 12402 37998 12414 38050
rect 14690 37998 14702 38050
rect 14754 37998 14766 38050
rect 15026 37998 15038 38050
rect 15090 37998 15102 38050
rect 15810 37998 15822 38050
rect 15874 37998 15886 38050
rect 16258 37998 16270 38050
rect 16322 37998 16334 38050
rect 8542 37986 8594 37998
rect 11118 37986 11170 37998
rect 16494 37986 16546 37998
rect 16718 38050 16770 38062
rect 16718 37986 16770 37998
rect 16830 38050 16882 38062
rect 16830 37986 16882 37998
rect 19854 38050 19906 38062
rect 19854 37986 19906 37998
rect 20302 38050 20354 38062
rect 20302 37986 20354 37998
rect 21198 38050 21250 38062
rect 21198 37986 21250 37998
rect 27694 38050 27746 38062
rect 43374 38050 43426 38062
rect 29362 37998 29374 38050
rect 29426 37998 29438 38050
rect 34850 37998 34862 38050
rect 34914 37998 34926 38050
rect 36194 37998 36206 38050
rect 36258 37998 36270 38050
rect 39218 37998 39230 38050
rect 39282 37998 39294 38050
rect 45266 37998 45278 38050
rect 45330 37998 45342 38050
rect 27694 37986 27746 37998
rect 43374 37986 43426 37998
rect 4174 37938 4226 37950
rect 7086 37938 7138 37950
rect 4498 37886 4510 37938
rect 4562 37886 4574 37938
rect 4174 37874 4226 37886
rect 7086 37874 7138 37886
rect 7534 37938 7586 37950
rect 7534 37874 7586 37886
rect 10334 37938 10386 37950
rect 10334 37874 10386 37886
rect 11230 37938 11282 37950
rect 13582 37938 13634 37950
rect 12450 37886 12462 37938
rect 12514 37886 12526 37938
rect 11230 37874 11282 37886
rect 13582 37874 13634 37886
rect 14366 37938 14418 37950
rect 14366 37874 14418 37886
rect 15710 37938 15762 37950
rect 15710 37874 15762 37886
rect 17502 37938 17554 37950
rect 17502 37874 17554 37886
rect 17950 37938 18002 37950
rect 17950 37874 18002 37886
rect 18062 37938 18114 37950
rect 18062 37874 18114 37886
rect 18510 37938 18562 37950
rect 18510 37874 18562 37886
rect 18734 37938 18786 37950
rect 18734 37874 18786 37886
rect 21646 37938 21698 37950
rect 21646 37874 21698 37886
rect 22654 37938 22706 37950
rect 22654 37874 22706 37886
rect 27358 37938 27410 37950
rect 27358 37874 27410 37886
rect 36430 37938 36482 37950
rect 36430 37874 36482 37886
rect 37214 37938 37266 37950
rect 37762 37886 37774 37938
rect 37826 37886 37838 37938
rect 38210 37886 38222 37938
rect 38274 37886 38286 37938
rect 40002 37886 40014 37938
rect 40066 37886 40078 37938
rect 43698 37886 43710 37938
rect 43762 37886 43774 37938
rect 44146 37886 44158 37938
rect 44210 37886 44222 37938
rect 46050 37886 46062 37938
rect 46114 37886 46126 37938
rect 37214 37874 37266 37886
rect 2606 37826 2658 37838
rect 2606 37762 2658 37774
rect 3614 37826 3666 37838
rect 3614 37762 3666 37774
rect 3726 37826 3778 37838
rect 3726 37762 3778 37774
rect 3950 37826 4002 37838
rect 3950 37762 4002 37774
rect 8766 37826 8818 37838
rect 13806 37826 13858 37838
rect 10658 37774 10670 37826
rect 10722 37774 10734 37826
rect 8766 37762 8818 37774
rect 13806 37762 13858 37774
rect 14030 37826 14082 37838
rect 14030 37762 14082 37774
rect 16606 37826 16658 37838
rect 16606 37762 16658 37774
rect 17726 37826 17778 37838
rect 17726 37762 17778 37774
rect 20750 37826 20802 37838
rect 20750 37762 20802 37774
rect 21758 37826 21810 37838
rect 21758 37762 21810 37774
rect 21870 37826 21922 37838
rect 21870 37762 21922 37774
rect 22318 37826 22370 37838
rect 22318 37762 22370 37774
rect 22766 37826 22818 37838
rect 22766 37762 22818 37774
rect 22990 37826 23042 37838
rect 22990 37762 23042 37774
rect 24670 37826 24722 37838
rect 24670 37762 24722 37774
rect 43038 37826 43090 37838
rect 43038 37762 43090 37774
rect 1344 37658 48608 37692
rect 1344 37606 19838 37658
rect 19890 37606 19942 37658
rect 19994 37606 20046 37658
rect 20098 37606 48608 37658
rect 1344 37572 48608 37606
rect 3614 37490 3666 37502
rect 3614 37426 3666 37438
rect 6078 37490 6130 37502
rect 6078 37426 6130 37438
rect 6190 37490 6242 37502
rect 15822 37490 15874 37502
rect 11106 37438 11118 37490
rect 11170 37438 11182 37490
rect 11778 37438 11790 37490
rect 11842 37438 11854 37490
rect 6190 37426 6242 37438
rect 15822 37426 15874 37438
rect 16046 37490 16098 37502
rect 16046 37426 16098 37438
rect 19518 37490 19570 37502
rect 19518 37426 19570 37438
rect 31054 37490 31106 37502
rect 39454 37490 39506 37502
rect 35410 37438 35422 37490
rect 35474 37438 35486 37490
rect 31054 37426 31106 37438
rect 39454 37426 39506 37438
rect 39902 37490 39954 37502
rect 39902 37426 39954 37438
rect 40350 37490 40402 37502
rect 40350 37426 40402 37438
rect 41022 37490 41074 37502
rect 41022 37426 41074 37438
rect 41694 37490 41746 37502
rect 41694 37426 41746 37438
rect 2046 37378 2098 37390
rect 2046 37314 2098 37326
rect 3054 37378 3106 37390
rect 3054 37314 3106 37326
rect 3838 37378 3890 37390
rect 3838 37314 3890 37326
rect 7310 37378 7362 37390
rect 7310 37314 7362 37326
rect 8206 37378 8258 37390
rect 14142 37378 14194 37390
rect 8978 37326 8990 37378
rect 9042 37326 9054 37378
rect 10098 37326 10110 37378
rect 10162 37326 10174 37378
rect 11666 37326 11678 37378
rect 11730 37326 11742 37378
rect 8206 37314 8258 37326
rect 14142 37314 14194 37326
rect 15710 37378 15762 37390
rect 17614 37378 17666 37390
rect 16370 37326 16382 37378
rect 16434 37326 16446 37378
rect 15710 37314 15762 37326
rect 17614 37314 17666 37326
rect 17726 37378 17778 37390
rect 17726 37314 17778 37326
rect 19406 37378 19458 37390
rect 23438 37378 23490 37390
rect 21634 37326 21646 37378
rect 21698 37326 21710 37378
rect 19406 37314 19458 37326
rect 23438 37314 23490 37326
rect 23550 37378 23602 37390
rect 23550 37314 23602 37326
rect 23774 37378 23826 37390
rect 23774 37314 23826 37326
rect 24222 37378 24274 37390
rect 24222 37314 24274 37326
rect 29150 37378 29202 37390
rect 37774 37378 37826 37390
rect 31602 37326 31614 37378
rect 31666 37326 31678 37378
rect 32162 37326 32174 37378
rect 32226 37326 32238 37378
rect 29150 37314 29202 37326
rect 37774 37314 37826 37326
rect 1710 37266 1762 37278
rect 1710 37202 1762 37214
rect 3950 37266 4002 37278
rect 5630 37266 5682 37278
rect 4610 37214 4622 37266
rect 4674 37214 4686 37266
rect 4834 37214 4846 37266
rect 4898 37214 4910 37266
rect 3950 37202 4002 37214
rect 5630 37202 5682 37214
rect 5966 37266 6018 37278
rect 5966 37202 6018 37214
rect 6638 37266 6690 37278
rect 6638 37202 6690 37214
rect 8094 37266 8146 37278
rect 9886 37266 9938 37278
rect 17390 37266 17442 37278
rect 8754 37214 8766 37266
rect 8818 37214 8830 37266
rect 10546 37214 10558 37266
rect 10610 37214 10622 37266
rect 10994 37214 11006 37266
rect 11058 37214 11070 37266
rect 11554 37214 11566 37266
rect 11618 37214 11630 37266
rect 13570 37214 13582 37266
rect 13634 37214 13646 37266
rect 16594 37214 16606 37266
rect 16658 37214 16670 37266
rect 8094 37202 8146 37214
rect 9886 37202 9938 37214
rect 17390 37202 17442 37214
rect 19070 37266 19122 37278
rect 24334 37266 24386 37278
rect 20178 37214 20190 37266
rect 20242 37214 20254 37266
rect 20514 37214 20526 37266
rect 20578 37214 20590 37266
rect 21074 37214 21086 37266
rect 21138 37214 21150 37266
rect 21522 37214 21534 37266
rect 21586 37214 21598 37266
rect 22418 37214 22430 37266
rect 22482 37214 22494 37266
rect 22978 37214 22990 37266
rect 23042 37214 23054 37266
rect 19070 37202 19122 37214
rect 24334 37202 24386 37214
rect 29486 37266 29538 37278
rect 29486 37202 29538 37214
rect 31390 37266 31442 37278
rect 31390 37202 31442 37214
rect 35758 37266 35810 37278
rect 37538 37214 37550 37266
rect 37602 37214 37614 37266
rect 41458 37214 41470 37266
rect 41522 37214 41534 37266
rect 44930 37214 44942 37266
rect 44994 37214 45006 37266
rect 45826 37214 45838 37266
rect 45890 37214 45902 37266
rect 35758 37202 35810 37214
rect 2494 37154 2546 37166
rect 2494 37090 2546 37102
rect 3502 37154 3554 37166
rect 7086 37154 7138 37166
rect 4722 37102 4734 37154
rect 4786 37102 4798 37154
rect 3502 37090 3554 37102
rect 7086 37090 7138 37102
rect 18286 37154 18338 37166
rect 18286 37090 18338 37102
rect 18622 37154 18674 37166
rect 36206 37154 36258 37166
rect 21858 37102 21870 37154
rect 21922 37102 21934 37154
rect 23426 37102 23438 37154
rect 23490 37102 23502 37154
rect 42018 37102 42030 37154
rect 42082 37102 42094 37154
rect 44146 37102 44158 37154
rect 44210 37102 44222 37154
rect 18622 37090 18674 37102
rect 36206 37090 36258 37102
rect 7422 37042 7474 37054
rect 6738 36990 6750 37042
rect 6802 37039 6814 37042
rect 6962 37039 6974 37042
rect 6802 36993 6974 37039
rect 6802 36990 6814 36993
rect 6962 36990 6974 36993
rect 7026 36990 7038 37042
rect 7422 36978 7474 36990
rect 8206 37042 8258 37054
rect 24222 37042 24274 37054
rect 18610 36990 18622 37042
rect 18674 37039 18686 37042
rect 19058 37039 19070 37042
rect 18674 36993 19070 37039
rect 18674 36990 18686 36993
rect 19058 36990 19070 36993
rect 19122 36990 19134 37042
rect 20850 36990 20862 37042
rect 20914 36990 20926 37042
rect 8206 36978 8258 36990
rect 24222 36978 24274 36990
rect 47966 37042 48018 37054
rect 47966 36978 48018 36990
rect 1344 36874 48608 36908
rect 1344 36822 4478 36874
rect 4530 36822 4582 36874
rect 4634 36822 4686 36874
rect 4738 36822 35198 36874
rect 35250 36822 35302 36874
rect 35354 36822 35406 36874
rect 35458 36822 48608 36874
rect 1344 36788 48608 36822
rect 12798 36706 12850 36718
rect 11554 36654 11566 36706
rect 11618 36654 11630 36706
rect 12798 36642 12850 36654
rect 41694 36706 41746 36718
rect 41694 36642 41746 36654
rect 43822 36706 43874 36718
rect 43822 36642 43874 36654
rect 4610 36568 4622 36620
rect 4674 36568 4686 36620
rect 5070 36594 5122 36606
rect 7422 36594 7474 36606
rect 6290 36542 6302 36594
rect 6354 36542 6366 36594
rect 5070 36530 5122 36542
rect 7422 36530 7474 36542
rect 13694 36594 13746 36606
rect 13694 36530 13746 36542
rect 14590 36594 14642 36606
rect 28030 36594 28082 36606
rect 22642 36542 22654 36594
rect 22706 36542 22718 36594
rect 26898 36542 26910 36594
rect 26962 36542 26974 36594
rect 29810 36542 29822 36594
rect 29874 36542 29886 36594
rect 35410 36542 35422 36594
rect 35474 36542 35486 36594
rect 37762 36542 37774 36594
rect 37826 36542 37838 36594
rect 39890 36542 39902 36594
rect 39954 36542 39966 36594
rect 14590 36530 14642 36542
rect 28030 36530 28082 36542
rect 7534 36482 7586 36494
rect 1810 36430 1822 36482
rect 1874 36430 1886 36482
rect 5954 36430 5966 36482
rect 6018 36430 6030 36482
rect 6626 36430 6638 36482
rect 6690 36430 6702 36482
rect 7534 36418 7586 36430
rect 9998 36482 10050 36494
rect 11006 36482 11058 36494
rect 10770 36430 10782 36482
rect 10834 36430 10846 36482
rect 9998 36418 10050 36430
rect 11006 36418 11058 36430
rect 11118 36482 11170 36494
rect 11118 36418 11170 36430
rect 12910 36482 12962 36494
rect 29262 36482 29314 36494
rect 36318 36482 36370 36494
rect 18498 36430 18510 36482
rect 18562 36430 18574 36482
rect 20738 36430 20750 36482
rect 20802 36430 20814 36482
rect 21410 36430 21422 36482
rect 21474 36430 21486 36482
rect 23202 36430 23214 36482
rect 23266 36430 23278 36482
rect 24098 36430 24110 36482
rect 24162 36430 24174 36482
rect 27458 36430 27470 36482
rect 27522 36430 27534 36482
rect 31602 36430 31614 36482
rect 31666 36430 31678 36482
rect 32610 36430 32622 36482
rect 32674 36430 32686 36482
rect 37090 36430 37102 36482
rect 37154 36430 37166 36482
rect 42466 36430 42478 36482
rect 42530 36430 42542 36482
rect 43138 36430 43150 36482
rect 43202 36430 43214 36482
rect 45042 36430 45054 36482
rect 45106 36430 45118 36482
rect 45602 36430 45614 36482
rect 45666 36430 45678 36482
rect 12910 36418 12962 36430
rect 29262 36418 29314 36430
rect 36318 36418 36370 36430
rect 9774 36370 9826 36382
rect 2482 36318 2494 36370
rect 2546 36318 2558 36370
rect 6178 36318 6190 36370
rect 6242 36318 6254 36370
rect 9774 36306 9826 36318
rect 9886 36370 9938 36382
rect 9886 36306 9938 36318
rect 12798 36370 12850 36382
rect 16606 36370 16658 36382
rect 19518 36370 19570 36382
rect 14914 36318 14926 36370
rect 14978 36318 14990 36370
rect 16370 36318 16382 36370
rect 16434 36318 16446 36370
rect 17042 36318 17054 36370
rect 17106 36318 17118 36370
rect 12798 36306 12850 36318
rect 16606 36306 16658 36318
rect 19518 36306 19570 36318
rect 22318 36370 22370 36382
rect 40350 36370 40402 36382
rect 24770 36318 24782 36370
rect 24834 36318 24846 36370
rect 33282 36318 33294 36370
rect 33346 36318 33358 36370
rect 22318 36306 22370 36318
rect 40350 36306 40402 36318
rect 40686 36370 40738 36382
rect 40686 36306 40738 36318
rect 41358 36370 41410 36382
rect 44158 36370 44210 36382
rect 42242 36318 42254 36370
rect 42306 36318 42318 36370
rect 43026 36318 43038 36370
rect 43090 36318 43102 36370
rect 41358 36306 41410 36318
rect 44158 36306 44210 36318
rect 44830 36370 44882 36382
rect 47394 36318 47406 36370
rect 47458 36318 47470 36370
rect 44830 36306 44882 36318
rect 7310 36258 7362 36270
rect 7310 36194 7362 36206
rect 7758 36258 7810 36270
rect 7758 36194 7810 36206
rect 8542 36258 8594 36270
rect 8542 36194 8594 36206
rect 8878 36258 8930 36270
rect 8878 36194 8930 36206
rect 9438 36258 9490 36270
rect 12350 36258 12402 36270
rect 10434 36206 10446 36258
rect 10498 36206 10510 36258
rect 9438 36194 9490 36206
rect 12350 36194 12402 36206
rect 13806 36258 13858 36270
rect 21758 36258 21810 36270
rect 17154 36206 17166 36258
rect 17218 36206 17230 36258
rect 13806 36194 13858 36206
rect 21758 36194 21810 36206
rect 21870 36258 21922 36270
rect 21870 36194 21922 36206
rect 21982 36258 22034 36270
rect 35758 36258 35810 36270
rect 27234 36206 27246 36258
rect 27298 36206 27310 36258
rect 21982 36194 22034 36206
rect 35758 36194 35810 36206
rect 1344 36090 48608 36124
rect 1344 36038 19838 36090
rect 19890 36038 19942 36090
rect 19994 36038 20046 36090
rect 20098 36038 48608 36090
rect 1344 36004 48608 36038
rect 2270 35922 2322 35934
rect 2270 35858 2322 35870
rect 2382 35922 2434 35934
rect 2382 35858 2434 35870
rect 5630 35922 5682 35934
rect 5630 35858 5682 35870
rect 5854 35922 5906 35934
rect 5854 35858 5906 35870
rect 6862 35922 6914 35934
rect 6862 35858 6914 35870
rect 9774 35922 9826 35934
rect 9774 35858 9826 35870
rect 11678 35922 11730 35934
rect 11678 35858 11730 35870
rect 19294 35922 19346 35934
rect 24334 35922 24386 35934
rect 19954 35870 19966 35922
rect 20018 35870 20030 35922
rect 19294 35858 19346 35870
rect 24334 35858 24386 35870
rect 24558 35922 24610 35934
rect 24558 35858 24610 35870
rect 25342 35922 25394 35934
rect 25342 35858 25394 35870
rect 31278 35922 31330 35934
rect 31278 35858 31330 35870
rect 33294 35922 33346 35934
rect 33294 35858 33346 35870
rect 33742 35922 33794 35934
rect 33742 35858 33794 35870
rect 37886 35922 37938 35934
rect 37886 35858 37938 35870
rect 40126 35922 40178 35934
rect 40126 35858 40178 35870
rect 41246 35922 41298 35934
rect 41246 35858 41298 35870
rect 41694 35922 41746 35934
rect 41694 35858 41746 35870
rect 8094 35810 8146 35822
rect 4834 35758 4846 35810
rect 4898 35758 4910 35810
rect 8094 35746 8146 35758
rect 10222 35810 10274 35822
rect 10222 35746 10274 35758
rect 10894 35810 10946 35822
rect 16046 35810 16098 35822
rect 11330 35758 11342 35810
rect 11394 35758 11406 35810
rect 13458 35758 13470 35810
rect 13522 35758 13534 35810
rect 14690 35758 14702 35810
rect 14754 35758 14766 35810
rect 10894 35746 10946 35758
rect 16046 35746 16098 35758
rect 17614 35810 17666 35822
rect 17614 35746 17666 35758
rect 17726 35810 17778 35822
rect 17726 35746 17778 35758
rect 19406 35810 19458 35822
rect 24222 35810 24274 35822
rect 20514 35758 20526 35810
rect 20578 35758 20590 35810
rect 22978 35758 22990 35810
rect 23042 35758 23054 35810
rect 19406 35746 19458 35758
rect 24222 35746 24274 35758
rect 26014 35810 26066 35822
rect 26338 35758 26350 35810
rect 26402 35758 26414 35810
rect 28690 35758 28702 35810
rect 28754 35758 28766 35810
rect 31938 35758 31950 35810
rect 32002 35758 32014 35810
rect 32386 35758 32398 35810
rect 32450 35758 32462 35810
rect 35298 35758 35310 35810
rect 35362 35758 35374 35810
rect 35522 35758 35534 35810
rect 35586 35758 35598 35810
rect 38770 35758 38782 35810
rect 38834 35758 38846 35810
rect 45714 35758 45726 35810
rect 45778 35758 45790 35810
rect 26014 35746 26066 35758
rect 2494 35698 2546 35710
rect 2494 35634 2546 35646
rect 2942 35698 2994 35710
rect 2942 35634 2994 35646
rect 3390 35698 3442 35710
rect 3390 35634 3442 35646
rect 3726 35698 3778 35710
rect 3726 35634 3778 35646
rect 5742 35698 5794 35710
rect 6638 35698 6690 35710
rect 6066 35646 6078 35698
rect 6130 35646 6142 35698
rect 6402 35646 6414 35698
rect 6466 35646 6478 35698
rect 5742 35634 5794 35646
rect 6638 35634 6690 35646
rect 6974 35698 7026 35710
rect 6974 35634 7026 35646
rect 7646 35698 7698 35710
rect 7646 35634 7698 35646
rect 7870 35698 7922 35710
rect 7870 35634 7922 35646
rect 8430 35698 8482 35710
rect 8430 35634 8482 35646
rect 8654 35698 8706 35710
rect 8654 35634 8706 35646
rect 9662 35698 9714 35710
rect 9662 35634 9714 35646
rect 9998 35698 10050 35710
rect 16718 35698 16770 35710
rect 12002 35646 12014 35698
rect 12066 35646 12078 35698
rect 15026 35646 15038 35698
rect 15090 35646 15102 35698
rect 9998 35634 10050 35646
rect 16158 35642 16210 35654
rect 16370 35646 16382 35698
rect 16434 35646 16446 35698
rect 1934 35586 1986 35598
rect 7982 35586 8034 35598
rect 16718 35634 16770 35646
rect 17950 35698 18002 35710
rect 18734 35698 18786 35710
rect 31614 35698 31666 35710
rect 18274 35646 18286 35698
rect 18338 35646 18350 35698
rect 20402 35646 20414 35698
rect 20466 35646 20478 35698
rect 22194 35646 22206 35698
rect 22258 35646 22270 35698
rect 23538 35646 23550 35698
rect 23602 35646 23614 35698
rect 26226 35646 26238 35698
rect 26290 35646 26302 35698
rect 26674 35646 26686 35698
rect 26738 35646 26750 35698
rect 27346 35646 27358 35698
rect 27410 35646 27422 35698
rect 28018 35646 28030 35698
rect 28082 35646 28094 35698
rect 17950 35634 18002 35646
rect 18734 35634 18786 35646
rect 31614 35634 31666 35646
rect 34078 35698 34130 35710
rect 34078 35634 34130 35646
rect 34638 35698 34690 35710
rect 34638 35634 34690 35646
rect 34974 35698 35026 35710
rect 34974 35634 35026 35646
rect 38222 35698 38274 35710
rect 38994 35646 39006 35698
rect 39058 35646 39070 35698
rect 44594 35646 44606 35698
rect 44658 35646 44670 35698
rect 45042 35646 45054 35698
rect 45106 35646 45118 35698
rect 38222 35634 38274 35646
rect 4498 35534 4510 35586
rect 4562 35534 4574 35586
rect 13682 35534 13694 35586
rect 13746 35534 13758 35586
rect 16158 35578 16210 35590
rect 30818 35534 30830 35586
rect 30882 35534 30894 35586
rect 47842 35534 47854 35586
rect 47906 35534 47918 35586
rect 1934 35522 1986 35534
rect 7982 35522 8034 35534
rect 3278 35474 3330 35486
rect 10782 35474 10834 35486
rect 16830 35474 16882 35486
rect 43598 35474 43650 35486
rect 8978 35422 8990 35474
rect 9042 35422 9054 35474
rect 15586 35422 15598 35474
rect 15650 35422 15662 35474
rect 41234 35422 41246 35474
rect 41298 35471 41310 35474
rect 41794 35471 41806 35474
rect 41298 35425 41806 35471
rect 41298 35422 41310 35425
rect 41794 35422 41806 35425
rect 41858 35422 41870 35474
rect 3278 35410 3330 35422
rect 10782 35410 10834 35422
rect 16830 35410 16882 35422
rect 43598 35410 43650 35422
rect 1344 35306 48608 35340
rect 1344 35254 4478 35306
rect 4530 35254 4582 35306
rect 4634 35254 4686 35306
rect 4738 35254 35198 35306
rect 35250 35254 35302 35306
rect 35354 35254 35406 35306
rect 35458 35254 48608 35306
rect 1344 35220 48608 35254
rect 5854 35138 5906 35150
rect 5854 35074 5906 35086
rect 8094 35138 8146 35150
rect 8094 35074 8146 35086
rect 25902 35138 25954 35150
rect 25902 35074 25954 35086
rect 2270 35026 2322 35038
rect 2270 34962 2322 34974
rect 3950 35026 4002 35038
rect 3950 34962 4002 34974
rect 5070 35026 5122 35038
rect 5070 34962 5122 34974
rect 5630 35026 5682 35038
rect 5630 34962 5682 34974
rect 7646 35026 7698 35038
rect 7646 34962 7698 34974
rect 8654 35026 8706 35038
rect 14254 35026 14306 35038
rect 17278 35026 17330 35038
rect 21422 35026 21474 35038
rect 32846 35026 32898 35038
rect 41806 35026 41858 35038
rect 12002 34974 12014 35026
rect 12066 34974 12078 35026
rect 14914 34974 14926 35026
rect 14978 34974 14990 35026
rect 17714 34974 17726 35026
rect 17778 34974 17790 35026
rect 22866 34974 22878 35026
rect 22930 34974 22942 35026
rect 32050 34974 32062 35026
rect 32114 34974 32126 35026
rect 39778 34974 39790 35026
rect 39842 34974 39854 35026
rect 8654 34962 8706 34974
rect 14254 34962 14306 34974
rect 17278 34962 17330 34974
rect 21422 34962 21474 34974
rect 32846 34962 32898 34974
rect 41806 34962 41858 34974
rect 8206 34914 8258 34926
rect 1810 34862 1822 34914
rect 1874 34862 1886 34914
rect 2706 34862 2718 34914
rect 2770 34862 2782 34914
rect 8206 34850 8258 34862
rect 9438 34914 9490 34926
rect 12910 34914 12962 34926
rect 9650 34862 9662 34914
rect 9714 34862 9726 34914
rect 10098 34862 10110 34914
rect 10162 34862 10174 34914
rect 10882 34862 10894 34914
rect 10946 34862 10958 34914
rect 11330 34862 11342 34914
rect 11394 34862 11406 34914
rect 12226 34862 12238 34914
rect 12290 34862 12302 34914
rect 9438 34850 9490 34862
rect 12910 34850 12962 34862
rect 13806 34914 13858 34926
rect 13806 34850 13858 34862
rect 14030 34914 14082 34926
rect 15710 34914 15762 34926
rect 15250 34862 15262 34914
rect 15314 34862 15326 34914
rect 14030 34850 14082 34862
rect 15710 34850 15762 34862
rect 16382 34914 16434 34926
rect 16382 34850 16434 34862
rect 16606 34914 16658 34926
rect 18510 34914 18562 34926
rect 17938 34862 17950 34914
rect 18002 34862 18014 34914
rect 16606 34850 16658 34862
rect 18510 34850 18562 34862
rect 19070 34914 19122 34926
rect 19070 34850 19122 34862
rect 19630 34914 19682 34926
rect 21310 34914 21362 34926
rect 26126 34914 26178 34926
rect 20066 34862 20078 34914
rect 20130 34862 20142 34914
rect 21746 34862 21758 34914
rect 21810 34862 21822 34914
rect 22082 34862 22094 34914
rect 22146 34862 22158 34914
rect 22978 34862 22990 34914
rect 23042 34862 23054 34914
rect 19630 34850 19682 34862
rect 21310 34850 21362 34862
rect 26126 34850 26178 34862
rect 26910 34914 26962 34926
rect 41134 34914 41186 34926
rect 29138 34862 29150 34914
rect 29202 34862 29214 34914
rect 33506 34862 33518 34914
rect 33570 34862 33582 34914
rect 34626 34862 34638 34914
rect 34690 34862 34702 34914
rect 37538 34862 37550 34914
rect 37602 34862 37614 34914
rect 26910 34850 26962 34862
rect 41134 34850 41186 34862
rect 42814 34914 42866 34926
rect 42814 34850 42866 34862
rect 43150 34914 43202 34926
rect 43922 34862 43934 34914
rect 43986 34862 43998 34914
rect 45826 34862 45838 34914
rect 45890 34862 45902 34914
rect 43150 34850 43202 34862
rect 3278 34802 3330 34814
rect 3278 34738 3330 34750
rect 3390 34802 3442 34814
rect 7422 34802 7474 34814
rect 7186 34750 7198 34802
rect 7250 34750 7262 34802
rect 3390 34738 3442 34750
rect 7422 34738 7474 34750
rect 7534 34802 7586 34814
rect 7534 34738 7586 34750
rect 8990 34802 9042 34814
rect 11678 34802 11730 34814
rect 10210 34750 10222 34802
rect 10274 34750 10286 34802
rect 8990 34738 9042 34750
rect 11678 34738 11730 34750
rect 13582 34802 13634 34814
rect 15486 34802 15538 34814
rect 15138 34750 15150 34802
rect 15202 34750 15214 34802
rect 13582 34738 13634 34750
rect 15486 34738 15538 34750
rect 16046 34802 16098 34814
rect 16046 34738 16098 34750
rect 19518 34802 19570 34814
rect 19518 34738 19570 34750
rect 21534 34802 21586 34814
rect 21534 34738 21586 34750
rect 22542 34802 22594 34814
rect 22542 34738 22594 34750
rect 24670 34802 24722 34814
rect 26686 34802 26738 34814
rect 44942 34802 44994 34814
rect 26450 34750 26462 34802
rect 26514 34750 26526 34802
rect 29922 34750 29934 34802
rect 29986 34750 29998 34802
rect 33394 34750 33406 34802
rect 33458 34750 33470 34802
rect 43810 34750 43822 34802
rect 43874 34750 43886 34802
rect 47170 34750 47182 34802
rect 47234 34750 47246 34802
rect 24670 34738 24722 34750
rect 26686 34738 26738 34750
rect 44942 34738 44994 34750
rect 2942 34690 2994 34702
rect 2942 34626 2994 34638
rect 3614 34690 3666 34702
rect 3614 34626 3666 34638
rect 3838 34690 3890 34702
rect 3838 34626 3890 34638
rect 4734 34690 4786 34702
rect 6638 34690 6690 34702
rect 6178 34638 6190 34690
rect 6242 34638 6254 34690
rect 4734 34626 4786 34638
rect 6638 34626 6690 34638
rect 7758 34690 7810 34702
rect 7758 34626 7810 34638
rect 9214 34690 9266 34702
rect 9214 34626 9266 34638
rect 9326 34690 9378 34702
rect 9326 34626 9378 34638
rect 14702 34690 14754 34702
rect 14702 34626 14754 34638
rect 16382 34690 16434 34702
rect 16382 34626 16434 34638
rect 18958 34690 19010 34702
rect 18958 34626 19010 34638
rect 19182 34690 19234 34702
rect 19182 34626 19234 34638
rect 24110 34690 24162 34702
rect 24110 34626 24162 34638
rect 24782 34690 24834 34702
rect 24782 34626 24834 34638
rect 25006 34690 25058 34702
rect 25006 34626 25058 34638
rect 25342 34690 25394 34702
rect 25342 34626 25394 34638
rect 32510 34690 32562 34702
rect 32510 34626 32562 34638
rect 34862 34690 34914 34702
rect 34862 34626 34914 34638
rect 37102 34690 37154 34702
rect 37102 34626 37154 34638
rect 40910 34690 40962 34702
rect 40910 34626 40962 34638
rect 41470 34690 41522 34702
rect 41470 34626 41522 34638
rect 42366 34690 42418 34702
rect 42366 34626 42418 34638
rect 45278 34690 45330 34702
rect 45278 34626 45330 34638
rect 1344 34522 48608 34556
rect 1344 34470 19838 34522
rect 19890 34470 19942 34522
rect 19994 34470 20046 34522
rect 20098 34470 48608 34522
rect 1344 34436 48608 34470
rect 2942 34354 2994 34366
rect 2594 34302 2606 34354
rect 2658 34302 2670 34354
rect 2942 34290 2994 34302
rect 3614 34354 3666 34366
rect 3614 34290 3666 34302
rect 4734 34354 4786 34366
rect 4734 34290 4786 34302
rect 6414 34354 6466 34366
rect 6414 34290 6466 34302
rect 6750 34354 6802 34366
rect 6750 34290 6802 34302
rect 10446 34354 10498 34366
rect 32062 34354 32114 34366
rect 13234 34302 13246 34354
rect 13298 34302 13310 34354
rect 10446 34290 10498 34302
rect 32062 34290 32114 34302
rect 45166 34354 45218 34366
rect 45166 34290 45218 34302
rect 3502 34242 3554 34254
rect 3502 34178 3554 34190
rect 3726 34242 3778 34254
rect 3726 34178 3778 34190
rect 6862 34242 6914 34254
rect 6862 34178 6914 34190
rect 8206 34242 8258 34254
rect 8206 34178 8258 34190
rect 8766 34242 8818 34254
rect 8766 34178 8818 34190
rect 8878 34242 8930 34254
rect 8878 34178 8930 34190
rect 9550 34242 9602 34254
rect 13582 34242 13634 34254
rect 12450 34190 12462 34242
rect 12514 34190 12526 34242
rect 9550 34178 9602 34190
rect 13582 34178 13634 34190
rect 15598 34242 15650 34254
rect 28814 34242 28866 34254
rect 18946 34190 18958 34242
rect 19010 34190 19022 34242
rect 21074 34190 21086 34242
rect 21138 34190 21150 34242
rect 21634 34190 21646 34242
rect 21698 34190 21710 34242
rect 15598 34178 15650 34190
rect 28814 34178 28866 34190
rect 32398 34242 32450 34254
rect 44158 34242 44210 34254
rect 36082 34190 36094 34242
rect 36146 34190 36158 34242
rect 41682 34190 41694 34242
rect 41746 34190 41758 34242
rect 32398 34178 32450 34190
rect 44158 34178 44210 34190
rect 1710 34130 1762 34142
rect 1710 34066 1762 34078
rect 3390 34130 3442 34142
rect 7982 34130 8034 34142
rect 4162 34078 4174 34130
rect 4226 34078 4238 34130
rect 5058 34078 5070 34130
rect 5122 34078 5134 34130
rect 3390 34066 3442 34078
rect 7982 34066 8034 34078
rect 8318 34130 8370 34142
rect 10222 34130 10274 34142
rect 12798 34130 12850 34142
rect 17950 34130 18002 34142
rect 20750 34130 20802 34142
rect 24110 34130 24162 34142
rect 9986 34078 9998 34130
rect 10050 34078 10062 34130
rect 10658 34078 10670 34130
rect 10722 34078 10734 34130
rect 11442 34078 11454 34130
rect 11506 34078 11518 34130
rect 12002 34078 12014 34130
rect 12066 34078 12078 34130
rect 12562 34078 12574 34130
rect 12626 34078 12638 34130
rect 13010 34078 13022 34130
rect 13074 34078 13086 34130
rect 15026 34078 15038 34130
rect 15090 34078 15102 34130
rect 19170 34078 19182 34130
rect 19234 34078 19246 34130
rect 19842 34078 19854 34130
rect 19906 34078 19918 34130
rect 21858 34078 21870 34130
rect 21922 34078 21934 34130
rect 22978 34078 22990 34130
rect 23042 34078 23054 34130
rect 8318 34066 8370 34078
rect 10222 34066 10274 34078
rect 12798 34066 12850 34078
rect 17950 34066 18002 34078
rect 20750 34066 20802 34078
rect 24110 34066 24162 34078
rect 24334 34130 24386 34142
rect 24334 34066 24386 34078
rect 24782 34130 24834 34142
rect 25218 34078 25230 34130
rect 25282 34078 25294 34130
rect 28578 34078 28590 34130
rect 28642 34078 28654 34130
rect 29362 34078 29374 34130
rect 29426 34078 29438 34130
rect 33170 34078 33182 34130
rect 33234 34078 33246 34130
rect 36866 34078 36878 34130
rect 36930 34078 36942 34130
rect 37426 34078 37438 34130
rect 37490 34078 37502 34130
rect 40898 34078 40910 34130
rect 40962 34078 40974 34130
rect 44594 34078 44606 34130
rect 44658 34078 44670 34130
rect 47954 34078 47966 34130
rect 48018 34078 48030 34130
rect 24782 34066 24834 34078
rect 2270 34018 2322 34030
rect 2270 33954 2322 33966
rect 5518 34018 5570 34030
rect 7310 34018 7362 34030
rect 5954 33966 5966 34018
rect 6018 33966 6030 34018
rect 5518 33954 5570 33966
rect 7310 33954 7362 33966
rect 7758 34018 7810 34030
rect 7758 33954 7810 33966
rect 9662 34018 9714 34030
rect 17390 34018 17442 34030
rect 10546 33966 10558 34018
rect 10610 33966 10622 34018
rect 9662 33954 9714 33966
rect 17390 33954 17442 33966
rect 20526 34018 20578 34030
rect 20526 33954 20578 33966
rect 22318 34018 22370 34030
rect 23774 34018 23826 34030
rect 23090 33966 23102 34018
rect 23154 33966 23166 34018
rect 22318 33954 22370 33966
rect 23774 33954 23826 33966
rect 24222 34018 24274 34030
rect 26002 33966 26014 34018
rect 26066 33966 26078 34018
rect 28130 33966 28142 34018
rect 28194 33966 28206 34018
rect 30258 33966 30270 34018
rect 30322 33966 30334 34018
rect 33506 33966 33518 34018
rect 33570 33966 33582 34018
rect 33954 33966 33966 34018
rect 34018 33966 34030 34018
rect 38098 33966 38110 34018
rect 38162 33966 38174 34018
rect 40226 33966 40238 34018
rect 40290 33966 40302 34018
rect 43810 33966 43822 34018
rect 43874 33966 43886 34018
rect 24222 33954 24274 33966
rect 8878 33906 8930 33918
rect 7186 33854 7198 33906
rect 7250 33903 7262 33906
rect 7858 33903 7870 33906
rect 7250 33857 7870 33903
rect 7250 33854 7262 33857
rect 7858 33854 7870 33857
rect 7922 33854 7934 33906
rect 46274 33854 46286 33906
rect 46338 33854 46350 33906
rect 8878 33842 8930 33854
rect 1344 33738 48608 33772
rect 1344 33686 4478 33738
rect 4530 33686 4582 33738
rect 4634 33686 4686 33738
rect 4738 33686 35198 33738
rect 35250 33686 35302 33738
rect 35354 33686 35406 33738
rect 35458 33686 48608 33738
rect 1344 33652 48608 33686
rect 3838 33570 3890 33582
rect 3838 33506 3890 33518
rect 34862 33570 34914 33582
rect 34862 33506 34914 33518
rect 3614 33458 3666 33470
rect 3614 33394 3666 33406
rect 4174 33458 4226 33470
rect 21310 33458 21362 33470
rect 9874 33406 9886 33458
rect 9938 33406 9950 33458
rect 17714 33406 17726 33458
rect 17778 33406 17790 33458
rect 19730 33406 19742 33458
rect 19794 33406 19806 33458
rect 4174 33394 4226 33406
rect 21310 33394 21362 33406
rect 24334 33458 24386 33470
rect 33406 33458 33458 33470
rect 29922 33406 29934 33458
rect 29986 33406 29998 33458
rect 32050 33406 32062 33458
rect 32114 33406 32126 33458
rect 24334 33394 24386 33406
rect 33406 33394 33458 33406
rect 45054 33458 45106 33470
rect 46050 33406 46062 33458
rect 46114 33406 46126 33458
rect 48178 33406 48190 33458
rect 48242 33406 48254 33458
rect 45054 33394 45106 33406
rect 3278 33346 3330 33358
rect 2818 33294 2830 33346
rect 2882 33294 2894 33346
rect 3278 33282 3330 33294
rect 4846 33346 4898 33358
rect 11790 33346 11842 33358
rect 6626 33294 6638 33346
rect 6690 33294 6702 33346
rect 7522 33294 7534 33346
rect 7586 33294 7598 33346
rect 8530 33294 8542 33346
rect 8594 33294 8606 33346
rect 9986 33294 9998 33346
rect 10050 33294 10062 33346
rect 10322 33294 10334 33346
rect 10386 33294 10398 33346
rect 11106 33294 11118 33346
rect 11170 33294 11182 33346
rect 4846 33282 4898 33294
rect 11790 33282 11842 33294
rect 12350 33346 12402 33358
rect 22206 33346 22258 33358
rect 14018 33294 14030 33346
rect 14082 33294 14094 33346
rect 15698 33294 15710 33346
rect 15762 33294 15774 33346
rect 16258 33294 16270 33346
rect 16322 33294 16334 33346
rect 16818 33294 16830 33346
rect 16882 33294 16894 33346
rect 18498 33294 18510 33346
rect 18562 33294 18574 33346
rect 19282 33294 19294 33346
rect 19346 33294 19358 33346
rect 21746 33294 21758 33346
rect 21810 33294 21822 33346
rect 12350 33282 12402 33294
rect 22206 33282 22258 33294
rect 23102 33346 23154 33358
rect 23102 33282 23154 33294
rect 23214 33346 23266 33358
rect 23214 33282 23266 33294
rect 23662 33346 23714 33358
rect 26350 33346 26402 33358
rect 32958 33346 33010 33358
rect 23874 33294 23886 33346
rect 23938 33294 23950 33346
rect 29250 33294 29262 33346
rect 29314 33294 29326 33346
rect 23662 33282 23714 33294
rect 26350 33282 26402 33294
rect 32958 33282 33010 33294
rect 35198 33346 35250 33358
rect 35746 33294 35758 33346
rect 35810 33294 35822 33346
rect 37538 33294 37550 33346
rect 37602 33294 37614 33346
rect 40674 33294 40686 33346
rect 40738 33294 40750 33346
rect 41682 33294 41694 33346
rect 41746 33294 41758 33346
rect 45378 33294 45390 33346
rect 45442 33294 45454 33346
rect 35198 33282 35250 33294
rect 1710 33234 1762 33246
rect 12910 33234 12962 33246
rect 14814 33234 14866 33246
rect 24222 33234 24274 33246
rect 32398 33234 32450 33246
rect 6514 33182 6526 33234
rect 6578 33182 6590 33234
rect 9538 33182 9550 33234
rect 9602 33182 9614 33234
rect 11554 33182 11566 33234
rect 11618 33182 11630 33234
rect 1710 33170 1762 33182
rect 12238 33178 12290 33190
rect 2046 33122 2098 33134
rect 2046 33058 2098 33070
rect 4510 33122 4562 33134
rect 8766 33122 8818 33134
rect 8082 33070 8094 33122
rect 8146 33070 8158 33122
rect 4510 33058 4562 33070
rect 8766 33058 8818 33070
rect 11678 33122 11730 33134
rect 11678 33058 11730 33070
rect 12014 33122 12066 33134
rect 14130 33182 14142 33234
rect 14194 33182 14206 33234
rect 15586 33182 15598 33234
rect 15650 33182 15662 33234
rect 26002 33182 26014 33234
rect 26066 33182 26078 33234
rect 35970 33182 35982 33234
rect 36034 33182 36046 33234
rect 39330 33182 39342 33234
rect 39394 33182 39406 33234
rect 43474 33182 43486 33234
rect 43538 33182 43550 33234
rect 12910 33170 12962 33182
rect 14814 33170 14866 33182
rect 24222 33170 24274 33182
rect 32398 33170 32450 33182
rect 12238 33114 12290 33126
rect 12574 33122 12626 33134
rect 12014 33058 12066 33070
rect 12574 33058 12626 33070
rect 12798 33122 12850 33134
rect 12798 33058 12850 33070
rect 13694 33122 13746 33134
rect 13694 33058 13746 33070
rect 22990 33122 23042 33134
rect 22990 33058 23042 33070
rect 24446 33122 24498 33134
rect 24446 33058 24498 33070
rect 24894 33122 24946 33134
rect 24894 33058 24946 33070
rect 25342 33122 25394 33134
rect 25342 33058 25394 33070
rect 28590 33122 28642 33134
rect 28590 33058 28642 33070
rect 37214 33122 37266 33134
rect 37214 33058 37266 33070
rect 40462 33122 40514 33134
rect 40462 33058 40514 33070
rect 1344 32954 48608 32988
rect 1344 32902 19838 32954
rect 19890 32902 19942 32954
rect 19994 32902 20046 32954
rect 20098 32902 48608 32954
rect 1344 32868 48608 32902
rect 4510 32786 4562 32798
rect 4510 32722 4562 32734
rect 4734 32786 4786 32798
rect 4734 32722 4786 32734
rect 6190 32786 6242 32798
rect 6190 32722 6242 32734
rect 6302 32786 6354 32798
rect 6302 32722 6354 32734
rect 7646 32786 7698 32798
rect 7646 32722 7698 32734
rect 8094 32786 8146 32798
rect 8094 32722 8146 32734
rect 15710 32786 15762 32798
rect 15710 32722 15762 32734
rect 16718 32786 16770 32798
rect 16718 32722 16770 32734
rect 18958 32786 19010 32798
rect 31166 32786 31218 32798
rect 22754 32734 22766 32786
rect 22818 32734 22830 32786
rect 18958 32722 19010 32734
rect 31166 32722 31218 32734
rect 40238 32786 40290 32798
rect 40238 32722 40290 32734
rect 42254 32786 42306 32798
rect 42254 32722 42306 32734
rect 2830 32674 2882 32686
rect 2830 32610 2882 32622
rect 2942 32674 2994 32686
rect 2942 32610 2994 32622
rect 3054 32674 3106 32686
rect 3054 32610 3106 32622
rect 3950 32674 4002 32686
rect 3950 32610 4002 32622
rect 10334 32674 10386 32686
rect 10334 32610 10386 32622
rect 10670 32674 10722 32686
rect 10670 32610 10722 32622
rect 15822 32674 15874 32686
rect 15822 32610 15874 32622
rect 17502 32674 17554 32686
rect 17502 32610 17554 32622
rect 21982 32674 22034 32686
rect 21982 32610 22034 32622
rect 23214 32674 23266 32686
rect 23214 32610 23266 32622
rect 23886 32674 23938 32686
rect 23886 32610 23938 32622
rect 23998 32674 24050 32686
rect 23998 32610 24050 32622
rect 26238 32674 26290 32686
rect 26238 32610 26290 32622
rect 29822 32674 29874 32686
rect 36990 32674 37042 32686
rect 32274 32622 32286 32674
rect 32338 32622 32350 32674
rect 29822 32610 29874 32622
rect 36990 32610 37042 32622
rect 38670 32674 38722 32686
rect 39106 32622 39118 32674
rect 39170 32622 39182 32674
rect 39666 32622 39678 32674
rect 39730 32622 39742 32674
rect 41346 32622 41358 32674
rect 41410 32622 41422 32674
rect 41570 32622 41582 32674
rect 41634 32622 41646 32674
rect 38670 32610 38722 32622
rect 3838 32562 3890 32574
rect 1810 32510 1822 32562
rect 1874 32510 1886 32562
rect 3838 32498 3890 32510
rect 4174 32562 4226 32574
rect 4174 32498 4226 32510
rect 4398 32562 4450 32574
rect 4398 32498 4450 32510
rect 5742 32562 5794 32574
rect 5742 32498 5794 32510
rect 6414 32562 6466 32574
rect 6414 32498 6466 32510
rect 7870 32562 7922 32574
rect 15486 32562 15538 32574
rect 9986 32510 9998 32562
rect 10050 32510 10062 32562
rect 11778 32510 11790 32562
rect 11842 32510 11854 32562
rect 13234 32510 13246 32562
rect 13298 32510 13310 32562
rect 13906 32510 13918 32562
rect 13970 32510 13982 32562
rect 15026 32510 15038 32562
rect 15090 32510 15102 32562
rect 7870 32498 7922 32510
rect 15486 32498 15538 32510
rect 16158 32562 16210 32574
rect 16158 32498 16210 32510
rect 19630 32562 19682 32574
rect 19630 32498 19682 32510
rect 22094 32562 22146 32574
rect 22094 32498 22146 32510
rect 23326 32562 23378 32574
rect 23326 32498 23378 32510
rect 23438 32562 23490 32574
rect 23438 32498 23490 32510
rect 24222 32562 24274 32574
rect 24222 32498 24274 32510
rect 26574 32562 26626 32574
rect 31502 32562 31554 32574
rect 37326 32562 37378 32574
rect 39902 32562 39954 32574
rect 29586 32510 29598 32562
rect 29650 32510 29662 32562
rect 32162 32510 32174 32562
rect 32226 32510 32238 32562
rect 38434 32510 38446 32562
rect 38498 32510 38510 32562
rect 42690 32510 42702 32562
rect 42754 32510 42766 32562
rect 45602 32510 45614 32562
rect 45666 32510 45678 32562
rect 26574 32498 26626 32510
rect 31502 32498 31554 32510
rect 37326 32498 37378 32510
rect 39902 32498 39954 32510
rect 2270 32450 2322 32462
rect 2270 32386 2322 32398
rect 5070 32450 5122 32462
rect 5070 32386 5122 32398
rect 5630 32450 5682 32462
rect 5630 32386 5682 32398
rect 6974 32450 7026 32462
rect 6974 32386 7026 32398
rect 7310 32450 7362 32462
rect 7310 32386 7362 32398
rect 7758 32450 7810 32462
rect 7758 32386 7810 32398
rect 8990 32450 9042 32462
rect 8990 32386 9042 32398
rect 9662 32450 9714 32462
rect 18062 32450 18114 32462
rect 15138 32398 15150 32450
rect 15202 32398 15214 32450
rect 9662 32386 9714 32398
rect 18062 32386 18114 32398
rect 18398 32450 18450 32462
rect 18398 32386 18450 32398
rect 20190 32450 20242 32462
rect 20190 32386 20242 32398
rect 20974 32450 21026 32462
rect 20974 32386 21026 32398
rect 21310 32450 21362 32462
rect 21310 32386 21362 32398
rect 24558 32450 24610 32462
rect 24558 32386 24610 32398
rect 17390 32338 17442 32350
rect 3490 32286 3502 32338
rect 3554 32286 3566 32338
rect 17390 32274 17442 32286
rect 21982 32338 22034 32350
rect 21982 32274 22034 32286
rect 41918 32338 41970 32350
rect 41918 32274 41970 32286
rect 45054 32338 45106 32350
rect 47058 32286 47070 32338
rect 47122 32286 47134 32338
rect 45054 32274 45106 32286
rect 1344 32170 48608 32204
rect 1344 32118 4478 32170
rect 4530 32118 4582 32170
rect 4634 32118 4686 32170
rect 4738 32118 35198 32170
rect 35250 32118 35302 32170
rect 35354 32118 35406 32170
rect 35458 32118 48608 32170
rect 1344 32084 48608 32118
rect 8878 32002 8930 32014
rect 8878 31938 8930 31950
rect 11454 32002 11506 32014
rect 11454 31938 11506 31950
rect 37662 32002 37714 32014
rect 37662 31938 37714 31950
rect 9102 31890 9154 31902
rect 2146 31838 2158 31890
rect 2210 31838 2222 31890
rect 3378 31838 3390 31890
rect 3442 31838 3454 31890
rect 6626 31838 6638 31890
rect 6690 31838 6702 31890
rect 9102 31826 9154 31838
rect 9326 31890 9378 31902
rect 9326 31826 9378 31838
rect 11902 31890 11954 31902
rect 11902 31826 11954 31838
rect 21422 31890 21474 31902
rect 24210 31838 24222 31890
rect 24274 31838 24286 31890
rect 27906 31838 27918 31890
rect 27970 31838 27982 31890
rect 29922 31838 29934 31890
rect 29986 31838 29998 31890
rect 32050 31838 32062 31890
rect 32114 31838 32126 31890
rect 35298 31838 35310 31890
rect 35362 31838 35374 31890
rect 40002 31838 40014 31890
rect 40066 31838 40078 31890
rect 42130 31838 42142 31890
rect 42194 31838 42206 31890
rect 47730 31838 47742 31890
rect 47794 31838 47806 31890
rect 21422 31826 21474 31838
rect 1710 31778 1762 31790
rect 4510 31778 4562 31790
rect 3714 31726 3726 31778
rect 3778 31726 3790 31778
rect 4050 31726 4062 31778
rect 4114 31726 4126 31778
rect 1710 31714 1762 31726
rect 4510 31714 4562 31726
rect 4846 31778 4898 31790
rect 4846 31714 4898 31726
rect 5854 31778 5906 31790
rect 6974 31778 7026 31790
rect 6402 31726 6414 31778
rect 6466 31726 6478 31778
rect 5854 31714 5906 31726
rect 6974 31714 7026 31726
rect 8206 31778 8258 31790
rect 8206 31714 8258 31726
rect 9550 31778 9602 31790
rect 9550 31714 9602 31726
rect 9774 31778 9826 31790
rect 12126 31778 12178 31790
rect 10210 31726 10222 31778
rect 10274 31726 10286 31778
rect 10994 31726 11006 31778
rect 11058 31726 11070 31778
rect 11554 31726 11566 31778
rect 11618 31726 11630 31778
rect 9774 31714 9826 31726
rect 12126 31714 12178 31726
rect 12686 31778 12738 31790
rect 12686 31714 12738 31726
rect 12798 31778 12850 31790
rect 12798 31714 12850 31726
rect 14702 31778 14754 31790
rect 14702 31714 14754 31726
rect 16718 31778 16770 31790
rect 16718 31714 16770 31726
rect 17166 31778 17218 31790
rect 17166 31714 17218 31726
rect 19630 31778 19682 31790
rect 20190 31778 20242 31790
rect 19842 31726 19854 31778
rect 19906 31726 19918 31778
rect 19630 31714 19682 31726
rect 20190 31714 20242 31726
rect 20302 31778 20354 31790
rect 20302 31714 20354 31726
rect 20414 31778 20466 31790
rect 20414 31714 20466 31726
rect 20638 31778 20690 31790
rect 23102 31778 23154 31790
rect 22194 31726 22206 31778
rect 22258 31726 22270 31778
rect 20638 31714 20690 31726
rect 23102 31714 23154 31726
rect 23214 31778 23266 31790
rect 37998 31778 38050 31790
rect 43822 31778 43874 31790
rect 24546 31726 24558 31778
rect 24610 31726 24622 31778
rect 24994 31726 25006 31778
rect 25058 31726 25070 31778
rect 25778 31726 25790 31778
rect 25842 31726 25854 31778
rect 29138 31726 29150 31778
rect 29202 31726 29214 31778
rect 32386 31726 32398 31778
rect 32450 31726 32462 31778
rect 39330 31726 39342 31778
rect 39394 31726 39406 31778
rect 43138 31726 43150 31778
rect 43202 31726 43214 31778
rect 45714 31726 45726 31778
rect 45778 31726 45790 31778
rect 23214 31714 23266 31726
rect 37998 31714 38050 31726
rect 43822 31714 43874 31726
rect 4734 31666 4786 31678
rect 3266 31614 3278 31666
rect 3330 31614 3342 31666
rect 4734 31602 4786 31614
rect 7534 31666 7586 31678
rect 17726 31666 17778 31678
rect 22766 31666 22818 31678
rect 44158 31666 44210 31678
rect 8530 31614 8542 31666
rect 8594 31614 8606 31666
rect 11442 31614 11454 31666
rect 11506 31614 11518 31666
rect 12450 31614 12462 31666
rect 12514 31614 12526 31666
rect 13906 31614 13918 31666
rect 13970 31614 13982 31666
rect 14242 31614 14254 31666
rect 14306 31614 14318 31666
rect 15138 31614 15150 31666
rect 15202 31614 15214 31666
rect 22418 31614 22430 31666
rect 22482 31614 22494 31666
rect 33170 31614 33182 31666
rect 33234 31614 33246 31666
rect 38210 31614 38222 31666
rect 38274 31614 38286 31666
rect 38770 31614 38782 31666
rect 38834 31614 38846 31666
rect 43250 31614 43262 31666
rect 43314 31614 43326 31666
rect 7534 31602 7586 31614
rect 17726 31602 17778 31614
rect 22766 31602 22818 31614
rect 44158 31602 44210 31614
rect 44830 31666 44882 31678
rect 44830 31602 44882 31614
rect 2830 31554 2882 31566
rect 2830 31490 2882 31502
rect 6638 31554 6690 31566
rect 6638 31490 6690 31502
rect 6862 31554 6914 31566
rect 6862 31490 6914 31502
rect 9662 31554 9714 31566
rect 19294 31554 19346 31566
rect 14578 31502 14590 31554
rect 14642 31502 14654 31554
rect 15250 31502 15262 31554
rect 15314 31502 15326 31554
rect 9662 31490 9714 31502
rect 19294 31490 19346 31502
rect 19406 31554 19458 31566
rect 19406 31490 19458 31502
rect 19518 31554 19570 31566
rect 19518 31490 19570 31502
rect 22990 31554 23042 31566
rect 22990 31490 23042 31502
rect 23774 31554 23826 31566
rect 23774 31490 23826 31502
rect 37214 31554 37266 31566
rect 37214 31490 37266 31502
rect 42702 31554 42754 31566
rect 42702 31490 42754 31502
rect 45166 31554 45218 31566
rect 45166 31490 45218 31502
rect 1344 31386 48608 31420
rect 1344 31334 19838 31386
rect 19890 31334 19942 31386
rect 19994 31334 20046 31386
rect 20098 31334 48608 31386
rect 1344 31300 48608 31334
rect 6078 31218 6130 31230
rect 6078 31154 6130 31166
rect 6526 31218 6578 31230
rect 6526 31154 6578 31166
rect 6750 31218 6802 31230
rect 10782 31218 10834 31230
rect 9538 31166 9550 31218
rect 9602 31166 9614 31218
rect 6750 31154 6802 31166
rect 10782 31154 10834 31166
rect 11118 31218 11170 31230
rect 11118 31154 11170 31166
rect 16718 31218 16770 31230
rect 22990 31218 23042 31230
rect 17714 31166 17726 31218
rect 17778 31166 17790 31218
rect 16718 31154 16770 31166
rect 22990 31154 23042 31166
rect 23550 31218 23602 31230
rect 23550 31154 23602 31166
rect 24558 31218 24610 31230
rect 24558 31154 24610 31166
rect 30718 31218 30770 31230
rect 30718 31154 30770 31166
rect 33406 31218 33458 31230
rect 41134 31218 41186 31230
rect 40002 31166 40014 31218
rect 40066 31166 40078 31218
rect 33406 31154 33458 31166
rect 41134 31154 41186 31166
rect 5294 31106 5346 31118
rect 2370 31054 2382 31106
rect 2434 31054 2446 31106
rect 3714 31054 3726 31106
rect 3778 31054 3790 31106
rect 5294 31042 5346 31054
rect 7086 31106 7138 31118
rect 7086 31042 7138 31054
rect 8878 31106 8930 31118
rect 8878 31042 8930 31054
rect 9774 31106 9826 31118
rect 14030 31106 14082 31118
rect 14590 31106 14642 31118
rect 13010 31054 13022 31106
rect 13074 31054 13086 31106
rect 14354 31054 14366 31106
rect 14418 31054 14430 31106
rect 9774 31042 9826 31054
rect 14030 31042 14082 31054
rect 14590 31042 14642 31054
rect 15598 31106 15650 31118
rect 29374 31106 29426 31118
rect 46062 31106 46114 31118
rect 22642 31054 22654 31106
rect 22706 31054 22718 31106
rect 31378 31054 31390 31106
rect 31442 31054 31454 31106
rect 31602 31054 31614 31106
rect 31666 31054 31678 31106
rect 34850 31054 34862 31106
rect 34914 31054 34926 31106
rect 35410 31054 35422 31106
rect 35474 31054 35486 31106
rect 36642 31054 36654 31106
rect 36706 31054 36718 31106
rect 41682 31054 41694 31106
rect 41746 31054 41758 31106
rect 42242 31054 42254 31106
rect 42306 31054 42318 31106
rect 44930 31054 44942 31106
rect 44994 31054 45006 31106
rect 47394 31054 47406 31106
rect 47458 31054 47470 31106
rect 47954 31054 47966 31106
rect 48018 31054 48030 31106
rect 15598 31042 15650 31054
rect 29374 31042 29426 31054
rect 46062 31042 46114 31054
rect 6414 30994 6466 31006
rect 4834 30942 4846 30994
rect 4898 30942 4910 30994
rect 5842 30942 5854 30994
rect 5906 30942 5918 30994
rect 6414 30930 6466 30942
rect 7982 30994 8034 31006
rect 7982 30930 8034 30942
rect 9550 30994 9602 31006
rect 9550 30930 9602 30942
rect 9998 30994 10050 31006
rect 9998 30930 10050 30942
rect 10110 30994 10162 31006
rect 14478 30994 14530 31006
rect 24446 30994 24498 31006
rect 11554 30942 11566 30994
rect 11618 30942 11630 30994
rect 11890 30942 11902 30994
rect 11954 30942 11966 30994
rect 15474 30942 15486 30994
rect 15538 30942 15550 30994
rect 16146 30942 16158 30994
rect 16210 30942 16222 30994
rect 16594 30942 16606 30994
rect 16658 30942 16670 30994
rect 17938 30942 17950 30994
rect 18002 30942 18014 30994
rect 18946 30942 18958 30994
rect 19010 30942 19022 30994
rect 21522 30942 21534 30994
rect 21586 30942 21598 30994
rect 21746 30942 21758 30994
rect 21810 30942 21822 30994
rect 10110 30930 10162 30942
rect 14478 30930 14530 30942
rect 24446 30930 24498 30942
rect 24782 30994 24834 31006
rect 29710 30994 29762 31006
rect 25330 30942 25342 30994
rect 25394 30942 25406 30994
rect 24782 30930 24834 30942
rect 29710 30930 29762 30942
rect 31054 30994 31106 31006
rect 31054 30930 31106 30942
rect 33742 30994 33794 31006
rect 33742 30930 33794 30942
rect 34302 30994 34354 31006
rect 34302 30930 34354 30942
rect 34638 30994 34690 31006
rect 41470 30994 41522 31006
rect 46398 30994 46450 31006
rect 35970 30942 35982 30994
rect 36034 30942 36046 30994
rect 40226 30942 40238 30994
rect 40290 30942 40302 30994
rect 45602 30942 45614 30994
rect 45666 30942 45678 30994
rect 34638 30930 34690 30942
rect 41470 30930 41522 30942
rect 46398 30930 46450 30942
rect 46846 30994 46898 31006
rect 46846 30930 46898 30942
rect 1934 30882 1986 30894
rect 1934 30818 1986 30830
rect 3950 30882 4002 30894
rect 8206 30882 8258 30894
rect 4946 30830 4958 30882
rect 5010 30830 5022 30882
rect 3950 30818 4002 30830
rect 8206 30818 8258 30830
rect 8430 30882 8482 30894
rect 21310 30882 21362 30894
rect 19506 30830 19518 30882
rect 19570 30830 19582 30882
rect 23986 30830 23998 30882
rect 24050 30830 24062 30882
rect 26002 30830 26014 30882
rect 26066 30830 26078 30882
rect 28130 30830 28142 30882
rect 28194 30830 28206 30882
rect 38770 30830 38782 30882
rect 38834 30830 38846 30882
rect 42802 30830 42814 30882
rect 42866 30830 42878 30882
rect 8430 30818 8482 30830
rect 21310 30818 21362 30830
rect 6974 30770 7026 30782
rect 6974 30706 7026 30718
rect 7310 30770 7362 30782
rect 7310 30706 7362 30718
rect 7758 30770 7810 30782
rect 7758 30706 7810 30718
rect 13694 30770 13746 30782
rect 13694 30706 13746 30718
rect 13806 30770 13858 30782
rect 13806 30706 13858 30718
rect 47182 30770 47234 30782
rect 47182 30706 47234 30718
rect 1344 30602 48608 30636
rect 1344 30550 4478 30602
rect 4530 30550 4582 30602
rect 4634 30550 4686 30602
rect 4738 30550 35198 30602
rect 35250 30550 35302 30602
rect 35354 30550 35406 30602
rect 35458 30550 48608 30602
rect 1344 30516 48608 30550
rect 12574 30434 12626 30446
rect 12574 30370 12626 30382
rect 19630 30434 19682 30446
rect 19630 30370 19682 30382
rect 20302 30434 20354 30446
rect 20302 30370 20354 30382
rect 5070 30322 5122 30334
rect 9662 30322 9714 30334
rect 13582 30322 13634 30334
rect 9426 30270 9438 30322
rect 9490 30270 9502 30322
rect 12898 30270 12910 30322
rect 12962 30270 12974 30322
rect 5070 30258 5122 30270
rect 9662 30258 9714 30270
rect 13582 30258 13634 30270
rect 14366 30322 14418 30334
rect 14366 30258 14418 30270
rect 16382 30322 16434 30334
rect 16382 30258 16434 30270
rect 17502 30322 17554 30334
rect 20638 30322 20690 30334
rect 34862 30322 34914 30334
rect 19394 30270 19406 30322
rect 19458 30270 19470 30322
rect 21746 30270 21758 30322
rect 21810 30270 21822 30322
rect 39890 30270 39902 30322
rect 39954 30270 39966 30322
rect 46050 30270 46062 30322
rect 46114 30270 46126 30322
rect 48178 30270 48190 30322
rect 48242 30270 48254 30322
rect 17502 30258 17554 30270
rect 20638 30258 20690 30270
rect 34862 30258 34914 30270
rect 7870 30210 7922 30222
rect 4274 30158 4286 30210
rect 4338 30158 4350 30210
rect 6402 30158 6414 30210
rect 6466 30158 6478 30210
rect 7870 30146 7922 30158
rect 8654 30210 8706 30222
rect 10558 30210 10610 30222
rect 8978 30158 8990 30210
rect 9042 30158 9054 30210
rect 8654 30146 8706 30158
rect 10558 30146 10610 30158
rect 11230 30210 11282 30222
rect 13470 30210 13522 30222
rect 11890 30158 11902 30210
rect 11954 30158 11966 30210
rect 11230 30146 11282 30158
rect 13470 30146 13522 30158
rect 13918 30210 13970 30222
rect 15710 30210 15762 30222
rect 15026 30158 15038 30210
rect 15090 30158 15102 30210
rect 13918 30146 13970 30158
rect 15710 30146 15762 30158
rect 16270 30210 16322 30222
rect 16270 30146 16322 30158
rect 17166 30210 17218 30222
rect 17166 30146 17218 30158
rect 18958 30210 19010 30222
rect 20750 30210 20802 30222
rect 22430 30210 22482 30222
rect 19954 30158 19966 30210
rect 20018 30158 20030 30210
rect 20514 30158 20526 30210
rect 20578 30158 20590 30210
rect 21858 30158 21870 30210
rect 21922 30158 21934 30210
rect 22194 30158 22206 30210
rect 22258 30158 22270 30210
rect 18958 30146 19010 30158
rect 20750 30146 20802 30158
rect 22430 30146 22482 30158
rect 22766 30210 22818 30222
rect 24110 30210 24162 30222
rect 23202 30158 23214 30210
rect 23266 30158 23278 30210
rect 22766 30146 22818 30158
rect 24110 30146 24162 30158
rect 24558 30210 24610 30222
rect 35634 30158 35646 30210
rect 35698 30158 35710 30210
rect 37090 30158 37102 30210
rect 37154 30158 37166 30210
rect 45378 30158 45390 30210
rect 45442 30158 45454 30210
rect 24558 30146 24610 30158
rect 8766 30098 8818 30110
rect 2482 30046 2494 30098
rect 2546 30046 2558 30098
rect 5954 30046 5966 30098
rect 6018 30046 6030 30098
rect 7634 30046 7646 30098
rect 7698 30046 7710 30098
rect 8766 30034 8818 30046
rect 11006 30098 11058 30110
rect 11006 30034 11058 30046
rect 13806 30098 13858 30110
rect 16046 30098 16098 30110
rect 14466 30046 14478 30098
rect 14530 30046 14542 30098
rect 14802 30046 14814 30098
rect 14866 30046 14878 30098
rect 13806 30034 13858 30046
rect 16046 30034 16098 30046
rect 16494 30098 16546 30110
rect 16494 30034 16546 30046
rect 21646 30098 21698 30110
rect 21646 30034 21698 30046
rect 23438 30098 23490 30110
rect 26798 30098 26850 30110
rect 23762 30046 23774 30098
rect 23826 30046 23838 30098
rect 23438 30034 23490 30046
rect 26798 30034 26850 30046
rect 30158 30098 30210 30110
rect 41246 30098 41298 30110
rect 35410 30046 35422 30098
rect 35474 30046 35486 30098
rect 37762 30046 37774 30098
rect 37826 30046 37838 30098
rect 30158 30034 30210 30046
rect 41246 30034 41298 30046
rect 10334 29986 10386 29998
rect 8194 29934 8206 29986
rect 8258 29934 8270 29986
rect 10334 29922 10386 29934
rect 10894 29986 10946 29998
rect 12798 29986 12850 29998
rect 12114 29934 12126 29986
rect 12178 29934 12190 29986
rect 10894 29922 10946 29934
rect 12798 29922 12850 29934
rect 15374 29986 15426 29998
rect 15374 29922 15426 29934
rect 15598 29986 15650 29998
rect 15598 29922 15650 29934
rect 16606 29986 16658 29998
rect 16606 29922 16658 29934
rect 18062 29986 18114 29998
rect 18062 29922 18114 29934
rect 18398 29986 18450 29998
rect 18398 29922 18450 29934
rect 19406 29986 19458 29998
rect 19406 29922 19458 29934
rect 21422 29986 21474 29998
rect 21422 29922 21474 29934
rect 22654 29986 22706 29998
rect 22654 29922 22706 29934
rect 26910 29986 26962 29998
rect 26910 29922 26962 29934
rect 27134 29986 27186 29998
rect 27134 29922 27186 29934
rect 29598 29986 29650 29998
rect 29598 29922 29650 29934
rect 34078 29986 34130 29998
rect 34078 29922 34130 29934
rect 34526 29986 34578 29998
rect 34526 29922 34578 29934
rect 41582 29986 41634 29998
rect 41582 29922 41634 29934
rect 44942 29986 44994 29998
rect 44942 29922 44994 29934
rect 1344 29818 48608 29852
rect 1344 29766 19838 29818
rect 19890 29766 19942 29818
rect 19994 29766 20046 29818
rect 20098 29766 48608 29818
rect 1344 29732 48608 29766
rect 9662 29650 9714 29662
rect 9662 29586 9714 29598
rect 11454 29650 11506 29662
rect 11454 29586 11506 29598
rect 11902 29650 11954 29662
rect 19070 29650 19122 29662
rect 18274 29598 18286 29650
rect 18338 29598 18350 29650
rect 11902 29586 11954 29598
rect 19070 29586 19122 29598
rect 19406 29650 19458 29662
rect 19406 29586 19458 29598
rect 20526 29650 20578 29662
rect 37774 29650 37826 29662
rect 22754 29598 22766 29650
rect 22818 29598 22830 29650
rect 26562 29598 26574 29650
rect 26626 29647 26638 29650
rect 26786 29647 26798 29650
rect 26626 29601 26798 29647
rect 26626 29598 26638 29601
rect 26786 29598 26798 29601
rect 26850 29598 26862 29650
rect 20526 29586 20578 29598
rect 37774 29586 37826 29598
rect 2718 29538 2770 29550
rect 2034 29486 2046 29538
rect 2098 29486 2110 29538
rect 2718 29474 2770 29486
rect 8318 29538 8370 29550
rect 8318 29474 8370 29486
rect 8878 29538 8930 29550
rect 16046 29538 16098 29550
rect 11106 29486 11118 29538
rect 11170 29486 11182 29538
rect 13010 29486 13022 29538
rect 13074 29486 13086 29538
rect 14242 29486 14254 29538
rect 14306 29486 14318 29538
rect 8878 29474 8930 29486
rect 16046 29474 16098 29486
rect 16382 29538 16434 29550
rect 16382 29474 16434 29486
rect 16830 29538 16882 29550
rect 16830 29474 16882 29486
rect 19518 29538 19570 29550
rect 27694 29538 27746 29550
rect 45278 29538 45330 29550
rect 22642 29486 22654 29538
rect 22706 29486 22718 29538
rect 24098 29486 24110 29538
rect 24162 29486 24174 29538
rect 26786 29486 26798 29538
rect 26850 29486 26862 29538
rect 27010 29486 27022 29538
rect 27074 29486 27086 29538
rect 29138 29486 29150 29538
rect 29202 29486 29214 29538
rect 39330 29486 39342 29538
rect 39394 29486 39406 29538
rect 41682 29486 41694 29538
rect 41746 29486 41758 29538
rect 19518 29474 19570 29486
rect 27694 29474 27746 29486
rect 45278 29474 45330 29486
rect 1710 29426 1762 29438
rect 1710 29362 1762 29374
rect 2494 29426 2546 29438
rect 2494 29362 2546 29374
rect 2606 29426 2658 29438
rect 8654 29426 8706 29438
rect 3154 29374 3166 29426
rect 3218 29374 3230 29426
rect 3490 29374 3502 29426
rect 3554 29374 3566 29426
rect 3826 29374 3838 29426
rect 3890 29374 3902 29426
rect 5394 29374 5406 29426
rect 5458 29374 5470 29426
rect 6738 29374 6750 29426
rect 6802 29374 6814 29426
rect 2606 29362 2658 29374
rect 8654 29362 8706 29374
rect 10782 29426 10834 29438
rect 17390 29426 17442 29438
rect 12450 29374 12462 29426
rect 12514 29374 12526 29426
rect 14018 29374 14030 29426
rect 14082 29374 14094 29426
rect 10782 29362 10834 29374
rect 17390 29362 17442 29374
rect 17950 29426 18002 29438
rect 38222 29426 38274 29438
rect 18498 29374 18510 29426
rect 18562 29374 18574 29426
rect 21746 29374 21758 29426
rect 21810 29374 21822 29426
rect 23762 29374 23774 29426
rect 23826 29374 23838 29426
rect 26562 29374 26574 29426
rect 26626 29374 26638 29426
rect 28466 29374 28478 29426
rect 28530 29374 28542 29426
rect 35970 29374 35982 29426
rect 36034 29374 36046 29426
rect 37538 29374 37550 29426
rect 37602 29374 37614 29426
rect 17950 29362 18002 29374
rect 38222 29362 38274 29374
rect 38558 29426 38610 29438
rect 39106 29374 39118 29426
rect 39170 29374 39182 29426
rect 41010 29374 41022 29426
rect 41074 29374 41086 29426
rect 45042 29374 45054 29426
rect 45106 29374 45118 29426
rect 45602 29374 45614 29426
rect 45666 29374 45678 29426
rect 38558 29362 38610 29374
rect 8430 29314 8482 29326
rect 6066 29262 6078 29314
rect 6130 29262 6142 29314
rect 6962 29262 6974 29314
rect 7026 29262 7038 29314
rect 8430 29250 8482 29262
rect 11790 29314 11842 29326
rect 18958 29314 19010 29326
rect 15026 29262 15038 29314
rect 15090 29262 15102 29314
rect 11790 29250 11842 29262
rect 18958 29250 19010 29262
rect 20078 29314 20130 29326
rect 39902 29314 39954 29326
rect 21298 29262 21310 29314
rect 21362 29262 21374 29314
rect 31266 29262 31278 29314
rect 31330 29262 31342 29314
rect 33058 29262 33070 29314
rect 33122 29262 33134 29314
rect 35186 29262 35198 29314
rect 35250 29262 35262 29314
rect 43810 29262 43822 29314
rect 43874 29262 43886 29314
rect 20078 29250 20130 29262
rect 39902 29250 39954 29262
rect 10110 29202 10162 29214
rect 10110 29138 10162 29150
rect 10334 29202 10386 29214
rect 10334 29138 10386 29150
rect 10558 29202 10610 29214
rect 10558 29138 10610 29150
rect 16718 29202 16770 29214
rect 16718 29138 16770 29150
rect 47966 29202 48018 29214
rect 47966 29138 48018 29150
rect 1344 29034 48608 29068
rect 1344 28982 4478 29034
rect 4530 28982 4582 29034
rect 4634 28982 4686 29034
rect 4738 28982 35198 29034
rect 35250 28982 35302 29034
rect 35354 28982 35406 29034
rect 35458 28982 48608 29034
rect 1344 28948 48608 28982
rect 5742 28866 5794 28878
rect 10446 28866 10498 28878
rect 7186 28814 7198 28866
rect 7250 28814 7262 28866
rect 5742 28802 5794 28814
rect 2718 28754 2770 28766
rect 7201 28751 7247 28814
rect 10446 28802 10498 28814
rect 25902 28866 25954 28878
rect 25902 28802 25954 28814
rect 30718 28866 30770 28878
rect 30718 28802 30770 28814
rect 35422 28866 35474 28878
rect 35422 28802 35474 28814
rect 41134 28866 41186 28878
rect 41134 28802 41186 28814
rect 41470 28866 41522 28878
rect 41470 28802 41522 28814
rect 43822 28866 43874 28878
rect 43822 28802 43874 28814
rect 19742 28754 19794 28766
rect 30270 28754 30322 28766
rect 7522 28751 7534 28754
rect 7201 28705 7534 28751
rect 7522 28702 7534 28705
rect 7586 28702 7598 28754
rect 12450 28702 12462 28754
rect 12514 28702 12526 28754
rect 13682 28702 13694 28754
rect 13746 28702 13758 28754
rect 17826 28702 17838 28754
rect 17890 28702 17902 28754
rect 20402 28702 20414 28754
rect 20466 28702 20478 28754
rect 29586 28702 29598 28754
rect 29650 28702 29662 28754
rect 2718 28690 2770 28702
rect 19742 28690 19794 28702
rect 30270 28690 30322 28702
rect 40686 28754 40738 28766
rect 40686 28690 40738 28702
rect 44158 28754 44210 28766
rect 47842 28702 47854 28754
rect 47906 28702 47918 28754
rect 44158 28690 44210 28702
rect 2158 28642 2210 28654
rect 2158 28578 2210 28590
rect 3054 28642 3106 28654
rect 5630 28642 5682 28654
rect 7534 28642 7586 28654
rect 4274 28590 4286 28642
rect 4338 28590 4350 28642
rect 4834 28590 4846 28642
rect 4898 28590 4910 28642
rect 6626 28590 6638 28642
rect 6690 28590 6702 28642
rect 6962 28590 6974 28642
rect 7026 28590 7038 28642
rect 3054 28578 3106 28590
rect 5630 28578 5682 28590
rect 7534 28578 7586 28590
rect 7982 28642 8034 28654
rect 7982 28578 8034 28590
rect 8094 28642 8146 28654
rect 9998 28642 10050 28654
rect 11230 28642 11282 28654
rect 17054 28642 17106 28654
rect 9762 28590 9774 28642
rect 9826 28590 9838 28642
rect 10546 28590 10558 28642
rect 10610 28590 10622 28642
rect 11778 28590 11790 28642
rect 11842 28590 11854 28642
rect 12338 28590 12350 28642
rect 12402 28590 12414 28642
rect 16034 28590 16046 28642
rect 16098 28590 16110 28642
rect 8094 28578 8146 28590
rect 9998 28578 10050 28590
rect 11230 28578 11282 28590
rect 17054 28578 17106 28590
rect 17390 28642 17442 28654
rect 17390 28578 17442 28590
rect 18958 28642 19010 28654
rect 23438 28642 23490 28654
rect 20178 28590 20190 28642
rect 20242 28590 20254 28642
rect 23090 28590 23102 28642
rect 23154 28590 23166 28642
rect 18958 28578 19010 28590
rect 23438 28578 23490 28590
rect 25790 28642 25842 28654
rect 31054 28642 31106 28654
rect 26226 28590 26238 28642
rect 26290 28590 26302 28642
rect 29250 28590 29262 28642
rect 29314 28590 29326 28642
rect 31826 28590 31838 28642
rect 31890 28590 31902 28642
rect 33170 28590 33182 28642
rect 33234 28590 33246 28642
rect 35858 28590 35870 28642
rect 35922 28590 35934 28642
rect 37762 28590 37774 28642
rect 37826 28590 37838 28642
rect 41906 28590 41918 28642
rect 41970 28590 41982 28642
rect 45042 28590 45054 28642
rect 45106 28590 45118 28642
rect 45602 28590 45614 28642
rect 45666 28590 45678 28642
rect 25790 28578 25842 28590
rect 31054 28578 31106 28590
rect 6190 28530 6242 28542
rect 3378 28478 3390 28530
rect 3442 28478 3454 28530
rect 4386 28478 4398 28530
rect 4450 28478 4462 28530
rect 6190 28466 6242 28478
rect 6414 28530 6466 28542
rect 6414 28466 6466 28478
rect 8206 28530 8258 28542
rect 8206 28466 8258 28478
rect 8766 28530 8818 28542
rect 20750 28530 20802 28542
rect 23998 28530 24050 28542
rect 27470 28530 27522 28542
rect 33406 28530 33458 28542
rect 12562 28478 12574 28530
rect 12626 28478 12638 28530
rect 16706 28478 16718 28530
rect 16770 28478 16782 28530
rect 21298 28478 21310 28530
rect 21362 28478 21374 28530
rect 26450 28478 26462 28530
rect 26514 28478 26526 28530
rect 26898 28478 26910 28530
rect 26962 28478 26974 28530
rect 31602 28478 31614 28530
rect 31666 28478 31678 28530
rect 36194 28478 36206 28530
rect 36258 28478 36270 28530
rect 37538 28478 37550 28530
rect 37602 28478 37614 28530
rect 39330 28478 39342 28530
rect 39394 28478 39406 28530
rect 42242 28478 42254 28530
rect 42306 28478 42318 28530
rect 43250 28478 43262 28530
rect 43314 28478 43326 28530
rect 43474 28478 43486 28530
rect 43538 28478 43550 28530
rect 8766 28466 8818 28478
rect 20750 28466 20802 28478
rect 23998 28466 24050 28478
rect 27470 28466 27522 28478
rect 33406 28466 33458 28478
rect 1934 28418 1986 28430
rect 6302 28418 6354 28430
rect 4946 28366 4958 28418
rect 5010 28366 5022 28418
rect 1934 28354 1986 28366
rect 6302 28354 6354 28366
rect 11678 28418 11730 28430
rect 11678 28354 11730 28366
rect 18398 28418 18450 28430
rect 35086 28418 35138 28430
rect 21522 28366 21534 28418
rect 21586 28366 21598 28418
rect 18398 28354 18450 28366
rect 35086 28354 35138 28366
rect 39678 28418 39730 28430
rect 39678 28354 39730 28366
rect 44830 28418 44882 28430
rect 44830 28354 44882 28366
rect 1344 28250 48608 28284
rect 1344 28198 19838 28250
rect 19890 28198 19942 28250
rect 19994 28198 20046 28250
rect 20098 28198 48608 28250
rect 1344 28164 48608 28198
rect 5182 28082 5234 28094
rect 5182 28018 5234 28030
rect 7758 28082 7810 28094
rect 7758 28018 7810 28030
rect 8430 28082 8482 28094
rect 8430 28018 8482 28030
rect 9438 28082 9490 28094
rect 9438 28018 9490 28030
rect 11566 28082 11618 28094
rect 11566 28018 11618 28030
rect 15038 28082 15090 28094
rect 15038 28018 15090 28030
rect 17502 28082 17554 28094
rect 26574 28082 26626 28094
rect 17826 28030 17838 28082
rect 17890 28030 17902 28082
rect 17502 28018 17554 28030
rect 26574 28018 26626 28030
rect 26686 28082 26738 28094
rect 42254 28082 42306 28094
rect 41570 28030 41582 28082
rect 41634 28030 41646 28082
rect 26686 28018 26738 28030
rect 42254 28018 42306 28030
rect 46062 28082 46114 28094
rect 46062 28018 46114 28030
rect 47630 28082 47682 28094
rect 47630 28018 47682 28030
rect 8094 27970 8146 27982
rect 15710 27970 15762 27982
rect 11218 27918 11230 27970
rect 11282 27918 11294 27970
rect 8094 27906 8146 27918
rect 15710 27906 15762 27918
rect 16606 27970 16658 27982
rect 16606 27906 16658 27918
rect 22206 27970 22258 27982
rect 22206 27906 22258 27918
rect 27134 27970 27186 27982
rect 43362 27918 43374 27970
rect 43426 27918 43438 27970
rect 46610 27918 46622 27970
rect 46674 27918 46686 27970
rect 27134 27906 27186 27918
rect 4958 27858 5010 27870
rect 1810 27806 1822 27858
rect 1874 27806 1886 27858
rect 4958 27794 5010 27806
rect 5630 27858 5682 27870
rect 7086 27858 7138 27870
rect 6626 27806 6638 27858
rect 6690 27806 6702 27858
rect 5630 27794 5682 27806
rect 7086 27794 7138 27806
rect 7198 27858 7250 27870
rect 14814 27858 14866 27870
rect 18398 27858 18450 27870
rect 22990 27858 23042 27870
rect 10098 27806 10110 27858
rect 10162 27806 10174 27858
rect 10434 27806 10446 27858
rect 10498 27806 10510 27858
rect 12450 27806 12462 27858
rect 12514 27806 12526 27858
rect 15362 27806 15374 27858
rect 15426 27806 15438 27858
rect 21298 27806 21310 27858
rect 21362 27806 21374 27858
rect 22754 27806 22766 27858
rect 22818 27806 22830 27858
rect 7198 27794 7250 27806
rect 14814 27794 14866 27806
rect 18398 27794 18450 27806
rect 22990 27794 23042 27806
rect 23438 27858 23490 27870
rect 41246 27858 41298 27870
rect 47294 27858 47346 27870
rect 24434 27806 24446 27858
rect 24498 27806 24510 27858
rect 27346 27806 27358 27858
rect 27410 27806 27422 27858
rect 29474 27806 29486 27858
rect 29538 27806 29550 27858
rect 33618 27806 33630 27858
rect 33682 27806 33694 27858
rect 37426 27806 37438 27858
rect 37490 27806 37502 27858
rect 42690 27806 42702 27858
rect 42754 27806 42766 27858
rect 46498 27806 46510 27858
rect 46562 27806 46574 27858
rect 23438 27794 23490 27806
rect 41246 27794 41298 27806
rect 47294 27794 47346 27806
rect 5070 27746 5122 27758
rect 8990 27746 9042 27758
rect 14926 27746 14978 27758
rect 2482 27694 2494 27746
rect 2546 27694 2558 27746
rect 4610 27694 4622 27746
rect 4674 27694 4686 27746
rect 6290 27694 6302 27746
rect 6354 27694 6366 27746
rect 9762 27694 9774 27746
rect 9826 27694 9838 27746
rect 13794 27694 13806 27746
rect 13858 27694 13870 27746
rect 5070 27682 5122 27694
rect 8990 27682 9042 27694
rect 14926 27682 14978 27694
rect 16046 27746 16098 27758
rect 23998 27746 24050 27758
rect 18834 27694 18846 27746
rect 18898 27694 18910 27746
rect 20290 27694 20302 27746
rect 20354 27694 20366 27746
rect 30258 27694 30270 27746
rect 30322 27694 30334 27746
rect 32386 27694 32398 27746
rect 32450 27694 32462 27746
rect 34402 27694 34414 27746
rect 34466 27694 34478 27746
rect 36530 27694 36542 27746
rect 36594 27694 36606 27746
rect 38210 27694 38222 27746
rect 38274 27694 38286 27746
rect 40338 27694 40350 27746
rect 40402 27694 40414 27746
rect 45490 27694 45502 27746
rect 45554 27694 45566 27746
rect 16046 27682 16098 27694
rect 23998 27682 24050 27694
rect 15822 27634 15874 27646
rect 15822 27570 15874 27582
rect 16158 27634 16210 27646
rect 16158 27570 16210 27582
rect 16718 27634 16770 27646
rect 16718 27570 16770 27582
rect 26462 27634 26514 27646
rect 26462 27570 26514 27582
rect 1344 27466 48608 27500
rect 1344 27414 4478 27466
rect 4530 27414 4582 27466
rect 4634 27414 4686 27466
rect 4738 27414 35198 27466
rect 35250 27414 35302 27466
rect 35354 27414 35406 27466
rect 35458 27414 48608 27466
rect 1344 27380 48608 27414
rect 12238 27298 12290 27310
rect 12238 27234 12290 27246
rect 31390 27298 31442 27310
rect 31390 27234 31442 27246
rect 2270 27186 2322 27198
rect 2270 27122 2322 27134
rect 5742 27186 5794 27198
rect 5742 27122 5794 27134
rect 6862 27186 6914 27198
rect 10222 27186 10274 27198
rect 9538 27134 9550 27186
rect 9602 27134 9614 27186
rect 6862 27122 6914 27134
rect 10222 27122 10274 27134
rect 11118 27186 11170 27198
rect 11118 27122 11170 27134
rect 13470 27186 13522 27198
rect 13470 27122 13522 27134
rect 15038 27186 15090 27198
rect 15038 27122 15090 27134
rect 20750 27186 20802 27198
rect 20750 27122 20802 27134
rect 23886 27186 23938 27198
rect 38334 27186 38386 27198
rect 26450 27134 26462 27186
rect 26514 27134 26526 27186
rect 28578 27134 28590 27186
rect 28642 27134 28654 27186
rect 40002 27134 40014 27186
rect 40066 27134 40078 27186
rect 46050 27134 46062 27186
rect 46114 27134 46126 27186
rect 48178 27134 48190 27186
rect 48242 27134 48254 27186
rect 23886 27122 23938 27134
rect 38334 27122 38386 27134
rect 4174 27074 4226 27086
rect 2930 27022 2942 27074
rect 2994 27022 3006 27074
rect 4174 27010 4226 27022
rect 4510 27074 4562 27086
rect 4510 27010 4562 27022
rect 5182 27074 5234 27086
rect 8318 27074 8370 27086
rect 6290 27022 6302 27074
rect 6354 27022 6366 27074
rect 7858 27022 7870 27074
rect 7922 27022 7934 27074
rect 5182 27010 5234 27022
rect 8318 27010 8370 27022
rect 8654 27074 8706 27086
rect 10558 27074 10610 27086
rect 9090 27022 9102 27074
rect 9154 27022 9166 27074
rect 8654 27010 8706 27022
rect 10558 27010 10610 27022
rect 11790 27074 11842 27086
rect 12910 27074 12962 27086
rect 15374 27074 15426 27086
rect 11890 27022 11902 27074
rect 11954 27022 11966 27074
rect 13682 27022 13694 27074
rect 13746 27022 13758 27074
rect 13906 27022 13918 27074
rect 13970 27022 13982 27074
rect 11790 27010 11842 27022
rect 12910 27010 12962 27022
rect 15374 27010 15426 27022
rect 15822 27074 15874 27086
rect 22990 27074 23042 27086
rect 18050 27022 18062 27074
rect 18114 27022 18126 27074
rect 19170 27022 19182 27074
rect 19234 27022 19246 27074
rect 20178 27022 20190 27074
rect 20242 27022 20254 27074
rect 20514 27022 20526 27074
rect 20578 27022 20590 27074
rect 15822 27010 15874 27022
rect 22990 27010 23042 27022
rect 23326 27074 23378 27086
rect 34750 27074 34802 27086
rect 25666 27022 25678 27074
rect 25730 27022 25742 27074
rect 23326 27010 23378 27022
rect 34750 27010 34802 27022
rect 37774 27074 37826 27086
rect 45378 27022 45390 27074
rect 45442 27022 45454 27074
rect 37774 27010 37826 27022
rect 1710 26962 1762 26974
rect 3502 26962 3554 26974
rect 3154 26910 3166 26962
rect 3218 26910 3230 26962
rect 1710 26898 1762 26910
rect 3502 26898 3554 26910
rect 3726 26962 3778 26974
rect 3726 26898 3778 26910
rect 4734 26962 4786 26974
rect 4734 26898 4786 26910
rect 5854 26962 5906 26974
rect 5854 26898 5906 26910
rect 5966 26962 6018 26974
rect 5966 26898 6018 26910
rect 6974 26962 7026 26974
rect 6974 26898 7026 26910
rect 7198 26962 7250 26974
rect 15710 26962 15762 26974
rect 8082 26910 8094 26962
rect 8146 26910 8158 26962
rect 12562 26910 12574 26962
rect 12626 26910 12638 26962
rect 7198 26898 7250 26910
rect 15710 26898 15762 26910
rect 16494 26962 16546 26974
rect 16494 26898 16546 26910
rect 16830 26962 16882 26974
rect 16830 26898 16882 26910
rect 17166 26962 17218 26974
rect 17166 26898 17218 26910
rect 17502 26962 17554 26974
rect 18734 26962 18786 26974
rect 17826 26910 17838 26962
rect 17890 26910 17902 26962
rect 17502 26898 17554 26910
rect 18734 26898 18786 26910
rect 21422 26962 21474 26974
rect 21422 26898 21474 26910
rect 21758 26962 21810 26974
rect 22430 26962 22482 26974
rect 22082 26910 22094 26962
rect 22146 26910 22158 26962
rect 21758 26898 21810 26910
rect 22430 26898 22482 26910
rect 24558 26962 24610 26974
rect 24558 26898 24610 26910
rect 30270 26962 30322 26974
rect 30270 26898 30322 26910
rect 30606 26962 30658 26974
rect 30606 26898 30658 26910
rect 31054 26962 31106 26974
rect 34414 26962 34466 26974
rect 31602 26910 31614 26962
rect 31666 26910 31678 26962
rect 32162 26910 32174 26962
rect 32226 26910 32238 26962
rect 31054 26898 31106 26910
rect 34414 26898 34466 26910
rect 39678 26962 39730 26974
rect 39678 26898 39730 26910
rect 39902 26962 39954 26974
rect 43922 26910 43934 26962
rect 43986 26910 43998 26962
rect 39902 26898 39954 26910
rect 3614 26850 3666 26862
rect 3614 26786 3666 26798
rect 4622 26850 4674 26862
rect 4622 26786 4674 26798
rect 5630 26850 5682 26862
rect 5630 26786 5682 26798
rect 6750 26850 6802 26862
rect 6750 26786 6802 26798
rect 11566 26850 11618 26862
rect 11566 26786 11618 26798
rect 11678 26850 11730 26862
rect 11678 26786 11730 26798
rect 15486 26850 15538 26862
rect 15486 26786 15538 26798
rect 18398 26850 18450 26862
rect 18398 26786 18450 26798
rect 18622 26850 18674 26862
rect 18622 26786 18674 26798
rect 19406 26850 19458 26862
rect 19406 26786 19458 26798
rect 24222 26850 24274 26862
rect 24222 26786 24274 26798
rect 44270 26850 44322 26862
rect 44270 26786 44322 26798
rect 1344 26682 48608 26716
rect 1344 26630 19838 26682
rect 19890 26630 19942 26682
rect 19994 26630 20046 26682
rect 20098 26630 48608 26682
rect 1344 26596 48608 26630
rect 2158 26514 2210 26526
rect 4734 26514 4786 26526
rect 4162 26462 4174 26514
rect 4226 26462 4238 26514
rect 2158 26450 2210 26462
rect 4734 26450 4786 26462
rect 4958 26514 5010 26526
rect 4958 26450 5010 26462
rect 5518 26514 5570 26526
rect 10558 26514 10610 26526
rect 8978 26462 8990 26514
rect 9042 26462 9054 26514
rect 5518 26450 5570 26462
rect 10558 26450 10610 26462
rect 11790 26514 11842 26526
rect 15822 26514 15874 26526
rect 12898 26462 12910 26514
rect 12962 26462 12974 26514
rect 11790 26450 11842 26462
rect 15822 26450 15874 26462
rect 16830 26514 16882 26526
rect 26686 26514 26738 26526
rect 22418 26462 22430 26514
rect 22482 26462 22494 26514
rect 16830 26450 16882 26462
rect 26686 26450 26738 26462
rect 39678 26514 39730 26526
rect 39678 26450 39730 26462
rect 5070 26402 5122 26414
rect 11342 26402 11394 26414
rect 7858 26350 7870 26402
rect 7922 26350 7934 26402
rect 5070 26338 5122 26350
rect 11342 26338 11394 26350
rect 12350 26402 12402 26414
rect 12350 26338 12402 26350
rect 16046 26402 16098 26414
rect 16046 26338 16098 26350
rect 17614 26402 17666 26414
rect 17614 26338 17666 26350
rect 18062 26402 18114 26414
rect 18062 26338 18114 26350
rect 18286 26402 18338 26414
rect 18286 26338 18338 26350
rect 18510 26402 18562 26414
rect 19954 26350 19966 26402
rect 20018 26350 20030 26402
rect 24546 26350 24558 26402
rect 24610 26350 24622 26402
rect 27794 26350 27806 26402
rect 27858 26350 27870 26402
rect 18510 26338 18562 26350
rect 2382 26290 2434 26302
rect 5854 26290 5906 26302
rect 8654 26290 8706 26302
rect 3378 26238 3390 26290
rect 3442 26238 3454 26290
rect 4386 26238 4398 26290
rect 4450 26238 4462 26290
rect 6962 26238 6974 26290
rect 7026 26238 7038 26290
rect 8082 26238 8094 26290
rect 8146 26238 8158 26290
rect 2382 26226 2434 26238
rect 5854 26226 5906 26238
rect 8654 26226 8706 26238
rect 9550 26290 9602 26302
rect 9550 26226 9602 26238
rect 9886 26290 9938 26302
rect 9886 26226 9938 26238
rect 9998 26290 10050 26302
rect 9998 26226 10050 26238
rect 10110 26290 10162 26302
rect 11566 26290 11618 26302
rect 10770 26238 10782 26290
rect 10834 26238 10846 26290
rect 10110 26226 10162 26238
rect 11566 26226 11618 26238
rect 11902 26290 11954 26302
rect 11902 26226 11954 26238
rect 12574 26290 12626 26302
rect 14926 26290 14978 26302
rect 13794 26238 13806 26290
rect 13858 26238 13870 26290
rect 12574 26226 12626 26238
rect 14926 26226 14978 26238
rect 15150 26290 15202 26302
rect 15150 26226 15202 26238
rect 15486 26290 15538 26302
rect 15486 26226 15538 26238
rect 15598 26290 15650 26302
rect 15598 26226 15650 26238
rect 16158 26290 16210 26302
rect 16158 26226 16210 26238
rect 17502 26290 17554 26302
rect 17502 26226 17554 26238
rect 17838 26290 17890 26302
rect 39454 26290 39506 26302
rect 19282 26238 19294 26290
rect 19346 26238 19358 26290
rect 22642 26238 22654 26290
rect 22706 26238 22718 26290
rect 24434 26238 24446 26290
rect 24498 26238 24510 26290
rect 27458 26238 27470 26290
rect 27522 26238 27534 26290
rect 33058 26238 33070 26290
rect 33122 26238 33134 26290
rect 39218 26238 39230 26290
rect 39282 26238 39294 26290
rect 17838 26226 17890 26238
rect 39454 26226 39506 26238
rect 39790 26290 39842 26302
rect 39790 26226 39842 26238
rect 40014 26290 40066 26302
rect 44706 26238 44718 26290
rect 44770 26238 44782 26290
rect 45602 26238 45614 26290
rect 45666 26238 45678 26290
rect 40014 26226 40066 26238
rect 2942 26178 2994 26190
rect 2942 26114 2994 26126
rect 3838 26178 3890 26190
rect 14254 26178 14306 26190
rect 7746 26126 7758 26178
rect 7810 26126 7822 26178
rect 11778 26126 11790 26178
rect 11842 26126 11854 26178
rect 13682 26126 13694 26178
rect 13746 26126 13758 26178
rect 3838 26114 3890 26126
rect 14254 26114 14306 26126
rect 15262 26178 15314 26190
rect 40910 26178 40962 26190
rect 22082 26126 22094 26178
rect 22146 26126 22158 26178
rect 33842 26126 33854 26178
rect 33906 26126 33918 26178
rect 35970 26126 35982 26178
rect 36034 26126 36046 26178
rect 36306 26126 36318 26178
rect 36370 26126 36382 26178
rect 38434 26126 38446 26178
rect 38498 26126 38510 26178
rect 41906 26126 41918 26178
rect 41970 26126 41982 26178
rect 44034 26126 44046 26178
rect 44098 26126 44110 26178
rect 15262 26114 15314 26126
rect 40910 26114 40962 26126
rect 6078 26066 6130 26078
rect 6078 26002 6130 26014
rect 6302 26066 6354 26078
rect 6302 26002 6354 26014
rect 6750 26066 6802 26078
rect 6750 26002 6802 26014
rect 10446 26066 10498 26078
rect 10446 26002 10498 26014
rect 18398 26066 18450 26078
rect 18398 26002 18450 26014
rect 23438 26066 23490 26078
rect 23438 26002 23490 26014
rect 23774 26066 23826 26078
rect 23774 26002 23826 26014
rect 27022 26066 27074 26078
rect 27022 26002 27074 26014
rect 41134 26066 41186 26078
rect 47966 26066 48018 26078
rect 41458 26014 41470 26066
rect 41522 26014 41534 26066
rect 41134 26002 41186 26014
rect 47966 26002 48018 26014
rect 1344 25898 48608 25932
rect 1344 25846 4478 25898
rect 4530 25846 4582 25898
rect 4634 25846 4686 25898
rect 4738 25846 35198 25898
rect 35250 25846 35302 25898
rect 35354 25846 35406 25898
rect 35458 25846 48608 25898
rect 1344 25812 48608 25846
rect 8878 25730 8930 25742
rect 8878 25666 8930 25678
rect 13470 25730 13522 25742
rect 13470 25666 13522 25678
rect 5182 25618 5234 25630
rect 13582 25618 13634 25630
rect 22318 25618 22370 25630
rect 37662 25618 37714 25630
rect 2482 25566 2494 25618
rect 2546 25566 2558 25618
rect 4610 25566 4622 25618
rect 4674 25566 4686 25618
rect 7298 25566 7310 25618
rect 7362 25566 7374 25618
rect 12450 25566 12462 25618
rect 12514 25566 12526 25618
rect 14242 25566 14254 25618
rect 14306 25566 14318 25618
rect 16370 25566 16382 25618
rect 16434 25566 16446 25618
rect 18162 25566 18174 25618
rect 18226 25566 18238 25618
rect 23986 25566 23998 25618
rect 24050 25566 24062 25618
rect 26114 25566 26126 25618
rect 26178 25566 26190 25618
rect 32162 25566 32174 25618
rect 32226 25566 32238 25618
rect 35186 25566 35198 25618
rect 35250 25566 35262 25618
rect 5182 25554 5234 25566
rect 13582 25554 13634 25566
rect 22318 25554 22370 25566
rect 37662 25554 37714 25566
rect 39454 25618 39506 25630
rect 40562 25566 40574 25618
rect 40626 25566 40638 25618
rect 48178 25566 48190 25618
rect 48242 25566 48254 25618
rect 39454 25554 39506 25566
rect 7870 25506 7922 25518
rect 10110 25506 10162 25518
rect 1810 25454 1822 25506
rect 1874 25454 1886 25506
rect 7186 25454 7198 25506
rect 7250 25454 7262 25506
rect 8082 25454 8094 25506
rect 8146 25454 8158 25506
rect 7870 25442 7922 25454
rect 10110 25442 10162 25454
rect 10446 25506 10498 25518
rect 17838 25506 17890 25518
rect 10658 25454 10670 25506
rect 10722 25454 10734 25506
rect 12002 25454 12014 25506
rect 12066 25454 12078 25506
rect 12786 25454 12798 25506
rect 12850 25454 12862 25506
rect 17042 25454 17054 25506
rect 17106 25454 17118 25506
rect 10446 25442 10498 25454
rect 17838 25442 17890 25454
rect 18734 25506 18786 25518
rect 18734 25442 18786 25454
rect 19854 25506 19906 25518
rect 21422 25506 21474 25518
rect 35646 25506 35698 25518
rect 20626 25454 20638 25506
rect 20690 25454 20702 25506
rect 23202 25454 23214 25506
rect 23266 25454 23278 25506
rect 29362 25454 29374 25506
rect 29426 25454 29438 25506
rect 19854 25442 19906 25454
rect 21422 25442 21474 25454
rect 35646 25442 35698 25454
rect 38110 25506 38162 25518
rect 38110 25442 38162 25454
rect 38334 25506 38386 25518
rect 38334 25442 38386 25454
rect 38670 25506 38722 25518
rect 38670 25442 38722 25454
rect 39566 25506 39618 25518
rect 39566 25442 39618 25454
rect 39790 25506 39842 25518
rect 43038 25506 43090 25518
rect 40002 25454 40014 25506
rect 40066 25454 40078 25506
rect 40226 25454 40238 25506
rect 40290 25454 40302 25506
rect 40786 25454 40798 25506
rect 40850 25454 40862 25506
rect 41794 25454 41806 25506
rect 41858 25454 41870 25506
rect 42354 25454 42366 25506
rect 42418 25454 42430 25506
rect 39790 25442 39842 25454
rect 43038 25442 43090 25454
rect 43598 25506 43650 25518
rect 45378 25454 45390 25506
rect 45442 25454 45454 25506
rect 43598 25442 43650 25454
rect 9774 25394 9826 25406
rect 19518 25394 19570 25406
rect 26462 25394 26514 25406
rect 33742 25394 33794 25406
rect 11890 25342 11902 25394
rect 11954 25342 11966 25394
rect 12450 25342 12462 25394
rect 12514 25342 12526 25394
rect 20402 25342 20414 25394
rect 20466 25342 20478 25394
rect 30034 25342 30046 25394
rect 30098 25342 30110 25394
rect 9774 25330 9826 25342
rect 19518 25330 19570 25342
rect 26462 25330 26514 25342
rect 33742 25330 33794 25342
rect 34078 25394 34130 25406
rect 34078 25330 34130 25342
rect 37550 25394 37602 25406
rect 37550 25330 37602 25342
rect 37774 25394 37826 25406
rect 37774 25330 37826 25342
rect 39342 25394 39394 25406
rect 43486 25394 43538 25406
rect 40674 25342 40686 25394
rect 40738 25342 40750 25394
rect 41346 25342 41358 25394
rect 41410 25342 41422 25394
rect 46050 25342 46062 25394
rect 46114 25342 46126 25394
rect 39342 25330 39394 25342
rect 43486 25330 43538 25342
rect 10110 25282 10162 25294
rect 10110 25218 10162 25230
rect 17614 25282 17666 25294
rect 17614 25218 17666 25230
rect 18174 25282 18226 25294
rect 18174 25218 18226 25230
rect 18398 25282 18450 25294
rect 18398 25218 18450 25230
rect 18846 25282 18898 25294
rect 18846 25218 18898 25230
rect 19070 25282 19122 25294
rect 19070 25218 19122 25230
rect 26798 25282 26850 25294
rect 26798 25218 26850 25230
rect 38446 25282 38498 25294
rect 38446 25218 38498 25230
rect 43374 25282 43426 25294
rect 43374 25218 43426 25230
rect 1344 25114 48608 25148
rect 1344 25062 19838 25114
rect 19890 25062 19942 25114
rect 19994 25062 20046 25114
rect 20098 25062 48608 25114
rect 1344 25028 48608 25062
rect 1710 24946 1762 24958
rect 1710 24882 1762 24894
rect 3838 24946 3890 24958
rect 15486 24946 15538 24958
rect 13234 24894 13246 24946
rect 13298 24894 13310 24946
rect 3838 24882 3890 24894
rect 15486 24882 15538 24894
rect 16718 24946 16770 24958
rect 16718 24882 16770 24894
rect 17614 24946 17666 24958
rect 19070 24946 19122 24958
rect 18162 24894 18174 24946
rect 18226 24894 18238 24946
rect 17614 24882 17666 24894
rect 19070 24882 19122 24894
rect 19406 24946 19458 24958
rect 19406 24882 19458 24894
rect 30942 24946 30994 24958
rect 30942 24882 30994 24894
rect 31278 24946 31330 24958
rect 31278 24882 31330 24894
rect 34526 24946 34578 24958
rect 43262 24946 43314 24958
rect 39218 24894 39230 24946
rect 39282 24894 39294 24946
rect 34526 24882 34578 24894
rect 43262 24882 43314 24894
rect 44606 24946 44658 24958
rect 45266 24894 45278 24946
rect 45330 24894 45342 24946
rect 44606 24882 44658 24894
rect 15038 24834 15090 24846
rect 2034 24782 2046 24834
rect 2098 24782 2110 24834
rect 7858 24782 7870 24834
rect 7922 24782 7934 24834
rect 10770 24782 10782 24834
rect 10834 24782 10846 24834
rect 11330 24782 11342 24834
rect 11394 24782 11406 24834
rect 12226 24782 12238 24834
rect 12290 24782 12302 24834
rect 13122 24782 13134 24834
rect 13186 24782 13198 24834
rect 15038 24770 15090 24782
rect 16158 24834 16210 24846
rect 22990 24834 23042 24846
rect 44942 24834 44994 24846
rect 21298 24782 21310 24834
rect 21362 24782 21374 24834
rect 28690 24782 28702 24834
rect 28754 24782 28766 24834
rect 35410 24782 35422 24834
rect 35474 24782 35486 24834
rect 16158 24770 16210 24782
rect 22990 24770 23042 24782
rect 44942 24770 44994 24782
rect 2382 24722 2434 24734
rect 2382 24658 2434 24670
rect 2942 24722 2994 24734
rect 2942 24658 2994 24670
rect 5630 24722 5682 24734
rect 5630 24658 5682 24670
rect 6974 24722 7026 24734
rect 16046 24722 16098 24734
rect 7746 24670 7758 24722
rect 7810 24670 7822 24722
rect 8306 24670 8318 24722
rect 8370 24670 8382 24722
rect 8978 24670 8990 24722
rect 9042 24670 9054 24722
rect 9538 24670 9550 24722
rect 9602 24670 9614 24722
rect 10882 24670 10894 24722
rect 10946 24670 10958 24722
rect 11442 24670 11454 24722
rect 11506 24670 11518 24722
rect 12450 24670 12462 24722
rect 12514 24670 12526 24722
rect 13010 24670 13022 24722
rect 13074 24670 13086 24722
rect 13906 24670 13918 24722
rect 13970 24670 13982 24722
rect 6974 24658 7026 24670
rect 16046 24658 16098 24670
rect 16382 24722 16434 24734
rect 16382 24658 16434 24670
rect 16606 24722 16658 24734
rect 16606 24658 16658 24670
rect 16942 24722 16994 24734
rect 16942 24658 16994 24670
rect 17838 24722 17890 24734
rect 23326 24722 23378 24734
rect 20402 24670 20414 24722
rect 20466 24670 20478 24722
rect 20738 24670 20750 24722
rect 20802 24670 20814 24722
rect 17838 24658 17890 24670
rect 23326 24658 23378 24670
rect 24670 24722 24722 24734
rect 30830 24722 30882 24734
rect 25218 24670 25230 24722
rect 25282 24670 25294 24722
rect 24670 24658 24722 24670
rect 30830 24658 30882 24670
rect 31054 24722 31106 24734
rect 38670 24722 38722 24734
rect 35634 24670 35646 24722
rect 35698 24670 35710 24722
rect 31054 24658 31106 24670
rect 38670 24658 38722 24670
rect 42478 24722 42530 24734
rect 42478 24658 42530 24670
rect 42702 24722 42754 24734
rect 44370 24670 44382 24722
rect 44434 24670 44446 24722
rect 48066 24670 48078 24722
rect 48130 24670 48142 24722
rect 42702 24658 42754 24670
rect 4174 24610 4226 24622
rect 4174 24546 4226 24558
rect 4622 24610 4674 24622
rect 4622 24546 4674 24558
rect 5070 24610 5122 24622
rect 5070 24546 5122 24558
rect 6078 24610 6130 24622
rect 6078 24546 6130 24558
rect 6302 24610 6354 24622
rect 6302 24546 6354 24558
rect 6750 24610 6802 24622
rect 21870 24610 21922 24622
rect 11666 24558 11678 24610
rect 11730 24558 11742 24610
rect 6750 24546 6802 24558
rect 21870 24546 21922 24558
rect 38446 24610 38498 24622
rect 38446 24546 38498 24558
rect 39678 24610 39730 24622
rect 39678 24546 39730 24558
rect 40238 24610 40290 24622
rect 40238 24546 40290 24558
rect 41022 24610 41074 24622
rect 43362 24558 43374 24610
rect 43426 24558 43438 24610
rect 46946 24558 46958 24610
rect 47010 24558 47022 24610
rect 41022 24546 41074 24558
rect 6526 24498 6578 24510
rect 4162 24446 4174 24498
rect 4226 24495 4238 24498
rect 5058 24495 5070 24498
rect 4226 24449 5070 24495
rect 4226 24446 4238 24449
rect 5058 24446 5070 24449
rect 5122 24446 5134 24498
rect 6526 24434 6578 24446
rect 7422 24498 7474 24510
rect 7422 24434 7474 24446
rect 34862 24498 34914 24510
rect 34862 24434 34914 24446
rect 38894 24498 38946 24510
rect 43038 24498 43090 24510
rect 39666 24446 39678 24498
rect 39730 24495 39742 24498
rect 40226 24495 40238 24498
rect 39730 24449 40238 24495
rect 39730 24446 39742 24449
rect 40226 24446 40238 24449
rect 40290 24446 40302 24498
rect 42130 24446 42142 24498
rect 42194 24446 42206 24498
rect 38894 24434 38946 24446
rect 43038 24434 43090 24446
rect 1344 24330 48608 24364
rect 1344 24278 4478 24330
rect 4530 24278 4582 24330
rect 4634 24278 4686 24330
rect 4738 24278 35198 24330
rect 35250 24278 35302 24330
rect 35354 24278 35406 24330
rect 35458 24278 48608 24330
rect 1344 24244 48608 24278
rect 19854 24162 19906 24174
rect 12786 24110 12798 24162
rect 12850 24159 12862 24162
rect 13010 24159 13022 24162
rect 12850 24113 13022 24159
rect 12850 24110 12862 24113
rect 13010 24110 13022 24113
rect 13074 24110 13086 24162
rect 19854 24098 19906 24110
rect 5182 24050 5234 24062
rect 12574 24050 12626 24062
rect 2482 23998 2494 24050
rect 2546 23998 2558 24050
rect 4610 23998 4622 24050
rect 4674 23998 4686 24050
rect 11218 23998 11230 24050
rect 11282 23998 11294 24050
rect 5182 23986 5234 23998
rect 12574 23986 12626 23998
rect 13022 24050 13074 24062
rect 29262 24050 29314 24062
rect 43710 24050 43762 24062
rect 23202 23998 23214 24050
rect 23266 23998 23278 24050
rect 25330 23998 25342 24050
rect 25394 23998 25406 24050
rect 25666 23998 25678 24050
rect 25730 23998 25742 24050
rect 27794 23998 27806 24050
rect 27858 23998 27870 24050
rect 33730 23998 33742 24050
rect 33794 23998 33806 24050
rect 13022 23986 13074 23998
rect 29262 23986 29314 23998
rect 43710 23986 43762 23998
rect 47966 24050 48018 24062
rect 47966 23986 48018 23998
rect 8878 23938 8930 23950
rect 29038 23938 29090 23950
rect 1810 23886 1822 23938
rect 1874 23886 1886 23938
rect 6738 23886 6750 23938
rect 6802 23886 6814 23938
rect 13682 23886 13694 23938
rect 13746 23886 13758 23938
rect 14466 23886 14478 23938
rect 14530 23886 14542 23938
rect 15250 23886 15262 23938
rect 15314 23886 15326 23938
rect 16034 23886 16046 23938
rect 16098 23886 16110 23938
rect 16818 23886 16830 23938
rect 16882 23886 16894 23938
rect 17266 23886 17278 23938
rect 17330 23886 17342 23938
rect 18050 23886 18062 23938
rect 18114 23886 18126 23938
rect 20290 23886 20302 23938
rect 20354 23886 20366 23938
rect 22418 23886 22430 23938
rect 22482 23886 22494 23938
rect 28578 23886 28590 23938
rect 28642 23886 28654 23938
rect 8878 23874 8930 23886
rect 29038 23874 29090 23886
rect 29486 23938 29538 23950
rect 29486 23874 29538 23886
rect 29598 23938 29650 23950
rect 29598 23874 29650 23886
rect 30606 23938 30658 23950
rect 38894 23938 38946 23950
rect 42590 23938 42642 23950
rect 30818 23886 30830 23938
rect 30882 23886 30894 23938
rect 37090 23886 37102 23938
rect 37154 23886 37166 23938
rect 39890 23886 39902 23938
rect 39954 23886 39966 23938
rect 40450 23886 40462 23938
rect 40514 23886 40526 23938
rect 41682 23886 41694 23938
rect 41746 23886 41758 23938
rect 30606 23874 30658 23886
rect 38894 23874 38946 23886
rect 42590 23874 42642 23886
rect 42926 23938 42978 23950
rect 42926 23874 42978 23886
rect 43262 23938 43314 23950
rect 45154 23886 45166 23938
rect 45218 23886 45230 23938
rect 45602 23886 45614 23938
rect 45666 23886 45678 23938
rect 43262 23874 43314 23886
rect 9998 23826 10050 23838
rect 17838 23826 17890 23838
rect 6850 23774 6862 23826
rect 6914 23774 6926 23826
rect 13570 23774 13582 23826
rect 13634 23774 13646 23826
rect 14242 23774 14254 23826
rect 14306 23774 14318 23826
rect 16146 23774 16158 23826
rect 16210 23774 16222 23826
rect 9998 23762 10050 23774
rect 17838 23762 17890 23774
rect 18286 23826 18338 23838
rect 18286 23762 18338 23774
rect 19070 23826 19122 23838
rect 19070 23762 19122 23774
rect 19518 23826 19570 23838
rect 30270 23826 30322 23838
rect 20626 23774 20638 23826
rect 20690 23774 20702 23826
rect 19518 23762 19570 23774
rect 30270 23762 30322 23774
rect 30382 23826 30434 23838
rect 43598 23826 43650 23838
rect 31602 23774 31614 23826
rect 31666 23774 31678 23826
rect 35970 23774 35982 23826
rect 36034 23774 36046 23826
rect 37314 23774 37326 23826
rect 37378 23774 37390 23826
rect 37986 23774 37998 23826
rect 38050 23774 38062 23826
rect 40002 23774 40014 23826
rect 40066 23774 40078 23826
rect 40674 23774 40686 23826
rect 40738 23774 40750 23826
rect 30382 23762 30434 23774
rect 43598 23762 43650 23774
rect 43822 23826 43874 23838
rect 43822 23762 43874 23774
rect 44942 23826 44994 23838
rect 44942 23762 44994 23774
rect 6078 23714 6130 23726
rect 6078 23650 6130 23662
rect 6526 23714 6578 23726
rect 11678 23714 11730 23726
rect 17390 23714 17442 23726
rect 8418 23662 8430 23714
rect 8482 23662 8494 23714
rect 14354 23662 14366 23714
rect 14418 23662 14430 23714
rect 6526 23650 6578 23662
rect 11678 23650 11730 23662
rect 17390 23650 17442 23662
rect 18398 23714 18450 23726
rect 18398 23650 18450 23662
rect 18734 23714 18786 23726
rect 18734 23650 18786 23662
rect 35646 23714 35698 23726
rect 35646 23650 35698 23662
rect 37662 23714 37714 23726
rect 37662 23650 37714 23662
rect 38334 23714 38386 23726
rect 42926 23714 42978 23726
rect 40562 23662 40574 23714
rect 40626 23662 40638 23714
rect 38334 23650 38386 23662
rect 42926 23650 42978 23662
rect 1344 23546 48608 23580
rect 1344 23494 19838 23546
rect 19890 23494 19942 23546
rect 19994 23494 20046 23546
rect 20098 23494 48608 23546
rect 1344 23460 48608 23494
rect 1710 23378 1762 23390
rect 1710 23314 1762 23326
rect 2942 23378 2994 23390
rect 2942 23314 2994 23326
rect 4510 23378 4562 23390
rect 4510 23314 4562 23326
rect 7982 23378 8034 23390
rect 7982 23314 8034 23326
rect 8206 23378 8258 23390
rect 8206 23314 8258 23326
rect 8990 23378 9042 23390
rect 13918 23378 13970 23390
rect 12562 23326 12574 23378
rect 12626 23326 12638 23378
rect 8990 23314 9042 23326
rect 13918 23314 13970 23326
rect 15710 23378 15762 23390
rect 17614 23378 17666 23390
rect 16818 23326 16830 23378
rect 16882 23326 16894 23378
rect 15710 23314 15762 23326
rect 17614 23314 17666 23326
rect 23326 23378 23378 23390
rect 23326 23314 23378 23326
rect 25678 23378 25730 23390
rect 25678 23314 25730 23326
rect 26462 23378 26514 23390
rect 26462 23314 26514 23326
rect 29374 23378 29426 23390
rect 29374 23314 29426 23326
rect 30942 23378 30994 23390
rect 30942 23314 30994 23326
rect 31166 23378 31218 23390
rect 31166 23314 31218 23326
rect 35198 23378 35250 23390
rect 35198 23314 35250 23326
rect 39006 23378 39058 23390
rect 41806 23378 41858 23390
rect 39330 23326 39342 23378
rect 39394 23326 39406 23378
rect 39006 23314 39058 23326
rect 41806 23314 41858 23326
rect 46510 23378 46562 23390
rect 46510 23314 46562 23326
rect 22878 23266 22930 23278
rect 25454 23266 25506 23278
rect 29486 23266 29538 23278
rect 2034 23214 2046 23266
rect 2098 23214 2110 23266
rect 8642 23214 8654 23266
rect 8706 23214 8718 23266
rect 10882 23214 10894 23266
rect 10946 23214 10958 23266
rect 13010 23214 13022 23266
rect 13074 23214 13086 23266
rect 14130 23214 14142 23266
rect 14194 23214 14206 23266
rect 18834 23214 18846 23266
rect 18898 23214 18910 23266
rect 24322 23214 24334 23266
rect 24386 23214 24398 23266
rect 27570 23214 27582 23266
rect 27634 23214 27646 23266
rect 22878 23202 22930 23214
rect 25454 23202 25506 23214
rect 29486 23202 29538 23214
rect 31054 23266 31106 23278
rect 31054 23202 31106 23214
rect 31726 23266 31778 23278
rect 31726 23202 31778 23214
rect 31950 23266 32002 23278
rect 31950 23202 32002 23214
rect 32062 23266 32114 23278
rect 39678 23266 39730 23278
rect 36306 23214 36318 23266
rect 36370 23214 36382 23266
rect 38658 23214 38670 23266
rect 38722 23214 38734 23266
rect 32062 23202 32114 23214
rect 39678 23202 39730 23214
rect 42030 23266 42082 23278
rect 42030 23202 42082 23214
rect 42366 23266 42418 23278
rect 43586 23214 43598 23266
rect 43650 23214 43662 23266
rect 47058 23214 47070 23266
rect 47122 23214 47134 23266
rect 47394 23214 47406 23266
rect 47458 23214 47470 23266
rect 42366 23202 42418 23214
rect 8318 23154 8370 23166
rect 4834 23102 4846 23154
rect 4898 23102 4910 23154
rect 8318 23090 8370 23102
rect 9662 23154 9714 23166
rect 9662 23090 9714 23102
rect 9886 23154 9938 23166
rect 9886 23090 9938 23102
rect 10110 23154 10162 23166
rect 10110 23090 10162 23102
rect 10558 23154 10610 23166
rect 13246 23154 13298 23166
rect 11442 23102 11454 23154
rect 11506 23102 11518 23154
rect 11778 23102 11790 23154
rect 11842 23102 11854 23154
rect 12226 23102 12238 23154
rect 12290 23102 12302 23154
rect 10558 23090 10610 23102
rect 13246 23090 13298 23102
rect 14478 23154 14530 23166
rect 14478 23090 14530 23102
rect 14926 23154 14978 23166
rect 22318 23154 22370 23166
rect 25678 23154 25730 23166
rect 16594 23102 16606 23154
rect 16658 23102 16670 23154
rect 18050 23102 18062 23154
rect 18114 23102 18126 23154
rect 24210 23102 24222 23154
rect 24274 23102 24286 23154
rect 14926 23090 14978 23102
rect 22318 23090 22370 23102
rect 25678 23090 25730 23102
rect 26014 23154 26066 23166
rect 26014 23090 26066 23102
rect 26798 23154 26850 23166
rect 29038 23154 29090 23166
rect 27458 23102 27470 23154
rect 27522 23102 27534 23154
rect 26798 23090 26850 23102
rect 29038 23090 29090 23102
rect 29710 23154 29762 23166
rect 29710 23090 29762 23102
rect 31614 23154 31666 23166
rect 31614 23090 31666 23102
rect 35534 23154 35586 23166
rect 46846 23154 46898 23166
rect 35970 23102 35982 23154
rect 36034 23102 36046 23154
rect 38434 23102 38446 23154
rect 38498 23102 38510 23154
rect 40002 23102 40014 23154
rect 40066 23102 40078 23154
rect 41234 23102 41246 23154
rect 41298 23102 41310 23154
rect 42914 23102 42926 23154
rect 42978 23102 42990 23154
rect 35534 23090 35586 23102
rect 46846 23090 46898 23102
rect 2606 23042 2658 23054
rect 2606 22978 2658 22990
rect 3502 23042 3554 23054
rect 3502 22978 3554 22990
rect 3950 23042 4002 23054
rect 16158 23042 16210 23054
rect 37998 23042 38050 23054
rect 5506 22990 5518 23042
rect 5570 22990 5582 23042
rect 7634 22990 7646 23042
rect 7698 22990 7710 23042
rect 9762 22990 9774 23042
rect 9826 22990 9838 23042
rect 20962 22990 20974 23042
rect 21026 22990 21038 23042
rect 3950 22978 4002 22990
rect 16158 22978 16210 22990
rect 37998 22978 38050 22990
rect 39790 23042 39842 23054
rect 48190 23042 48242 23054
rect 45714 22990 45726 23042
rect 45778 22990 45790 23042
rect 39790 22978 39842 22990
rect 48190 22978 48242 22990
rect 10334 22930 10386 22942
rect 23662 22930 23714 22942
rect 2594 22878 2606 22930
rect 2658 22927 2670 22930
rect 3154 22927 3166 22930
rect 2658 22881 3166 22927
rect 2658 22878 2670 22881
rect 3154 22878 3166 22881
rect 3218 22878 3230 22930
rect 3490 22878 3502 22930
rect 3554 22927 3566 22930
rect 4498 22927 4510 22930
rect 3554 22881 4510 22927
rect 3554 22878 3566 22881
rect 4498 22878 4510 22881
rect 4562 22878 4574 22930
rect 15586 22878 15598 22930
rect 15650 22927 15662 22930
rect 16146 22927 16158 22930
rect 15650 22881 16158 22927
rect 15650 22878 15662 22881
rect 16146 22878 16158 22881
rect 16210 22878 16222 22930
rect 10334 22866 10386 22878
rect 23662 22866 23714 22878
rect 40910 22930 40962 22942
rect 40910 22866 40962 22878
rect 41246 22930 41298 22942
rect 41246 22866 41298 22878
rect 1344 22762 48608 22796
rect 1344 22710 4478 22762
rect 4530 22710 4582 22762
rect 4634 22710 4686 22762
rect 4738 22710 35198 22762
rect 35250 22710 35302 22762
rect 35354 22710 35406 22762
rect 35458 22710 48608 22762
rect 1344 22676 48608 22710
rect 7422 22594 7474 22606
rect 35198 22594 35250 22606
rect 10658 22542 10670 22594
rect 10722 22591 10734 22594
rect 10882 22591 10894 22594
rect 10722 22545 10894 22591
rect 10722 22542 10734 22545
rect 10882 22542 10894 22545
rect 10946 22542 10958 22594
rect 12002 22542 12014 22594
rect 12066 22591 12078 22594
rect 12226 22591 12238 22594
rect 12066 22545 12238 22591
rect 12066 22542 12078 22545
rect 12226 22542 12238 22545
rect 12290 22542 12302 22594
rect 22306 22542 22318 22594
rect 22370 22542 22382 22594
rect 7422 22530 7474 22542
rect 5854 22482 5906 22494
rect 2482 22430 2494 22482
rect 2546 22430 2558 22482
rect 4610 22430 4622 22482
rect 4674 22430 4686 22482
rect 5854 22418 5906 22430
rect 6414 22482 6466 22494
rect 6414 22418 6466 22430
rect 7310 22482 7362 22494
rect 7310 22418 7362 22430
rect 10222 22482 10274 22494
rect 10222 22418 10274 22430
rect 10894 22482 10946 22494
rect 10894 22418 10946 22430
rect 11342 22482 11394 22494
rect 11342 22418 11394 22430
rect 11902 22482 11954 22494
rect 11902 22418 11954 22430
rect 12350 22482 12402 22494
rect 12350 22418 12402 22430
rect 12798 22482 12850 22494
rect 12798 22418 12850 22430
rect 14478 22482 14530 22494
rect 19070 22482 19122 22494
rect 17826 22430 17838 22482
rect 17890 22430 17902 22482
rect 14478 22418 14530 22430
rect 19070 22418 19122 22430
rect 6526 22370 6578 22382
rect 9214 22370 9266 22382
rect 1810 22318 1822 22370
rect 1874 22318 1886 22370
rect 6738 22318 6750 22370
rect 6802 22318 6814 22370
rect 7970 22318 7982 22370
rect 8034 22318 8046 22370
rect 6526 22306 6578 22318
rect 9214 22306 9266 22318
rect 10446 22370 10498 22382
rect 10446 22306 10498 22318
rect 14030 22370 14082 22382
rect 22094 22370 22146 22382
rect 14802 22318 14814 22370
rect 14866 22318 14878 22370
rect 14030 22306 14082 22318
rect 22094 22306 22146 22318
rect 6078 22258 6130 22270
rect 6078 22194 6130 22206
rect 8766 22258 8818 22270
rect 8766 22194 8818 22206
rect 8878 22258 8930 22270
rect 8878 22194 8930 22206
rect 9326 22258 9378 22270
rect 9326 22194 9378 22206
rect 9774 22258 9826 22270
rect 9774 22194 9826 22206
rect 9998 22258 10050 22270
rect 9998 22194 10050 22206
rect 13470 22258 13522 22270
rect 13470 22194 13522 22206
rect 13694 22258 13746 22270
rect 21758 22258 21810 22270
rect 15586 22206 15598 22258
rect 15650 22206 15662 22258
rect 13694 22194 13746 22206
rect 21758 22194 21810 22206
rect 5070 22146 5122 22158
rect 5070 22082 5122 22094
rect 6302 22146 6354 22158
rect 9550 22146 9602 22158
rect 7746 22094 7758 22146
rect 7810 22094 7822 22146
rect 6302 22082 6354 22094
rect 9550 22082 9602 22094
rect 12910 22146 12962 22158
rect 12910 22082 12962 22094
rect 13806 22146 13858 22158
rect 13806 22082 13858 22094
rect 21982 22146 22034 22158
rect 22321 22146 22367 22542
rect 35198 22530 35250 22542
rect 32734 22482 32786 22494
rect 22754 22430 22766 22482
rect 22818 22430 22830 22482
rect 28130 22430 28142 22482
rect 28194 22430 28206 22482
rect 32050 22430 32062 22482
rect 32114 22430 32126 22482
rect 32734 22418 32786 22430
rect 44382 22482 44434 22494
rect 44382 22418 44434 22430
rect 45054 22482 45106 22494
rect 48178 22430 48190 22482
rect 48242 22430 48254 22482
rect 45054 22418 45106 22430
rect 38782 22370 38834 22382
rect 25218 22318 25230 22370
rect 25282 22318 25294 22370
rect 29250 22318 29262 22370
rect 29314 22318 29326 22370
rect 34066 22318 34078 22370
rect 34130 22318 34142 22370
rect 35970 22318 35982 22370
rect 36034 22318 36046 22370
rect 38782 22306 38834 22318
rect 39342 22370 39394 22382
rect 42590 22370 42642 22382
rect 39890 22318 39902 22370
rect 39954 22318 39966 22370
rect 40562 22318 40574 22370
rect 40626 22318 40638 22370
rect 41794 22318 41806 22370
rect 41858 22318 41870 22370
rect 39342 22306 39394 22318
rect 42590 22306 42642 22318
rect 42814 22370 42866 22382
rect 42814 22306 42866 22318
rect 43150 22370 43202 22382
rect 43150 22306 43202 22318
rect 43486 22370 43538 22382
rect 45378 22318 45390 22370
rect 45442 22318 45454 22370
rect 43486 22306 43538 22318
rect 22542 22258 22594 22270
rect 22542 22194 22594 22206
rect 23662 22258 23714 22270
rect 39118 22258 39170 22270
rect 43710 22258 43762 22270
rect 26002 22206 26014 22258
rect 26066 22206 26078 22258
rect 29922 22206 29934 22258
rect 29986 22206 29998 22258
rect 35746 22206 35758 22258
rect 35810 22206 35822 22258
rect 39778 22206 39790 22258
rect 39842 22206 39854 22258
rect 40786 22206 40798 22258
rect 40850 22206 40862 22258
rect 42242 22206 42254 22258
rect 42306 22206 42318 22258
rect 46050 22206 46062 22258
rect 46114 22206 46126 22258
rect 23662 22194 23714 22206
rect 39118 22194 39170 22206
rect 43710 22194 43762 22206
rect 22766 22146 22818 22158
rect 22306 22094 22318 22146
rect 22370 22094 22382 22146
rect 21982 22082 22034 22094
rect 22766 22082 22818 22094
rect 22990 22146 23042 22158
rect 22990 22082 23042 22094
rect 23326 22146 23378 22158
rect 23326 22082 23378 22094
rect 24222 22146 24274 22158
rect 24222 22082 24274 22094
rect 34302 22146 34354 22158
rect 34302 22082 34354 22094
rect 34862 22146 34914 22158
rect 34862 22082 34914 22094
rect 37102 22146 37154 22158
rect 37102 22082 37154 22094
rect 37550 22146 37602 22158
rect 37550 22082 37602 22094
rect 38110 22146 38162 22158
rect 39006 22146 39058 22158
rect 38434 22094 38446 22146
rect 38498 22094 38510 22146
rect 38110 22082 38162 22094
rect 39006 22082 39058 22094
rect 42030 22146 42082 22158
rect 42030 22082 42082 22094
rect 43598 22146 43650 22158
rect 43598 22082 43650 22094
rect 1344 21978 48608 22012
rect 1344 21926 19838 21978
rect 19890 21926 19942 21978
rect 19994 21926 20046 21978
rect 20098 21926 48608 21978
rect 1344 21892 48608 21926
rect 5630 21810 5682 21822
rect 5630 21746 5682 21758
rect 6302 21810 6354 21822
rect 6302 21746 6354 21758
rect 6974 21810 7026 21822
rect 6974 21746 7026 21758
rect 7982 21810 8034 21822
rect 7982 21746 8034 21758
rect 8654 21810 8706 21822
rect 8654 21746 8706 21758
rect 10110 21810 10162 21822
rect 10110 21746 10162 21758
rect 15934 21810 15986 21822
rect 26126 21810 26178 21822
rect 20626 21758 20638 21810
rect 20690 21758 20702 21810
rect 22194 21758 22206 21810
rect 22258 21758 22270 21810
rect 22866 21758 22878 21810
rect 22930 21758 22942 21810
rect 15934 21746 15986 21758
rect 26126 21746 26178 21758
rect 26238 21810 26290 21822
rect 26238 21746 26290 21758
rect 27918 21810 27970 21822
rect 29598 21810 29650 21822
rect 29138 21758 29150 21810
rect 29202 21758 29214 21810
rect 27918 21746 27970 21758
rect 29598 21746 29650 21758
rect 29710 21810 29762 21822
rect 29710 21746 29762 21758
rect 30718 21810 30770 21822
rect 30718 21746 30770 21758
rect 31390 21810 31442 21822
rect 42142 21810 42194 21822
rect 39218 21758 39230 21810
rect 39282 21758 39294 21810
rect 41794 21758 41806 21810
rect 41858 21758 41870 21810
rect 31390 21746 31442 21758
rect 42142 21746 42194 21758
rect 7646 21698 7698 21710
rect 7410 21646 7422 21698
rect 7474 21646 7486 21698
rect 7646 21634 7698 21646
rect 7758 21698 7810 21710
rect 21758 21698 21810 21710
rect 8306 21646 8318 21698
rect 8370 21646 8382 21698
rect 12898 21646 12910 21698
rect 12962 21646 12974 21698
rect 7758 21634 7810 21646
rect 21758 21634 21810 21646
rect 32062 21698 32114 21710
rect 32062 21634 32114 21646
rect 32174 21698 32226 21710
rect 42478 21698 42530 21710
rect 37538 21646 37550 21698
rect 37602 21646 37614 21698
rect 38994 21646 39006 21698
rect 39058 21646 39070 21698
rect 40002 21646 40014 21698
rect 40066 21646 40078 21698
rect 45378 21646 45390 21698
rect 45442 21646 45454 21698
rect 47506 21646 47518 21698
rect 47570 21646 47582 21698
rect 48066 21646 48078 21698
rect 48130 21646 48142 21698
rect 32174 21634 32226 21646
rect 42478 21634 42530 21646
rect 5742 21586 5794 21598
rect 1810 21534 1822 21586
rect 1874 21534 1886 21586
rect 5742 21522 5794 21534
rect 6190 21586 6242 21598
rect 6190 21522 6242 21534
rect 6414 21586 6466 21598
rect 6414 21522 6466 21534
rect 10334 21586 10386 21598
rect 10334 21522 10386 21534
rect 10894 21586 10946 21598
rect 15486 21586 15538 21598
rect 21646 21586 21698 21598
rect 26350 21586 26402 21598
rect 11330 21534 11342 21586
rect 11394 21534 11406 21586
rect 12226 21534 12238 21586
rect 12290 21534 12302 21586
rect 17490 21534 17502 21586
rect 17554 21534 17566 21586
rect 20850 21534 20862 21586
rect 20914 21534 20926 21586
rect 21410 21534 21422 21586
rect 21474 21534 21486 21586
rect 23090 21534 23102 21586
rect 23154 21534 23166 21586
rect 23426 21534 23438 21586
rect 23490 21534 23502 21586
rect 10894 21522 10946 21534
rect 15486 21522 15538 21534
rect 21646 21522 21698 21534
rect 26350 21522 26402 21534
rect 26798 21586 26850 21598
rect 26798 21522 26850 21534
rect 27694 21586 27746 21598
rect 27694 21522 27746 21534
rect 28030 21586 28082 21598
rect 29486 21586 29538 21598
rect 28914 21534 28926 21586
rect 28978 21534 28990 21586
rect 28030 21522 28082 21534
rect 29486 21522 29538 21534
rect 30158 21586 30210 21598
rect 30158 21522 30210 21534
rect 30494 21586 30546 21598
rect 30494 21522 30546 21534
rect 30830 21586 30882 21598
rect 30830 21522 30882 21534
rect 31166 21586 31218 21598
rect 31166 21522 31218 21534
rect 31838 21586 31890 21598
rect 40910 21586 40962 21598
rect 42814 21586 42866 21598
rect 47294 21586 47346 21598
rect 33058 21534 33070 21586
rect 33122 21534 33134 21586
rect 37874 21534 37886 21586
rect 37938 21534 37950 21586
rect 39218 21534 39230 21586
rect 39282 21534 39294 21586
rect 39890 21534 39902 21586
rect 39954 21534 39966 21586
rect 41346 21534 41358 21586
rect 41410 21534 41422 21586
rect 46050 21534 46062 21586
rect 46114 21534 46126 21586
rect 31838 21522 31890 21534
rect 40910 21522 40962 21534
rect 42814 21522 42866 21534
rect 47294 21522 47346 21534
rect 5182 21474 5234 21486
rect 11790 21474 11842 21486
rect 16494 21474 16546 21486
rect 31278 21474 31330 21486
rect 36990 21474 37042 21486
rect 2482 21422 2494 21474
rect 2546 21422 2558 21474
rect 4610 21422 4622 21474
rect 4674 21422 4686 21474
rect 7634 21422 7646 21474
rect 7698 21422 7710 21474
rect 15026 21422 15038 21474
rect 15090 21422 15102 21474
rect 18162 21422 18174 21474
rect 18226 21422 18238 21474
rect 20290 21422 20302 21474
rect 20354 21422 20366 21474
rect 22978 21422 22990 21474
rect 23042 21422 23054 21474
rect 35186 21422 35198 21474
rect 35250 21422 35262 21474
rect 43250 21422 43262 21474
rect 43314 21422 43326 21474
rect 5182 21410 5234 21422
rect 11790 21410 11842 21422
rect 16494 21410 16546 21422
rect 31278 21410 31330 21422
rect 36990 21410 37042 21422
rect 32174 21362 32226 21374
rect 16146 21310 16158 21362
rect 16210 21359 16222 21362
rect 16370 21359 16382 21362
rect 16210 21313 16382 21359
rect 16210 21310 16222 21313
rect 16370 21310 16382 21313
rect 16434 21310 16446 21362
rect 32174 21298 32226 21310
rect 37214 21362 37266 21374
rect 37214 21298 37266 21310
rect 46958 21362 47010 21374
rect 46958 21298 47010 21310
rect 1344 21194 48608 21228
rect 1344 21142 4478 21194
rect 4530 21142 4582 21194
rect 4634 21142 4686 21194
rect 4738 21142 35198 21194
rect 35250 21142 35302 21194
rect 35354 21142 35406 21194
rect 35458 21142 48608 21194
rect 1344 21108 48608 21142
rect 7310 21026 7362 21038
rect 13582 21026 13634 21038
rect 9986 21023 9998 21026
rect 7310 20962 7362 20974
rect 9441 20977 9998 21023
rect 5070 20914 5122 20926
rect 7982 20914 8034 20926
rect 1698 20862 1710 20914
rect 1762 20862 1774 20914
rect 6066 20862 6078 20914
rect 6130 20862 6142 20914
rect 5070 20850 5122 20862
rect 7982 20850 8034 20862
rect 6526 20802 6578 20814
rect 8878 20802 8930 20814
rect 4498 20750 4510 20802
rect 4562 20750 4574 20802
rect 6738 20750 6750 20802
rect 6802 20750 6814 20802
rect 7858 20750 7870 20802
rect 7922 20750 7934 20802
rect 6526 20738 6578 20750
rect 8878 20738 8930 20750
rect 9214 20802 9266 20814
rect 9441 20802 9487 20977
rect 9986 20974 9998 20977
rect 10050 20974 10062 21026
rect 13582 20962 13634 20974
rect 15038 21026 15090 21038
rect 34750 21026 34802 21038
rect 23650 20974 23662 21026
rect 23714 20974 23726 21026
rect 15038 20962 15090 20974
rect 34750 20962 34802 20974
rect 35086 21026 35138 21038
rect 35086 20962 35138 20974
rect 47966 21026 48018 21038
rect 47966 20962 48018 20974
rect 9886 20914 9938 20926
rect 9886 20850 9938 20862
rect 10334 20914 10386 20926
rect 10334 20850 10386 20862
rect 11006 20914 11058 20926
rect 11006 20850 11058 20862
rect 11342 20914 11394 20926
rect 11342 20850 11394 20862
rect 12798 20914 12850 20926
rect 12798 20850 12850 20862
rect 22430 20914 22482 20926
rect 22430 20850 22482 20862
rect 23998 20914 24050 20926
rect 36430 20914 36482 20926
rect 32162 20862 32174 20914
rect 32226 20862 32238 20914
rect 34290 20862 34302 20914
rect 34354 20862 34366 20914
rect 37650 20862 37662 20914
rect 37714 20862 37726 20914
rect 39106 20862 39118 20914
rect 39170 20862 39182 20914
rect 41234 20862 41246 20914
rect 41298 20862 41310 20914
rect 43586 20862 43598 20914
rect 43650 20862 43662 20914
rect 23998 20850 24050 20862
rect 36430 20850 36482 20862
rect 11790 20802 11842 20814
rect 9426 20750 9438 20802
rect 9490 20750 9502 20802
rect 11554 20750 11566 20802
rect 11618 20750 11630 20802
rect 9214 20738 9266 20750
rect 11790 20738 11842 20750
rect 12126 20802 12178 20814
rect 13470 20802 13522 20814
rect 12338 20750 12350 20802
rect 12402 20750 12414 20802
rect 12126 20738 12178 20750
rect 13470 20738 13522 20750
rect 13918 20802 13970 20814
rect 16158 20802 16210 20814
rect 14466 20750 14478 20802
rect 14530 20750 14542 20802
rect 14690 20750 14702 20802
rect 14754 20750 14766 20802
rect 13918 20738 13970 20750
rect 16158 20738 16210 20750
rect 16270 20802 16322 20814
rect 16270 20738 16322 20750
rect 21422 20802 21474 20814
rect 21422 20738 21474 20750
rect 21982 20802 22034 20814
rect 21982 20738 22034 20750
rect 22990 20802 23042 20814
rect 22990 20738 23042 20750
rect 23102 20802 23154 20814
rect 23102 20738 23154 20750
rect 23214 20802 23266 20814
rect 23214 20738 23266 20750
rect 25902 20802 25954 20814
rect 25902 20738 25954 20750
rect 26350 20802 26402 20814
rect 31490 20750 31502 20802
rect 31554 20750 31566 20802
rect 35858 20750 35870 20802
rect 35922 20750 35934 20802
rect 38322 20750 38334 20802
rect 38386 20750 38398 20802
rect 42018 20750 42030 20802
rect 42082 20750 42094 20802
rect 42802 20750 42814 20802
rect 42866 20750 42878 20802
rect 43698 20750 43710 20802
rect 43762 20750 43774 20802
rect 45042 20750 45054 20802
rect 45106 20750 45118 20802
rect 45602 20750 45614 20802
rect 45666 20750 45678 20802
rect 26350 20738 26402 20750
rect 10558 20690 10610 20702
rect 3826 20638 3838 20690
rect 3890 20638 3902 20690
rect 10558 20626 10610 20638
rect 10670 20690 10722 20702
rect 10670 20626 10722 20638
rect 14142 20690 14194 20702
rect 14142 20626 14194 20638
rect 15374 20690 15426 20702
rect 16718 20690 16770 20702
rect 15474 20638 15486 20690
rect 15538 20687 15550 20690
rect 15922 20687 15934 20690
rect 15538 20641 15934 20687
rect 15538 20638 15550 20641
rect 15922 20638 15934 20641
rect 15986 20638 15998 20690
rect 15374 20626 15426 20638
rect 16718 20626 16770 20638
rect 24110 20690 24162 20702
rect 26574 20690 26626 20702
rect 25442 20638 25454 20690
rect 25506 20638 25518 20690
rect 24110 20626 24162 20638
rect 26574 20626 26626 20638
rect 28366 20690 28418 20702
rect 37214 20690 37266 20702
rect 45278 20690 45330 20702
rect 30706 20638 30718 20690
rect 30770 20638 30782 20690
rect 35746 20638 35758 20690
rect 35810 20638 35822 20690
rect 42914 20638 42926 20690
rect 42978 20638 42990 20690
rect 43810 20638 43822 20690
rect 43874 20638 43886 20690
rect 28366 20626 28418 20638
rect 37214 20626 37266 20638
rect 45278 20626 45330 20638
rect 8766 20578 8818 20590
rect 8766 20514 8818 20526
rect 9102 20578 9154 20590
rect 9102 20514 9154 20526
rect 10894 20578 10946 20590
rect 10894 20514 10946 20526
rect 11566 20578 11618 20590
rect 11566 20514 11618 20526
rect 13694 20578 13746 20590
rect 13694 20514 13746 20526
rect 14926 20578 14978 20590
rect 14926 20514 14978 20526
rect 15262 20578 15314 20590
rect 15262 20514 15314 20526
rect 16382 20578 16434 20590
rect 16382 20514 16434 20526
rect 16494 20578 16546 20590
rect 16494 20514 16546 20526
rect 17278 20578 17330 20590
rect 17278 20514 17330 20526
rect 24782 20578 24834 20590
rect 24782 20514 24834 20526
rect 25118 20578 25170 20590
rect 25118 20514 25170 20526
rect 26126 20578 26178 20590
rect 26126 20514 26178 20526
rect 28030 20578 28082 20590
rect 28030 20514 28082 20526
rect 31054 20578 31106 20590
rect 31054 20514 31106 20526
rect 1344 20410 48608 20444
rect 1344 20358 19838 20410
rect 19890 20358 19942 20410
rect 19994 20358 20046 20410
rect 20098 20358 48608 20410
rect 1344 20324 48608 20358
rect 16046 20242 16098 20254
rect 15698 20190 15710 20242
rect 15762 20190 15774 20242
rect 16046 20178 16098 20190
rect 31950 20242 32002 20254
rect 31950 20178 32002 20190
rect 33182 20242 33234 20254
rect 42130 20190 42142 20242
rect 42194 20190 42206 20242
rect 33182 20178 33234 20190
rect 2158 20130 2210 20142
rect 2158 20066 2210 20078
rect 2830 20130 2882 20142
rect 2830 20066 2882 20078
rect 3278 20130 3330 20142
rect 3278 20066 3330 20078
rect 3614 20130 3666 20142
rect 3614 20066 3666 20078
rect 4174 20130 4226 20142
rect 4174 20066 4226 20078
rect 4734 20130 4786 20142
rect 4734 20066 4786 20078
rect 7982 20130 8034 20142
rect 7982 20066 8034 20078
rect 8990 20130 9042 20142
rect 16830 20130 16882 20142
rect 16594 20078 16606 20130
rect 16658 20078 16670 20130
rect 8990 20066 9042 20078
rect 16830 20066 16882 20078
rect 18398 20130 18450 20142
rect 28814 20130 28866 20142
rect 20962 20078 20974 20130
rect 21026 20078 21038 20130
rect 21522 20078 21534 20130
rect 21586 20078 21598 20130
rect 18398 20066 18450 20078
rect 28814 20066 28866 20078
rect 30158 20130 30210 20142
rect 41246 20130 41298 20142
rect 35298 20078 35310 20130
rect 35362 20078 35374 20130
rect 30158 20066 30210 20078
rect 41246 20066 41298 20078
rect 43710 20130 43762 20142
rect 45054 20130 45106 20142
rect 44370 20078 44382 20130
rect 44434 20078 44446 20130
rect 43710 20066 43762 20078
rect 45054 20066 45106 20078
rect 5406 20018 5458 20030
rect 8542 20018 8594 20030
rect 4386 19966 4398 20018
rect 4450 19966 4462 20018
rect 5618 19966 5630 20018
rect 5682 19966 5694 20018
rect 6850 19966 6862 20018
rect 6914 19966 6926 20018
rect 8306 19966 8318 20018
rect 8370 19966 8382 20018
rect 5406 19954 5458 19966
rect 8542 19954 8594 19966
rect 8766 20018 8818 20030
rect 12686 20018 12738 20030
rect 13918 20018 13970 20030
rect 9538 19966 9550 20018
rect 9602 19966 9614 20018
rect 11106 19966 11118 20018
rect 11170 19966 11182 20018
rect 11330 19966 11342 20018
rect 11394 19966 11406 20018
rect 11890 19966 11902 20018
rect 11954 19966 11966 20018
rect 12786 19966 12798 20018
rect 12850 19966 12862 20018
rect 13682 19966 13694 20018
rect 13746 19966 13758 20018
rect 8766 19954 8818 19966
rect 12686 19954 12738 19966
rect 13918 19954 13970 19966
rect 14030 20018 14082 20030
rect 14030 19954 14082 19966
rect 15150 20018 15202 20030
rect 18734 20018 18786 20030
rect 28926 20018 28978 20030
rect 16034 19966 16046 20018
rect 16098 19966 16110 20018
rect 25554 19966 25566 20018
rect 25618 19966 25630 20018
rect 15150 19954 15202 19966
rect 18734 19954 18786 19966
rect 28926 19954 28978 19966
rect 30046 20018 30098 20030
rect 30046 19954 30098 19966
rect 30382 20018 30434 20030
rect 30382 19954 30434 19966
rect 31614 20018 31666 20030
rect 31614 19954 31666 19966
rect 31838 20018 31890 20030
rect 31838 19954 31890 19966
rect 32174 20018 32226 20030
rect 40910 20018 40962 20030
rect 34626 19966 34638 20018
rect 34690 19966 34702 20018
rect 37762 19966 37774 20018
rect 37826 19966 37838 20018
rect 32174 19954 32226 19966
rect 40910 19954 40962 19966
rect 41582 20018 41634 20030
rect 41582 19954 41634 19966
rect 41806 20018 41858 20030
rect 41806 19954 41858 19966
rect 42478 20018 42530 20030
rect 42478 19954 42530 19966
rect 43038 20018 43090 20030
rect 44046 20018 44098 20030
rect 43474 19966 43486 20018
rect 43538 19966 43550 20018
rect 45378 19966 45390 20018
rect 45442 19966 45454 20018
rect 43038 19954 43090 19966
rect 44046 19954 44098 19966
rect 4958 19906 5010 19918
rect 7422 19906 7474 19918
rect 4050 19854 4062 19906
rect 4114 19854 4126 19906
rect 5730 19854 5742 19906
rect 5794 19854 5806 19906
rect 6402 19854 6414 19906
rect 6466 19854 6478 19906
rect 4958 19842 5010 19854
rect 7422 19842 7474 19854
rect 8654 19906 8706 19918
rect 8654 19842 8706 19854
rect 10110 19906 10162 19918
rect 15374 19906 15426 19918
rect 30830 19906 30882 19918
rect 11778 19854 11790 19906
rect 11842 19854 11854 19906
rect 26226 19854 26238 19906
rect 26290 19854 26302 19906
rect 28354 19854 28366 19906
rect 28418 19854 28430 19906
rect 37426 19854 37438 19906
rect 37490 19854 37502 19906
rect 40114 19854 40126 19906
rect 40178 19854 40190 19906
rect 46050 19854 46062 19906
rect 46114 19854 46126 19906
rect 48178 19854 48190 19906
rect 48242 19854 48254 19906
rect 10110 19842 10162 19854
rect 15374 19842 15426 19854
rect 30830 19842 30882 19854
rect 3726 19794 3778 19806
rect 3726 19730 3778 19742
rect 5070 19794 5122 19806
rect 5070 19730 5122 19742
rect 9886 19794 9938 19806
rect 20414 19794 20466 19806
rect 13346 19742 13358 19794
rect 13410 19742 13422 19794
rect 14466 19742 14478 19794
rect 14530 19742 14542 19794
rect 16258 19742 16270 19794
rect 16322 19742 16334 19794
rect 9886 19730 9938 19742
rect 20414 19730 20466 19742
rect 20750 19794 20802 19806
rect 20750 19730 20802 19742
rect 28814 19794 28866 19806
rect 30594 19742 30606 19794
rect 30658 19791 30670 19794
rect 30818 19791 30830 19794
rect 30658 19745 30830 19791
rect 30658 19742 30670 19745
rect 30818 19742 30830 19745
rect 30882 19742 30894 19794
rect 28814 19730 28866 19742
rect 1344 19626 48608 19660
rect 1344 19574 4478 19626
rect 4530 19574 4582 19626
rect 4634 19574 4686 19626
rect 4738 19574 35198 19626
rect 35250 19574 35302 19626
rect 35354 19574 35406 19626
rect 35458 19574 48608 19626
rect 1344 19540 48608 19574
rect 4846 19458 4898 19470
rect 2034 19406 2046 19458
rect 2098 19455 2110 19458
rect 2930 19455 2942 19458
rect 2098 19409 2942 19455
rect 2098 19406 2110 19409
rect 2930 19406 2942 19409
rect 2994 19406 3006 19458
rect 4846 19394 4898 19406
rect 11230 19458 11282 19470
rect 14254 19458 14306 19470
rect 42366 19458 42418 19470
rect 11778 19406 11790 19458
rect 11842 19455 11854 19458
rect 12226 19455 12238 19458
rect 11842 19409 12238 19455
rect 11842 19406 11854 19409
rect 12226 19406 12238 19409
rect 12290 19406 12302 19458
rect 15250 19406 15262 19458
rect 15314 19406 15326 19458
rect 11230 19394 11282 19406
rect 14254 19394 14306 19406
rect 42366 19394 42418 19406
rect 47966 19458 48018 19470
rect 47966 19394 48018 19406
rect 2158 19346 2210 19358
rect 2158 19282 2210 19294
rect 2494 19346 2546 19358
rect 2494 19282 2546 19294
rect 2942 19346 2994 19358
rect 2942 19282 2994 19294
rect 3502 19346 3554 19358
rect 3502 19282 3554 19294
rect 5854 19346 5906 19358
rect 5854 19282 5906 19294
rect 6302 19346 6354 19358
rect 6302 19282 6354 19294
rect 7086 19346 7138 19358
rect 7086 19282 7138 19294
rect 8766 19346 8818 19358
rect 8766 19282 8818 19294
rect 10110 19346 10162 19358
rect 11790 19346 11842 19358
rect 10770 19294 10782 19346
rect 10834 19294 10846 19346
rect 10110 19282 10162 19294
rect 11790 19282 11842 19294
rect 13022 19346 13074 19358
rect 13022 19282 13074 19294
rect 15822 19346 15874 19358
rect 26462 19346 26514 19358
rect 16706 19294 16718 19346
rect 16770 19294 16782 19346
rect 18610 19294 18622 19346
rect 18674 19294 18686 19346
rect 20738 19294 20750 19346
rect 20802 19294 20814 19346
rect 25554 19294 25566 19346
rect 25618 19294 25630 19346
rect 15822 19282 15874 19294
rect 26462 19282 26514 19294
rect 30158 19346 30210 19358
rect 30158 19282 30210 19294
rect 32174 19346 32226 19358
rect 41022 19346 41074 19358
rect 33954 19294 33966 19346
rect 34018 19294 34030 19346
rect 35970 19294 35982 19346
rect 36034 19294 36046 19346
rect 39890 19294 39902 19346
rect 39954 19294 39966 19346
rect 32174 19282 32226 19294
rect 41022 19282 41074 19294
rect 42926 19346 42978 19358
rect 42926 19282 42978 19294
rect 43374 19346 43426 19358
rect 44942 19346 44994 19358
rect 43810 19294 43822 19346
rect 43874 19294 43886 19346
rect 43374 19282 43426 19294
rect 44942 19282 44994 19294
rect 3726 19234 3778 19246
rect 3726 19170 3778 19182
rect 3950 19234 4002 19246
rect 3950 19170 4002 19182
rect 4398 19234 4450 19246
rect 4398 19170 4450 19182
rect 4958 19234 5010 19246
rect 4958 19170 5010 19182
rect 8094 19234 8146 19246
rect 8094 19170 8146 19182
rect 8206 19234 8258 19246
rect 8206 19170 8258 19182
rect 8430 19234 8482 19246
rect 8430 19170 8482 19182
rect 8990 19234 9042 19246
rect 12238 19234 12290 19246
rect 10434 19182 10446 19234
rect 10498 19182 10510 19234
rect 8990 19170 9042 19182
rect 12238 19170 12290 19182
rect 13918 19234 13970 19246
rect 13918 19170 13970 19182
rect 14142 19234 14194 19246
rect 14142 19170 14194 19182
rect 14366 19234 14418 19246
rect 14366 19170 14418 19182
rect 14702 19234 14754 19246
rect 14702 19170 14754 19182
rect 14926 19234 14978 19246
rect 14926 19170 14978 19182
rect 16494 19234 16546 19246
rect 16494 19170 16546 19182
rect 17278 19234 17330 19246
rect 21310 19234 21362 19246
rect 26350 19234 26402 19246
rect 17826 19182 17838 19234
rect 17890 19182 17902 19234
rect 22642 19182 22654 19234
rect 22706 19182 22718 19234
rect 17278 19170 17330 19182
rect 21310 19170 21362 19182
rect 26350 19170 26402 19182
rect 26574 19234 26626 19246
rect 26574 19170 26626 19182
rect 27022 19234 27074 19246
rect 27022 19170 27074 19182
rect 29486 19234 29538 19246
rect 29486 19170 29538 19182
rect 29934 19234 29986 19246
rect 29934 19170 29986 19182
rect 30270 19234 30322 19246
rect 30270 19170 30322 19182
rect 30830 19234 30882 19246
rect 30830 19170 30882 19182
rect 31278 19234 31330 19246
rect 32286 19234 32338 19246
rect 31826 19182 31838 19234
rect 31890 19182 31902 19234
rect 31278 19170 31330 19182
rect 32286 19170 32338 19182
rect 32398 19234 32450 19246
rect 32398 19170 32450 19182
rect 33182 19234 33234 19246
rect 33182 19170 33234 19182
rect 33294 19234 33346 19246
rect 34414 19234 34466 19246
rect 41694 19234 41746 19246
rect 33506 19182 33518 19234
rect 33570 19182 33582 19234
rect 33842 19182 33854 19234
rect 33906 19182 33918 19234
rect 37538 19182 37550 19234
rect 37602 19182 37614 19234
rect 33294 19170 33346 19182
rect 34414 19170 34466 19182
rect 41694 19170 41746 19182
rect 42030 19234 42082 19246
rect 42030 19170 42082 19182
rect 44718 19234 44770 19246
rect 45602 19182 45614 19234
rect 45666 19182 45678 19234
rect 44718 19170 44770 19182
rect 8654 19122 8706 19134
rect 8654 19058 8706 19070
rect 9326 19122 9378 19134
rect 9326 19058 9378 19070
rect 11342 19122 11394 19134
rect 11342 19058 11394 19070
rect 13694 19122 13746 19134
rect 13694 19058 13746 19070
rect 16270 19122 16322 19134
rect 16270 19058 16322 19070
rect 16830 19122 16882 19134
rect 16830 19058 16882 19070
rect 17390 19122 17442 19134
rect 29150 19122 29202 19134
rect 23426 19070 23438 19122
rect 23490 19070 23502 19122
rect 17390 19058 17442 19070
rect 29150 19058 29202 19070
rect 29262 19122 29314 19134
rect 29262 19058 29314 19070
rect 29710 19122 29762 19134
rect 29710 19058 29762 19070
rect 30606 19122 30658 19134
rect 30606 19058 30658 19070
rect 32846 19122 32898 19134
rect 32846 19058 32898 19070
rect 34862 19122 34914 19134
rect 34862 19058 34914 19070
rect 35422 19122 35474 19134
rect 35422 19058 35474 19070
rect 41358 19122 41410 19134
rect 41358 19058 41410 19070
rect 42254 19122 42306 19134
rect 42254 19058 42306 19070
rect 4174 19010 4226 19022
rect 4174 18946 4226 18958
rect 4286 19010 4338 19022
rect 4286 18946 4338 18958
rect 7422 19010 7474 19022
rect 7422 18946 7474 18958
rect 9214 19010 9266 19022
rect 9214 18946 9266 18958
rect 16718 19010 16770 19022
rect 16718 18946 16770 18958
rect 17614 19010 17666 19022
rect 17614 18946 17666 18958
rect 21646 19010 21698 19022
rect 21646 18946 21698 18958
rect 26126 19010 26178 19022
rect 26126 18946 26178 18958
rect 28590 19010 28642 19022
rect 28590 18946 28642 18958
rect 30942 19010 30994 19022
rect 30942 18946 30994 18958
rect 32062 19010 32114 19022
rect 32062 18946 32114 18958
rect 33070 19010 33122 19022
rect 33070 18946 33122 18958
rect 34078 19010 34130 19022
rect 34078 18946 34130 18958
rect 34302 19010 34354 19022
rect 34302 18946 34354 18958
rect 36430 19010 36482 19022
rect 36430 18946 36482 18958
rect 37214 19010 37266 19022
rect 37214 18946 37266 18958
rect 40462 19010 40514 19022
rect 40462 18946 40514 18958
rect 41694 19010 41746 19022
rect 41694 18946 41746 18958
rect 42366 19010 42418 19022
rect 42366 18946 42418 18958
rect 44270 19010 44322 19022
rect 44270 18946 44322 18958
rect 45054 19010 45106 19022
rect 45054 18946 45106 18958
rect 45278 19010 45330 19022
rect 45278 18946 45330 18958
rect 1344 18842 48608 18876
rect 1344 18790 19838 18842
rect 19890 18790 19942 18842
rect 19994 18790 20046 18842
rect 20098 18790 48608 18842
rect 1344 18756 48608 18790
rect 5294 18674 5346 18686
rect 5294 18610 5346 18622
rect 7422 18674 7474 18686
rect 7422 18610 7474 18622
rect 10222 18674 10274 18686
rect 5070 18562 5122 18574
rect 7746 18566 7758 18618
rect 7810 18566 7822 18618
rect 10222 18610 10274 18622
rect 12126 18674 12178 18686
rect 12126 18610 12178 18622
rect 16046 18674 16098 18686
rect 16046 18610 16098 18622
rect 18622 18674 18674 18686
rect 18622 18610 18674 18622
rect 25454 18674 25506 18686
rect 25454 18610 25506 18622
rect 29710 18674 29762 18686
rect 29710 18610 29762 18622
rect 30382 18674 30434 18686
rect 30382 18610 30434 18622
rect 31278 18674 31330 18686
rect 31278 18610 31330 18622
rect 31950 18674 32002 18686
rect 31950 18610 32002 18622
rect 32174 18674 32226 18686
rect 32174 18610 32226 18622
rect 39006 18674 39058 18686
rect 39006 18610 39058 18622
rect 40462 18674 40514 18686
rect 40462 18610 40514 18622
rect 42702 18674 42754 18686
rect 42702 18610 42754 18622
rect 43710 18674 43762 18686
rect 43710 18610 43762 18622
rect 45614 18674 45666 18686
rect 45614 18610 45666 18622
rect 46510 18674 46562 18686
rect 46510 18610 46562 18622
rect 47182 18674 47234 18686
rect 47182 18610 47234 18622
rect 11118 18562 11170 18574
rect 7074 18510 7086 18562
rect 7138 18510 7150 18562
rect 10770 18510 10782 18562
rect 10834 18510 10846 18562
rect 5070 18498 5122 18510
rect 11118 18498 11170 18510
rect 11454 18562 11506 18574
rect 13246 18562 13298 18574
rect 12898 18510 12910 18562
rect 12962 18510 12974 18562
rect 11454 18498 11506 18510
rect 13246 18498 13298 18510
rect 13470 18562 13522 18574
rect 13470 18498 13522 18510
rect 14590 18562 14642 18574
rect 14590 18498 14642 18510
rect 16606 18562 16658 18574
rect 25902 18562 25954 18574
rect 19506 18510 19518 18562
rect 19570 18510 19582 18562
rect 21746 18510 21758 18562
rect 21810 18510 21822 18562
rect 16606 18498 16658 18510
rect 25902 18498 25954 18510
rect 26574 18562 26626 18574
rect 28366 18562 28418 18574
rect 27234 18510 27246 18562
rect 27298 18510 27310 18562
rect 26574 18498 26626 18510
rect 28366 18498 28418 18510
rect 28478 18562 28530 18574
rect 28478 18498 28530 18510
rect 29934 18562 29986 18574
rect 29934 18498 29986 18510
rect 30158 18562 30210 18574
rect 30158 18498 30210 18510
rect 31166 18562 31218 18574
rect 45838 18562 45890 18574
rect 36418 18510 36430 18562
rect 36482 18510 36494 18562
rect 31166 18498 31218 18510
rect 45838 18498 45890 18510
rect 47854 18562 47906 18574
rect 47854 18498 47906 18510
rect 5518 18450 5570 18462
rect 9774 18450 9826 18462
rect 12574 18450 12626 18462
rect 18958 18450 19010 18462
rect 24222 18450 24274 18462
rect 1810 18398 1822 18450
rect 1874 18398 1886 18450
rect 7970 18398 7982 18450
rect 8034 18398 8046 18450
rect 11890 18398 11902 18450
rect 11954 18398 11966 18450
rect 13682 18398 13694 18450
rect 13746 18398 13758 18450
rect 16258 18398 16270 18450
rect 16322 18398 16334 18450
rect 19618 18398 19630 18450
rect 19682 18398 19694 18450
rect 21074 18398 21086 18450
rect 21138 18398 21150 18450
rect 5518 18386 5570 18398
rect 9774 18386 9826 18398
rect 12574 18386 12626 18398
rect 18958 18386 19010 18398
rect 24222 18386 24274 18398
rect 25342 18450 25394 18462
rect 25342 18386 25394 18398
rect 25678 18450 25730 18462
rect 25678 18386 25730 18398
rect 26350 18450 26402 18462
rect 26350 18386 26402 18398
rect 27022 18450 27074 18462
rect 27022 18386 27074 18398
rect 27582 18450 27634 18462
rect 27582 18386 27634 18398
rect 28142 18450 28194 18462
rect 31502 18450 31554 18462
rect 30594 18398 30606 18450
rect 30658 18398 30670 18450
rect 28142 18386 28194 18398
rect 31502 18386 31554 18398
rect 31838 18450 31890 18462
rect 36094 18450 36146 18462
rect 38446 18450 38498 18462
rect 39902 18450 39954 18462
rect 32386 18398 32398 18450
rect 32450 18398 32462 18450
rect 35298 18398 35310 18450
rect 35362 18398 35374 18450
rect 37090 18398 37102 18450
rect 37154 18398 37166 18450
rect 37874 18398 37886 18450
rect 37938 18398 37950 18450
rect 39442 18398 39454 18450
rect 39506 18398 39518 18450
rect 39666 18398 39678 18450
rect 39730 18398 39742 18450
rect 31838 18386 31890 18398
rect 36094 18386 36146 18398
rect 38446 18386 38498 18398
rect 39902 18386 39954 18398
rect 40350 18450 40402 18462
rect 42142 18450 42194 18462
rect 41794 18398 41806 18450
rect 41858 18398 41870 18450
rect 40350 18386 40402 18398
rect 42142 18386 42194 18398
rect 42590 18450 42642 18462
rect 42590 18386 42642 18398
rect 43262 18450 43314 18462
rect 43262 18386 43314 18398
rect 43486 18450 43538 18462
rect 43486 18386 43538 18398
rect 43934 18450 43986 18462
rect 47518 18450 47570 18462
rect 44818 18398 44830 18450
rect 44882 18398 44894 18450
rect 46050 18398 46062 18450
rect 46114 18398 46126 18450
rect 46722 18398 46734 18450
rect 46786 18398 46798 18450
rect 43934 18386 43986 18398
rect 47518 18386 47570 18398
rect 48190 18450 48242 18462
rect 48190 18386 48242 18398
rect 5182 18338 5234 18350
rect 2482 18286 2494 18338
rect 2546 18286 2558 18338
rect 4610 18286 4622 18338
rect 4674 18286 4686 18338
rect 5182 18274 5234 18286
rect 6190 18338 6242 18350
rect 6190 18274 6242 18286
rect 6750 18338 6802 18350
rect 6750 18274 6802 18286
rect 9102 18338 9154 18350
rect 9102 18274 9154 18286
rect 11566 18338 11618 18350
rect 11566 18274 11618 18286
rect 13582 18338 13634 18350
rect 13582 18274 13634 18286
rect 14702 18338 14754 18350
rect 14702 18274 14754 18286
rect 17502 18338 17554 18350
rect 24334 18338 24386 18350
rect 23874 18286 23886 18338
rect 23938 18286 23950 18338
rect 17502 18274 17554 18286
rect 24334 18274 24386 18286
rect 25566 18338 25618 18350
rect 25566 18274 25618 18286
rect 26798 18338 26850 18350
rect 26798 18274 26850 18286
rect 30270 18338 30322 18350
rect 40126 18338 40178 18350
rect 32274 18286 32286 18338
rect 32338 18286 32350 18338
rect 34066 18286 34078 18338
rect 34130 18286 34142 18338
rect 37538 18286 37550 18338
rect 37602 18286 37614 18338
rect 30270 18274 30322 18286
rect 40126 18274 40178 18286
rect 42254 18338 42306 18350
rect 42254 18274 42306 18286
rect 44046 18338 44098 18350
rect 45278 18338 45330 18350
rect 46398 18338 46450 18350
rect 44370 18286 44382 18338
rect 44434 18286 44446 18338
rect 45714 18286 45726 18338
rect 45778 18286 45790 18338
rect 44046 18274 44098 18286
rect 45278 18274 45330 18286
rect 46398 18274 46450 18286
rect 5742 18226 5794 18238
rect 12238 18226 12290 18238
rect 9874 18174 9886 18226
rect 9938 18223 9950 18226
rect 10322 18223 10334 18226
rect 9938 18177 10334 18223
rect 9938 18174 9950 18177
rect 10322 18174 10334 18177
rect 10386 18174 10398 18226
rect 5742 18162 5794 18174
rect 12238 18162 12290 18174
rect 14814 18226 14866 18238
rect 14814 18162 14866 18174
rect 16270 18226 16322 18238
rect 42702 18226 42754 18238
rect 37090 18174 37102 18226
rect 37154 18174 37166 18226
rect 16270 18162 16322 18174
rect 42702 18162 42754 18174
rect 1344 18058 48608 18092
rect 1344 18006 4478 18058
rect 4530 18006 4582 18058
rect 4634 18006 4686 18058
rect 4738 18006 35198 18058
rect 35250 18006 35302 18058
rect 35354 18006 35406 18058
rect 35458 18006 48608 18058
rect 1344 17972 48608 18006
rect 8990 17890 9042 17902
rect 7186 17838 7198 17890
rect 7250 17838 7262 17890
rect 38658 17838 38670 17890
rect 38722 17838 38734 17890
rect 8990 17826 9042 17838
rect 1934 17778 1986 17790
rect 13582 17778 13634 17790
rect 30830 17778 30882 17790
rect 7074 17726 7086 17778
rect 7138 17726 7150 17778
rect 9538 17726 9550 17778
rect 9602 17726 9614 17778
rect 14690 17726 14702 17778
rect 14754 17726 14766 17778
rect 16818 17726 16830 17778
rect 16882 17726 16894 17778
rect 20066 17726 20078 17778
rect 20130 17726 20142 17778
rect 28578 17726 28590 17778
rect 28642 17726 28654 17778
rect 1934 17714 1986 17726
rect 13582 17714 13634 17726
rect 30830 17714 30882 17726
rect 31278 17778 31330 17790
rect 31278 17714 31330 17726
rect 36430 17778 36482 17790
rect 42702 17778 42754 17790
rect 40450 17726 40462 17778
rect 40514 17726 40526 17778
rect 36430 17714 36482 17726
rect 42702 17714 42754 17726
rect 43486 17778 43538 17790
rect 43486 17714 43538 17726
rect 44158 17778 44210 17790
rect 44158 17714 44210 17726
rect 44942 17778 44994 17790
rect 48178 17726 48190 17778
rect 48242 17726 48254 17778
rect 44942 17714 44994 17726
rect 5630 17666 5682 17678
rect 8654 17666 8706 17678
rect 3826 17614 3838 17666
rect 3890 17614 3902 17666
rect 6402 17614 6414 17666
rect 6466 17614 6478 17666
rect 5630 17602 5682 17614
rect 8654 17602 8706 17614
rect 9774 17666 9826 17678
rect 11678 17666 11730 17678
rect 9874 17614 9886 17666
rect 9938 17614 9950 17666
rect 11442 17614 11454 17666
rect 11506 17614 11518 17666
rect 9774 17602 9826 17614
rect 11678 17602 11730 17614
rect 12238 17666 12290 17678
rect 12238 17602 12290 17614
rect 12686 17666 12738 17678
rect 29822 17666 29874 17678
rect 14018 17614 14030 17666
rect 14082 17614 14094 17666
rect 19730 17614 19742 17666
rect 19794 17614 19806 17666
rect 21858 17614 21870 17666
rect 21922 17614 21934 17666
rect 25778 17614 25790 17666
rect 25842 17614 25854 17666
rect 29586 17614 29598 17666
rect 29650 17614 29662 17666
rect 12686 17602 12738 17614
rect 29822 17602 29874 17614
rect 30046 17666 30098 17678
rect 30046 17602 30098 17614
rect 30158 17666 30210 17678
rect 30158 17602 30210 17614
rect 31838 17666 31890 17678
rect 31838 17602 31890 17614
rect 32174 17666 32226 17678
rect 32174 17602 32226 17614
rect 32286 17666 32338 17678
rect 32286 17602 32338 17614
rect 32510 17666 32562 17678
rect 35982 17666 36034 17678
rect 41918 17666 41970 17678
rect 35186 17614 35198 17666
rect 35250 17614 35262 17666
rect 37090 17614 37102 17666
rect 37154 17614 37166 17666
rect 38210 17614 38222 17666
rect 38274 17614 38286 17666
rect 39218 17614 39230 17666
rect 39282 17614 39294 17666
rect 40338 17614 40350 17666
rect 40402 17614 40414 17666
rect 32510 17602 32562 17614
rect 35982 17602 36034 17614
rect 41918 17602 41970 17614
rect 42030 17666 42082 17678
rect 42030 17602 42082 17614
rect 43598 17666 43650 17678
rect 45378 17614 45390 17666
rect 45442 17614 45454 17666
rect 43598 17602 43650 17614
rect 5854 17554 5906 17566
rect 4722 17502 4734 17554
rect 4786 17502 4798 17554
rect 5854 17490 5906 17502
rect 5966 17554 6018 17566
rect 5966 17490 6018 17502
rect 6750 17554 6802 17566
rect 6750 17490 6802 17502
rect 8206 17554 8258 17566
rect 8206 17490 8258 17502
rect 8878 17554 8930 17566
rect 8878 17490 8930 17502
rect 12910 17554 12962 17566
rect 18958 17554 19010 17566
rect 32958 17554 33010 17566
rect 42366 17554 42418 17566
rect 17826 17502 17838 17554
rect 17890 17502 17902 17554
rect 26450 17502 26462 17554
rect 26514 17502 26526 17554
rect 33506 17502 33518 17554
rect 33570 17502 33582 17554
rect 34290 17502 34302 17554
rect 34354 17502 34366 17554
rect 35634 17502 35646 17554
rect 35698 17502 35710 17554
rect 12910 17490 12962 17502
rect 18958 17490 19010 17502
rect 32958 17490 33010 17502
rect 42366 17490 42418 17502
rect 42814 17554 42866 17566
rect 46050 17502 46062 17554
rect 46114 17502 46126 17554
rect 42814 17490 42866 17502
rect 5070 17442 5122 17454
rect 5070 17378 5122 17390
rect 5742 17442 5794 17454
rect 11566 17442 11618 17454
rect 10098 17390 10110 17442
rect 10162 17390 10174 17442
rect 5742 17378 5794 17390
rect 11566 17378 11618 17390
rect 12574 17442 12626 17454
rect 12574 17378 12626 17390
rect 17502 17442 17554 17454
rect 17502 17378 17554 17390
rect 18286 17442 18338 17454
rect 18286 17378 18338 17390
rect 19294 17442 19346 17454
rect 19294 17378 19346 17390
rect 22094 17442 22146 17454
rect 22094 17378 22146 17390
rect 22542 17442 22594 17454
rect 22542 17378 22594 17390
rect 29934 17442 29986 17454
rect 29934 17378 29986 17390
rect 32622 17442 32674 17454
rect 32622 17378 32674 17390
rect 32846 17442 32898 17454
rect 32846 17378 32898 17390
rect 33854 17442 33906 17454
rect 33854 17378 33906 17390
rect 34638 17442 34690 17454
rect 34638 17378 34690 17390
rect 34974 17442 35026 17454
rect 34974 17378 35026 17390
rect 42142 17442 42194 17454
rect 42142 17378 42194 17390
rect 44046 17442 44098 17454
rect 44046 17378 44098 17390
rect 44270 17442 44322 17454
rect 44270 17378 44322 17390
rect 1344 17274 48608 17308
rect 1344 17222 19838 17274
rect 19890 17222 19942 17274
rect 19994 17222 20046 17274
rect 20098 17222 48608 17274
rect 1344 17188 48608 17222
rect 3278 17106 3330 17118
rect 3278 17042 3330 17054
rect 4286 17106 4338 17118
rect 4286 17042 4338 17054
rect 5070 17106 5122 17118
rect 5070 17042 5122 17054
rect 5742 17106 5794 17118
rect 5742 17042 5794 17054
rect 6638 17106 6690 17118
rect 6638 17042 6690 17054
rect 7422 17106 7474 17118
rect 7422 17042 7474 17054
rect 7646 17106 7698 17118
rect 7646 17042 7698 17054
rect 8542 17106 8594 17118
rect 8542 17042 8594 17054
rect 9886 17106 9938 17118
rect 15822 17106 15874 17118
rect 23774 17106 23826 17118
rect 14466 17054 14478 17106
rect 14530 17054 14542 17106
rect 16594 17054 16606 17106
rect 16658 17054 16670 17106
rect 9886 17042 9938 17054
rect 15822 17042 15874 17054
rect 23774 17042 23826 17054
rect 24222 17106 24274 17118
rect 24222 17042 24274 17054
rect 25230 17106 25282 17118
rect 29486 17106 29538 17118
rect 25554 17054 25566 17106
rect 25618 17054 25630 17106
rect 25230 17042 25282 17054
rect 29486 17042 29538 17054
rect 31390 17106 31442 17118
rect 31390 17042 31442 17054
rect 31726 17106 31778 17118
rect 35422 17106 35474 17118
rect 33282 17054 33294 17106
rect 33346 17054 33358 17106
rect 31726 17042 31778 17054
rect 35422 17042 35474 17054
rect 38670 17106 38722 17118
rect 38670 17042 38722 17054
rect 40238 17106 40290 17118
rect 40238 17042 40290 17054
rect 41358 17106 41410 17118
rect 46062 17106 46114 17118
rect 43698 17054 43710 17106
rect 43762 17054 43774 17106
rect 41358 17042 41410 17054
rect 46062 17042 46114 17054
rect 4958 16994 5010 17006
rect 4958 16930 5010 16942
rect 5294 16994 5346 17006
rect 14926 16994 14978 17006
rect 26574 16994 26626 17006
rect 6066 16942 6078 16994
rect 6130 16942 6142 16994
rect 9538 16942 9550 16994
rect 9602 16942 9614 16994
rect 11218 16942 11230 16994
rect 11282 16942 11294 16994
rect 13794 16942 13806 16994
rect 13858 16942 13870 16994
rect 19506 16942 19518 16994
rect 19570 16942 19582 16994
rect 5294 16930 5346 16942
rect 14926 16930 14978 16942
rect 26574 16930 26626 16942
rect 26910 16994 26962 17006
rect 26910 16930 26962 16942
rect 28926 16994 28978 17006
rect 28926 16930 28978 16942
rect 29262 16994 29314 17006
rect 29262 16930 29314 16942
rect 30270 16994 30322 17006
rect 30270 16930 30322 16942
rect 30494 16994 30546 17006
rect 30494 16930 30546 16942
rect 31502 16994 31554 17006
rect 31502 16930 31554 16942
rect 31950 16994 32002 17006
rect 39006 16994 39058 17006
rect 42814 16994 42866 17006
rect 44270 16994 44322 17006
rect 33058 16942 33070 16994
rect 33122 16942 33134 16994
rect 34962 16942 34974 16994
rect 35026 16942 35038 16994
rect 36530 16942 36542 16994
rect 36594 16942 36606 16994
rect 36866 16942 36878 16994
rect 36930 16942 36942 16994
rect 39890 16942 39902 16994
rect 39954 16942 39966 16994
rect 43250 16942 43262 16994
rect 43314 16942 43326 16994
rect 31950 16930 32002 16942
rect 39006 16930 39058 16942
rect 42814 16930 42866 16942
rect 44270 16930 44322 16942
rect 46958 16994 47010 17006
rect 46958 16930 47010 16942
rect 47518 16994 47570 17006
rect 47518 16930 47570 16942
rect 47630 16994 47682 17006
rect 47630 16930 47682 16942
rect 48078 16994 48130 17006
rect 48078 16930 48130 16942
rect 2830 16882 2882 16894
rect 4510 16882 4562 16894
rect 4162 16830 4174 16882
rect 4226 16830 4238 16882
rect 2830 16818 2882 16830
rect 4510 16818 4562 16830
rect 8094 16882 8146 16894
rect 16270 16882 16322 16894
rect 17950 16882 18002 16894
rect 22318 16882 22370 16894
rect 10322 16830 10334 16882
rect 10386 16830 10398 16882
rect 12114 16830 12126 16882
rect 12178 16830 12190 16882
rect 14130 16830 14142 16882
rect 14194 16830 14206 16882
rect 17490 16830 17502 16882
rect 17554 16830 17566 16882
rect 18722 16830 18734 16882
rect 18786 16830 18798 16882
rect 8094 16818 8146 16830
rect 16270 16818 16322 16830
rect 17950 16818 18002 16830
rect 22318 16818 22370 16830
rect 22542 16882 22594 16894
rect 22542 16818 22594 16830
rect 23214 16882 23266 16894
rect 23214 16818 23266 16830
rect 26350 16882 26402 16894
rect 26350 16818 26402 16830
rect 26798 16882 26850 16894
rect 26798 16818 26850 16830
rect 29486 16882 29538 16894
rect 29486 16818 29538 16830
rect 29822 16882 29874 16894
rect 39230 16882 39282 16894
rect 40910 16882 40962 16894
rect 33506 16830 33518 16882
rect 33570 16830 33582 16882
rect 34178 16830 34190 16882
rect 34242 16830 34254 16882
rect 34402 16830 34414 16882
rect 34466 16830 34478 16882
rect 36194 16830 36206 16882
rect 36258 16830 36270 16882
rect 37202 16830 37214 16882
rect 37266 16830 37278 16882
rect 37762 16830 37774 16882
rect 37826 16830 37838 16882
rect 39554 16830 39566 16882
rect 39618 16830 39630 16882
rect 29822 16818 29874 16830
rect 39230 16818 39282 16830
rect 40910 16818 40962 16830
rect 41134 16882 41186 16894
rect 41134 16818 41186 16830
rect 42702 16882 42754 16894
rect 45726 16882 45778 16894
rect 43810 16830 43822 16882
rect 43874 16830 43886 16882
rect 44818 16830 44830 16882
rect 44882 16830 44894 16882
rect 42702 16818 42754 16830
rect 45726 16818 45778 16830
rect 46174 16882 46226 16894
rect 46174 16818 46226 16830
rect 46286 16882 46338 16894
rect 46286 16818 46338 16830
rect 47294 16882 47346 16894
rect 47294 16818 47346 16830
rect 3166 16770 3218 16782
rect 7534 16770 7586 16782
rect 4386 16718 4398 16770
rect 4450 16718 4462 16770
rect 3166 16706 3218 16718
rect 7534 16706 7586 16718
rect 7870 16770 7922 16782
rect 7870 16706 7922 16718
rect 16046 16770 16098 16782
rect 31614 16770 31666 16782
rect 21634 16718 21646 16770
rect 21698 16718 21710 16770
rect 30146 16718 30158 16770
rect 30210 16718 30222 16770
rect 16046 16706 16098 16718
rect 31614 16706 31666 16718
rect 38110 16770 38162 16782
rect 38110 16706 38162 16718
rect 38222 16770 38274 16782
rect 38222 16706 38274 16718
rect 39118 16770 39170 16782
rect 39118 16706 39170 16718
rect 41022 16770 41074 16782
rect 41022 16706 41074 16718
rect 41806 16770 41858 16782
rect 45502 16770 45554 16782
rect 44706 16718 44718 16770
rect 44770 16718 44782 16770
rect 41806 16706 41858 16718
rect 45502 16706 45554 16718
rect 46846 16770 46898 16782
rect 46846 16706 46898 16718
rect 3614 16658 3666 16670
rect 3614 16594 3666 16606
rect 3838 16658 3890 16670
rect 26126 16658 26178 16670
rect 22866 16606 22878 16658
rect 22930 16606 22942 16658
rect 3838 16594 3890 16606
rect 26126 16594 26178 16606
rect 41918 16658 41970 16670
rect 41918 16594 41970 16606
rect 42142 16658 42194 16670
rect 42142 16594 42194 16606
rect 42254 16658 42306 16670
rect 42254 16594 42306 16606
rect 42814 16658 42866 16670
rect 42814 16594 42866 16606
rect 46734 16658 46786 16670
rect 46734 16594 46786 16606
rect 1344 16490 48608 16524
rect 1344 16438 4478 16490
rect 4530 16438 4582 16490
rect 4634 16438 4686 16490
rect 4738 16438 35198 16490
rect 35250 16438 35302 16490
rect 35354 16438 35406 16490
rect 35458 16438 48608 16490
rect 1344 16404 48608 16438
rect 7198 16322 7250 16334
rect 7198 16258 7250 16270
rect 11902 16322 11954 16334
rect 11902 16258 11954 16270
rect 18958 16322 19010 16334
rect 18958 16258 19010 16270
rect 19294 16322 19346 16334
rect 19294 16258 19346 16270
rect 34862 16322 34914 16334
rect 38670 16322 38722 16334
rect 37650 16270 37662 16322
rect 37714 16270 37726 16322
rect 34862 16258 34914 16270
rect 38670 16258 38722 16270
rect 39230 16322 39282 16334
rect 39230 16258 39282 16270
rect 40686 16322 40738 16334
rect 40686 16258 40738 16270
rect 43374 16322 43426 16334
rect 44930 16270 44942 16322
rect 44994 16270 45006 16322
rect 43374 16258 43426 16270
rect 5070 16210 5122 16222
rect 1698 16158 1710 16210
rect 1762 16158 1774 16210
rect 3826 16158 3838 16210
rect 3890 16158 3902 16210
rect 5070 16146 5122 16158
rect 5854 16210 5906 16222
rect 5854 16146 5906 16158
rect 6190 16210 6242 16222
rect 6190 16146 6242 16158
rect 7646 16210 7698 16222
rect 20750 16210 20802 16222
rect 25902 16210 25954 16222
rect 14578 16158 14590 16210
rect 14642 16158 14654 16210
rect 21746 16158 21758 16210
rect 21810 16158 21822 16210
rect 7646 16146 7698 16158
rect 20750 16146 20802 16158
rect 25902 16146 25954 16158
rect 27918 16210 27970 16222
rect 27918 16146 27970 16158
rect 29262 16210 29314 16222
rect 29262 16146 29314 16158
rect 30158 16210 30210 16222
rect 30158 16146 30210 16158
rect 33854 16210 33906 16222
rect 33854 16146 33906 16158
rect 35646 16210 35698 16222
rect 35646 16146 35698 16158
rect 43038 16210 43090 16222
rect 43038 16146 43090 16158
rect 44382 16210 44434 16222
rect 46958 16210 47010 16222
rect 46386 16158 46398 16210
rect 46450 16158 46462 16210
rect 44382 16146 44434 16158
rect 46958 16146 47010 16158
rect 7422 16098 7474 16110
rect 4610 16046 4622 16098
rect 4674 16046 4686 16098
rect 7422 16034 7474 16046
rect 8094 16098 8146 16110
rect 8094 16034 8146 16046
rect 9998 16098 10050 16110
rect 9998 16034 10050 16046
rect 12238 16098 12290 16110
rect 12238 16034 12290 16046
rect 12686 16098 12738 16110
rect 16942 16098 16994 16110
rect 23886 16098 23938 16110
rect 14018 16046 14030 16098
rect 14082 16046 14094 16098
rect 20066 16046 20078 16098
rect 20130 16046 20142 16098
rect 22418 16046 22430 16098
rect 22482 16046 22494 16098
rect 23650 16046 23662 16098
rect 23714 16046 23726 16098
rect 12686 16034 12738 16046
rect 16942 16034 16994 16046
rect 23886 16034 23938 16046
rect 24670 16098 24722 16110
rect 28254 16098 28306 16110
rect 25666 16046 25678 16098
rect 25730 16046 25742 16098
rect 24670 16034 24722 16046
rect 28254 16034 28306 16046
rect 29038 16098 29090 16110
rect 29038 16034 29090 16046
rect 29710 16098 29762 16110
rect 29710 16034 29762 16046
rect 31726 16098 31778 16110
rect 35198 16098 35250 16110
rect 31938 16046 31950 16098
rect 32002 16046 32014 16098
rect 34290 16046 34302 16098
rect 34354 16046 34366 16098
rect 31726 16034 31778 16046
rect 35198 16034 35250 16046
rect 35534 16098 35586 16110
rect 35534 16034 35586 16046
rect 36206 16098 36258 16110
rect 37998 16098 38050 16110
rect 37202 16046 37214 16098
rect 37266 16046 37278 16098
rect 37650 16046 37662 16098
rect 37714 16046 37726 16098
rect 36206 16034 36258 16046
rect 37998 16034 38050 16046
rect 39454 16098 39506 16110
rect 39454 16034 39506 16046
rect 40350 16098 40402 16110
rect 40350 16034 40402 16046
rect 40798 16098 40850 16110
rect 41582 16098 41634 16110
rect 41346 16046 41358 16098
rect 41410 16046 41422 16098
rect 40798 16034 40850 16046
rect 41582 16034 41634 16046
rect 45166 16098 45218 16110
rect 45166 16034 45218 16046
rect 45614 16098 45666 16110
rect 45614 16034 45666 16046
rect 45950 16098 46002 16110
rect 45950 16034 46002 16046
rect 9886 15986 9938 15998
rect 9886 15922 9938 15934
rect 12014 15986 12066 15998
rect 12014 15922 12066 15934
rect 12910 15986 12962 15998
rect 24334 15986 24386 15998
rect 17266 15934 17278 15986
rect 17330 15934 17342 15986
rect 19954 15934 19966 15986
rect 20018 15934 20030 15986
rect 22194 15934 22206 15986
rect 22258 15934 22270 15986
rect 23202 15934 23214 15986
rect 23266 15934 23278 15986
rect 12910 15922 12962 15934
rect 24334 15922 24386 15934
rect 26014 15986 26066 15998
rect 29486 15986 29538 15998
rect 28578 15934 28590 15986
rect 28642 15934 28654 15986
rect 26014 15922 26066 15934
rect 29486 15922 29538 15934
rect 30046 15986 30098 15998
rect 30046 15922 30098 15934
rect 30270 15986 30322 15998
rect 30270 15922 30322 15934
rect 31614 15986 31666 15998
rect 38334 15986 38386 15998
rect 34514 15934 34526 15986
rect 34578 15934 34590 15986
rect 31614 15922 31666 15934
rect 38334 15922 38386 15934
rect 38894 15986 38946 15998
rect 38894 15922 38946 15934
rect 40014 15986 40066 15998
rect 40014 15922 40066 15934
rect 41470 15986 41522 15998
rect 41470 15922 41522 15934
rect 42142 15986 42194 15998
rect 42142 15922 42194 15934
rect 42478 15986 42530 15998
rect 42478 15922 42530 15934
rect 43710 15986 43762 15998
rect 43710 15922 43762 15934
rect 47294 15986 47346 15998
rect 47294 15922 47346 15934
rect 7870 15874 7922 15886
rect 7870 15810 7922 15822
rect 7982 15874 8034 15886
rect 7982 15810 8034 15822
rect 11902 15874 11954 15886
rect 11902 15810 11954 15822
rect 12574 15874 12626 15886
rect 12574 15810 12626 15822
rect 16494 15874 16546 15886
rect 16494 15810 16546 15822
rect 21310 15874 21362 15886
rect 21310 15810 21362 15822
rect 22878 15874 22930 15886
rect 22878 15810 22930 15822
rect 23998 15874 24050 15886
rect 23998 15810 24050 15822
rect 24110 15874 24162 15886
rect 34974 15874 35026 15886
rect 24994 15822 25006 15874
rect 25058 15822 25070 15874
rect 31154 15822 31166 15874
rect 31218 15822 31230 15874
rect 24110 15810 24162 15822
rect 34974 15810 35026 15822
rect 35758 15874 35810 15886
rect 35758 15810 35810 15822
rect 38222 15874 38274 15886
rect 38222 15810 38274 15822
rect 39566 15874 39618 15886
rect 39566 15810 39618 15822
rect 40238 15874 40290 15886
rect 40238 15810 40290 15822
rect 41134 15874 41186 15886
rect 41134 15810 41186 15822
rect 42030 15874 42082 15886
rect 42030 15810 42082 15822
rect 42254 15874 42306 15886
rect 42254 15810 42306 15822
rect 43486 15874 43538 15886
rect 43486 15810 43538 15822
rect 47854 15874 47906 15886
rect 47854 15810 47906 15822
rect 1344 15706 48608 15740
rect 1344 15654 19838 15706
rect 19890 15654 19942 15706
rect 19994 15654 20046 15706
rect 20098 15654 48608 15706
rect 1344 15620 48608 15654
rect 4734 15538 4786 15550
rect 4734 15474 4786 15486
rect 4958 15538 5010 15550
rect 12238 15538 12290 15550
rect 10994 15486 11006 15538
rect 11058 15486 11070 15538
rect 4958 15474 5010 15486
rect 12238 15474 12290 15486
rect 24446 15538 24498 15550
rect 24446 15474 24498 15486
rect 27918 15538 27970 15550
rect 27918 15474 27970 15486
rect 28814 15538 28866 15550
rect 34526 15538 34578 15550
rect 36654 15538 36706 15550
rect 33058 15486 33070 15538
rect 33122 15486 33134 15538
rect 34850 15486 34862 15538
rect 34914 15486 34926 15538
rect 35858 15486 35870 15538
rect 35922 15486 35934 15538
rect 28814 15474 28866 15486
rect 34526 15474 34578 15486
rect 36654 15474 36706 15486
rect 37774 15538 37826 15550
rect 37774 15474 37826 15486
rect 37998 15538 38050 15550
rect 37998 15474 38050 15486
rect 40014 15538 40066 15550
rect 40014 15474 40066 15486
rect 41470 15538 41522 15550
rect 41470 15474 41522 15486
rect 41694 15538 41746 15550
rect 41694 15474 41746 15486
rect 43486 15538 43538 15550
rect 43486 15474 43538 15486
rect 7086 15426 7138 15438
rect 5618 15374 5630 15426
rect 5682 15374 5694 15426
rect 7086 15362 7138 15374
rect 9550 15426 9602 15438
rect 16382 15426 16434 15438
rect 13234 15374 13246 15426
rect 13298 15374 13310 15426
rect 9550 15362 9602 15374
rect 16382 15362 16434 15374
rect 16606 15426 16658 15438
rect 25342 15426 25394 15438
rect 17714 15374 17726 15426
rect 17778 15374 17790 15426
rect 19394 15374 19406 15426
rect 19458 15374 19470 15426
rect 16606 15362 16658 15374
rect 25342 15362 25394 15374
rect 27694 15426 27746 15438
rect 27694 15362 27746 15374
rect 31614 15426 31666 15438
rect 31614 15362 31666 15374
rect 31726 15426 31778 15438
rect 31726 15362 31778 15374
rect 36318 15426 36370 15438
rect 36318 15362 36370 15374
rect 37550 15426 37602 15438
rect 37550 15362 37602 15374
rect 39678 15426 39730 15438
rect 39678 15362 39730 15374
rect 39790 15426 39842 15438
rect 39790 15362 39842 15374
rect 40238 15426 40290 15438
rect 40238 15362 40290 15374
rect 40350 15426 40402 15438
rect 40350 15362 40402 15374
rect 41246 15426 41298 15438
rect 41246 15362 41298 15374
rect 44830 15426 44882 15438
rect 44830 15362 44882 15374
rect 47406 15426 47458 15438
rect 47406 15362 47458 15374
rect 5406 15314 5458 15326
rect 5406 15250 5458 15262
rect 6862 15314 6914 15326
rect 7534 15314 7586 15326
rect 11342 15314 11394 15326
rect 7186 15262 7198 15314
rect 7250 15262 7262 15314
rect 10770 15262 10782 15314
rect 10834 15262 10846 15314
rect 6862 15250 6914 15262
rect 7534 15250 7586 15262
rect 11342 15250 11394 15262
rect 11790 15314 11842 15326
rect 17390 15314 17442 15326
rect 24110 15314 24162 15326
rect 11790 15250 11842 15262
rect 12562 15250 12574 15302
rect 12626 15250 12638 15302
rect 19282 15262 19294 15314
rect 19346 15262 19358 15314
rect 21298 15262 21310 15314
rect 21362 15262 21374 15314
rect 17390 15250 17442 15262
rect 24110 15250 24162 15262
rect 24222 15314 24274 15326
rect 26126 15314 26178 15326
rect 27582 15314 27634 15326
rect 35534 15314 35586 15326
rect 24658 15262 24670 15314
rect 24722 15262 24734 15314
rect 26562 15262 26574 15314
rect 26626 15262 26638 15314
rect 31938 15262 31950 15314
rect 32002 15262 32014 15314
rect 33282 15262 33294 15314
rect 33346 15262 33358 15314
rect 34290 15262 34302 15314
rect 34354 15262 34366 15314
rect 35074 15262 35086 15314
rect 35138 15262 35150 15314
rect 24222 15250 24274 15262
rect 26126 15250 26178 15262
rect 27582 15250 27634 15262
rect 35534 15250 35586 15262
rect 36542 15314 36594 15326
rect 36542 15250 36594 15262
rect 36878 15314 36930 15326
rect 41582 15314 41634 15326
rect 43822 15314 43874 15326
rect 39106 15262 39118 15314
rect 39170 15262 39182 15314
rect 41906 15262 41918 15314
rect 41970 15262 41982 15314
rect 45938 15262 45950 15314
rect 46002 15262 46014 15314
rect 46386 15262 46398 15314
rect 46450 15262 46462 15314
rect 36878 15250 36930 15262
rect 41582 15250 41634 15262
rect 43822 15250 43874 15262
rect 4846 15202 4898 15214
rect 4846 15138 4898 15150
rect 5966 15202 6018 15214
rect 5966 15138 6018 15150
rect 6974 15202 7026 15214
rect 6974 15138 7026 15150
rect 9662 15202 9714 15214
rect 9662 15138 9714 15150
rect 10222 15202 10274 15214
rect 10222 15138 10274 15150
rect 11566 15202 11618 15214
rect 15822 15202 15874 15214
rect 18622 15202 18674 15214
rect 29822 15202 29874 15214
rect 42366 15202 42418 15214
rect 15362 15150 15374 15202
rect 15426 15150 15438 15202
rect 16258 15150 16270 15202
rect 16322 15150 16334 15202
rect 21858 15150 21870 15202
rect 21922 15150 21934 15202
rect 24434 15150 24446 15202
rect 24498 15150 24510 15202
rect 26674 15150 26686 15202
rect 26738 15150 26750 15202
rect 38770 15150 38782 15202
rect 38834 15150 38846 15202
rect 11566 15138 11618 15150
rect 15822 15138 15874 15150
rect 18622 15138 18674 15150
rect 29822 15138 29874 15150
rect 42366 15138 42418 15150
rect 42814 15202 42866 15214
rect 44594 15150 44606 15202
rect 44658 15150 44670 15202
rect 42814 15138 42866 15150
rect 18286 15090 18338 15102
rect 38110 15090 38162 15102
rect 31154 15038 31166 15090
rect 31218 15038 31230 15090
rect 18286 15026 18338 15038
rect 38110 15026 38162 15038
rect 39678 15090 39730 15102
rect 39678 15026 39730 15038
rect 1344 14922 48608 14956
rect 1344 14870 4478 14922
rect 4530 14870 4582 14922
rect 4634 14870 4686 14922
rect 4738 14870 35198 14922
rect 35250 14870 35302 14922
rect 35354 14870 35406 14922
rect 35458 14870 48608 14922
rect 1344 14836 48608 14870
rect 26574 14754 26626 14766
rect 21746 14702 21758 14754
rect 21810 14702 21822 14754
rect 26574 14690 26626 14702
rect 34414 14754 34466 14766
rect 34414 14690 34466 14702
rect 38110 14754 38162 14766
rect 38110 14690 38162 14702
rect 41582 14754 41634 14766
rect 41582 14690 41634 14702
rect 10782 14642 10834 14654
rect 2482 14590 2494 14642
rect 2546 14590 2558 14642
rect 4610 14590 4622 14642
rect 4674 14590 4686 14642
rect 7858 14590 7870 14642
rect 7922 14590 7934 14642
rect 9986 14590 9998 14642
rect 10050 14590 10062 14642
rect 10782 14578 10834 14590
rect 12014 14642 12066 14654
rect 28590 14642 28642 14654
rect 40574 14642 40626 14654
rect 13906 14590 13918 14642
rect 13970 14590 13982 14642
rect 20066 14590 20078 14642
rect 20130 14590 20142 14642
rect 21970 14590 21982 14642
rect 22034 14590 22046 14642
rect 23650 14590 23662 14642
rect 23714 14590 23726 14642
rect 26226 14590 26238 14642
rect 26290 14590 26302 14642
rect 35298 14590 35310 14642
rect 35362 14590 35374 14642
rect 12014 14578 12066 14590
rect 28590 14578 28642 14590
rect 40574 14578 40626 14590
rect 43486 14642 43538 14654
rect 43486 14578 43538 14590
rect 44942 14642 44994 14654
rect 46050 14590 46062 14642
rect 46114 14590 46126 14642
rect 48178 14590 48190 14642
rect 48242 14590 48254 14642
rect 44942 14578 44994 14590
rect 10446 14530 10498 14542
rect 1810 14478 1822 14530
rect 1874 14478 1886 14530
rect 7186 14478 7198 14530
rect 7250 14478 7262 14530
rect 10446 14466 10498 14478
rect 10670 14530 10722 14542
rect 10670 14466 10722 14478
rect 12238 14530 12290 14542
rect 12238 14466 12290 14478
rect 12910 14530 12962 14542
rect 16606 14530 16658 14542
rect 16258 14478 16270 14530
rect 16322 14478 16334 14530
rect 12910 14466 12962 14478
rect 16606 14466 16658 14478
rect 16942 14530 16994 14542
rect 26014 14530 26066 14542
rect 37886 14530 37938 14542
rect 40014 14530 40066 14542
rect 17266 14478 17278 14530
rect 17330 14478 17342 14530
rect 20626 14478 20638 14530
rect 20690 14478 20702 14530
rect 21858 14478 21870 14530
rect 21922 14478 21934 14530
rect 22194 14478 22206 14530
rect 22258 14478 22270 14530
rect 23538 14478 23550 14530
rect 23602 14478 23614 14530
rect 24322 14478 24334 14530
rect 24386 14478 24398 14530
rect 24994 14478 25006 14530
rect 25058 14478 25070 14530
rect 29474 14478 29486 14530
rect 29538 14478 29550 14530
rect 30146 14478 30158 14530
rect 30210 14478 30222 14530
rect 35634 14478 35646 14530
rect 35698 14478 35710 14530
rect 35970 14478 35982 14530
rect 36034 14478 36046 14530
rect 38994 14478 39006 14530
rect 39058 14478 39070 14530
rect 16942 14466 16994 14478
rect 26014 14466 26066 14478
rect 37886 14466 37938 14478
rect 40014 14466 40066 14478
rect 40686 14530 40738 14542
rect 40686 14466 40738 14478
rect 41022 14530 41074 14542
rect 41022 14466 41074 14478
rect 41470 14530 41522 14542
rect 41470 14466 41522 14478
rect 41694 14530 41746 14542
rect 43026 14478 43038 14530
rect 43090 14478 43102 14530
rect 44258 14478 44270 14530
rect 44322 14478 44334 14530
rect 45266 14478 45278 14530
rect 45330 14478 45342 14530
rect 41694 14466 41746 14478
rect 10334 14418 10386 14430
rect 20414 14418 20466 14430
rect 17938 14366 17950 14418
rect 18002 14366 18014 14418
rect 10334 14354 10386 14366
rect 20414 14354 20466 14366
rect 23998 14418 24050 14430
rect 23998 14354 24050 14366
rect 25678 14418 25730 14430
rect 25678 14354 25730 14366
rect 27246 14418 27298 14430
rect 31166 14418 31218 14430
rect 30370 14366 30382 14418
rect 30434 14366 30446 14418
rect 27246 14354 27298 14366
rect 31166 14354 31218 14366
rect 31278 14418 31330 14430
rect 31278 14354 31330 14366
rect 34302 14418 34354 14430
rect 34302 14354 34354 14366
rect 37214 14418 37266 14430
rect 37214 14354 37266 14366
rect 37550 14418 37602 14430
rect 43474 14366 43486 14418
rect 43538 14366 43550 14418
rect 43810 14366 43822 14418
rect 43874 14366 43886 14418
rect 37550 14354 37602 14366
rect 5070 14306 5122 14318
rect 5070 14242 5122 14254
rect 12686 14306 12738 14318
rect 12686 14242 12738 14254
rect 12798 14306 12850 14318
rect 12798 14242 12850 14254
rect 16718 14306 16770 14318
rect 16718 14242 16770 14254
rect 24558 14306 24610 14318
rect 24558 14242 24610 14254
rect 24670 14306 24722 14318
rect 24670 14242 24722 14254
rect 24782 14306 24834 14318
rect 24782 14242 24834 14254
rect 25790 14306 25842 14318
rect 25790 14242 25842 14254
rect 26350 14306 26402 14318
rect 26350 14242 26402 14254
rect 27022 14306 27074 14318
rect 27022 14242 27074 14254
rect 27358 14306 27410 14318
rect 27358 14242 27410 14254
rect 27470 14306 27522 14318
rect 27470 14242 27522 14254
rect 28030 14306 28082 14318
rect 39790 14306 39842 14318
rect 29698 14254 29710 14306
rect 29762 14254 29774 14306
rect 30706 14254 30718 14306
rect 30770 14254 30782 14306
rect 35858 14254 35870 14306
rect 35922 14254 35934 14306
rect 38434 14254 38446 14306
rect 38498 14254 38510 14306
rect 38770 14254 38782 14306
rect 38834 14254 38846 14306
rect 39442 14254 39454 14306
rect 39506 14254 39518 14306
rect 28030 14242 28082 14254
rect 39790 14242 39842 14254
rect 40462 14306 40514 14318
rect 40462 14242 40514 14254
rect 41246 14306 41298 14318
rect 42366 14306 42418 14318
rect 42018 14254 42030 14306
rect 42082 14254 42094 14306
rect 41246 14242 41298 14254
rect 42366 14242 42418 14254
rect 1344 14138 48608 14172
rect 1344 14086 19838 14138
rect 19890 14086 19942 14138
rect 19994 14086 20046 14138
rect 20098 14086 48608 14138
rect 1344 14052 48608 14086
rect 4622 13970 4674 13982
rect 4622 13906 4674 13918
rect 9662 13970 9714 13982
rect 11454 13970 11506 13982
rect 10770 13918 10782 13970
rect 10834 13918 10846 13970
rect 9662 13906 9714 13918
rect 11454 13906 11506 13918
rect 12798 13970 12850 13982
rect 12798 13906 12850 13918
rect 12910 13970 12962 13982
rect 12910 13906 12962 13918
rect 13470 13970 13522 13982
rect 13470 13906 13522 13918
rect 17502 13970 17554 13982
rect 17502 13906 17554 13918
rect 17950 13970 18002 13982
rect 17950 13906 18002 13918
rect 18734 13970 18786 13982
rect 18734 13906 18786 13918
rect 23550 13970 23602 13982
rect 23550 13906 23602 13918
rect 25342 13970 25394 13982
rect 25342 13906 25394 13918
rect 26126 13970 26178 13982
rect 30942 13970 30994 13982
rect 27906 13918 27918 13970
rect 27970 13918 27982 13970
rect 26126 13906 26178 13918
rect 30942 13906 30994 13918
rect 31054 13970 31106 13982
rect 47070 13970 47122 13982
rect 37874 13918 37886 13970
rect 37938 13918 37950 13970
rect 31054 13906 31106 13918
rect 47070 13906 47122 13918
rect 18286 13858 18338 13870
rect 6514 13806 6526 13858
rect 6578 13806 6590 13858
rect 14466 13806 14478 13858
rect 14530 13806 14542 13858
rect 18286 13794 18338 13806
rect 23326 13858 23378 13870
rect 23326 13794 23378 13806
rect 24446 13858 24498 13870
rect 24446 13794 24498 13806
rect 24670 13858 24722 13870
rect 24670 13794 24722 13806
rect 27022 13858 27074 13870
rect 31166 13858 31218 13870
rect 29250 13806 29262 13858
rect 29314 13806 29326 13858
rect 27022 13794 27074 13806
rect 31166 13794 31218 13806
rect 31278 13858 31330 13870
rect 37202 13806 37214 13858
rect 37266 13806 37278 13858
rect 42242 13806 42254 13858
rect 42306 13806 42318 13858
rect 43698 13806 43710 13858
rect 43762 13806 43774 13858
rect 31278 13794 31330 13806
rect 4846 13746 4898 13758
rect 4846 13682 4898 13694
rect 5070 13746 5122 13758
rect 9998 13746 10050 13758
rect 5842 13694 5854 13746
rect 5906 13694 5918 13746
rect 5070 13682 5122 13694
rect 9998 13682 10050 13694
rect 10222 13746 10274 13758
rect 10222 13682 10274 13694
rect 10446 13746 10498 13758
rect 10446 13682 10498 13694
rect 12238 13746 12290 13758
rect 12238 13682 12290 13694
rect 12686 13746 12738 13758
rect 23774 13746 23826 13758
rect 26910 13746 26962 13758
rect 13794 13694 13806 13746
rect 13858 13694 13870 13746
rect 22530 13694 22542 13746
rect 22594 13694 22606 13746
rect 23986 13694 23998 13746
rect 24050 13694 24062 13746
rect 12686 13682 12738 13694
rect 23774 13682 23826 13694
rect 26910 13682 26962 13694
rect 27470 13746 27522 13758
rect 33406 13746 33458 13758
rect 29586 13694 29598 13746
rect 29650 13694 29662 13746
rect 30706 13694 30718 13746
rect 30770 13694 30782 13746
rect 31714 13694 31726 13746
rect 31778 13694 31790 13746
rect 27470 13682 27522 13694
rect 33406 13682 33458 13694
rect 33966 13746 34018 13758
rect 34862 13746 34914 13758
rect 47742 13746 47794 13758
rect 34402 13694 34414 13746
rect 34466 13694 34478 13746
rect 35410 13694 35422 13746
rect 35474 13694 35486 13746
rect 35858 13694 35870 13746
rect 35922 13694 35934 13746
rect 36866 13694 36878 13746
rect 36930 13694 36942 13746
rect 38546 13694 38558 13746
rect 38610 13694 38622 13746
rect 40002 13694 40014 13746
rect 40066 13694 40078 13746
rect 40786 13694 40798 13746
rect 40850 13694 40862 13746
rect 41570 13694 41582 13746
rect 41634 13694 41646 13746
rect 42130 13694 42142 13746
rect 42194 13694 42206 13746
rect 43362 13694 43374 13746
rect 43426 13694 43438 13746
rect 46274 13694 46286 13746
rect 46338 13694 46350 13746
rect 46722 13694 46734 13746
rect 46786 13694 46798 13746
rect 33966 13682 34018 13694
rect 34862 13682 34914 13694
rect 47742 13682 47794 13694
rect 4734 13634 4786 13646
rect 12014 13634 12066 13646
rect 19182 13634 19234 13646
rect 8642 13582 8654 13634
rect 8706 13582 8718 13634
rect 16594 13582 16606 13634
rect 16658 13582 16670 13634
rect 4734 13570 4786 13582
rect 12014 13570 12066 13582
rect 19182 13570 19234 13582
rect 19630 13634 19682 13646
rect 22990 13634 23042 13646
rect 21410 13582 21422 13634
rect 21474 13582 21486 13634
rect 19630 13570 19682 13582
rect 22990 13570 23042 13582
rect 23662 13634 23714 13646
rect 28478 13634 28530 13646
rect 24434 13582 24446 13634
rect 24498 13582 24510 13634
rect 23662 13570 23714 13582
rect 28478 13570 28530 13582
rect 28926 13634 28978 13646
rect 42702 13634 42754 13646
rect 47966 13634 48018 13646
rect 30034 13582 30046 13634
rect 30098 13582 30110 13634
rect 43922 13582 43934 13634
rect 43986 13582 43998 13634
rect 28926 13570 28978 13582
rect 42702 13570 42754 13582
rect 47966 13570 48018 13582
rect 5294 13522 5346 13534
rect 5294 13458 5346 13470
rect 19406 13522 19458 13534
rect 26686 13522 26738 13534
rect 22754 13470 22766 13522
rect 22818 13519 22830 13522
rect 22978 13519 22990 13522
rect 22818 13473 22990 13519
rect 22818 13470 22830 13473
rect 22978 13470 22990 13473
rect 23042 13470 23054 13522
rect 19406 13458 19458 13470
rect 26686 13458 26738 13470
rect 27246 13522 27298 13534
rect 27246 13458 27298 13470
rect 28254 13522 28306 13534
rect 47518 13522 47570 13534
rect 35858 13470 35870 13522
rect 35922 13470 35934 13522
rect 28254 13458 28306 13470
rect 47518 13458 47570 13470
rect 1344 13354 48608 13388
rect 1344 13302 4478 13354
rect 4530 13302 4582 13354
rect 4634 13302 4686 13354
rect 4738 13302 35198 13354
rect 35250 13302 35302 13354
rect 35354 13302 35406 13354
rect 35458 13302 48608 13354
rect 1344 13268 48608 13302
rect 13694 13186 13746 13198
rect 13694 13122 13746 13134
rect 20078 13186 20130 13198
rect 20078 13122 20130 13134
rect 24782 13186 24834 13198
rect 24782 13122 24834 13134
rect 27022 13186 27074 13198
rect 27022 13122 27074 13134
rect 27246 13186 27298 13198
rect 27246 13122 27298 13134
rect 35422 13186 35474 13198
rect 40686 13186 40738 13198
rect 44158 13186 44210 13198
rect 40338 13134 40350 13186
rect 40402 13134 40414 13186
rect 42690 13134 42702 13186
rect 42754 13134 42766 13186
rect 35422 13122 35474 13134
rect 40686 13122 40738 13134
rect 44158 13122 44210 13134
rect 6638 13074 6690 13086
rect 2482 13022 2494 13074
rect 2546 13022 2558 13074
rect 4610 13022 4622 13074
rect 4674 13022 4686 13074
rect 6638 13010 6690 13022
rect 10446 13074 10498 13086
rect 10446 13010 10498 13022
rect 11454 13074 11506 13086
rect 11454 13010 11506 13022
rect 13022 13074 13074 13086
rect 13022 13010 13074 13022
rect 13470 13074 13522 13086
rect 19630 13074 19682 13086
rect 28702 13074 28754 13086
rect 17714 13022 17726 13074
rect 17778 13022 17790 13074
rect 24322 13022 24334 13074
rect 24386 13022 24398 13074
rect 13470 13010 13522 13022
rect 19630 13010 19682 13022
rect 28702 13010 28754 13022
rect 29486 13074 29538 13086
rect 34190 13074 34242 13086
rect 31602 13022 31614 13074
rect 31666 13022 31678 13074
rect 33730 13022 33742 13074
rect 33794 13022 33806 13074
rect 29486 13010 29538 13022
rect 34190 13010 34242 13022
rect 34526 13074 34578 13086
rect 34526 13010 34578 13022
rect 36430 13074 36482 13086
rect 39666 13022 39678 13074
rect 39730 13022 39742 13074
rect 41458 13022 41470 13074
rect 41522 13022 41534 13074
rect 48178 13022 48190 13074
rect 48242 13022 48254 13074
rect 36430 13010 36482 13022
rect 4958 12962 5010 12974
rect 5854 12962 5906 12974
rect 1810 12910 1822 12962
rect 1874 12910 1886 12962
rect 5618 12910 5630 12962
rect 5682 12910 5694 12962
rect 4958 12898 5010 12910
rect 5854 12898 5906 12910
rect 6078 12962 6130 12974
rect 6078 12898 6130 12910
rect 8878 12962 8930 12974
rect 10110 12962 10162 12974
rect 26798 12962 26850 12974
rect 9202 12910 9214 12962
rect 9266 12910 9278 12962
rect 9986 12910 9998 12962
rect 10050 12910 10062 12962
rect 10322 12910 10334 12962
rect 10386 12910 10398 12962
rect 10994 12910 11006 12962
rect 11058 12910 11070 12962
rect 14802 12910 14814 12962
rect 14866 12910 14878 12962
rect 21298 12910 21310 12962
rect 21362 12910 21374 12962
rect 8878 12898 8930 12910
rect 10110 12898 10162 12910
rect 26798 12898 26850 12910
rect 27470 12962 27522 12974
rect 27470 12898 27522 12910
rect 30046 12962 30098 12974
rect 30046 12898 30098 12910
rect 30606 12962 30658 12974
rect 34750 12962 34802 12974
rect 30818 12910 30830 12962
rect 30882 12910 30894 12962
rect 30606 12898 30658 12910
rect 34750 12898 34802 12910
rect 34974 12962 35026 12974
rect 34974 12898 35026 12910
rect 35646 12962 35698 12974
rect 35646 12898 35698 12910
rect 36094 12962 36146 12974
rect 40910 12962 40962 12974
rect 37650 12910 37662 12962
rect 37714 12910 37726 12962
rect 38882 12910 38894 12962
rect 38946 12910 38958 12962
rect 40002 12910 40014 12962
rect 40066 12910 40078 12962
rect 36094 12898 36146 12910
rect 40910 12898 40962 12910
rect 41246 12962 41298 12974
rect 41246 12898 41298 12910
rect 43598 12962 43650 12974
rect 43598 12898 43650 12910
rect 44382 12962 44434 12974
rect 44382 12898 44434 12910
rect 44830 12962 44882 12974
rect 45266 12910 45278 12962
rect 45330 12910 45342 12962
rect 44830 12898 44882 12910
rect 5070 12850 5122 12862
rect 5070 12786 5122 12798
rect 9438 12850 9490 12862
rect 9438 12786 9490 12798
rect 10558 12850 10610 12862
rect 10558 12786 10610 12798
rect 14366 12850 14418 12862
rect 14366 12786 14418 12798
rect 14478 12850 14530 12862
rect 20078 12850 20130 12862
rect 15586 12798 15598 12850
rect 15650 12798 15662 12850
rect 14478 12786 14530 12798
rect 20078 12786 20130 12798
rect 20190 12850 20242 12862
rect 25006 12850 25058 12862
rect 29598 12850 29650 12862
rect 22082 12798 22094 12850
rect 22146 12798 22158 12850
rect 26450 12798 26462 12850
rect 26514 12798 26526 12850
rect 20190 12786 20242 12798
rect 25006 12786 25058 12798
rect 29598 12786 29650 12798
rect 30270 12850 30322 12862
rect 30270 12786 30322 12798
rect 30382 12850 30434 12862
rect 30382 12786 30434 12798
rect 41582 12850 41634 12862
rect 44942 12850 44994 12862
rect 41682 12798 41694 12850
rect 41746 12798 41758 12850
rect 42578 12798 42590 12850
rect 42642 12798 42654 12850
rect 46050 12798 46062 12850
rect 46114 12798 46126 12850
rect 41582 12786 41634 12798
rect 44942 12786 44994 12798
rect 5742 12738 5794 12750
rect 5742 12674 5794 12686
rect 9550 12738 9602 12750
rect 18174 12738 18226 12750
rect 14018 12686 14030 12738
rect 14082 12686 14094 12738
rect 9550 12674 9602 12686
rect 18174 12674 18226 12686
rect 19182 12738 19234 12750
rect 19182 12674 19234 12686
rect 20638 12738 20690 12750
rect 20638 12674 20690 12686
rect 24894 12738 24946 12750
rect 24894 12674 24946 12686
rect 26126 12738 26178 12750
rect 26126 12674 26178 12686
rect 27918 12738 27970 12750
rect 27918 12674 27970 12686
rect 29374 12738 29426 12750
rect 29374 12674 29426 12686
rect 41470 12738 41522 12750
rect 41470 12674 41522 12686
rect 1344 12570 48608 12604
rect 1344 12518 19838 12570
rect 19890 12518 19942 12570
rect 19994 12518 20046 12570
rect 20098 12518 48608 12570
rect 1344 12484 48608 12518
rect 3166 12402 3218 12414
rect 3166 12338 3218 12350
rect 4286 12402 4338 12414
rect 4286 12338 4338 12350
rect 11118 12402 11170 12414
rect 11118 12338 11170 12350
rect 13134 12402 13186 12414
rect 13134 12338 13186 12350
rect 14478 12402 14530 12414
rect 16718 12402 16770 12414
rect 20078 12402 20130 12414
rect 15586 12350 15598 12402
rect 15650 12350 15662 12402
rect 18610 12350 18622 12402
rect 18674 12350 18686 12402
rect 14478 12338 14530 12350
rect 16718 12338 16770 12350
rect 20078 12338 20130 12350
rect 22766 12402 22818 12414
rect 22766 12338 22818 12350
rect 23998 12402 24050 12414
rect 34638 12402 34690 12414
rect 29362 12350 29374 12402
rect 29426 12350 29438 12402
rect 23998 12338 24050 12350
rect 34638 12338 34690 12350
rect 47966 12402 48018 12414
rect 47966 12338 48018 12350
rect 5406 12290 5458 12302
rect 9662 12290 9714 12302
rect 6850 12238 6862 12290
rect 6914 12238 6926 12290
rect 5406 12226 5458 12238
rect 9662 12226 9714 12238
rect 11230 12290 11282 12302
rect 11230 12226 11282 12238
rect 15150 12290 15202 12302
rect 19518 12290 19570 12302
rect 15362 12238 15374 12290
rect 15426 12238 15438 12290
rect 15150 12226 15202 12238
rect 19518 12226 19570 12238
rect 22990 12290 23042 12302
rect 22990 12226 23042 12238
rect 23438 12290 23490 12302
rect 23438 12226 23490 12238
rect 24222 12290 24274 12302
rect 24222 12226 24274 12238
rect 27246 12290 27298 12302
rect 27246 12226 27298 12238
rect 29262 12290 29314 12302
rect 29262 12226 29314 12238
rect 31838 12290 31890 12302
rect 31838 12226 31890 12238
rect 31950 12290 32002 12302
rect 31950 12226 32002 12238
rect 35982 12290 36034 12302
rect 35982 12226 36034 12238
rect 37102 12290 37154 12302
rect 40350 12290 40402 12302
rect 39890 12238 39902 12290
rect 39954 12238 39966 12290
rect 37102 12226 37154 12238
rect 40350 12226 40402 12238
rect 41918 12290 41970 12302
rect 47406 12290 47458 12302
rect 43250 12238 43262 12290
rect 43314 12238 43326 12290
rect 41918 12226 41970 12238
rect 47406 12226 47458 12238
rect 3390 12178 3442 12190
rect 3390 12114 3442 12126
rect 3614 12178 3666 12190
rect 3614 12114 3666 12126
rect 3838 12178 3890 12190
rect 3838 12114 3890 12126
rect 4510 12178 4562 12190
rect 4510 12114 4562 12126
rect 4734 12178 4786 12190
rect 4734 12114 4786 12126
rect 4958 12178 5010 12190
rect 4958 12114 5010 12126
rect 5294 12178 5346 12190
rect 18958 12178 19010 12190
rect 6178 12126 6190 12178
rect 6242 12126 6254 12178
rect 10322 12126 10334 12178
rect 10386 12126 10398 12178
rect 15922 12126 15934 12178
rect 15986 12126 15998 12178
rect 18162 12126 18174 12178
rect 18226 12126 18238 12178
rect 18722 12126 18734 12178
rect 18786 12126 18798 12178
rect 5294 12114 5346 12126
rect 18958 12114 19010 12126
rect 19294 12178 19346 12190
rect 19294 12114 19346 12126
rect 26686 12178 26738 12190
rect 26686 12114 26738 12126
rect 28702 12178 28754 12190
rect 28702 12114 28754 12126
rect 30942 12178 30994 12190
rect 30942 12114 30994 12126
rect 31166 12178 31218 12190
rect 31166 12114 31218 12126
rect 31502 12178 31554 12190
rect 37326 12178 37378 12190
rect 35522 12126 35534 12178
rect 35586 12126 35598 12178
rect 31502 12114 31554 12126
rect 37326 12114 37378 12126
rect 37774 12178 37826 12190
rect 37774 12114 37826 12126
rect 37998 12178 38050 12190
rect 41470 12178 41522 12190
rect 38770 12126 38782 12178
rect 38834 12126 38846 12178
rect 39330 12126 39342 12178
rect 39394 12126 39406 12178
rect 37998 12114 38050 12126
rect 41470 12114 41522 12126
rect 42814 12178 42866 12190
rect 46846 12178 46898 12190
rect 43138 12126 43150 12178
rect 43202 12126 43214 12178
rect 44034 12126 44046 12178
rect 44098 12126 44110 12178
rect 44482 12126 44494 12178
rect 44546 12126 44558 12178
rect 42814 12114 42866 12126
rect 46846 12114 46898 12126
rect 3278 12066 3330 12078
rect 3278 12002 3330 12014
rect 4398 12066 4450 12078
rect 12126 12066 12178 12078
rect 8978 12014 8990 12066
rect 9042 12014 9054 12066
rect 10658 12014 10670 12066
rect 10722 12014 10734 12066
rect 4398 12002 4450 12014
rect 12126 12002 12178 12014
rect 14030 12066 14082 12078
rect 14030 12002 14082 12014
rect 16606 12066 16658 12078
rect 16606 12002 16658 12014
rect 18510 12066 18562 12078
rect 24110 12066 24162 12078
rect 19506 12014 19518 12066
rect 19570 12014 19582 12066
rect 22642 12014 22654 12066
rect 22706 12014 22718 12066
rect 18510 12002 18562 12014
rect 24110 12002 24162 12014
rect 31054 12066 31106 12078
rect 31054 12002 31106 12014
rect 32622 12066 32674 12078
rect 32622 12002 32674 12014
rect 33294 12066 33346 12078
rect 33294 12002 33346 12014
rect 33742 12066 33794 12078
rect 33742 12002 33794 12014
rect 34302 12066 34354 12078
rect 34302 12002 34354 12014
rect 35086 12066 35138 12078
rect 38446 12066 38498 12078
rect 42254 12066 42306 12078
rect 36642 12014 36654 12066
rect 36706 12014 36718 12066
rect 39442 12014 39454 12066
rect 39506 12014 39518 12066
rect 41010 12014 41022 12066
rect 41074 12014 41086 12066
rect 35086 12002 35138 12014
rect 38446 12002 38498 12014
rect 42254 12002 42306 12014
rect 45950 12066 46002 12078
rect 45950 12002 46002 12014
rect 46286 12066 46338 12078
rect 46286 12002 46338 12014
rect 16494 11954 16546 11966
rect 9426 11902 9438 11954
rect 9490 11951 9502 11954
rect 9762 11951 9774 11954
rect 9490 11905 9774 11951
rect 9490 11902 9502 11905
rect 9762 11902 9774 11905
rect 9826 11902 9838 11954
rect 15698 11902 15710 11954
rect 15762 11902 15774 11954
rect 16494 11890 16546 11902
rect 31950 11954 32002 11966
rect 38222 11954 38274 11966
rect 34178 11902 34190 11954
rect 34242 11951 34254 11954
rect 34962 11951 34974 11954
rect 34242 11905 34974 11951
rect 34242 11902 34254 11905
rect 34962 11902 34974 11905
rect 35026 11902 35038 11954
rect 31950 11890 32002 11902
rect 38222 11890 38274 11902
rect 40238 11954 40290 11966
rect 40238 11890 40290 11902
rect 45838 11954 45890 11966
rect 45838 11890 45890 11902
rect 1344 11786 48608 11820
rect 1344 11734 4478 11786
rect 4530 11734 4582 11786
rect 4634 11734 4686 11786
rect 4738 11734 35198 11786
rect 35250 11734 35302 11786
rect 35354 11734 35406 11786
rect 35458 11734 48608 11786
rect 1344 11700 48608 11734
rect 9998 11618 10050 11630
rect 9998 11554 10050 11566
rect 11006 11618 11058 11630
rect 11006 11554 11058 11566
rect 30046 11618 30098 11630
rect 30046 11554 30098 11566
rect 37102 11618 37154 11630
rect 37102 11554 37154 11566
rect 39902 11618 39954 11630
rect 39902 11554 39954 11566
rect 6414 11506 6466 11518
rect 2482 11454 2494 11506
rect 2546 11454 2558 11506
rect 4610 11454 4622 11506
rect 4674 11454 4686 11506
rect 6414 11442 6466 11454
rect 9326 11506 9378 11518
rect 28142 11506 28194 11518
rect 35086 11506 35138 11518
rect 12786 11454 12798 11506
rect 12850 11454 12862 11506
rect 13794 11454 13806 11506
rect 13858 11454 13870 11506
rect 18610 11454 18622 11506
rect 18674 11454 18686 11506
rect 20738 11454 20750 11506
rect 20802 11454 20814 11506
rect 24098 11454 24110 11506
rect 24162 11454 24174 11506
rect 26226 11454 26238 11506
rect 26290 11454 26302 11506
rect 32498 11454 32510 11506
rect 32562 11454 32574 11506
rect 34626 11454 34638 11506
rect 34690 11454 34702 11506
rect 9326 11442 9378 11454
rect 28142 11442 28194 11454
rect 35086 11442 35138 11454
rect 36206 11506 36258 11518
rect 36206 11442 36258 11454
rect 36990 11506 37042 11518
rect 37986 11454 37998 11506
rect 38050 11454 38062 11506
rect 40674 11454 40686 11506
rect 40738 11454 40750 11506
rect 47730 11454 47742 11506
rect 47794 11454 47806 11506
rect 36990 11442 37042 11454
rect 4958 11394 5010 11406
rect 1810 11342 1822 11394
rect 1874 11342 1886 11394
rect 4958 11330 5010 11342
rect 5630 11394 5682 11406
rect 5630 11330 5682 11342
rect 7758 11394 7810 11406
rect 7758 11330 7810 11342
rect 7982 11394 8034 11406
rect 10222 11394 10274 11406
rect 8754 11342 8766 11394
rect 8818 11342 8830 11394
rect 9762 11342 9774 11394
rect 9826 11342 9838 11394
rect 7982 11330 8034 11342
rect 10222 11330 10274 11342
rect 11230 11394 11282 11406
rect 11230 11330 11282 11342
rect 11678 11394 11730 11406
rect 13470 11394 13522 11406
rect 28478 11394 28530 11406
rect 12226 11342 12238 11394
rect 12290 11342 12302 11394
rect 12898 11342 12910 11394
rect 12962 11342 12974 11394
rect 17938 11342 17950 11394
rect 18002 11342 18014 11394
rect 23314 11342 23326 11394
rect 23378 11342 23390 11394
rect 11678 11330 11730 11342
rect 13470 11330 13522 11342
rect 28478 11330 28530 11342
rect 29038 11394 29090 11406
rect 30606 11394 30658 11406
rect 29362 11342 29374 11394
rect 29426 11342 29438 11394
rect 29038 11330 29090 11342
rect 30606 11330 30658 11342
rect 31054 11394 31106 11406
rect 39678 11394 39730 11406
rect 31826 11342 31838 11394
rect 31890 11342 31902 11394
rect 43586 11342 43598 11394
rect 43650 11342 43662 11394
rect 44818 11342 44830 11394
rect 44882 11342 44894 11394
rect 31054 11330 31106 11342
rect 39678 11330 39730 11342
rect 5070 11282 5122 11294
rect 10334 11282 10386 11294
rect 5954 11230 5966 11282
rect 6018 11230 6030 11282
rect 8978 11230 8990 11282
rect 9042 11230 9054 11282
rect 5070 11218 5122 11230
rect 10334 11218 10386 11230
rect 12686 11282 12738 11294
rect 12686 11218 12738 11230
rect 13694 11282 13746 11294
rect 13694 11218 13746 11230
rect 29598 11282 29650 11294
rect 29598 11218 29650 11230
rect 29710 11282 29762 11294
rect 30046 11282 30098 11294
rect 29710 11218 29762 11230
rect 29934 11226 29986 11238
rect 7870 11170 7922 11182
rect 7870 11106 7922 11118
rect 8206 11170 8258 11182
rect 8206 11106 8258 11118
rect 9438 11170 9490 11182
rect 11790 11170 11842 11182
rect 10658 11118 10670 11170
rect 10722 11118 10734 11170
rect 9438 11106 9490 11118
rect 11790 11106 11842 11118
rect 12014 11170 12066 11182
rect 12014 11106 12066 11118
rect 12462 11170 12514 11182
rect 12462 11106 12514 11118
rect 14366 11170 14418 11182
rect 14366 11106 14418 11118
rect 21422 11170 21474 11182
rect 21422 11106 21474 11118
rect 22990 11170 23042 11182
rect 22990 11106 23042 11118
rect 28590 11170 28642 11182
rect 30046 11218 30098 11230
rect 31278 11282 31330 11294
rect 31278 11218 31330 11230
rect 37550 11282 37602 11294
rect 40238 11282 40290 11294
rect 38994 11230 39006 11282
rect 39058 11230 39070 11282
rect 42802 11230 42814 11282
rect 42866 11230 42878 11282
rect 45602 11230 45614 11282
rect 45666 11230 45678 11282
rect 37550 11218 37602 11230
rect 40238 11218 40290 11230
rect 29934 11162 29986 11174
rect 30830 11170 30882 11182
rect 28590 11106 28642 11118
rect 30830 11106 30882 11118
rect 35870 11170 35922 11182
rect 35870 11106 35922 11118
rect 40014 11170 40066 11182
rect 40014 11106 40066 11118
rect 44270 11170 44322 11182
rect 44270 11106 44322 11118
rect 48190 11170 48242 11182
rect 48190 11106 48242 11118
rect 1344 11002 48608 11036
rect 1344 10950 19838 11002
rect 19890 10950 19942 11002
rect 19994 10950 20046 11002
rect 20098 10950 48608 11002
rect 1344 10916 48608 10950
rect 8206 10834 8258 10846
rect 8206 10770 8258 10782
rect 8430 10834 8482 10846
rect 8430 10770 8482 10782
rect 9662 10834 9714 10846
rect 9662 10770 9714 10782
rect 15038 10834 15090 10846
rect 15038 10770 15090 10782
rect 16382 10834 16434 10846
rect 16382 10770 16434 10782
rect 16942 10834 16994 10846
rect 16942 10770 16994 10782
rect 17502 10834 17554 10846
rect 17502 10770 17554 10782
rect 31726 10834 31778 10846
rect 31726 10770 31778 10782
rect 40238 10834 40290 10846
rect 40238 10770 40290 10782
rect 41134 10834 41186 10846
rect 41134 10770 41186 10782
rect 41358 10834 41410 10846
rect 41358 10770 41410 10782
rect 41470 10834 41522 10846
rect 41470 10770 41522 10782
rect 41582 10834 41634 10846
rect 42702 10834 42754 10846
rect 41906 10782 41918 10834
rect 41970 10782 41982 10834
rect 41582 10770 41634 10782
rect 42702 10770 42754 10782
rect 45054 10834 45106 10846
rect 46174 10834 46226 10846
rect 45826 10782 45838 10834
rect 45890 10782 45902 10834
rect 45054 10770 45106 10782
rect 46174 10770 46226 10782
rect 6302 10722 6354 10734
rect 6302 10658 6354 10670
rect 6638 10722 6690 10734
rect 6638 10658 6690 10670
rect 9886 10722 9938 10734
rect 9886 10658 9938 10670
rect 10110 10722 10162 10734
rect 29038 10722 29090 10734
rect 13794 10670 13806 10722
rect 13858 10670 13870 10722
rect 26002 10670 26014 10722
rect 26066 10670 26078 10722
rect 10110 10658 10162 10670
rect 29038 10658 29090 10670
rect 29374 10722 29426 10734
rect 29374 10658 29426 10670
rect 30606 10722 30658 10734
rect 39678 10722 39730 10734
rect 33842 10670 33854 10722
rect 33906 10670 33918 10722
rect 37090 10670 37102 10722
rect 37154 10670 37166 10722
rect 30606 10658 30658 10670
rect 39678 10658 39730 10670
rect 43374 10722 43426 10734
rect 43374 10658 43426 10670
rect 43934 10722 43986 10734
rect 43934 10658 43986 10670
rect 44270 10722 44322 10734
rect 46846 10722 46898 10734
rect 46498 10670 46510 10722
rect 46562 10670 46574 10722
rect 47170 10670 47182 10722
rect 47234 10670 47246 10722
rect 44270 10658 44322 10670
rect 46846 10658 46898 10670
rect 4958 10610 5010 10622
rect 4958 10546 5010 10558
rect 5182 10610 5234 10622
rect 5182 10546 5234 10558
rect 8878 10610 8930 10622
rect 8878 10546 8930 10558
rect 9438 10610 9490 10622
rect 9438 10546 9490 10558
rect 10558 10610 10610 10622
rect 10558 10546 10610 10558
rect 10894 10610 10946 10622
rect 28478 10610 28530 10622
rect 14578 10558 14590 10610
rect 14642 10558 14654 10610
rect 20514 10558 20526 10610
rect 20578 10558 20590 10610
rect 25218 10558 25230 10610
rect 25282 10558 25294 10610
rect 10894 10546 10946 10558
rect 28478 10546 28530 10558
rect 28702 10610 28754 10622
rect 30830 10610 30882 10622
rect 29586 10558 29598 10610
rect 29650 10558 29662 10610
rect 28702 10546 28754 10558
rect 30830 10546 30882 10558
rect 31166 10610 31218 10622
rect 31166 10546 31218 10558
rect 31502 10610 31554 10622
rect 43486 10610 43538 10622
rect 33170 10558 33182 10610
rect 33234 10558 33246 10610
rect 36306 10558 36318 10610
rect 36370 10558 36382 10610
rect 42130 10558 42142 10610
rect 42194 10558 42206 10610
rect 31502 10546 31554 10558
rect 43486 10546 43538 10558
rect 43710 10610 43762 10622
rect 43710 10546 43762 10558
rect 44606 10610 44658 10622
rect 44818 10558 44830 10610
rect 44882 10558 44894 10610
rect 47394 10558 47406 10610
rect 47458 10558 47470 10610
rect 44606 10546 44658 10558
rect 7534 10498 7586 10510
rect 7534 10434 7586 10446
rect 8318 10498 8370 10510
rect 8318 10434 8370 10446
rect 10782 10498 10834 10510
rect 15486 10498 15538 10510
rect 24670 10498 24722 10510
rect 28590 10498 28642 10510
rect 11666 10446 11678 10498
rect 11730 10446 11742 10498
rect 15922 10446 15934 10498
rect 15986 10446 15998 10498
rect 21186 10446 21198 10498
rect 21250 10446 21262 10498
rect 23314 10446 23326 10498
rect 23378 10446 23390 10498
rect 28130 10446 28142 10498
rect 28194 10446 28206 10498
rect 10782 10434 10834 10446
rect 15486 10434 15538 10446
rect 24670 10434 24722 10446
rect 28590 10434 28642 10446
rect 30158 10498 30210 10510
rect 30158 10434 30210 10446
rect 31054 10498 31106 10510
rect 31054 10434 31106 10446
rect 32510 10498 32562 10510
rect 40350 10498 40402 10510
rect 35970 10446 35982 10498
rect 36034 10446 36046 10498
rect 39218 10446 39230 10498
rect 39282 10446 39294 10498
rect 32510 10434 32562 10446
rect 40350 10434 40402 10446
rect 45390 10498 45442 10510
rect 45390 10434 45442 10446
rect 47966 10498 48018 10510
rect 47966 10434 48018 10446
rect 4846 10386 4898 10398
rect 4846 10322 4898 10334
rect 5294 10386 5346 10398
rect 5294 10322 5346 10334
rect 10446 10386 10498 10398
rect 10446 10322 10498 10334
rect 31838 10386 31890 10398
rect 31838 10322 31890 10334
rect 39566 10386 39618 10398
rect 45502 10386 45554 10398
rect 44818 10334 44830 10386
rect 44882 10334 44894 10386
rect 39566 10322 39618 10334
rect 45502 10322 45554 10334
rect 47854 10386 47906 10398
rect 47854 10322 47906 10334
rect 1344 10218 48608 10252
rect 1344 10166 4478 10218
rect 4530 10166 4582 10218
rect 4634 10166 4686 10218
rect 4738 10166 35198 10218
rect 35250 10166 35302 10218
rect 35354 10166 35406 10218
rect 35458 10166 48608 10218
rect 1344 10132 48608 10166
rect 10334 10050 10386 10062
rect 10334 9986 10386 9998
rect 10446 10050 10498 10062
rect 10446 9986 10498 9998
rect 30382 10050 30434 10062
rect 30382 9986 30434 9998
rect 35534 10050 35586 10062
rect 35534 9986 35586 9998
rect 9214 9938 9266 9950
rect 34078 9938 34130 9950
rect 1698 9886 1710 9938
rect 1762 9886 1774 9938
rect 3826 9886 3838 9938
rect 3890 9886 3902 9938
rect 16482 9886 16494 9938
rect 16546 9886 16558 9938
rect 19730 9886 19742 9938
rect 19794 9886 19806 9938
rect 23202 9886 23214 9938
rect 23266 9886 23278 9938
rect 25330 9886 25342 9938
rect 25394 9886 25406 9938
rect 25666 9886 25678 9938
rect 25730 9886 25742 9938
rect 27794 9886 27806 9938
rect 27858 9886 27870 9938
rect 30034 9886 30046 9938
rect 30098 9886 30110 9938
rect 31490 9886 31502 9938
rect 31554 9886 31566 9938
rect 33618 9886 33630 9938
rect 33682 9886 33694 9938
rect 9214 9874 9266 9886
rect 34078 9874 34130 9886
rect 37438 9938 37490 9950
rect 37438 9874 37490 9886
rect 37886 9938 37938 9950
rect 41010 9886 41022 9938
rect 41074 9886 41086 9938
rect 44258 9886 44270 9938
rect 44322 9886 44334 9938
rect 37886 9874 37938 9886
rect 5070 9826 5122 9838
rect 4610 9774 4622 9826
rect 4674 9774 4686 9826
rect 5070 9762 5122 9774
rect 6190 9826 6242 9838
rect 6190 9762 6242 9774
rect 6414 9826 6466 9838
rect 6974 9826 7026 9838
rect 6626 9774 6638 9826
rect 6690 9774 6702 9826
rect 6414 9762 6466 9774
rect 6974 9762 7026 9774
rect 7870 9826 7922 9838
rect 7870 9762 7922 9774
rect 7982 9826 8034 9838
rect 7982 9762 8034 9774
rect 9998 9826 10050 9838
rect 9998 9762 10050 9774
rect 10670 9826 10722 9838
rect 10670 9762 10722 9774
rect 10894 9826 10946 9838
rect 29038 9826 29090 9838
rect 12898 9774 12910 9826
rect 12962 9774 12974 9826
rect 13570 9774 13582 9826
rect 13634 9774 13646 9826
rect 16930 9774 16942 9826
rect 16994 9774 17006 9826
rect 22418 9774 22430 9826
rect 22482 9774 22494 9826
rect 28578 9774 28590 9826
rect 28642 9774 28654 9826
rect 10894 9762 10946 9774
rect 29038 9762 29090 9774
rect 29374 9826 29426 9838
rect 30706 9774 30718 9826
rect 30770 9774 30782 9826
rect 36306 9774 36318 9826
rect 36370 9774 36382 9826
rect 38098 9774 38110 9826
rect 38162 9774 38174 9826
rect 41346 9774 41358 9826
rect 41410 9774 41422 9826
rect 47842 9774 47854 9826
rect 47906 9774 47918 9826
rect 29374 9762 29426 9774
rect 7310 9714 7362 9726
rect 7310 9650 7362 9662
rect 7534 9714 7586 9726
rect 7534 9650 7586 9662
rect 11006 9714 11058 9726
rect 11006 9650 11058 9662
rect 11342 9714 11394 9726
rect 11342 9650 11394 9662
rect 11678 9714 11730 9726
rect 11678 9650 11730 9662
rect 12574 9714 12626 9726
rect 30158 9714 30210 9726
rect 44942 9714 44994 9726
rect 14354 9662 14366 9714
rect 14418 9662 14430 9714
rect 17602 9662 17614 9714
rect 17666 9662 17678 9714
rect 36082 9662 36094 9714
rect 36146 9662 36158 9714
rect 38882 9662 38894 9714
rect 38946 9662 38958 9714
rect 42130 9662 42142 9714
rect 42194 9662 42206 9714
rect 12574 9650 12626 9662
rect 30158 9650 30210 9662
rect 44942 9650 44994 9662
rect 6526 9602 6578 9614
rect 6526 9538 6578 9550
rect 7086 9602 7138 9614
rect 7086 9538 7138 9550
rect 7646 9602 7698 9614
rect 7646 9538 7698 9550
rect 12238 9602 12290 9614
rect 12238 9538 12290 9550
rect 12686 9602 12738 9614
rect 12686 9538 12738 9550
rect 20190 9602 20242 9614
rect 20190 9538 20242 9550
rect 22094 9602 22146 9614
rect 22094 9538 22146 9550
rect 29262 9602 29314 9614
rect 29262 9538 29314 9550
rect 34862 9602 34914 9614
rect 34862 9538 34914 9550
rect 35198 9602 35250 9614
rect 35198 9538 35250 9550
rect 45054 9602 45106 9614
rect 45054 9538 45106 9550
rect 45278 9602 45330 9614
rect 45278 9538 45330 9550
rect 47182 9602 47234 9614
rect 47182 9538 47234 9550
rect 1344 9434 48608 9468
rect 1344 9382 19838 9434
rect 19890 9382 19942 9434
rect 19994 9382 20046 9434
rect 20098 9382 48608 9434
rect 1344 9348 48608 9382
rect 3838 9266 3890 9278
rect 3838 9202 3890 9214
rect 4958 9266 5010 9278
rect 4958 9202 5010 9214
rect 15038 9266 15090 9278
rect 15038 9202 15090 9214
rect 17502 9266 17554 9278
rect 17502 9202 17554 9214
rect 17950 9266 18002 9278
rect 17950 9202 18002 9214
rect 18846 9266 18898 9278
rect 18846 9202 18898 9214
rect 29150 9266 29202 9278
rect 29150 9202 29202 9214
rect 33294 9266 33346 9278
rect 33294 9202 33346 9214
rect 34302 9266 34354 9278
rect 34302 9202 34354 9214
rect 34638 9266 34690 9278
rect 34638 9202 34690 9214
rect 38222 9266 38274 9278
rect 38222 9202 38274 9214
rect 38558 9266 38610 9278
rect 38558 9202 38610 9214
rect 38782 9266 38834 9278
rect 38782 9202 38834 9214
rect 41582 9266 41634 9278
rect 41582 9202 41634 9214
rect 41918 9266 41970 9278
rect 41918 9202 41970 9214
rect 4622 9154 4674 9166
rect 4622 9090 4674 9102
rect 5742 9154 5794 9166
rect 10670 9154 10722 9166
rect 6850 9102 6862 9154
rect 6914 9102 6926 9154
rect 5742 9090 5794 9102
rect 10670 9090 10722 9102
rect 18398 9154 18450 9166
rect 28030 9154 28082 9166
rect 27570 9102 27582 9154
rect 27634 9102 27646 9154
rect 18398 9090 18450 9102
rect 28030 9090 28082 9102
rect 28142 9154 28194 9166
rect 28142 9090 28194 9102
rect 33518 9154 33570 9166
rect 33518 9090 33570 9102
rect 37326 9154 37378 9166
rect 37326 9090 37378 9102
rect 42478 9154 42530 9166
rect 42478 9090 42530 9102
rect 43822 9154 43874 9166
rect 43822 9090 43874 9102
rect 44270 9154 44322 9166
rect 44270 9090 44322 9102
rect 4174 9042 4226 9054
rect 5294 9042 5346 9054
rect 14926 9042 14978 9054
rect 16382 9042 16434 9054
rect 35198 9042 35250 9054
rect 3938 8990 3950 9042
rect 4002 8990 4014 9042
rect 4386 8990 4398 9042
rect 4450 8990 4462 9042
rect 4946 8990 4958 9042
rect 5010 8990 5022 9042
rect 5506 8990 5518 9042
rect 5570 8990 5582 9042
rect 6178 8990 6190 9042
rect 6242 8990 6254 9042
rect 10434 8990 10446 9042
rect 10498 8990 10510 9042
rect 14578 8990 14590 9042
rect 14642 8990 14654 9042
rect 15138 8990 15150 9042
rect 15202 8990 15214 9042
rect 15698 8990 15710 9042
rect 15762 8990 15774 9042
rect 16594 8990 16606 9042
rect 16658 8990 16670 9042
rect 19618 8990 19630 9042
rect 19682 8990 19694 9042
rect 20178 8990 20190 9042
rect 20242 8990 20254 9042
rect 4174 8978 4226 8990
rect 5294 8978 5346 8990
rect 14926 8978 14978 8990
rect 16382 8978 16434 8990
rect 35198 8978 35250 8990
rect 36430 9042 36482 9054
rect 36430 8978 36482 8990
rect 36878 9042 36930 9054
rect 36878 8978 36930 8990
rect 39118 9042 39170 9054
rect 39118 8978 39170 8990
rect 41470 9042 41522 9054
rect 41470 8978 41522 8990
rect 41694 9042 41746 9054
rect 41694 8978 41746 8990
rect 44158 9042 44210 9054
rect 44158 8978 44210 8990
rect 44494 9042 44546 9054
rect 44494 8978 44546 8990
rect 44718 9042 44770 9054
rect 44718 8978 44770 8990
rect 44942 9042 44994 9054
rect 45826 8990 45838 9042
rect 45890 8990 45902 9042
rect 44942 8978 44994 8990
rect 9998 8930 10050 8942
rect 8978 8878 8990 8930
rect 9042 8878 9054 8930
rect 9998 8866 10050 8878
rect 11454 8930 11506 8942
rect 22990 8930 23042 8942
rect 28702 8930 28754 8942
rect 11666 8878 11678 8930
rect 11730 8878 11742 8930
rect 13794 8878 13806 8930
rect 13858 8878 13870 8930
rect 22530 8878 22542 8930
rect 22594 8878 22606 8930
rect 26226 8878 26238 8930
rect 26290 8878 26302 8930
rect 11454 8866 11506 8878
rect 22990 8866 23042 8878
rect 28702 8866 28754 8878
rect 29934 8930 29986 8942
rect 29934 8866 29986 8878
rect 30382 8930 30434 8942
rect 30382 8866 30434 8878
rect 30830 8930 30882 8942
rect 30830 8866 30882 8878
rect 31278 8930 31330 8942
rect 31278 8866 31330 8878
rect 31726 8930 31778 8942
rect 31726 8866 31778 8878
rect 32510 8930 32562 8942
rect 32510 8866 32562 8878
rect 35758 8930 35810 8942
rect 35758 8866 35810 8878
rect 36206 8930 36258 8942
rect 36206 8866 36258 8878
rect 37886 8930 37938 8942
rect 37886 8866 37938 8878
rect 38894 8930 38946 8942
rect 38894 8866 38946 8878
rect 39454 8930 39506 8942
rect 39454 8866 39506 8878
rect 40014 8930 40066 8942
rect 40014 8866 40066 8878
rect 40350 8930 40402 8942
rect 40350 8866 40402 8878
rect 41134 8930 41186 8942
rect 41134 8866 41186 8878
rect 42814 8930 42866 8942
rect 42814 8866 42866 8878
rect 43262 8930 43314 8942
rect 43262 8866 43314 8878
rect 16270 8818 16322 8830
rect 15474 8766 15486 8818
rect 15538 8766 15550 8818
rect 16270 8754 16322 8766
rect 28142 8818 28194 8830
rect 33182 8818 33234 8830
rect 30370 8766 30382 8818
rect 30434 8815 30446 8818
rect 30818 8815 30830 8818
rect 30434 8769 30830 8815
rect 30434 8766 30446 8769
rect 30818 8766 30830 8769
rect 30882 8766 30894 8818
rect 28142 8754 28194 8766
rect 33182 8754 33234 8766
rect 36654 8818 36706 8830
rect 42926 8818 42978 8830
rect 39442 8766 39454 8818
rect 39506 8815 39518 8818
rect 40338 8815 40350 8818
rect 39506 8769 40350 8815
rect 39506 8766 39518 8769
rect 40338 8766 40350 8769
rect 40402 8766 40414 8818
rect 36654 8754 36706 8766
rect 42926 8754 42978 8766
rect 43374 8818 43426 8830
rect 43374 8754 43426 8766
rect 43710 8818 43762 8830
rect 47966 8818 48018 8830
rect 45266 8766 45278 8818
rect 45330 8766 45342 8818
rect 43710 8754 43762 8766
rect 47966 8754 48018 8766
rect 1344 8650 48608 8684
rect 1344 8598 4478 8650
rect 4530 8598 4582 8650
rect 4634 8598 4686 8650
rect 4738 8598 35198 8650
rect 35250 8598 35302 8650
rect 35354 8598 35406 8650
rect 35458 8598 48608 8650
rect 1344 8564 48608 8598
rect 10770 8430 10782 8482
rect 10834 8430 10846 8482
rect 13682 8430 13694 8482
rect 13746 8430 13758 8482
rect 4958 8370 5010 8382
rect 2482 8318 2494 8370
rect 2546 8318 2558 8370
rect 4610 8318 4622 8370
rect 4674 8318 4686 8370
rect 4958 8306 5010 8318
rect 5742 8370 5794 8382
rect 5742 8306 5794 8318
rect 11454 8370 11506 8382
rect 11454 8306 11506 8318
rect 13022 8370 13074 8382
rect 13022 8306 13074 8318
rect 15150 8370 15202 8382
rect 15150 8306 15202 8318
rect 17950 8370 18002 8382
rect 17950 8306 18002 8318
rect 19966 8370 20018 8382
rect 22430 8370 22482 8382
rect 28702 8370 28754 8382
rect 20290 8318 20302 8370
rect 20354 8318 20366 8370
rect 25666 8318 25678 8370
rect 25730 8318 25742 8370
rect 19966 8306 20018 8318
rect 22430 8306 22482 8318
rect 28702 8306 28754 8318
rect 33966 8370 34018 8382
rect 33966 8306 34018 8318
rect 34414 8370 34466 8382
rect 38334 8370 38386 8382
rect 35298 8318 35310 8370
rect 35362 8318 35374 8370
rect 34414 8306 34466 8318
rect 38334 8306 38386 8318
rect 44158 8370 44210 8382
rect 44158 8306 44210 8318
rect 47966 8370 48018 8382
rect 47966 8306 48018 8318
rect 9438 8258 9490 8270
rect 19742 8258 19794 8270
rect 1810 8206 1822 8258
rect 1874 8206 1886 8258
rect 10322 8206 10334 8258
rect 10386 8206 10398 8258
rect 10770 8206 10782 8258
rect 10834 8206 10846 8258
rect 13458 8206 13470 8258
rect 13522 8206 13534 8258
rect 16818 8206 16830 8258
rect 16882 8206 16894 8258
rect 19394 8206 19406 8258
rect 19458 8206 19470 8258
rect 9438 8194 9490 8206
rect 19742 8194 19794 8206
rect 21982 8258 22034 8270
rect 35646 8258 35698 8270
rect 36542 8258 36594 8270
rect 40014 8258 40066 8270
rect 22754 8206 22766 8258
rect 22818 8206 22830 8258
rect 30930 8206 30942 8258
rect 30994 8206 31006 8258
rect 31602 8206 31614 8258
rect 31666 8206 31678 8258
rect 33170 8206 33182 8258
rect 33234 8206 33246 8258
rect 35858 8206 35870 8258
rect 35922 8206 35934 8258
rect 38770 8206 38782 8258
rect 38834 8206 38846 8258
rect 40450 8206 40462 8258
rect 40514 8206 40526 8258
rect 41346 8206 41358 8258
rect 41410 8206 41422 8258
rect 45042 8206 45054 8258
rect 45106 8206 45118 8258
rect 45938 8206 45950 8258
rect 46002 8206 46014 8258
rect 21982 8194 22034 8206
rect 35646 8194 35698 8206
rect 36542 8194 36594 8206
rect 40014 8194 40066 8206
rect 12238 8146 12290 8158
rect 14254 8146 14306 8158
rect 14018 8094 14030 8146
rect 14082 8094 14094 8146
rect 12238 8082 12290 8094
rect 14254 8082 14306 8094
rect 15598 8146 15650 8158
rect 21646 8146 21698 8158
rect 27134 8146 27186 8158
rect 19282 8094 19294 8146
rect 19346 8094 19358 8146
rect 23538 8094 23550 8146
rect 23602 8094 23614 8146
rect 15598 8082 15650 8094
rect 21646 8082 21698 8094
rect 27134 8082 27186 8094
rect 27582 8146 27634 8158
rect 27582 8082 27634 8094
rect 27806 8146 27858 8158
rect 27806 8082 27858 8094
rect 29822 8146 29874 8158
rect 39342 8146 39394 8158
rect 37314 8094 37326 8146
rect 37378 8094 37390 8146
rect 29822 8082 29874 8094
rect 39342 8082 39394 8094
rect 39678 8146 39730 8158
rect 39678 8082 39730 8094
rect 40686 8146 40738 8158
rect 42366 8146 42418 8158
rect 41906 8094 41918 8146
rect 41970 8094 41982 8146
rect 40686 8082 40738 8094
rect 42366 8082 42418 8094
rect 42478 8146 42530 8158
rect 42478 8082 42530 8094
rect 42926 8146 42978 8158
rect 43934 8146 43986 8158
rect 43810 8094 43822 8146
rect 43874 8094 43886 8146
rect 45266 8094 45278 8146
rect 45330 8094 45342 8146
rect 42926 8082 42978 8094
rect 43934 8082 43986 8094
rect 5070 8034 5122 8046
rect 5070 7970 5122 7982
rect 8878 8034 8930 8046
rect 8878 7970 8930 7982
rect 9774 8034 9826 8046
rect 9774 7970 9826 7982
rect 12014 8034 12066 8046
rect 12014 7970 12066 7982
rect 12350 8034 12402 8046
rect 14702 8034 14754 8046
rect 13906 7982 13918 8034
rect 13970 7982 13982 8034
rect 12350 7970 12402 7982
rect 14702 7970 14754 7982
rect 15486 8034 15538 8046
rect 15486 7970 15538 7982
rect 16270 8034 16322 8046
rect 17502 8034 17554 8046
rect 17042 7982 17054 8034
rect 17106 7982 17118 8034
rect 16270 7970 16322 7982
rect 17502 7970 17554 7982
rect 18398 8034 18450 8046
rect 20862 8034 20914 8046
rect 18834 7982 18846 8034
rect 18898 7982 18910 8034
rect 18398 7970 18450 7982
rect 20862 7970 20914 7982
rect 27694 8034 27746 8046
rect 27694 7970 27746 7982
rect 29486 8034 29538 8046
rect 29486 7970 29538 7982
rect 29934 8034 29986 8046
rect 29934 7970 29986 7982
rect 30046 8034 30098 8046
rect 30046 7970 30098 7982
rect 30718 8034 30770 8046
rect 30718 7970 30770 7982
rect 31390 8034 31442 8046
rect 31390 7970 31442 7982
rect 32174 8034 32226 8046
rect 32174 7970 32226 7982
rect 32622 8034 32674 8046
rect 32622 7970 32674 7982
rect 33406 8034 33458 8046
rect 33406 7970 33458 7982
rect 34974 8034 35026 8046
rect 34974 7970 35026 7982
rect 36990 8034 37042 8046
rect 36990 7970 37042 7982
rect 37774 8034 37826 8046
rect 40126 8034 40178 8046
rect 42142 8034 42194 8046
rect 38994 7982 39006 8034
rect 39058 7982 39070 8034
rect 40786 7982 40798 8034
rect 40850 7982 40862 8034
rect 37774 7970 37826 7982
rect 40126 7970 40178 7982
rect 42142 7970 42194 7982
rect 42814 8034 42866 8046
rect 42814 7970 42866 7982
rect 44046 8034 44098 8046
rect 44046 7970 44098 7982
rect 44270 8034 44322 8046
rect 44270 7970 44322 7982
rect 1344 7866 48608 7900
rect 1344 7814 19838 7866
rect 19890 7814 19942 7866
rect 19994 7814 20046 7866
rect 20098 7814 48608 7866
rect 1344 7780 48608 7814
rect 6638 7698 6690 7710
rect 6638 7634 6690 7646
rect 7086 7698 7138 7710
rect 20078 7698 20130 7710
rect 19394 7646 19406 7698
rect 19458 7646 19470 7698
rect 7086 7634 7138 7646
rect 20078 7634 20130 7646
rect 26014 7698 26066 7710
rect 26014 7634 26066 7646
rect 27918 7698 27970 7710
rect 27918 7634 27970 7646
rect 32174 7698 32226 7710
rect 32174 7634 32226 7646
rect 37214 7698 37266 7710
rect 37214 7634 37266 7646
rect 38222 7698 38274 7710
rect 45266 7646 45278 7698
rect 45330 7646 45342 7698
rect 38222 7634 38274 7646
rect 13246 7586 13298 7598
rect 4050 7534 4062 7586
rect 4114 7534 4126 7586
rect 13246 7522 13298 7534
rect 19070 7586 19122 7598
rect 19070 7522 19122 7534
rect 19742 7586 19794 7598
rect 27134 7586 27186 7598
rect 40910 7586 40962 7598
rect 21410 7534 21422 7586
rect 21474 7534 21486 7586
rect 21970 7534 21982 7586
rect 22034 7534 22046 7586
rect 26338 7534 26350 7586
rect 26402 7534 26414 7586
rect 36754 7534 36766 7586
rect 36818 7534 36830 7586
rect 39890 7534 39902 7586
rect 39954 7534 39966 7586
rect 42130 7534 42142 7586
rect 42194 7534 42206 7586
rect 19742 7522 19794 7534
rect 27134 7522 27186 7534
rect 40910 7522 40962 7534
rect 6526 7474 6578 7486
rect 13134 7474 13186 7486
rect 17950 7474 18002 7486
rect 3266 7422 3278 7474
rect 3330 7422 3342 7474
rect 9874 7422 9886 7474
rect 9938 7422 9950 7474
rect 13682 7422 13694 7474
rect 13746 7422 13758 7474
rect 6526 7410 6578 7422
rect 13134 7410 13186 7422
rect 17950 7410 18002 7422
rect 21198 7474 21250 7486
rect 36430 7474 36482 7486
rect 44718 7474 44770 7486
rect 26562 7422 26574 7474
rect 26626 7422 26638 7474
rect 27458 7422 27470 7474
rect 27522 7422 27534 7474
rect 28354 7422 28366 7474
rect 28418 7422 28430 7474
rect 28914 7422 28926 7474
rect 28978 7422 28990 7474
rect 35410 7422 35422 7474
rect 35474 7422 35486 7474
rect 35970 7422 35982 7474
rect 36034 7422 36046 7474
rect 38434 7422 38446 7474
rect 38498 7422 38510 7474
rect 39554 7422 39566 7474
rect 39618 7422 39630 7474
rect 41458 7422 41470 7474
rect 41522 7422 41534 7474
rect 21198 7410 21250 7422
rect 36430 7410 36482 7422
rect 44718 7410 44770 7422
rect 44942 7474 44994 7486
rect 45714 7422 45726 7474
rect 45778 7422 45790 7474
rect 44942 7410 44994 7422
rect 7534 7362 7586 7374
rect 6178 7310 6190 7362
rect 6242 7310 6254 7362
rect 7534 7298 7586 7310
rect 8654 7362 8706 7374
rect 8654 7298 8706 7310
rect 9102 7362 9154 7374
rect 18398 7362 18450 7374
rect 10658 7310 10670 7362
rect 10722 7310 10734 7362
rect 12786 7310 12798 7362
rect 12850 7310 12862 7362
rect 14466 7310 14478 7362
rect 14530 7310 14542 7362
rect 16594 7310 16606 7362
rect 16658 7310 16670 7362
rect 17490 7310 17502 7362
rect 17554 7310 17566 7362
rect 9102 7298 9154 7310
rect 18398 7298 18450 7310
rect 18958 7362 19010 7374
rect 18958 7298 19010 7310
rect 20190 7362 20242 7374
rect 20190 7298 20242 7310
rect 22766 7362 22818 7374
rect 22766 7298 22818 7310
rect 23550 7362 23602 7374
rect 23550 7298 23602 7310
rect 24446 7362 24498 7374
rect 31614 7362 31666 7374
rect 37662 7362 37714 7374
rect 40350 7362 40402 7374
rect 47966 7362 48018 7374
rect 31266 7310 31278 7362
rect 31330 7310 31342 7362
rect 33058 7310 33070 7362
rect 33122 7310 33134 7362
rect 39330 7310 39342 7362
rect 39394 7310 39406 7362
rect 44258 7310 44270 7362
rect 44322 7310 44334 7362
rect 24446 7298 24498 7310
rect 31614 7298 31666 7310
rect 37662 7298 37714 7310
rect 40350 7298 40402 7310
rect 47966 7298 48018 7310
rect 7422 7250 7474 7262
rect 7422 7186 7474 7198
rect 13246 7250 13298 7262
rect 13246 7186 13298 7198
rect 20862 7250 20914 7262
rect 20862 7186 20914 7198
rect 22654 7250 22706 7262
rect 22654 7186 22706 7198
rect 27470 7250 27522 7262
rect 27470 7186 27522 7198
rect 31726 7250 31778 7262
rect 31726 7186 31778 7198
rect 40238 7250 40290 7262
rect 40238 7186 40290 7198
rect 41022 7250 41074 7262
rect 41022 7186 41074 7198
rect 1344 7082 48608 7116
rect 1344 7030 4478 7082
rect 4530 7030 4582 7082
rect 4634 7030 4686 7082
rect 4738 7030 35198 7082
rect 35250 7030 35302 7082
rect 35354 7030 35406 7082
rect 35458 7030 48608 7082
rect 1344 6996 48608 7030
rect 11566 6914 11618 6926
rect 11566 6850 11618 6862
rect 31054 6914 31106 6926
rect 31054 6850 31106 6862
rect 35310 6914 35362 6926
rect 35310 6850 35362 6862
rect 11678 6802 11730 6814
rect 32174 6802 32226 6814
rect 7186 6750 7198 6802
rect 7250 6750 7262 6802
rect 9314 6750 9326 6802
rect 9378 6750 9390 6802
rect 12114 6750 12126 6802
rect 12178 6750 12190 6802
rect 19842 6750 19854 6802
rect 19906 6750 19918 6802
rect 23202 6750 23214 6802
rect 23266 6750 23278 6802
rect 27794 6750 27806 6802
rect 27858 6750 27870 6802
rect 30706 6750 30718 6802
rect 30770 6750 30782 6802
rect 11678 6738 11730 6750
rect 32174 6738 32226 6750
rect 32958 6802 33010 6814
rect 38770 6750 38782 6802
rect 38834 6750 38846 6802
rect 39330 6750 39342 6802
rect 39394 6750 39406 6802
rect 43474 6750 43486 6802
rect 43538 6750 43550 6802
rect 48178 6750 48190 6802
rect 48242 6750 48254 6802
rect 32958 6738 33010 6750
rect 10222 6690 10274 6702
rect 6514 6638 6526 6690
rect 6578 6638 6590 6690
rect 9762 6638 9774 6690
rect 9826 6638 9838 6690
rect 10222 6626 10274 6638
rect 10670 6690 10722 6702
rect 10670 6626 10722 6638
rect 12910 6690 12962 6702
rect 21982 6690 22034 6702
rect 29486 6690 29538 6702
rect 13682 6638 13694 6690
rect 13746 6638 13758 6690
rect 17042 6638 17054 6690
rect 17106 6638 17118 6690
rect 23650 6638 23662 6690
rect 23714 6638 23726 6690
rect 24770 6638 24782 6690
rect 24834 6638 24846 6690
rect 25442 6638 25454 6690
rect 25506 6638 25518 6690
rect 12910 6626 12962 6638
rect 21982 6626 22034 6638
rect 29486 6626 29538 6638
rect 29710 6690 29762 6702
rect 29710 6626 29762 6638
rect 30382 6690 30434 6702
rect 30382 6626 30434 6638
rect 32286 6690 32338 6702
rect 34302 6690 34354 6702
rect 33282 6638 33294 6690
rect 33346 6638 33358 6690
rect 34066 6638 34078 6690
rect 34130 6638 34142 6690
rect 32286 6626 32338 6638
rect 34302 6626 34354 6638
rect 34638 6690 34690 6702
rect 34638 6626 34690 6638
rect 37886 6690 37938 6702
rect 37886 6626 37938 6638
rect 38222 6690 38274 6702
rect 38434 6638 38446 6690
rect 38498 6638 38510 6690
rect 39106 6638 39118 6690
rect 39170 6638 39182 6690
rect 40562 6638 40574 6690
rect 40626 6638 40638 6690
rect 45378 6638 45390 6690
rect 45442 6638 45454 6690
rect 46050 6638 46062 6690
rect 46114 6638 46126 6690
rect 38222 6626 38274 6638
rect 11006 6578 11058 6590
rect 12574 6578 12626 6590
rect 23102 6578 23154 6590
rect 12450 6526 12462 6578
rect 12514 6526 12526 6578
rect 17714 6526 17726 6578
rect 17778 6526 17790 6578
rect 11006 6514 11058 6526
rect 12574 6514 12626 6526
rect 23102 6514 23154 6526
rect 23214 6578 23266 6590
rect 23214 6514 23266 6526
rect 23998 6578 24050 6590
rect 23998 6514 24050 6526
rect 24334 6578 24386 6590
rect 35198 6578 35250 6590
rect 33058 6526 33070 6578
rect 33122 6526 33134 6578
rect 24334 6514 24386 6526
rect 35198 6514 35250 6526
rect 36318 6578 36370 6590
rect 36318 6514 36370 6526
rect 37326 6578 37378 6590
rect 37326 6514 37378 6526
rect 40126 6578 40178 6590
rect 43934 6578 43986 6590
rect 43698 6526 43710 6578
rect 43762 6526 43774 6578
rect 40126 6514 40178 6526
rect 43934 6514 43986 6526
rect 44270 6578 44322 6590
rect 44270 6514 44322 6526
rect 44942 6578 44994 6590
rect 44942 6514 44994 6526
rect 11118 6466 11170 6478
rect 11118 6402 11170 6414
rect 11342 6466 11394 6478
rect 11342 6402 11394 6414
rect 12686 6466 12738 6478
rect 12686 6402 12738 6414
rect 14702 6466 14754 6478
rect 14702 6402 14754 6414
rect 20302 6466 20354 6478
rect 20302 6402 20354 6414
rect 20750 6466 20802 6478
rect 20750 6402 20802 6414
rect 21422 6466 21474 6478
rect 21422 6402 21474 6414
rect 22206 6466 22258 6478
rect 22878 6466 22930 6478
rect 22530 6414 22542 6466
rect 22594 6414 22606 6466
rect 22206 6402 22258 6414
rect 22878 6402 22930 6414
rect 24110 6466 24162 6478
rect 24110 6402 24162 6414
rect 28702 6466 28754 6478
rect 28702 6402 28754 6414
rect 30158 6466 30210 6478
rect 30158 6402 30210 6414
rect 30270 6466 30322 6478
rect 30270 6402 30322 6414
rect 30830 6466 30882 6478
rect 30830 6402 30882 6414
rect 31838 6466 31890 6478
rect 31838 6402 31890 6414
rect 32062 6466 32114 6478
rect 32062 6402 32114 6414
rect 34526 6466 34578 6478
rect 34526 6402 34578 6414
rect 35758 6466 35810 6478
rect 35758 6402 35810 6414
rect 36430 6466 36482 6478
rect 36430 6402 36482 6414
rect 37438 6466 37490 6478
rect 37438 6402 37490 6414
rect 37662 6466 37714 6478
rect 37662 6402 37714 6414
rect 37998 6466 38050 6478
rect 37998 6402 38050 6414
rect 40238 6466 40290 6478
rect 40238 6402 40290 6414
rect 41582 6466 41634 6478
rect 41582 6402 41634 6414
rect 44046 6466 44098 6478
rect 44046 6402 44098 6414
rect 44830 6466 44882 6478
rect 44830 6402 44882 6414
rect 1344 6298 48608 6332
rect 1344 6246 19838 6298
rect 19890 6246 19942 6298
rect 19994 6246 20046 6298
rect 20098 6246 48608 6298
rect 1344 6212 48608 6246
rect 6302 6130 6354 6142
rect 6302 6066 6354 6078
rect 6638 6130 6690 6142
rect 6638 6066 6690 6078
rect 7422 6130 7474 6142
rect 7422 6066 7474 6078
rect 7534 6130 7586 6142
rect 7534 6066 7586 6078
rect 7646 6130 7698 6142
rect 7646 6066 7698 6078
rect 8654 6130 8706 6142
rect 12350 6130 12402 6142
rect 9762 6078 9774 6130
rect 9826 6078 9838 6130
rect 11442 6078 11454 6130
rect 11506 6078 11518 6130
rect 8654 6066 8706 6078
rect 12350 6066 12402 6078
rect 12910 6130 12962 6142
rect 12910 6066 12962 6078
rect 22542 6130 22594 6142
rect 26350 6130 26402 6142
rect 22754 6078 22766 6130
rect 22818 6078 22830 6130
rect 22542 6066 22594 6078
rect 26350 6066 26402 6078
rect 27470 6130 27522 6142
rect 27470 6066 27522 6078
rect 27694 6130 27746 6142
rect 27694 6066 27746 6078
rect 29486 6130 29538 6142
rect 29486 6066 29538 6078
rect 33182 6130 33234 6142
rect 33182 6066 33234 6078
rect 33294 6130 33346 6142
rect 46958 6130 47010 6142
rect 39442 6078 39454 6130
rect 39506 6078 39518 6130
rect 33294 6066 33346 6078
rect 46958 6066 47010 6078
rect 1710 6018 1762 6030
rect 1710 5954 1762 5966
rect 7758 6018 7810 6030
rect 7758 5954 7810 5966
rect 10782 6018 10834 6030
rect 10782 5954 10834 5966
rect 11902 6018 11954 6030
rect 11902 5954 11954 5966
rect 13134 6018 13186 6030
rect 17502 6018 17554 6030
rect 13570 5966 13582 6018
rect 13634 5966 13646 6018
rect 13134 5954 13186 5966
rect 17502 5954 17554 5966
rect 19294 6018 19346 6030
rect 19294 5954 19346 5966
rect 20078 6018 20130 6030
rect 23102 6018 23154 6030
rect 21634 5966 21646 6018
rect 21698 5966 21710 6018
rect 20078 5954 20130 5966
rect 23102 5954 23154 5966
rect 23886 6018 23938 6030
rect 23886 5954 23938 5966
rect 25790 6018 25842 6030
rect 25790 5954 25842 5966
rect 28926 6018 28978 6030
rect 28926 5954 28978 5966
rect 30382 6018 30434 6030
rect 30382 5954 30434 5966
rect 31166 6018 31218 6030
rect 31166 5954 31218 5966
rect 31502 6018 31554 6030
rect 31502 5954 31554 5966
rect 32062 6018 32114 6030
rect 33406 6018 33458 6030
rect 32386 5966 32398 6018
rect 32450 5966 32462 6018
rect 32062 5954 32114 5966
rect 33406 5954 33458 5966
rect 33742 6018 33794 6030
rect 33742 5954 33794 5966
rect 33854 6018 33906 6030
rect 33854 5954 33906 5966
rect 34414 6018 34466 6030
rect 39790 6018 39842 6030
rect 36530 5966 36542 6018
rect 36594 5966 36606 6018
rect 34414 5954 34466 5966
rect 39790 5954 39842 5966
rect 40350 6018 40402 6030
rect 48190 6018 48242 6030
rect 47282 5966 47294 6018
rect 47346 5966 47358 6018
rect 40350 5954 40402 5966
rect 48190 5954 48242 5966
rect 7086 5906 7138 5918
rect 8542 5906 8594 5918
rect 10446 5906 10498 5918
rect 8194 5854 8206 5906
rect 8258 5854 8270 5906
rect 9986 5854 9998 5906
rect 10050 5854 10062 5906
rect 7086 5842 7138 5854
rect 8542 5842 8594 5854
rect 10446 5842 10498 5854
rect 11118 5906 11170 5918
rect 11118 5842 11170 5854
rect 11790 5906 11842 5918
rect 11790 5842 11842 5854
rect 12686 5906 12738 5918
rect 12686 5842 12738 5854
rect 13246 5906 13298 5918
rect 13246 5842 13298 5854
rect 13918 5906 13970 5918
rect 17614 5906 17666 5918
rect 16706 5854 16718 5906
rect 16770 5854 16782 5906
rect 13918 5842 13970 5854
rect 17614 5842 17666 5854
rect 17950 5906 18002 5918
rect 20526 5906 20578 5918
rect 19058 5854 19070 5906
rect 19122 5854 19134 5906
rect 19842 5854 19854 5906
rect 19906 5854 19918 5906
rect 17950 5842 18002 5854
rect 20526 5842 20578 5854
rect 20862 5906 20914 5918
rect 22206 5906 22258 5918
rect 21298 5854 21310 5906
rect 21362 5854 21374 5906
rect 20862 5842 20914 5854
rect 22206 5842 22258 5854
rect 22318 5906 22370 5918
rect 22318 5842 22370 5854
rect 22766 5906 22818 5918
rect 22766 5842 22818 5854
rect 23438 5906 23490 5918
rect 23438 5842 23490 5854
rect 23774 5906 23826 5918
rect 23774 5842 23826 5854
rect 26238 5906 26290 5918
rect 26238 5842 26290 5854
rect 26462 5906 26514 5918
rect 27022 5906 27074 5918
rect 26786 5854 26798 5906
rect 26850 5854 26862 5906
rect 26462 5842 26514 5854
rect 27022 5842 27074 5854
rect 27582 5906 27634 5918
rect 27582 5842 27634 5854
rect 28590 5906 28642 5918
rect 28590 5842 28642 5854
rect 29374 5906 29426 5918
rect 29374 5842 29426 5854
rect 29598 5906 29650 5918
rect 29598 5842 29650 5854
rect 30046 5906 30098 5918
rect 30046 5842 30098 5854
rect 30494 5906 30546 5918
rect 30494 5842 30546 5854
rect 34190 5906 34242 5918
rect 34190 5842 34242 5854
rect 34526 5906 34578 5918
rect 34526 5842 34578 5854
rect 35310 5906 35362 5918
rect 39118 5906 39170 5918
rect 35858 5854 35870 5906
rect 35922 5854 35934 5906
rect 35310 5842 35362 5854
rect 39118 5842 39170 5854
rect 39902 5906 39954 5918
rect 39902 5842 39954 5854
rect 40126 5906 40178 5918
rect 46734 5906 46786 5918
rect 47854 5906 47906 5918
rect 40898 5854 40910 5906
rect 40962 5854 40974 5906
rect 43810 5854 43822 5906
rect 43874 5854 43886 5906
rect 47170 5854 47182 5906
rect 47234 5854 47246 5906
rect 40126 5842 40178 5854
rect 46734 5842 46786 5854
rect 47854 5842 47906 5854
rect 5854 5794 5906 5806
rect 5854 5730 5906 5742
rect 6974 5794 7026 5806
rect 18062 5794 18114 5806
rect 14690 5742 14702 5794
rect 14754 5742 14766 5794
rect 6974 5730 7026 5742
rect 18062 5730 18114 5742
rect 18510 5794 18562 5806
rect 18510 5730 18562 5742
rect 24446 5794 24498 5806
rect 24446 5730 24498 5742
rect 25342 5794 25394 5806
rect 25342 5730 25394 5742
rect 28142 5794 28194 5806
rect 28142 5730 28194 5742
rect 34974 5794 35026 5806
rect 34974 5730 35026 5742
rect 35422 5794 35474 5806
rect 38658 5742 38670 5794
rect 38722 5742 38734 5794
rect 42018 5742 42030 5794
rect 42082 5742 42094 5794
rect 47058 5742 47070 5794
rect 47122 5742 47134 5794
rect 35422 5730 35474 5742
rect 8654 5682 8706 5694
rect 8654 5618 8706 5630
rect 11902 5682 11954 5694
rect 11902 5618 11954 5630
rect 17502 5682 17554 5694
rect 17502 5618 17554 5630
rect 18398 5682 18450 5694
rect 18398 5618 18450 5630
rect 23886 5682 23938 5694
rect 23886 5618 23938 5630
rect 25230 5682 25282 5694
rect 25230 5618 25282 5630
rect 25902 5682 25954 5694
rect 25902 5618 25954 5630
rect 29038 5682 29090 5694
rect 29038 5618 29090 5630
rect 30382 5682 30434 5694
rect 30382 5618 30434 5630
rect 33854 5682 33906 5694
rect 33854 5618 33906 5630
rect 34862 5682 34914 5694
rect 34862 5618 34914 5630
rect 44830 5682 44882 5694
rect 44830 5618 44882 5630
rect 1344 5514 48608 5548
rect 1344 5462 4478 5514
rect 4530 5462 4582 5514
rect 4634 5462 4686 5514
rect 4738 5462 35198 5514
rect 35250 5462 35302 5514
rect 35354 5462 35406 5514
rect 35458 5462 48608 5514
rect 1344 5428 48608 5462
rect 21534 5346 21586 5358
rect 21534 5282 21586 5294
rect 21982 5346 22034 5358
rect 21982 5282 22034 5294
rect 22094 5346 22146 5358
rect 22094 5282 22146 5294
rect 22430 5346 22482 5358
rect 22430 5282 22482 5294
rect 35198 5346 35250 5358
rect 35198 5282 35250 5294
rect 37662 5346 37714 5358
rect 37662 5282 37714 5294
rect 38894 5346 38946 5358
rect 38894 5282 38946 5294
rect 20078 5234 20130 5246
rect 10322 5182 10334 5234
rect 10386 5182 10398 5234
rect 15138 5182 15150 5234
rect 15202 5182 15214 5234
rect 16930 5182 16942 5234
rect 16994 5182 17006 5234
rect 19058 5182 19070 5234
rect 19122 5182 19134 5234
rect 20078 5170 20130 5182
rect 20750 5234 20802 5246
rect 20750 5170 20802 5182
rect 21422 5234 21474 5246
rect 26798 5234 26850 5246
rect 24210 5182 24222 5234
rect 24274 5182 24286 5234
rect 26338 5182 26350 5234
rect 26402 5182 26414 5234
rect 21422 5170 21474 5182
rect 26798 5170 26850 5182
rect 28590 5234 28642 5246
rect 36318 5234 36370 5246
rect 42702 5234 42754 5246
rect 29138 5182 29150 5234
rect 29202 5182 29214 5234
rect 32610 5182 32622 5234
rect 32674 5182 32686 5234
rect 34738 5182 34750 5234
rect 34802 5182 34814 5234
rect 40114 5182 40126 5234
rect 40178 5182 40190 5234
rect 42242 5182 42254 5234
rect 42306 5182 42318 5234
rect 28590 5170 28642 5182
rect 36318 5170 36370 5182
rect 42702 5170 42754 5182
rect 5630 5122 5682 5134
rect 5630 5058 5682 5070
rect 6414 5122 6466 5134
rect 10670 5122 10722 5134
rect 20190 5122 20242 5134
rect 6962 5070 6974 5122
rect 7026 5070 7038 5122
rect 7410 5070 7422 5122
rect 7474 5070 7486 5122
rect 8194 5070 8206 5122
rect 8258 5070 8270 5122
rect 11106 5070 11118 5122
rect 11170 5070 11182 5122
rect 11330 5070 11342 5122
rect 11394 5070 11406 5122
rect 12002 5070 12014 5122
rect 12066 5070 12078 5122
rect 12786 5070 12798 5122
rect 12850 5070 12862 5122
rect 13458 5070 13470 5122
rect 13522 5070 13534 5122
rect 13794 5070 13806 5122
rect 13858 5070 13870 5122
rect 14802 5070 14814 5122
rect 14866 5070 14878 5122
rect 15026 5070 15038 5122
rect 15090 5070 15102 5122
rect 16146 5070 16158 5122
rect 16210 5070 16222 5122
rect 6414 5058 6466 5070
rect 10670 5058 10722 5070
rect 20190 5058 20242 5070
rect 22318 5122 22370 5134
rect 26686 5122 26738 5134
rect 22866 5070 22878 5122
rect 22930 5070 22942 5122
rect 23538 5070 23550 5122
rect 23602 5070 23614 5122
rect 22318 5058 22370 5070
rect 26686 5058 26738 5070
rect 27246 5122 27298 5134
rect 30606 5122 30658 5134
rect 36430 5122 36482 5134
rect 37774 5122 37826 5134
rect 28018 5070 28030 5122
rect 28082 5070 28094 5122
rect 29250 5070 29262 5122
rect 29314 5070 29326 5122
rect 29474 5070 29486 5122
rect 29538 5070 29550 5122
rect 31042 5070 31054 5122
rect 31106 5070 31118 5122
rect 31938 5070 31950 5122
rect 32002 5070 32014 5122
rect 35634 5070 35646 5122
rect 35698 5070 35710 5122
rect 37090 5070 37102 5122
rect 37154 5070 37166 5122
rect 27246 5058 27298 5070
rect 30606 5058 30658 5070
rect 36430 5058 36482 5070
rect 37774 5058 37826 5070
rect 38110 5122 38162 5134
rect 42590 5122 42642 5134
rect 43710 5122 43762 5134
rect 39442 5070 39454 5122
rect 39506 5070 39518 5122
rect 43250 5070 43262 5122
rect 43314 5070 43326 5122
rect 38110 5058 38162 5070
rect 42590 5058 42642 5070
rect 43710 5058 43762 5070
rect 44270 5122 44322 5134
rect 45042 5070 45054 5122
rect 45106 5070 45118 5122
rect 47954 5070 47966 5122
rect 48018 5070 48030 5122
rect 44270 5058 44322 5070
rect 5070 5010 5122 5022
rect 5070 4946 5122 4958
rect 6526 5010 6578 5022
rect 6526 4946 6578 4958
rect 6638 5010 6690 5022
rect 6638 4946 6690 4958
rect 10894 5010 10946 5022
rect 12574 5010 12626 5022
rect 11778 4958 11790 5010
rect 11842 4958 11854 5010
rect 10894 4946 10946 4958
rect 12574 4946 12626 4958
rect 15262 5010 15314 5022
rect 15262 4946 15314 4958
rect 19406 5010 19458 5022
rect 19406 4946 19458 4958
rect 19742 5010 19794 5022
rect 29710 5010 29762 5022
rect 23090 4958 23102 5010
rect 23154 4958 23166 5010
rect 27794 4958 27806 5010
rect 27858 4958 27870 5010
rect 19742 4946 19794 4958
rect 29710 4946 29762 4958
rect 35310 5010 35362 5022
rect 35310 4946 35362 4958
rect 36094 5010 36146 5022
rect 36094 4946 36146 4958
rect 37326 5010 37378 5022
rect 37326 4946 37378 4958
rect 38782 5010 38834 5022
rect 38782 4946 38834 4958
rect 42926 5010 42978 5022
rect 42926 4946 42978 4958
rect 47742 5010 47794 5022
rect 47742 4946 47794 4958
rect 1710 4898 1762 4910
rect 1710 4834 1762 4846
rect 5742 4898 5794 4910
rect 5742 4834 5794 4846
rect 6302 4898 6354 4910
rect 6302 4834 6354 4846
rect 10782 4898 10834 4910
rect 10782 4834 10834 4846
rect 14030 4898 14082 4910
rect 14030 4834 14082 4846
rect 14142 4898 14194 4910
rect 14142 4834 14194 4846
rect 14254 4898 14306 4910
rect 14254 4834 14306 4846
rect 15486 4898 15538 4910
rect 15486 4834 15538 4846
rect 28478 4898 28530 4910
rect 28478 4834 28530 4846
rect 29934 4898 29986 4910
rect 35198 4898 35250 4910
rect 30258 4846 30270 4898
rect 30322 4846 30334 4898
rect 31266 4846 31278 4898
rect 31330 4846 31342 4898
rect 29934 4834 29986 4846
rect 35198 4834 35250 4846
rect 36206 4898 36258 4910
rect 36206 4834 36258 4846
rect 38222 4898 38274 4910
rect 38222 4834 38274 4846
rect 38894 4898 38946 4910
rect 38894 4834 38946 4846
rect 42814 4898 42866 4910
rect 42814 4834 42866 4846
rect 45838 4898 45890 4910
rect 45838 4834 45890 4846
rect 1344 4730 48608 4764
rect 1344 4678 19838 4730
rect 19890 4678 19942 4730
rect 19994 4678 20046 4730
rect 20098 4678 48608 4730
rect 1344 4644 48608 4678
rect 7534 4562 7586 4574
rect 4050 4510 4062 4562
rect 4114 4510 4126 4562
rect 7534 4498 7586 4510
rect 8094 4562 8146 4574
rect 8094 4498 8146 4510
rect 8542 4562 8594 4574
rect 8542 4498 8594 4510
rect 17950 4562 18002 4574
rect 17950 4498 18002 4510
rect 18062 4562 18114 4574
rect 18062 4498 18114 4510
rect 21982 4562 22034 4574
rect 21982 4498 22034 4510
rect 22094 4562 22146 4574
rect 22094 4498 22146 4510
rect 22206 4562 22258 4574
rect 22206 4498 22258 4510
rect 23438 4562 23490 4574
rect 23438 4498 23490 4510
rect 24110 4562 24162 4574
rect 24110 4498 24162 4510
rect 24558 4562 24610 4574
rect 24558 4498 24610 4510
rect 25790 4562 25842 4574
rect 25790 4498 25842 4510
rect 26014 4562 26066 4574
rect 26014 4498 26066 4510
rect 33070 4562 33122 4574
rect 33070 4498 33122 4510
rect 34078 4562 34130 4574
rect 34078 4498 34130 4510
rect 34302 4562 34354 4574
rect 34302 4498 34354 4510
rect 34638 4562 34690 4574
rect 34638 4498 34690 4510
rect 36094 4562 36146 4574
rect 36094 4498 36146 4510
rect 36318 4562 36370 4574
rect 36318 4498 36370 4510
rect 40238 4562 40290 4574
rect 40238 4498 40290 4510
rect 40462 4562 40514 4574
rect 40462 4498 40514 4510
rect 43934 4562 43986 4574
rect 43934 4498 43986 4510
rect 44158 4562 44210 4574
rect 44158 4498 44210 4510
rect 47630 4562 47682 4574
rect 47630 4498 47682 4510
rect 1710 4450 1762 4462
rect 8430 4450 8482 4462
rect 6290 4398 6302 4450
rect 6354 4398 6366 4450
rect 1710 4386 1762 4398
rect 8430 4386 8482 4398
rect 8878 4450 8930 4462
rect 8878 4386 8930 4398
rect 17838 4450 17890 4462
rect 22318 4450 22370 4462
rect 19394 4398 19406 4450
rect 19458 4398 19470 4450
rect 17838 4386 17890 4398
rect 22318 4386 22370 4398
rect 23774 4450 23826 4462
rect 23774 4386 23826 4398
rect 24670 4450 24722 4462
rect 24670 4386 24722 4398
rect 25678 4450 25730 4462
rect 33966 4450 34018 4462
rect 27458 4398 27470 4450
rect 27522 4398 27534 4450
rect 33842 4398 33854 4450
rect 33906 4398 33918 4450
rect 25678 4386 25730 4398
rect 33966 4386 34018 4398
rect 34974 4450 35026 4462
rect 34974 4386 35026 4398
rect 35982 4450 36034 4462
rect 40126 4450 40178 4462
rect 38770 4398 38782 4450
rect 38834 4398 38846 4450
rect 35982 4386 36034 4398
rect 40126 4386 40178 4398
rect 43822 4450 43874 4462
rect 45154 4398 45166 4450
rect 45218 4398 45230 4450
rect 43822 4386 43874 4398
rect 7422 4338 7474 4350
rect 18174 4338 18226 4350
rect 23102 4338 23154 4350
rect 7074 4286 7086 4338
rect 7138 4286 7150 4338
rect 9650 4286 9662 4338
rect 9714 4286 9726 4338
rect 12898 4286 12910 4338
rect 12962 4286 12974 4338
rect 16594 4286 16606 4338
rect 16658 4286 16670 4338
rect 17490 4286 17502 4338
rect 17554 4286 17566 4338
rect 18722 4286 18734 4338
rect 18786 4286 18798 4338
rect 22754 4286 22766 4338
rect 22818 4286 22830 4338
rect 25218 4286 25230 4338
rect 25282 4286 25294 4338
rect 26786 4286 26798 4338
rect 26850 4286 26862 4338
rect 29922 4286 29934 4338
rect 29986 4286 29998 4338
rect 35522 4286 35534 4338
rect 35586 4286 35598 4338
rect 39554 4286 39566 4338
rect 39618 4286 39630 4338
rect 41122 4286 41134 4338
rect 41186 4286 41198 4338
rect 44482 4286 44494 4338
rect 44546 4286 44558 4338
rect 47842 4286 47854 4338
rect 47906 4286 47918 4338
rect 7422 4274 7474 4286
rect 18174 4274 18226 4286
rect 23102 4274 23154 4286
rect 7982 4226 8034 4238
rect 7982 4162 8034 4174
rect 8990 4226 9042 4238
rect 33182 4226 33234 4238
rect 13682 4174 13694 4226
rect 13746 4174 13758 4226
rect 15810 4174 15822 4226
rect 15874 4174 15886 4226
rect 16258 4174 16270 4226
rect 16322 4174 16334 4226
rect 21522 4174 21534 4226
rect 21586 4174 21598 4226
rect 25666 4174 25678 4226
rect 25730 4174 25742 4226
rect 29586 4174 29598 4226
rect 29650 4174 29662 4226
rect 8990 4162 9042 4174
rect 33182 4162 33234 4174
rect 34190 4226 34242 4238
rect 35970 4174 35982 4226
rect 36034 4174 36046 4226
rect 36642 4174 36654 4226
rect 36706 4174 36718 4226
rect 42018 4174 42030 4226
rect 42082 4174 42094 4226
rect 47282 4174 47294 4226
rect 47346 4174 47358 4226
rect 34190 4162 34242 4174
rect 7534 4114 7586 4126
rect 7534 4050 7586 4062
rect 10670 4114 10722 4126
rect 10670 4050 10722 4062
rect 24558 4114 24610 4126
rect 24558 4050 24610 4062
rect 30942 4114 30994 4126
rect 30942 4050 30994 4062
rect 1344 3946 48608 3980
rect 1344 3894 4478 3946
rect 4530 3894 4582 3946
rect 4634 3894 4686 3946
rect 4738 3894 35198 3946
rect 35250 3894 35302 3946
rect 35354 3894 35406 3946
rect 35458 3894 48608 3946
rect 1344 3860 48608 3894
rect 6190 3778 6242 3790
rect 6190 3714 6242 3726
rect 6638 3778 6690 3790
rect 6638 3714 6690 3726
rect 4622 3666 4674 3678
rect 4622 3602 4674 3614
rect 5070 3666 5122 3678
rect 5070 3602 5122 3614
rect 5854 3666 5906 3678
rect 5854 3602 5906 3614
rect 6526 3666 6578 3678
rect 6526 3602 6578 3614
rect 16158 3666 16210 3678
rect 16158 3602 16210 3614
rect 18622 3666 18674 3678
rect 18622 3602 18674 3614
rect 22094 3666 22146 3678
rect 22094 3602 22146 3614
rect 29374 3666 29426 3678
rect 29374 3602 29426 3614
rect 33854 3666 33906 3678
rect 40798 3666 40850 3678
rect 36978 3614 36990 3666
rect 37042 3614 37054 3666
rect 33854 3602 33906 3614
rect 40798 3602 40850 3614
rect 44606 3666 44658 3678
rect 44606 3602 44658 3614
rect 48190 3666 48242 3678
rect 48190 3602 48242 3614
rect 4174 3554 4226 3566
rect 8430 3554 8482 3566
rect 13470 3554 13522 3566
rect 31278 3554 31330 3566
rect 42702 3554 42754 3566
rect 7186 3502 7198 3554
rect 7250 3502 7262 3554
rect 7858 3502 7870 3554
rect 7922 3502 7934 3554
rect 9538 3502 9550 3554
rect 9602 3502 9614 3554
rect 10434 3502 10446 3554
rect 10498 3502 10510 3554
rect 14242 3502 14254 3554
rect 14306 3502 14318 3554
rect 17042 3502 17054 3554
rect 17106 3502 17118 3554
rect 17714 3502 17726 3554
rect 17778 3502 17790 3554
rect 21074 3502 21086 3554
rect 21138 3502 21150 3554
rect 24658 3502 24670 3554
rect 24722 3502 24734 3554
rect 25442 3502 25454 3554
rect 25506 3502 25518 3554
rect 28578 3502 28590 3554
rect 28642 3502 28654 3554
rect 32274 3502 32286 3554
rect 32338 3502 32350 3554
rect 33282 3502 33294 3554
rect 33346 3502 33358 3554
rect 36194 3502 36206 3554
rect 36258 3502 36270 3554
rect 39106 3502 39118 3554
rect 39170 3502 39182 3554
rect 40002 3502 40014 3554
rect 40066 3502 40078 3554
rect 43698 3502 43710 3554
rect 43762 3502 43774 3554
rect 46722 3502 46734 3554
rect 46786 3502 46798 3554
rect 47618 3502 47630 3554
rect 47682 3502 47694 3554
rect 4174 3490 4226 3502
rect 8430 3490 8482 3502
rect 13470 3490 13522 3502
rect 31278 3490 31330 3502
rect 42702 3490 42754 3502
rect 6078 3442 6130 3454
rect 6078 3378 6130 3390
rect 6974 3442 7026 3454
rect 6974 3378 7026 3390
rect 7646 3442 7698 3454
rect 7646 3378 7698 3390
rect 8766 3442 8818 3454
rect 8766 3378 8818 3390
rect 9326 3442 9378 3454
rect 13134 3442 13186 3454
rect 11554 3390 11566 3442
rect 11618 3390 11630 3442
rect 9326 3378 9378 3390
rect 13134 3378 13186 3390
rect 17278 3442 17330 3454
rect 17278 3378 17330 3390
rect 24894 3442 24946 3454
rect 32510 3442 32562 3454
rect 26898 3390 26910 3442
rect 26962 3390 26974 3442
rect 31602 3390 31614 3442
rect 31666 3390 31678 3442
rect 24894 3378 24946 3390
rect 32510 3378 32562 3390
rect 35982 3442 36034 3454
rect 46510 3442 46562 3454
rect 43026 3390 43038 3442
rect 43090 3390 43102 3442
rect 35982 3378 36034 3390
rect 46510 3378 46562 3390
rect 47406 3442 47458 3454
rect 47406 3378 47458 3390
rect 48078 3442 48130 3454
rect 48078 3378 48130 3390
rect 1710 3330 1762 3342
rect 1710 3266 1762 3278
rect 2158 3330 2210 3342
rect 2158 3266 2210 3278
rect 1344 3162 48608 3196
rect 1344 3110 19838 3162
rect 19890 3110 19942 3162
rect 19994 3110 20046 3162
rect 20098 3110 48608 3162
rect 1344 3076 48608 3110
<< via1 >>
rect 4478 46230 4530 46282
rect 4582 46230 4634 46282
rect 4686 46230 4738 46282
rect 35198 46230 35250 46282
rect 35302 46230 35354 46282
rect 35406 46230 35458 46282
rect 29374 46062 29426 46114
rect 33182 46062 33234 46114
rect 36990 46062 37042 46114
rect 10670 45950 10722 46002
rect 17726 45950 17778 46002
rect 26910 45950 26962 46002
rect 13918 45838 13970 45890
rect 15262 45838 15314 45890
rect 16270 45838 16322 45890
rect 18398 45838 18450 45890
rect 19630 45838 19682 45890
rect 20078 45838 20130 45890
rect 23886 45838 23938 45890
rect 25454 45838 25506 45890
rect 28590 45838 28642 45890
rect 31502 45838 31554 45890
rect 32174 45838 32226 45890
rect 35982 45838 36034 45890
rect 39790 45838 39842 45890
rect 42926 45838 42978 45890
rect 44046 45838 44098 45890
rect 19406 45726 19458 45778
rect 24558 45726 24610 45778
rect 35422 45726 35474 45778
rect 39230 45726 39282 45778
rect 1710 45614 1762 45666
rect 8094 45614 8146 45666
rect 9550 45614 9602 45666
rect 11118 45614 11170 45666
rect 11678 45614 11730 45666
rect 12126 45614 12178 45666
rect 12574 45614 12626 45666
rect 13470 45614 13522 45666
rect 13694 45614 13746 45666
rect 14590 45614 14642 45666
rect 15038 45614 15090 45666
rect 15822 45614 15874 45666
rect 17166 45614 17218 45666
rect 18174 45614 18226 45666
rect 18734 45614 18786 45666
rect 20974 45614 21026 45666
rect 22990 45614 23042 45666
rect 24894 45614 24946 45666
rect 31278 45614 31330 45666
rect 35086 45614 35138 45666
rect 38894 45614 38946 45666
rect 40798 45614 40850 45666
rect 42702 45614 42754 45666
rect 44606 45614 44658 45666
rect 46846 45614 46898 45666
rect 47742 45614 47794 45666
rect 48190 45614 48242 45666
rect 19838 45446 19890 45498
rect 19942 45446 19994 45498
rect 20046 45446 20098 45498
rect 25342 45278 25394 45330
rect 30158 45278 30210 45330
rect 31278 45278 31330 45330
rect 46062 45278 46114 45330
rect 26462 45166 26514 45218
rect 29038 45166 29090 45218
rect 31950 45166 32002 45218
rect 32398 45166 32450 45218
rect 34638 45166 34690 45218
rect 37886 45166 37938 45218
rect 42590 45166 42642 45218
rect 48190 45166 48242 45218
rect 13246 45054 13298 45106
rect 13694 45054 13746 45106
rect 17614 45054 17666 45106
rect 20750 45054 20802 45106
rect 24446 45054 24498 45106
rect 25678 45054 25730 45106
rect 26350 45054 26402 45106
rect 29822 45054 29874 45106
rect 30382 45054 30434 45106
rect 33966 45054 34018 45106
rect 37102 45054 37154 45106
rect 41806 45054 41858 45106
rect 45054 45054 45106 45106
rect 7422 44942 7474 44994
rect 7982 44942 8034 44994
rect 8430 44942 8482 44994
rect 9102 44942 9154 44994
rect 9662 44942 9714 44994
rect 10110 44942 10162 44994
rect 10446 44942 10498 44994
rect 12574 44942 12626 44994
rect 14478 44942 14530 44994
rect 16606 44942 16658 44994
rect 18286 44942 18338 44994
rect 20414 44942 20466 44994
rect 21534 44942 21586 44994
rect 23662 44942 23714 44994
rect 24110 44942 24162 44994
rect 26910 44942 26962 44994
rect 33294 44942 33346 44994
rect 36766 44942 36818 44994
rect 40014 44942 40066 44994
rect 41134 44942 41186 44994
rect 41582 44942 41634 44994
rect 44718 44942 44770 44994
rect 7534 44830 7586 44882
rect 8430 44830 8482 44882
rect 31614 44830 31666 44882
rect 4478 44662 4530 44714
rect 4582 44662 4634 44714
rect 4686 44662 4738 44714
rect 35198 44662 35250 44714
rect 35302 44662 35354 44714
rect 35406 44662 35458 44714
rect 27358 44494 27410 44546
rect 27694 44494 27746 44546
rect 34526 44494 34578 44546
rect 42030 44494 42082 44546
rect 44942 44494 44994 44546
rect 11678 44382 11730 44434
rect 17390 44382 17442 44434
rect 20638 44382 20690 44434
rect 23102 44382 23154 44434
rect 25230 44382 25282 44434
rect 31054 44382 31106 44434
rect 33182 44382 33234 44434
rect 37102 44382 37154 44434
rect 40686 44382 40738 44434
rect 7422 44270 7474 44322
rect 7870 44270 7922 44322
rect 8094 44270 8146 44322
rect 8766 44270 8818 44322
rect 17838 44270 17890 44322
rect 21870 44270 21922 44322
rect 25902 44270 25954 44322
rect 28366 44270 28418 44322
rect 29934 44270 29986 44322
rect 30382 44270 30434 44322
rect 33742 44270 33794 44322
rect 37774 44270 37826 44322
rect 41022 44270 41074 44322
rect 44158 44270 44210 44322
rect 45278 44270 45330 44322
rect 45726 44270 45778 44322
rect 47182 44270 47234 44322
rect 8430 44158 8482 44210
rect 9550 44158 9602 44210
rect 12910 44158 12962 44210
rect 14702 44158 14754 44210
rect 16382 44158 16434 44210
rect 16494 44158 16546 44210
rect 18510 44158 18562 44210
rect 22094 44158 22146 44210
rect 22654 44158 22706 44210
rect 28478 44158 28530 44210
rect 38558 44158 38610 44210
rect 45838 44158 45890 44210
rect 47518 44158 47570 44210
rect 47966 44158 48018 44210
rect 4846 44046 4898 44098
rect 5854 44046 5906 44098
rect 6414 44046 6466 44098
rect 6862 44046 6914 44098
rect 7198 44046 7250 44098
rect 7310 44046 7362 44098
rect 8318 44046 8370 44098
rect 12014 44046 12066 44098
rect 12350 44046 12402 44098
rect 12574 44046 12626 44098
rect 12798 44046 12850 44098
rect 13694 44046 13746 44098
rect 14142 44046 14194 44098
rect 14366 44046 14418 44098
rect 14590 44046 14642 44098
rect 15486 44046 15538 44098
rect 15822 44046 15874 44098
rect 16158 44046 16210 44098
rect 17054 44046 17106 44098
rect 21534 44046 21586 44098
rect 26462 44046 26514 44098
rect 29374 44046 29426 44098
rect 43934 44046 43986 44098
rect 46846 44046 46898 44098
rect 19838 43878 19890 43930
rect 19942 43878 19994 43930
rect 20046 43878 20098 43930
rect 15598 43710 15650 43762
rect 21422 43710 21474 43762
rect 29150 43710 29202 43762
rect 45278 43710 45330 43762
rect 6862 43598 6914 43650
rect 11454 43598 11506 43650
rect 16494 43598 16546 43650
rect 18286 43598 18338 43650
rect 18622 43598 18674 43650
rect 19070 43598 19122 43650
rect 23662 43598 23714 43650
rect 25342 43598 25394 43650
rect 39006 43598 39058 43650
rect 39566 43598 39618 43650
rect 39902 43598 39954 43650
rect 40910 43598 40962 43650
rect 43934 43598 43986 43650
rect 6190 43486 6242 43538
rect 9998 43486 10050 43538
rect 10894 43486 10946 43538
rect 11342 43486 11394 43538
rect 11566 43486 11618 43538
rect 11902 43486 11954 43538
rect 12462 43486 12514 43538
rect 15710 43486 15762 43538
rect 16270 43486 16322 43538
rect 18958 43486 19010 43538
rect 19294 43486 19346 43538
rect 21646 43486 21698 43538
rect 22542 43486 22594 43538
rect 25902 43486 25954 43538
rect 29710 43486 29762 43538
rect 33294 43486 33346 43538
rect 35982 43486 36034 43538
rect 39342 43486 39394 43538
rect 41246 43486 41298 43538
rect 44606 43486 44658 43538
rect 45838 43486 45890 43538
rect 1822 43374 1874 43426
rect 2270 43374 2322 43426
rect 3950 43374 4002 43426
rect 4398 43374 4450 43426
rect 4846 43374 4898 43426
rect 5406 43374 5458 43426
rect 5854 43374 5906 43426
rect 8990 43374 9042 43426
rect 9550 43374 9602 43426
rect 10446 43374 10498 43426
rect 13134 43374 13186 43426
rect 15262 43374 15314 43426
rect 17502 43374 17554 43426
rect 17950 43374 18002 43426
rect 19742 43374 19794 43426
rect 20638 43374 20690 43426
rect 21086 43374 21138 43426
rect 26574 43374 26626 43426
rect 28702 43374 28754 43426
rect 30382 43374 30434 43426
rect 32510 43374 32562 43426
rect 34078 43374 34130 43426
rect 36990 43374 37042 43426
rect 41806 43374 41858 43426
rect 3838 43262 3890 43314
rect 4846 43262 4898 43314
rect 15934 43262 15986 43314
rect 47966 43262 48018 43314
rect 4478 43094 4530 43146
rect 4582 43094 4634 43146
rect 4686 43094 4738 43146
rect 35198 43094 35250 43146
rect 35302 43094 35354 43146
rect 35406 43094 35458 43146
rect 29598 42926 29650 42978
rect 32174 42926 32226 42978
rect 34526 42926 34578 42978
rect 37214 42926 37266 42978
rect 40126 42926 40178 42978
rect 42926 42926 42978 42978
rect 43262 42926 43314 42978
rect 10110 42814 10162 42866
rect 13694 42814 13746 42866
rect 14590 42814 14642 42866
rect 15710 42814 15762 42866
rect 19070 42814 19122 42866
rect 26126 42814 26178 42866
rect 46958 42814 47010 42866
rect 5630 42702 5682 42754
rect 9102 42702 9154 42754
rect 11006 42702 11058 42754
rect 11342 42702 11394 42754
rect 13806 42702 13858 42754
rect 14254 42702 14306 42754
rect 18622 42702 18674 42754
rect 19966 42702 20018 42754
rect 20414 42702 20466 42754
rect 23326 42702 23378 42754
rect 31166 42702 31218 42754
rect 36206 42702 36258 42754
rect 39342 42702 39394 42754
rect 42030 42702 42082 42754
rect 43710 42702 43762 42754
rect 48190 42702 48242 42754
rect 6414 42590 6466 42642
rect 9214 42590 9266 42642
rect 10222 42590 10274 42642
rect 11454 42590 11506 42642
rect 17838 42590 17890 42642
rect 19406 42590 19458 42642
rect 23998 42590 24050 42642
rect 27022 42590 27074 42642
rect 27358 42590 27410 42642
rect 29262 42590 29314 42642
rect 29934 42590 29986 42642
rect 30270 42590 30322 42642
rect 34750 42590 34802 42642
rect 35086 42590 35138 42642
rect 43822 42590 43874 42642
rect 45278 42590 45330 42642
rect 1822 42478 1874 42530
rect 2494 42478 2546 42530
rect 2942 42478 2994 42530
rect 3390 42478 3442 42530
rect 3950 42478 4002 42530
rect 4398 42478 4450 42530
rect 4846 42478 4898 42530
rect 8654 42478 8706 42530
rect 9438 42478 9490 42530
rect 13582 42478 13634 42530
rect 15038 42478 15090 42530
rect 18958 42478 19010 42530
rect 19182 42478 19234 42530
rect 26574 42478 26626 42530
rect 34190 42478 34242 42530
rect 36430 42478 36482 42530
rect 19838 42310 19890 42362
rect 19942 42310 19994 42362
rect 20046 42310 20098 42362
rect 7982 42142 8034 42194
rect 12462 42142 12514 42194
rect 15262 42142 15314 42194
rect 15598 42142 15650 42194
rect 24222 42142 24274 42194
rect 31278 42142 31330 42194
rect 48190 42142 48242 42194
rect 4846 42030 4898 42082
rect 5854 42030 5906 42082
rect 8878 42030 8930 42082
rect 11902 42030 11954 42082
rect 16606 42030 16658 42082
rect 18286 42030 18338 42082
rect 18958 42030 19010 42082
rect 26238 42030 26290 42082
rect 27694 42030 27746 42082
rect 30382 42030 30434 42082
rect 31614 42030 31666 42082
rect 1710 41918 1762 41970
rect 3838 41918 3890 41970
rect 4286 41918 4338 41970
rect 4622 41918 4674 41970
rect 6974 41918 7026 41970
rect 7422 41918 7474 41970
rect 10446 41918 10498 41970
rect 10670 41918 10722 41970
rect 13358 41918 13410 41970
rect 13582 41918 13634 41970
rect 13806 41918 13858 41970
rect 14030 41918 14082 41970
rect 14366 41918 14418 41970
rect 14926 41918 14978 41970
rect 15934 41918 15986 41970
rect 18510 41918 18562 41970
rect 20638 41918 20690 41970
rect 23774 41918 23826 41970
rect 24558 41918 24610 41970
rect 26350 41918 26402 41970
rect 27470 41918 27522 41970
rect 30718 41918 30770 41970
rect 32510 41918 32562 41970
rect 33182 41918 33234 41970
rect 36318 41918 36370 41970
rect 37102 41918 37154 41970
rect 39678 41918 39730 41970
rect 44494 41918 44546 41970
rect 44830 41918 44882 41970
rect 2270 41806 2322 41858
rect 3166 41806 3218 41858
rect 9774 41806 9826 41858
rect 11566 41806 11618 41858
rect 12910 41806 12962 41858
rect 16158 41806 16210 41858
rect 17502 41806 17554 41858
rect 20974 41806 21026 41858
rect 23102 41806 23154 41858
rect 25342 41806 25394 41858
rect 28814 41806 28866 41858
rect 30046 41806 30098 41858
rect 33854 41806 33906 41858
rect 35982 41806 36034 41858
rect 39230 41806 39282 41858
rect 40126 41806 40178 41858
rect 41022 41806 41074 41858
rect 41582 41806 41634 41858
rect 43710 41806 43762 41858
rect 45614 41806 45666 41858
rect 47742 41806 47794 41858
rect 10334 41694 10386 41746
rect 16718 41694 16770 41746
rect 25678 41694 25730 41746
rect 4478 41526 4530 41578
rect 4582 41526 4634 41578
rect 4686 41526 4738 41578
rect 35198 41526 35250 41578
rect 35302 41526 35354 41578
rect 35406 41526 35458 41578
rect 12686 41358 12738 41410
rect 16270 41358 16322 41410
rect 34638 41358 34690 41410
rect 37214 41358 37266 41410
rect 37550 41358 37602 41410
rect 5070 41246 5122 41298
rect 5854 41246 5906 41298
rect 15038 41246 15090 41298
rect 17278 41246 17330 41298
rect 18398 41246 18450 41298
rect 21758 41246 21810 41298
rect 24110 41246 24162 41298
rect 24894 41246 24946 41298
rect 25678 41246 25730 41298
rect 27806 41246 27858 41298
rect 30158 41246 30210 41298
rect 32286 41246 32338 41298
rect 32734 41246 32786 41298
rect 43934 41246 43986 41298
rect 47854 41246 47906 41298
rect 2158 41134 2210 41186
rect 5630 41134 5682 41186
rect 8766 41134 8818 41186
rect 9326 41134 9378 41186
rect 11006 41134 11058 41186
rect 12910 41134 12962 41186
rect 13806 41134 13858 41186
rect 14926 41134 14978 41186
rect 15710 41134 15762 41186
rect 16382 41134 16434 41186
rect 17054 41134 17106 41186
rect 17390 41134 17442 41186
rect 18510 41134 18562 41186
rect 19854 41134 19906 41186
rect 20414 41134 20466 41186
rect 21310 41134 21362 41186
rect 28590 41134 28642 41186
rect 29374 41134 29426 41186
rect 33630 41134 33682 41186
rect 35198 41134 35250 41186
rect 36206 41134 36258 41186
rect 38894 41134 38946 41186
rect 39230 41134 39282 41186
rect 39678 41134 39730 41186
rect 40798 41134 40850 41186
rect 41470 41134 41522 41186
rect 41806 41134 41858 41186
rect 45614 41134 45666 41186
rect 2942 41022 2994 41074
rect 7086 41022 7138 41074
rect 7982 41022 8034 41074
rect 9774 41022 9826 41074
rect 12126 41022 12178 41074
rect 12350 41022 12402 41074
rect 14254 41022 14306 41074
rect 15934 41022 15986 41074
rect 16830 41022 16882 41074
rect 18286 41022 18338 41074
rect 18846 41022 18898 41074
rect 19966 41022 20018 41074
rect 20302 41022 20354 41074
rect 22654 41022 22706 41074
rect 33854 41022 33906 41074
rect 34302 41022 34354 41074
rect 35422 41022 35474 41074
rect 37774 41022 37826 41074
rect 38222 41022 38274 41074
rect 39790 41022 39842 41074
rect 42030 41022 42082 41074
rect 42366 41022 42418 41074
rect 43150 41022 43202 41074
rect 44942 41022 44994 41074
rect 45278 41022 45330 41074
rect 1822 40910 1874 40962
rect 9326 40910 9378 40962
rect 12462 40910 12514 40962
rect 13582 40910 13634 40962
rect 16494 40910 16546 40962
rect 17950 40910 18002 40962
rect 19406 40910 19458 40962
rect 22990 40910 23042 40962
rect 36430 40910 36482 40962
rect 41022 40910 41074 40962
rect 43486 40910 43538 40962
rect 19838 40742 19890 40794
rect 19942 40742 19994 40794
rect 20046 40742 20098 40794
rect 6302 40574 6354 40626
rect 7198 40574 7250 40626
rect 15934 40574 15986 40626
rect 18286 40574 18338 40626
rect 19742 40574 19794 40626
rect 28254 40574 28306 40626
rect 30942 40574 30994 40626
rect 36318 40574 36370 40626
rect 43822 40574 43874 40626
rect 44606 40574 44658 40626
rect 5294 40462 5346 40514
rect 5966 40462 6018 40514
rect 10558 40462 10610 40514
rect 11902 40462 11954 40514
rect 13022 40462 13074 40514
rect 15486 40462 15538 40514
rect 16830 40462 16882 40514
rect 20414 40462 20466 40514
rect 20862 40462 20914 40514
rect 22318 40462 22370 40514
rect 23214 40462 23266 40514
rect 26462 40462 26514 40514
rect 27022 40462 27074 40514
rect 29262 40462 29314 40514
rect 31502 40462 31554 40514
rect 31950 40462 32002 40514
rect 35646 40462 35698 40514
rect 37438 40462 37490 40514
rect 41694 40462 41746 40514
rect 42030 40462 42082 40514
rect 42926 40462 42978 40514
rect 45278 40462 45330 40514
rect 1822 40350 1874 40402
rect 5070 40350 5122 40402
rect 8766 40350 8818 40402
rect 11006 40350 11058 40402
rect 11342 40350 11394 40402
rect 13694 40350 13746 40402
rect 14814 40350 14866 40402
rect 16718 40350 16770 40402
rect 18846 40350 18898 40402
rect 19182 40350 19234 40402
rect 20190 40350 20242 40402
rect 20638 40350 20690 40402
rect 20974 40350 21026 40402
rect 22766 40350 22818 40402
rect 23438 40350 23490 40402
rect 29150 40350 29202 40402
rect 29934 40350 29986 40402
rect 33182 40350 33234 40402
rect 33966 40350 34018 40402
rect 35198 40350 35250 40402
rect 36654 40350 36706 40402
rect 42702 40350 42754 40402
rect 45054 40350 45106 40402
rect 45614 40350 45666 40402
rect 2494 40238 2546 40290
rect 4622 40238 4674 40290
rect 6638 40238 6690 40290
rect 8094 40238 8146 40290
rect 9886 40238 9938 40290
rect 10110 40238 10162 40290
rect 10894 40238 10946 40290
rect 16046 40238 16098 40290
rect 17614 40238 17666 40290
rect 17950 40238 18002 40290
rect 19294 40238 19346 40290
rect 26238 40238 26290 40290
rect 31278 40238 31330 40290
rect 33518 40238 33570 40290
rect 34414 40238 34466 40290
rect 39566 40238 39618 40290
rect 40014 40238 40066 40290
rect 7646 40126 7698 40178
rect 8318 40126 8370 40178
rect 8542 40126 8594 40178
rect 9438 40126 9490 40178
rect 10334 40126 10386 40178
rect 16270 40126 16322 40178
rect 19518 40126 19570 40178
rect 19742 40126 19794 40178
rect 25902 40126 25954 40178
rect 28590 40126 28642 40178
rect 41022 40126 41074 40178
rect 41358 40126 41410 40178
rect 43486 40126 43538 40178
rect 47966 40126 48018 40178
rect 4478 39958 4530 40010
rect 4582 39958 4634 40010
rect 4686 39958 4738 40010
rect 35198 39958 35250 40010
rect 35302 39958 35354 40010
rect 35406 39958 35458 40010
rect 6302 39790 6354 39842
rect 7422 39790 7474 39842
rect 7646 39790 7698 39842
rect 7870 39790 7922 39842
rect 13470 39790 13522 39842
rect 16494 39790 16546 39842
rect 16830 39790 16882 39842
rect 17166 39790 17218 39842
rect 38334 39790 38386 39842
rect 38670 39790 38722 39842
rect 43038 39790 43090 39842
rect 43374 39790 43426 39842
rect 2270 39678 2322 39730
rect 3390 39678 3442 39730
rect 7198 39678 7250 39730
rect 18958 39678 19010 39730
rect 22990 39678 23042 39730
rect 26798 39678 26850 39730
rect 31614 39678 31666 39730
rect 34862 39678 34914 39730
rect 36430 39678 36482 39730
rect 37102 39678 37154 39730
rect 42030 39678 42082 39730
rect 46062 39678 46114 39730
rect 48190 39678 48242 39730
rect 1710 39566 1762 39618
rect 2606 39566 2658 39618
rect 3278 39566 3330 39618
rect 3838 39566 3890 39618
rect 4062 39566 4114 39618
rect 10334 39566 10386 39618
rect 12350 39566 12402 39618
rect 14254 39566 14306 39618
rect 15822 39566 15874 39618
rect 16046 39566 16098 39618
rect 17166 39566 17218 39618
rect 18398 39566 18450 39618
rect 18622 39566 18674 39618
rect 19854 39566 19906 39618
rect 20302 39566 20354 39618
rect 22094 39566 22146 39618
rect 22654 39566 22706 39618
rect 23438 39566 23490 39618
rect 23998 39566 24050 39618
rect 31950 39566 32002 39618
rect 39118 39566 39170 39618
rect 44158 39566 44210 39618
rect 45390 39566 45442 39618
rect 2942 39454 2994 39506
rect 4398 39454 4450 39506
rect 5966 39454 6018 39506
rect 6190 39454 6242 39506
rect 8542 39454 8594 39506
rect 11230 39454 11282 39506
rect 13918 39454 13970 39506
rect 14030 39454 14082 39506
rect 14702 39454 14754 39506
rect 15934 39454 15986 39506
rect 18846 39454 18898 39506
rect 19070 39454 19122 39506
rect 19406 39454 19458 39506
rect 24670 39454 24722 39506
rect 32734 39454 32786 39506
rect 35198 39454 35250 39506
rect 37774 39454 37826 39506
rect 38110 39454 38162 39506
rect 39902 39454 39954 39506
rect 43934 39454 43986 39506
rect 3502 39342 3554 39394
rect 4286 39342 4338 39394
rect 4846 39342 4898 39394
rect 6862 39342 6914 39394
rect 8318 39342 8370 39394
rect 9886 39342 9938 39394
rect 13022 39342 13074 39394
rect 14590 39342 14642 39394
rect 15262 39342 15314 39394
rect 18062 39342 18114 39394
rect 21422 39342 21474 39394
rect 27246 39342 27298 39394
rect 29262 39342 29314 39394
rect 35534 39342 35586 39394
rect 42478 39342 42530 39394
rect 45054 39342 45106 39394
rect 19838 39174 19890 39226
rect 19942 39174 19994 39226
rect 20046 39174 20098 39226
rect 6526 39006 6578 39058
rect 6750 39006 6802 39058
rect 8542 39006 8594 39058
rect 9998 39006 10050 39058
rect 10894 39006 10946 39058
rect 16046 39006 16098 39058
rect 20302 39006 20354 39058
rect 21646 39006 21698 39058
rect 21870 39006 21922 39058
rect 22654 39006 22706 39058
rect 22990 39006 23042 39058
rect 23662 39006 23714 39058
rect 25230 39006 25282 39058
rect 31838 39006 31890 39058
rect 33070 39006 33122 39058
rect 40238 39006 40290 39058
rect 40910 39006 40962 39058
rect 41694 39006 41746 39058
rect 5294 38894 5346 38946
rect 7982 38894 8034 38946
rect 11790 38894 11842 38946
rect 12238 38894 12290 38946
rect 18174 38894 18226 38946
rect 19518 38894 19570 38946
rect 20526 38894 20578 38946
rect 21198 38894 21250 38946
rect 21310 38894 21362 38946
rect 23326 38894 23378 38946
rect 25566 38894 25618 38946
rect 30382 38894 30434 38946
rect 31054 38894 31106 38946
rect 35086 38894 35138 38946
rect 39342 38894 39394 38946
rect 39566 38894 39618 38946
rect 43262 38894 43314 38946
rect 45950 38894 46002 38946
rect 47854 38894 47906 38946
rect 1822 38782 1874 38834
rect 5742 38782 5794 38834
rect 5854 38782 5906 38834
rect 6302 38782 6354 38834
rect 7086 38782 7138 38834
rect 7534 38782 7586 38834
rect 10446 38782 10498 38834
rect 13246 38782 13298 38834
rect 13806 38782 13858 38834
rect 14926 38782 14978 38834
rect 15486 38782 15538 38834
rect 21534 38782 21586 38834
rect 21982 38782 22034 38834
rect 26126 38782 26178 38834
rect 29822 38782 29874 38834
rect 30494 38782 30546 38834
rect 31278 38782 31330 38834
rect 33406 38782 33458 38834
rect 34078 38782 34130 38834
rect 34414 38782 34466 38834
rect 35198 38782 35250 38834
rect 35870 38782 35922 38834
rect 39902 38782 39954 38834
rect 41134 38782 41186 38834
rect 42478 38782 42530 38834
rect 46286 38782 46338 38834
rect 46734 38782 46786 38834
rect 47518 38782 47570 38834
rect 2494 38670 2546 38722
rect 4734 38670 4786 38722
rect 5182 38670 5234 38722
rect 6078 38670 6130 38722
rect 8990 38670 9042 38722
rect 11342 38670 11394 38722
rect 15598 38670 15650 38722
rect 16830 38670 16882 38722
rect 17838 38670 17890 38722
rect 19854 38670 19906 38722
rect 20190 38670 20242 38722
rect 24110 38670 24162 38722
rect 26910 38670 26962 38722
rect 29038 38670 29090 38722
rect 29486 38670 29538 38722
rect 36542 38670 36594 38722
rect 38670 38670 38722 38722
rect 42142 38670 42194 38722
rect 45390 38643 45442 38695
rect 47070 38670 47122 38722
rect 6862 38558 6914 38610
rect 11678 38558 11730 38610
rect 12350 38558 12402 38610
rect 13806 38558 13858 38610
rect 4478 38390 4530 38442
rect 4582 38390 4634 38442
rect 4686 38390 4738 38442
rect 35198 38390 35250 38442
rect 35302 38390 35354 38442
rect 35406 38390 35458 38442
rect 7758 38222 7810 38274
rect 20078 38222 20130 38274
rect 23662 38222 23714 38274
rect 24110 38222 24162 38274
rect 24334 38222 24386 38274
rect 37550 38222 37602 38274
rect 2270 38110 2322 38162
rect 2718 38110 2770 38162
rect 3614 38110 3666 38162
rect 4846 38110 4898 38162
rect 6190 38110 6242 38162
rect 7646 38110 7698 38162
rect 8318 38110 8370 38162
rect 8654 38110 8706 38162
rect 9886 38110 9938 38162
rect 12798 38110 12850 38162
rect 13694 38110 13746 38162
rect 17390 38110 17442 38162
rect 18622 38110 18674 38162
rect 19406 38110 19458 38162
rect 23662 38110 23714 38162
rect 24110 38110 24162 38162
rect 30046 38110 30098 38162
rect 32174 38110 32226 38162
rect 32622 38110 32674 38162
rect 34526 38110 34578 38162
rect 38894 38110 38946 38162
rect 42142 38110 42194 38162
rect 42590 38110 42642 38162
rect 44942 38110 44994 38162
rect 48190 38110 48242 38162
rect 1710 37998 1762 38050
rect 2830 37998 2882 38050
rect 3278 37998 3330 38050
rect 6526 37998 6578 38050
rect 8094 37998 8146 38050
rect 8542 37998 8594 38050
rect 9662 37998 9714 38050
rect 11118 37998 11170 38050
rect 11454 37998 11506 38050
rect 12014 37998 12066 38050
rect 12350 37998 12402 38050
rect 14702 37998 14754 38050
rect 15038 37998 15090 38050
rect 15822 37998 15874 38050
rect 16270 37998 16322 38050
rect 16494 37998 16546 38050
rect 16718 37998 16770 38050
rect 16830 37998 16882 38050
rect 19854 37998 19906 38050
rect 20302 37998 20354 38050
rect 21198 37998 21250 38050
rect 27694 37998 27746 38050
rect 29374 37998 29426 38050
rect 34862 37998 34914 38050
rect 36206 37998 36258 38050
rect 39230 37998 39282 38050
rect 43374 37998 43426 38050
rect 45278 37998 45330 38050
rect 4174 37886 4226 37938
rect 4510 37886 4562 37938
rect 7086 37886 7138 37938
rect 7534 37886 7586 37938
rect 10334 37886 10386 37938
rect 11230 37886 11282 37938
rect 12462 37886 12514 37938
rect 13582 37886 13634 37938
rect 14366 37886 14418 37938
rect 15710 37886 15762 37938
rect 17502 37886 17554 37938
rect 17950 37886 18002 37938
rect 18062 37886 18114 37938
rect 18510 37886 18562 37938
rect 18734 37886 18786 37938
rect 21646 37886 21698 37938
rect 22654 37886 22706 37938
rect 27358 37886 27410 37938
rect 36430 37886 36482 37938
rect 37214 37886 37266 37938
rect 37774 37886 37826 37938
rect 38222 37886 38274 37938
rect 40014 37886 40066 37938
rect 43710 37886 43762 37938
rect 44158 37886 44210 37938
rect 46062 37886 46114 37938
rect 2606 37774 2658 37826
rect 3614 37774 3666 37826
rect 3726 37774 3778 37826
rect 3950 37774 4002 37826
rect 8766 37774 8818 37826
rect 10670 37774 10722 37826
rect 13806 37774 13858 37826
rect 14030 37774 14082 37826
rect 16606 37774 16658 37826
rect 17726 37774 17778 37826
rect 20750 37774 20802 37826
rect 21758 37774 21810 37826
rect 21870 37774 21922 37826
rect 22318 37774 22370 37826
rect 22766 37774 22818 37826
rect 22990 37774 23042 37826
rect 24670 37774 24722 37826
rect 43038 37774 43090 37826
rect 19838 37606 19890 37658
rect 19942 37606 19994 37658
rect 20046 37606 20098 37658
rect 3614 37438 3666 37490
rect 6078 37438 6130 37490
rect 6190 37438 6242 37490
rect 11118 37438 11170 37490
rect 11790 37438 11842 37490
rect 15822 37438 15874 37490
rect 16046 37438 16098 37490
rect 19518 37438 19570 37490
rect 31054 37438 31106 37490
rect 35422 37438 35474 37490
rect 39454 37438 39506 37490
rect 39902 37438 39954 37490
rect 40350 37438 40402 37490
rect 41022 37438 41074 37490
rect 41694 37438 41746 37490
rect 2046 37326 2098 37378
rect 3054 37326 3106 37378
rect 3838 37326 3890 37378
rect 7310 37326 7362 37378
rect 8206 37326 8258 37378
rect 8990 37326 9042 37378
rect 10110 37326 10162 37378
rect 11678 37326 11730 37378
rect 14142 37326 14194 37378
rect 15710 37326 15762 37378
rect 16382 37326 16434 37378
rect 17614 37326 17666 37378
rect 17726 37326 17778 37378
rect 19406 37326 19458 37378
rect 21646 37326 21698 37378
rect 23438 37326 23490 37378
rect 23550 37326 23602 37378
rect 23774 37326 23826 37378
rect 24222 37326 24274 37378
rect 29150 37326 29202 37378
rect 31614 37326 31666 37378
rect 32174 37326 32226 37378
rect 37774 37326 37826 37378
rect 1710 37214 1762 37266
rect 3950 37214 4002 37266
rect 4622 37214 4674 37266
rect 4846 37214 4898 37266
rect 5630 37214 5682 37266
rect 5966 37214 6018 37266
rect 6638 37214 6690 37266
rect 8094 37214 8146 37266
rect 8766 37214 8818 37266
rect 9886 37214 9938 37266
rect 10558 37214 10610 37266
rect 11006 37214 11058 37266
rect 11566 37214 11618 37266
rect 13582 37214 13634 37266
rect 16606 37214 16658 37266
rect 17390 37214 17442 37266
rect 19070 37214 19122 37266
rect 20190 37214 20242 37266
rect 20526 37214 20578 37266
rect 21086 37214 21138 37266
rect 21534 37214 21586 37266
rect 22430 37214 22482 37266
rect 22990 37214 23042 37266
rect 24334 37214 24386 37266
rect 29486 37214 29538 37266
rect 31390 37214 31442 37266
rect 35758 37214 35810 37266
rect 37550 37214 37602 37266
rect 41470 37214 41522 37266
rect 44942 37214 44994 37266
rect 45838 37214 45890 37266
rect 2494 37102 2546 37154
rect 3502 37102 3554 37154
rect 4734 37102 4786 37154
rect 7086 37102 7138 37154
rect 18286 37102 18338 37154
rect 18622 37102 18674 37154
rect 21870 37102 21922 37154
rect 23438 37102 23490 37154
rect 36206 37102 36258 37154
rect 42030 37102 42082 37154
rect 44158 37102 44210 37154
rect 6750 36990 6802 37042
rect 6974 36990 7026 37042
rect 7422 36990 7474 37042
rect 8206 36990 8258 37042
rect 18622 36990 18674 37042
rect 19070 36990 19122 37042
rect 20862 36990 20914 37042
rect 24222 36990 24274 37042
rect 47966 36990 48018 37042
rect 4478 36822 4530 36874
rect 4582 36822 4634 36874
rect 4686 36822 4738 36874
rect 35198 36822 35250 36874
rect 35302 36822 35354 36874
rect 35406 36822 35458 36874
rect 11566 36654 11618 36706
rect 12798 36654 12850 36706
rect 41694 36654 41746 36706
rect 43822 36654 43874 36706
rect 4622 36568 4674 36620
rect 5070 36542 5122 36594
rect 6302 36542 6354 36594
rect 7422 36542 7474 36594
rect 13694 36542 13746 36594
rect 14590 36542 14642 36594
rect 22654 36542 22706 36594
rect 26910 36542 26962 36594
rect 28030 36542 28082 36594
rect 29822 36542 29874 36594
rect 35422 36542 35474 36594
rect 37774 36542 37826 36594
rect 39902 36542 39954 36594
rect 1822 36430 1874 36482
rect 5966 36430 6018 36482
rect 6638 36430 6690 36482
rect 7534 36430 7586 36482
rect 9998 36430 10050 36482
rect 10782 36430 10834 36482
rect 11006 36430 11058 36482
rect 11118 36430 11170 36482
rect 12910 36430 12962 36482
rect 18510 36430 18562 36482
rect 20750 36430 20802 36482
rect 21422 36430 21474 36482
rect 23214 36430 23266 36482
rect 24110 36430 24162 36482
rect 27470 36430 27522 36482
rect 29262 36430 29314 36482
rect 31614 36430 31666 36482
rect 32622 36430 32674 36482
rect 36318 36430 36370 36482
rect 37102 36430 37154 36482
rect 42478 36430 42530 36482
rect 43150 36430 43202 36482
rect 45054 36430 45106 36482
rect 45614 36430 45666 36482
rect 2494 36318 2546 36370
rect 6190 36318 6242 36370
rect 9774 36318 9826 36370
rect 9886 36318 9938 36370
rect 12798 36318 12850 36370
rect 14926 36318 14978 36370
rect 16382 36318 16434 36370
rect 16606 36318 16658 36370
rect 17054 36318 17106 36370
rect 19518 36318 19570 36370
rect 22318 36318 22370 36370
rect 24782 36318 24834 36370
rect 33294 36318 33346 36370
rect 40350 36318 40402 36370
rect 40686 36318 40738 36370
rect 41358 36318 41410 36370
rect 42254 36318 42306 36370
rect 43038 36318 43090 36370
rect 44158 36318 44210 36370
rect 44830 36318 44882 36370
rect 47406 36318 47458 36370
rect 7310 36206 7362 36258
rect 7758 36206 7810 36258
rect 8542 36206 8594 36258
rect 8878 36206 8930 36258
rect 9438 36206 9490 36258
rect 10446 36206 10498 36258
rect 12350 36206 12402 36258
rect 13806 36206 13858 36258
rect 17166 36206 17218 36258
rect 21758 36206 21810 36258
rect 21870 36206 21922 36258
rect 21982 36206 22034 36258
rect 27246 36206 27298 36258
rect 35758 36206 35810 36258
rect 19838 36038 19890 36090
rect 19942 36038 19994 36090
rect 20046 36038 20098 36090
rect 2270 35870 2322 35922
rect 2382 35870 2434 35922
rect 5630 35870 5682 35922
rect 5854 35870 5906 35922
rect 6862 35870 6914 35922
rect 9774 35870 9826 35922
rect 11678 35870 11730 35922
rect 19294 35870 19346 35922
rect 19966 35870 20018 35922
rect 24334 35870 24386 35922
rect 24558 35870 24610 35922
rect 25342 35870 25394 35922
rect 31278 35870 31330 35922
rect 33294 35870 33346 35922
rect 33742 35870 33794 35922
rect 37886 35870 37938 35922
rect 40126 35870 40178 35922
rect 41246 35870 41298 35922
rect 41694 35870 41746 35922
rect 4846 35758 4898 35810
rect 8094 35758 8146 35810
rect 10222 35758 10274 35810
rect 10894 35758 10946 35810
rect 11342 35758 11394 35810
rect 13470 35758 13522 35810
rect 14702 35758 14754 35810
rect 16046 35758 16098 35810
rect 17614 35758 17666 35810
rect 17726 35758 17778 35810
rect 19406 35758 19458 35810
rect 20526 35758 20578 35810
rect 22990 35758 23042 35810
rect 24222 35758 24274 35810
rect 26014 35758 26066 35810
rect 26350 35758 26402 35810
rect 28702 35758 28754 35810
rect 31950 35758 32002 35810
rect 32398 35758 32450 35810
rect 35310 35758 35362 35810
rect 35534 35758 35586 35810
rect 38782 35758 38834 35810
rect 45726 35758 45778 35810
rect 2494 35646 2546 35698
rect 2942 35646 2994 35698
rect 3390 35646 3442 35698
rect 3726 35646 3778 35698
rect 5742 35646 5794 35698
rect 6078 35646 6130 35698
rect 6414 35646 6466 35698
rect 6638 35646 6690 35698
rect 6974 35646 7026 35698
rect 7646 35646 7698 35698
rect 7870 35646 7922 35698
rect 8430 35646 8482 35698
rect 8654 35646 8706 35698
rect 9662 35646 9714 35698
rect 9998 35646 10050 35698
rect 12014 35646 12066 35698
rect 15038 35646 15090 35698
rect 16382 35646 16434 35698
rect 16718 35646 16770 35698
rect 16158 35590 16210 35642
rect 17950 35646 18002 35698
rect 18286 35646 18338 35698
rect 18734 35646 18786 35698
rect 20414 35646 20466 35698
rect 22206 35646 22258 35698
rect 23550 35646 23602 35698
rect 26238 35646 26290 35698
rect 26686 35646 26738 35698
rect 27358 35646 27410 35698
rect 28030 35646 28082 35698
rect 31614 35646 31666 35698
rect 34078 35646 34130 35698
rect 34638 35646 34690 35698
rect 34974 35646 35026 35698
rect 38222 35646 38274 35698
rect 39006 35646 39058 35698
rect 44606 35646 44658 35698
rect 45054 35646 45106 35698
rect 1934 35534 1986 35586
rect 4510 35534 4562 35586
rect 7982 35534 8034 35586
rect 13694 35534 13746 35586
rect 30830 35534 30882 35586
rect 47854 35534 47906 35586
rect 3278 35422 3330 35474
rect 8990 35422 9042 35474
rect 10782 35422 10834 35474
rect 15598 35422 15650 35474
rect 16830 35422 16882 35474
rect 41246 35422 41298 35474
rect 41806 35422 41858 35474
rect 43598 35422 43650 35474
rect 4478 35254 4530 35306
rect 4582 35254 4634 35306
rect 4686 35254 4738 35306
rect 35198 35254 35250 35306
rect 35302 35254 35354 35306
rect 35406 35254 35458 35306
rect 5854 35086 5906 35138
rect 8094 35086 8146 35138
rect 25902 35086 25954 35138
rect 2270 34974 2322 35026
rect 3950 34974 4002 35026
rect 5070 34974 5122 35026
rect 5630 34974 5682 35026
rect 7646 34974 7698 35026
rect 8654 34974 8706 35026
rect 12014 34974 12066 35026
rect 14254 34974 14306 35026
rect 14926 34974 14978 35026
rect 17278 34974 17330 35026
rect 17726 34974 17778 35026
rect 21422 34974 21474 35026
rect 22878 34974 22930 35026
rect 32062 34974 32114 35026
rect 32846 34974 32898 35026
rect 39790 34974 39842 35026
rect 41806 34974 41858 35026
rect 1822 34862 1874 34914
rect 2718 34862 2770 34914
rect 8206 34862 8258 34914
rect 9438 34862 9490 34914
rect 9662 34862 9714 34914
rect 10110 34862 10162 34914
rect 10894 34862 10946 34914
rect 11342 34862 11394 34914
rect 12238 34862 12290 34914
rect 12910 34862 12962 34914
rect 13806 34862 13858 34914
rect 14030 34862 14082 34914
rect 15262 34862 15314 34914
rect 15710 34862 15762 34914
rect 16382 34862 16434 34914
rect 16606 34862 16658 34914
rect 17950 34862 18002 34914
rect 18510 34862 18562 34914
rect 19070 34862 19122 34914
rect 19630 34862 19682 34914
rect 20078 34862 20130 34914
rect 21310 34862 21362 34914
rect 21758 34862 21810 34914
rect 22094 34862 22146 34914
rect 22990 34862 23042 34914
rect 26126 34862 26178 34914
rect 26910 34862 26962 34914
rect 29150 34862 29202 34914
rect 33518 34862 33570 34914
rect 34638 34862 34690 34914
rect 37550 34862 37602 34914
rect 41134 34862 41186 34914
rect 42814 34862 42866 34914
rect 43150 34862 43202 34914
rect 43934 34862 43986 34914
rect 45838 34862 45890 34914
rect 3278 34750 3330 34802
rect 3390 34750 3442 34802
rect 7198 34750 7250 34802
rect 7422 34750 7474 34802
rect 7534 34750 7586 34802
rect 8990 34750 9042 34802
rect 10222 34750 10274 34802
rect 11678 34750 11730 34802
rect 13582 34750 13634 34802
rect 15150 34750 15202 34802
rect 15486 34750 15538 34802
rect 16046 34750 16098 34802
rect 19518 34750 19570 34802
rect 21534 34750 21586 34802
rect 22542 34750 22594 34802
rect 24670 34750 24722 34802
rect 26462 34750 26514 34802
rect 26686 34750 26738 34802
rect 29934 34750 29986 34802
rect 33406 34750 33458 34802
rect 43822 34750 43874 34802
rect 44942 34750 44994 34802
rect 47182 34750 47234 34802
rect 2942 34638 2994 34690
rect 3614 34638 3666 34690
rect 3838 34638 3890 34690
rect 4734 34638 4786 34690
rect 6190 34638 6242 34690
rect 6638 34638 6690 34690
rect 7758 34638 7810 34690
rect 9214 34638 9266 34690
rect 9326 34638 9378 34690
rect 14702 34638 14754 34690
rect 16382 34638 16434 34690
rect 18958 34638 19010 34690
rect 19182 34638 19234 34690
rect 24110 34638 24162 34690
rect 24782 34638 24834 34690
rect 25006 34638 25058 34690
rect 25342 34638 25394 34690
rect 32510 34638 32562 34690
rect 34862 34638 34914 34690
rect 37102 34638 37154 34690
rect 40910 34638 40962 34690
rect 41470 34638 41522 34690
rect 42366 34638 42418 34690
rect 45278 34638 45330 34690
rect 19838 34470 19890 34522
rect 19942 34470 19994 34522
rect 20046 34470 20098 34522
rect 2606 34302 2658 34354
rect 2942 34302 2994 34354
rect 3614 34302 3666 34354
rect 4734 34302 4786 34354
rect 6414 34302 6466 34354
rect 6750 34302 6802 34354
rect 10446 34302 10498 34354
rect 13246 34302 13298 34354
rect 32062 34302 32114 34354
rect 45166 34302 45218 34354
rect 3502 34190 3554 34242
rect 3726 34190 3778 34242
rect 6862 34190 6914 34242
rect 8206 34190 8258 34242
rect 8766 34190 8818 34242
rect 8878 34190 8930 34242
rect 9550 34190 9602 34242
rect 12462 34190 12514 34242
rect 13582 34190 13634 34242
rect 15598 34190 15650 34242
rect 18958 34190 19010 34242
rect 21086 34190 21138 34242
rect 21646 34190 21698 34242
rect 28814 34190 28866 34242
rect 32398 34190 32450 34242
rect 36094 34190 36146 34242
rect 41694 34190 41746 34242
rect 44158 34190 44210 34242
rect 1710 34078 1762 34130
rect 3390 34078 3442 34130
rect 4174 34078 4226 34130
rect 5070 34078 5122 34130
rect 7982 34078 8034 34130
rect 8318 34078 8370 34130
rect 9998 34078 10050 34130
rect 10222 34078 10274 34130
rect 10670 34078 10722 34130
rect 11454 34078 11506 34130
rect 12014 34078 12066 34130
rect 12574 34078 12626 34130
rect 12798 34078 12850 34130
rect 13022 34078 13074 34130
rect 15038 34078 15090 34130
rect 17950 34078 18002 34130
rect 19182 34078 19234 34130
rect 19854 34078 19906 34130
rect 20750 34078 20802 34130
rect 21870 34078 21922 34130
rect 22990 34078 23042 34130
rect 24110 34078 24162 34130
rect 24334 34078 24386 34130
rect 24782 34078 24834 34130
rect 25230 34078 25282 34130
rect 28590 34078 28642 34130
rect 29374 34078 29426 34130
rect 33182 34078 33234 34130
rect 36878 34078 36930 34130
rect 37438 34078 37490 34130
rect 40910 34078 40962 34130
rect 44606 34078 44658 34130
rect 47966 34078 48018 34130
rect 2270 33966 2322 34018
rect 5518 33966 5570 34018
rect 5966 33966 6018 34018
rect 7310 33966 7362 34018
rect 7758 33966 7810 34018
rect 9662 33966 9714 34018
rect 10558 33966 10610 34018
rect 17390 33966 17442 34018
rect 20526 33966 20578 34018
rect 22318 33966 22370 34018
rect 23102 33966 23154 34018
rect 23774 33966 23826 34018
rect 24222 33966 24274 34018
rect 26014 33966 26066 34018
rect 28142 33966 28194 34018
rect 30270 33966 30322 34018
rect 33518 33966 33570 34018
rect 33966 33966 34018 34018
rect 38110 33966 38162 34018
rect 40238 33966 40290 34018
rect 43822 33966 43874 34018
rect 7198 33854 7250 33906
rect 7870 33854 7922 33906
rect 8878 33854 8930 33906
rect 46286 33854 46338 33906
rect 4478 33686 4530 33738
rect 4582 33686 4634 33738
rect 4686 33686 4738 33738
rect 35198 33686 35250 33738
rect 35302 33686 35354 33738
rect 35406 33686 35458 33738
rect 3838 33518 3890 33570
rect 34862 33518 34914 33570
rect 3614 33406 3666 33458
rect 4174 33406 4226 33458
rect 9886 33406 9938 33458
rect 17726 33406 17778 33458
rect 19742 33406 19794 33458
rect 21310 33406 21362 33458
rect 24334 33406 24386 33458
rect 29934 33406 29986 33458
rect 32062 33406 32114 33458
rect 33406 33406 33458 33458
rect 45054 33406 45106 33458
rect 46062 33406 46114 33458
rect 48190 33406 48242 33458
rect 2830 33294 2882 33346
rect 3278 33294 3330 33346
rect 4846 33294 4898 33346
rect 6638 33294 6690 33346
rect 7534 33294 7586 33346
rect 8542 33294 8594 33346
rect 9998 33294 10050 33346
rect 10334 33294 10386 33346
rect 11118 33294 11170 33346
rect 11790 33294 11842 33346
rect 12350 33294 12402 33346
rect 14030 33294 14082 33346
rect 15710 33294 15762 33346
rect 16270 33294 16322 33346
rect 16830 33294 16882 33346
rect 18510 33294 18562 33346
rect 19294 33294 19346 33346
rect 21758 33294 21810 33346
rect 22206 33294 22258 33346
rect 23102 33294 23154 33346
rect 23214 33294 23266 33346
rect 23662 33294 23714 33346
rect 23886 33294 23938 33346
rect 26350 33294 26402 33346
rect 29262 33294 29314 33346
rect 32958 33294 33010 33346
rect 35198 33294 35250 33346
rect 35758 33294 35810 33346
rect 37550 33294 37602 33346
rect 40686 33294 40738 33346
rect 41694 33294 41746 33346
rect 45390 33294 45442 33346
rect 1710 33182 1762 33234
rect 6526 33182 6578 33234
rect 9550 33182 9602 33234
rect 11566 33182 11618 33234
rect 2046 33070 2098 33122
rect 4510 33070 4562 33122
rect 8094 33070 8146 33122
rect 8766 33070 8818 33122
rect 11678 33070 11730 33122
rect 12014 33070 12066 33122
rect 12238 33126 12290 33178
rect 12910 33182 12962 33234
rect 14142 33182 14194 33234
rect 14814 33182 14866 33234
rect 15598 33182 15650 33234
rect 24222 33182 24274 33234
rect 26014 33182 26066 33234
rect 32398 33182 32450 33234
rect 35982 33182 36034 33234
rect 39342 33182 39394 33234
rect 43486 33182 43538 33234
rect 12574 33070 12626 33122
rect 12798 33070 12850 33122
rect 13694 33070 13746 33122
rect 22990 33070 23042 33122
rect 24446 33070 24498 33122
rect 24894 33070 24946 33122
rect 25342 33070 25394 33122
rect 28590 33070 28642 33122
rect 37214 33070 37266 33122
rect 40462 33070 40514 33122
rect 19838 32902 19890 32954
rect 19942 32902 19994 32954
rect 20046 32902 20098 32954
rect 4510 32734 4562 32786
rect 4734 32734 4786 32786
rect 6190 32734 6242 32786
rect 6302 32734 6354 32786
rect 7646 32734 7698 32786
rect 8094 32734 8146 32786
rect 15710 32734 15762 32786
rect 16718 32734 16770 32786
rect 18958 32734 19010 32786
rect 22766 32734 22818 32786
rect 31166 32734 31218 32786
rect 40238 32734 40290 32786
rect 42254 32734 42306 32786
rect 2830 32622 2882 32674
rect 2942 32622 2994 32674
rect 3054 32622 3106 32674
rect 3950 32622 4002 32674
rect 10334 32622 10386 32674
rect 10670 32622 10722 32674
rect 15822 32622 15874 32674
rect 17502 32622 17554 32674
rect 21982 32622 22034 32674
rect 23214 32622 23266 32674
rect 23886 32622 23938 32674
rect 23998 32622 24050 32674
rect 26238 32622 26290 32674
rect 29822 32622 29874 32674
rect 32286 32622 32338 32674
rect 36990 32622 37042 32674
rect 38670 32622 38722 32674
rect 39118 32622 39170 32674
rect 39678 32622 39730 32674
rect 41358 32622 41410 32674
rect 41582 32622 41634 32674
rect 1822 32510 1874 32562
rect 3838 32510 3890 32562
rect 4174 32510 4226 32562
rect 4398 32510 4450 32562
rect 5742 32510 5794 32562
rect 6414 32510 6466 32562
rect 7870 32510 7922 32562
rect 9998 32510 10050 32562
rect 11790 32510 11842 32562
rect 13246 32510 13298 32562
rect 13918 32510 13970 32562
rect 15038 32510 15090 32562
rect 15486 32510 15538 32562
rect 16158 32510 16210 32562
rect 19630 32510 19682 32562
rect 22094 32510 22146 32562
rect 23326 32510 23378 32562
rect 23438 32510 23490 32562
rect 24222 32510 24274 32562
rect 26574 32510 26626 32562
rect 29598 32510 29650 32562
rect 31502 32510 31554 32562
rect 32174 32510 32226 32562
rect 37326 32510 37378 32562
rect 38446 32510 38498 32562
rect 39902 32510 39954 32562
rect 42702 32510 42754 32562
rect 45614 32510 45666 32562
rect 2270 32398 2322 32450
rect 5070 32398 5122 32450
rect 5630 32398 5682 32450
rect 6974 32398 7026 32450
rect 7310 32398 7362 32450
rect 7758 32398 7810 32450
rect 8990 32398 9042 32450
rect 9662 32398 9714 32450
rect 15150 32398 15202 32450
rect 18062 32398 18114 32450
rect 18398 32398 18450 32450
rect 20190 32398 20242 32450
rect 20974 32398 21026 32450
rect 21310 32398 21362 32450
rect 24558 32398 24610 32450
rect 3502 32286 3554 32338
rect 17390 32286 17442 32338
rect 21982 32286 22034 32338
rect 41918 32286 41970 32338
rect 45054 32286 45106 32338
rect 47070 32286 47122 32338
rect 4478 32118 4530 32170
rect 4582 32118 4634 32170
rect 4686 32118 4738 32170
rect 35198 32118 35250 32170
rect 35302 32118 35354 32170
rect 35406 32118 35458 32170
rect 8878 31950 8930 32002
rect 11454 31950 11506 32002
rect 37662 31950 37714 32002
rect 2158 31838 2210 31890
rect 3390 31838 3442 31890
rect 6638 31838 6690 31890
rect 9102 31838 9154 31890
rect 9326 31838 9378 31890
rect 11902 31838 11954 31890
rect 21422 31838 21474 31890
rect 24222 31838 24274 31890
rect 27918 31838 27970 31890
rect 29934 31838 29986 31890
rect 32062 31838 32114 31890
rect 35310 31838 35362 31890
rect 40014 31838 40066 31890
rect 42142 31838 42194 31890
rect 47742 31838 47794 31890
rect 1710 31726 1762 31778
rect 3726 31726 3778 31778
rect 4062 31726 4114 31778
rect 4510 31726 4562 31778
rect 4846 31726 4898 31778
rect 5854 31726 5906 31778
rect 6414 31726 6466 31778
rect 6974 31726 7026 31778
rect 8206 31726 8258 31778
rect 9550 31726 9602 31778
rect 9774 31726 9826 31778
rect 10222 31726 10274 31778
rect 11006 31726 11058 31778
rect 11566 31726 11618 31778
rect 12126 31726 12178 31778
rect 12686 31726 12738 31778
rect 12798 31726 12850 31778
rect 14702 31726 14754 31778
rect 16718 31726 16770 31778
rect 17166 31726 17218 31778
rect 19630 31726 19682 31778
rect 19854 31726 19906 31778
rect 20190 31726 20242 31778
rect 20302 31726 20354 31778
rect 20414 31726 20466 31778
rect 20638 31726 20690 31778
rect 22206 31726 22258 31778
rect 23102 31726 23154 31778
rect 23214 31726 23266 31778
rect 24558 31726 24610 31778
rect 25006 31726 25058 31778
rect 25790 31726 25842 31778
rect 29150 31726 29202 31778
rect 32398 31726 32450 31778
rect 37998 31726 38050 31778
rect 39342 31726 39394 31778
rect 43150 31726 43202 31778
rect 43822 31726 43874 31778
rect 45726 31726 45778 31778
rect 3278 31614 3330 31666
rect 4734 31614 4786 31666
rect 7534 31614 7586 31666
rect 8542 31614 8594 31666
rect 11454 31614 11506 31666
rect 12462 31614 12514 31666
rect 13918 31614 13970 31666
rect 14254 31614 14306 31666
rect 15150 31614 15202 31666
rect 17726 31614 17778 31666
rect 22430 31614 22482 31666
rect 22766 31614 22818 31666
rect 33182 31614 33234 31666
rect 38222 31614 38274 31666
rect 38782 31614 38834 31666
rect 43262 31614 43314 31666
rect 44158 31614 44210 31666
rect 44830 31614 44882 31666
rect 2830 31502 2882 31554
rect 6638 31502 6690 31554
rect 6862 31502 6914 31554
rect 9662 31502 9714 31554
rect 14590 31502 14642 31554
rect 15262 31502 15314 31554
rect 19294 31502 19346 31554
rect 19406 31502 19458 31554
rect 19518 31502 19570 31554
rect 22990 31502 23042 31554
rect 23774 31502 23826 31554
rect 37214 31502 37266 31554
rect 42702 31502 42754 31554
rect 45166 31502 45218 31554
rect 19838 31334 19890 31386
rect 19942 31334 19994 31386
rect 20046 31334 20098 31386
rect 6078 31166 6130 31218
rect 6526 31166 6578 31218
rect 6750 31166 6802 31218
rect 9550 31166 9602 31218
rect 10782 31166 10834 31218
rect 11118 31166 11170 31218
rect 16718 31166 16770 31218
rect 17726 31166 17778 31218
rect 22990 31166 23042 31218
rect 23550 31166 23602 31218
rect 24558 31166 24610 31218
rect 30718 31166 30770 31218
rect 33406 31166 33458 31218
rect 40014 31166 40066 31218
rect 41134 31166 41186 31218
rect 2382 31054 2434 31106
rect 3726 31054 3778 31106
rect 5294 31054 5346 31106
rect 7086 31054 7138 31106
rect 8878 31054 8930 31106
rect 9774 31054 9826 31106
rect 13022 31054 13074 31106
rect 14030 31054 14082 31106
rect 14366 31054 14418 31106
rect 14590 31054 14642 31106
rect 15598 31054 15650 31106
rect 22654 31054 22706 31106
rect 29374 31054 29426 31106
rect 31390 31054 31442 31106
rect 31614 31054 31666 31106
rect 34862 31054 34914 31106
rect 35422 31054 35474 31106
rect 36654 31054 36706 31106
rect 41694 31054 41746 31106
rect 42254 31054 42306 31106
rect 44942 31054 44994 31106
rect 46062 31054 46114 31106
rect 47406 31054 47458 31106
rect 47966 31054 48018 31106
rect 4846 30942 4898 30994
rect 5854 30942 5906 30994
rect 6414 30942 6466 30994
rect 7982 30942 8034 30994
rect 9550 30942 9602 30994
rect 9998 30942 10050 30994
rect 10110 30942 10162 30994
rect 11566 30942 11618 30994
rect 11902 30942 11954 30994
rect 14478 30942 14530 30994
rect 15486 30942 15538 30994
rect 16158 30942 16210 30994
rect 16606 30942 16658 30994
rect 17950 30942 18002 30994
rect 18958 30942 19010 30994
rect 21534 30942 21586 30994
rect 21758 30942 21810 30994
rect 24446 30942 24498 30994
rect 24782 30942 24834 30994
rect 25342 30942 25394 30994
rect 29710 30942 29762 30994
rect 31054 30942 31106 30994
rect 33742 30942 33794 30994
rect 34302 30942 34354 30994
rect 34638 30942 34690 30994
rect 35982 30942 36034 30994
rect 40238 30942 40290 30994
rect 41470 30942 41522 30994
rect 45614 30942 45666 30994
rect 46398 30942 46450 30994
rect 46846 30942 46898 30994
rect 1934 30830 1986 30882
rect 3950 30830 4002 30882
rect 4958 30830 5010 30882
rect 8206 30830 8258 30882
rect 8430 30830 8482 30882
rect 19518 30830 19570 30882
rect 21310 30830 21362 30882
rect 23998 30830 24050 30882
rect 26014 30830 26066 30882
rect 28142 30830 28194 30882
rect 38782 30830 38834 30882
rect 42814 30830 42866 30882
rect 6974 30718 7026 30770
rect 7310 30718 7362 30770
rect 7758 30718 7810 30770
rect 13694 30718 13746 30770
rect 13806 30718 13858 30770
rect 47182 30718 47234 30770
rect 4478 30550 4530 30602
rect 4582 30550 4634 30602
rect 4686 30550 4738 30602
rect 35198 30550 35250 30602
rect 35302 30550 35354 30602
rect 35406 30550 35458 30602
rect 12574 30382 12626 30434
rect 19630 30382 19682 30434
rect 20302 30382 20354 30434
rect 5070 30270 5122 30322
rect 9438 30270 9490 30322
rect 9662 30270 9714 30322
rect 12910 30270 12962 30322
rect 13582 30270 13634 30322
rect 14366 30270 14418 30322
rect 16382 30270 16434 30322
rect 17502 30270 17554 30322
rect 19406 30270 19458 30322
rect 20638 30270 20690 30322
rect 21758 30270 21810 30322
rect 34862 30270 34914 30322
rect 39902 30270 39954 30322
rect 46062 30270 46114 30322
rect 48190 30270 48242 30322
rect 4286 30158 4338 30210
rect 6414 30158 6466 30210
rect 7870 30158 7922 30210
rect 8654 30158 8706 30210
rect 8990 30158 9042 30210
rect 10558 30158 10610 30210
rect 11230 30158 11282 30210
rect 11902 30158 11954 30210
rect 13470 30158 13522 30210
rect 13918 30158 13970 30210
rect 15038 30158 15090 30210
rect 15710 30158 15762 30210
rect 16270 30158 16322 30210
rect 17166 30158 17218 30210
rect 18958 30158 19010 30210
rect 19966 30158 20018 30210
rect 20526 30158 20578 30210
rect 20750 30158 20802 30210
rect 21870 30158 21922 30210
rect 22206 30158 22258 30210
rect 22430 30158 22482 30210
rect 22766 30158 22818 30210
rect 23214 30158 23266 30210
rect 24110 30158 24162 30210
rect 24558 30158 24610 30210
rect 35646 30158 35698 30210
rect 37102 30158 37154 30210
rect 45390 30158 45442 30210
rect 2494 30046 2546 30098
rect 5966 30046 6018 30098
rect 7646 30046 7698 30098
rect 8766 30046 8818 30098
rect 11006 30046 11058 30098
rect 13806 30046 13858 30098
rect 14478 30046 14530 30098
rect 14814 30046 14866 30098
rect 16046 30046 16098 30098
rect 16494 30046 16546 30098
rect 21646 30046 21698 30098
rect 23438 30046 23490 30098
rect 23774 30046 23826 30098
rect 26798 30046 26850 30098
rect 30158 30046 30210 30098
rect 35422 30046 35474 30098
rect 37774 30046 37826 30098
rect 41246 30046 41298 30098
rect 8206 29934 8258 29986
rect 10334 29934 10386 29986
rect 10894 29934 10946 29986
rect 12126 29934 12178 29986
rect 12798 29934 12850 29986
rect 15374 29934 15426 29986
rect 15598 29934 15650 29986
rect 16606 29934 16658 29986
rect 18062 29934 18114 29986
rect 18398 29934 18450 29986
rect 19406 29934 19458 29986
rect 21422 29934 21474 29986
rect 22654 29934 22706 29986
rect 26910 29934 26962 29986
rect 27134 29934 27186 29986
rect 29598 29934 29650 29986
rect 34078 29934 34130 29986
rect 34526 29934 34578 29986
rect 41582 29934 41634 29986
rect 44942 29934 44994 29986
rect 19838 29766 19890 29818
rect 19942 29766 19994 29818
rect 20046 29766 20098 29818
rect 9662 29598 9714 29650
rect 11454 29598 11506 29650
rect 11902 29598 11954 29650
rect 18286 29598 18338 29650
rect 19070 29598 19122 29650
rect 19406 29598 19458 29650
rect 20526 29598 20578 29650
rect 22766 29598 22818 29650
rect 26574 29598 26626 29650
rect 26798 29598 26850 29650
rect 37774 29598 37826 29650
rect 2046 29486 2098 29538
rect 2718 29486 2770 29538
rect 8318 29486 8370 29538
rect 8878 29486 8930 29538
rect 11118 29486 11170 29538
rect 13022 29486 13074 29538
rect 14254 29486 14306 29538
rect 16046 29486 16098 29538
rect 16382 29486 16434 29538
rect 16830 29486 16882 29538
rect 19518 29486 19570 29538
rect 22654 29486 22706 29538
rect 24110 29486 24162 29538
rect 26798 29486 26850 29538
rect 27022 29486 27074 29538
rect 27694 29486 27746 29538
rect 29150 29486 29202 29538
rect 39342 29486 39394 29538
rect 41694 29486 41746 29538
rect 45278 29486 45330 29538
rect 1710 29374 1762 29426
rect 2494 29374 2546 29426
rect 2606 29374 2658 29426
rect 3166 29374 3218 29426
rect 3502 29374 3554 29426
rect 3838 29374 3890 29426
rect 5406 29374 5458 29426
rect 6750 29374 6802 29426
rect 8654 29374 8706 29426
rect 10782 29374 10834 29426
rect 12462 29374 12514 29426
rect 14030 29374 14082 29426
rect 17390 29374 17442 29426
rect 17950 29374 18002 29426
rect 18510 29374 18562 29426
rect 21758 29374 21810 29426
rect 23774 29374 23826 29426
rect 26574 29374 26626 29426
rect 28478 29374 28530 29426
rect 35982 29374 36034 29426
rect 37550 29374 37602 29426
rect 38222 29374 38274 29426
rect 38558 29374 38610 29426
rect 39118 29374 39170 29426
rect 41022 29374 41074 29426
rect 45054 29374 45106 29426
rect 45614 29374 45666 29426
rect 6078 29262 6130 29314
rect 6974 29262 7026 29314
rect 8430 29262 8482 29314
rect 11790 29262 11842 29314
rect 15038 29262 15090 29314
rect 18958 29262 19010 29314
rect 20078 29262 20130 29314
rect 21310 29262 21362 29314
rect 31278 29262 31330 29314
rect 33070 29262 33122 29314
rect 35198 29262 35250 29314
rect 39902 29262 39954 29314
rect 43822 29262 43874 29314
rect 10110 29150 10162 29202
rect 10334 29150 10386 29202
rect 10558 29150 10610 29202
rect 16718 29150 16770 29202
rect 47966 29150 48018 29202
rect 4478 28982 4530 29034
rect 4582 28982 4634 29034
rect 4686 28982 4738 29034
rect 35198 28982 35250 29034
rect 35302 28982 35354 29034
rect 35406 28982 35458 29034
rect 5742 28814 5794 28866
rect 7198 28814 7250 28866
rect 10446 28814 10498 28866
rect 2718 28702 2770 28754
rect 25902 28814 25954 28866
rect 30718 28814 30770 28866
rect 35422 28814 35474 28866
rect 41134 28814 41186 28866
rect 41470 28814 41522 28866
rect 43822 28814 43874 28866
rect 7534 28702 7586 28754
rect 12462 28702 12514 28754
rect 13694 28702 13746 28754
rect 17838 28702 17890 28754
rect 19742 28702 19794 28754
rect 20414 28702 20466 28754
rect 29598 28702 29650 28754
rect 30270 28702 30322 28754
rect 40686 28702 40738 28754
rect 44158 28702 44210 28754
rect 47854 28702 47906 28754
rect 2158 28590 2210 28642
rect 3054 28590 3106 28642
rect 4286 28590 4338 28642
rect 4846 28590 4898 28642
rect 5630 28590 5682 28642
rect 6638 28590 6690 28642
rect 6974 28590 7026 28642
rect 7534 28590 7586 28642
rect 7982 28590 8034 28642
rect 8094 28590 8146 28642
rect 9774 28590 9826 28642
rect 9998 28590 10050 28642
rect 10558 28590 10610 28642
rect 11230 28590 11282 28642
rect 11790 28590 11842 28642
rect 12350 28590 12402 28642
rect 16046 28590 16098 28642
rect 17054 28590 17106 28642
rect 17390 28590 17442 28642
rect 18958 28590 19010 28642
rect 20190 28590 20242 28642
rect 23102 28590 23154 28642
rect 23438 28590 23490 28642
rect 25790 28590 25842 28642
rect 26238 28590 26290 28642
rect 29262 28590 29314 28642
rect 31054 28590 31106 28642
rect 31838 28590 31890 28642
rect 33182 28590 33234 28642
rect 35870 28590 35922 28642
rect 37774 28590 37826 28642
rect 41918 28590 41970 28642
rect 45054 28590 45106 28642
rect 45614 28590 45666 28642
rect 3390 28478 3442 28530
rect 4398 28478 4450 28530
rect 6190 28478 6242 28530
rect 6414 28478 6466 28530
rect 8206 28478 8258 28530
rect 8766 28478 8818 28530
rect 12574 28478 12626 28530
rect 16718 28478 16770 28530
rect 20750 28478 20802 28530
rect 21310 28478 21362 28530
rect 23998 28478 24050 28530
rect 26462 28478 26514 28530
rect 26910 28478 26962 28530
rect 27470 28478 27522 28530
rect 31614 28478 31666 28530
rect 33406 28478 33458 28530
rect 36206 28478 36258 28530
rect 37550 28478 37602 28530
rect 39342 28478 39394 28530
rect 42254 28478 42306 28530
rect 43262 28478 43314 28530
rect 43486 28478 43538 28530
rect 1934 28366 1986 28418
rect 4958 28366 5010 28418
rect 6302 28366 6354 28418
rect 11678 28366 11730 28418
rect 18398 28366 18450 28418
rect 21534 28366 21586 28418
rect 35086 28366 35138 28418
rect 39678 28366 39730 28418
rect 44830 28366 44882 28418
rect 19838 28198 19890 28250
rect 19942 28198 19994 28250
rect 20046 28198 20098 28250
rect 5182 28030 5234 28082
rect 7758 28030 7810 28082
rect 8430 28030 8482 28082
rect 9438 28030 9490 28082
rect 11566 28030 11618 28082
rect 15038 28030 15090 28082
rect 17502 28030 17554 28082
rect 17838 28030 17890 28082
rect 26574 28030 26626 28082
rect 26686 28030 26738 28082
rect 41582 28030 41634 28082
rect 42254 28030 42306 28082
rect 46062 28030 46114 28082
rect 47630 28030 47682 28082
rect 8094 27918 8146 27970
rect 11230 27918 11282 27970
rect 15710 27918 15762 27970
rect 16606 27918 16658 27970
rect 22206 27918 22258 27970
rect 27134 27918 27186 27970
rect 43374 27918 43426 27970
rect 46622 27918 46674 27970
rect 1822 27806 1874 27858
rect 4958 27806 5010 27858
rect 5630 27806 5682 27858
rect 6638 27806 6690 27858
rect 7086 27806 7138 27858
rect 7198 27806 7250 27858
rect 10110 27806 10162 27858
rect 10446 27806 10498 27858
rect 12462 27806 12514 27858
rect 14814 27806 14866 27858
rect 15374 27806 15426 27858
rect 18398 27806 18450 27858
rect 21310 27806 21362 27858
rect 22766 27806 22818 27858
rect 22990 27806 23042 27858
rect 23438 27806 23490 27858
rect 24446 27806 24498 27858
rect 27358 27806 27410 27858
rect 29486 27806 29538 27858
rect 33630 27806 33682 27858
rect 37438 27806 37490 27858
rect 41246 27806 41298 27858
rect 42702 27806 42754 27858
rect 46510 27806 46562 27858
rect 47294 27806 47346 27858
rect 2494 27694 2546 27746
rect 4622 27694 4674 27746
rect 5070 27694 5122 27746
rect 6302 27694 6354 27746
rect 8990 27694 9042 27746
rect 9774 27694 9826 27746
rect 13806 27694 13858 27746
rect 14926 27694 14978 27746
rect 16046 27694 16098 27746
rect 18846 27694 18898 27746
rect 20302 27694 20354 27746
rect 23998 27694 24050 27746
rect 30270 27694 30322 27746
rect 32398 27694 32450 27746
rect 34414 27694 34466 27746
rect 36542 27694 36594 27746
rect 38222 27694 38274 27746
rect 40350 27694 40402 27746
rect 45502 27694 45554 27746
rect 15822 27582 15874 27634
rect 16158 27582 16210 27634
rect 16718 27582 16770 27634
rect 26462 27582 26514 27634
rect 4478 27414 4530 27466
rect 4582 27414 4634 27466
rect 4686 27414 4738 27466
rect 35198 27414 35250 27466
rect 35302 27414 35354 27466
rect 35406 27414 35458 27466
rect 12238 27246 12290 27298
rect 31390 27246 31442 27298
rect 2270 27134 2322 27186
rect 5742 27134 5794 27186
rect 6862 27134 6914 27186
rect 9550 27134 9602 27186
rect 10222 27134 10274 27186
rect 11118 27134 11170 27186
rect 13470 27134 13522 27186
rect 15038 27134 15090 27186
rect 20750 27134 20802 27186
rect 23886 27134 23938 27186
rect 26462 27134 26514 27186
rect 28590 27134 28642 27186
rect 38334 27134 38386 27186
rect 40014 27134 40066 27186
rect 46062 27134 46114 27186
rect 48190 27134 48242 27186
rect 2942 27022 2994 27074
rect 4174 27022 4226 27074
rect 4510 27022 4562 27074
rect 5182 27022 5234 27074
rect 6302 27022 6354 27074
rect 7870 27022 7922 27074
rect 8318 27022 8370 27074
rect 8654 27022 8706 27074
rect 9102 27022 9154 27074
rect 10558 27022 10610 27074
rect 11790 27022 11842 27074
rect 11902 27022 11954 27074
rect 12910 27022 12962 27074
rect 13694 27022 13746 27074
rect 13918 27022 13970 27074
rect 15374 27022 15426 27074
rect 15822 27022 15874 27074
rect 18062 27022 18114 27074
rect 19182 27022 19234 27074
rect 20190 27022 20242 27074
rect 20526 27022 20578 27074
rect 22990 27022 23042 27074
rect 23326 27022 23378 27074
rect 25678 27022 25730 27074
rect 34750 27022 34802 27074
rect 37774 27022 37826 27074
rect 45390 27022 45442 27074
rect 1710 26910 1762 26962
rect 3166 26910 3218 26962
rect 3502 26910 3554 26962
rect 3726 26910 3778 26962
rect 4734 26910 4786 26962
rect 5854 26910 5906 26962
rect 5966 26910 6018 26962
rect 6974 26910 7026 26962
rect 7198 26910 7250 26962
rect 8094 26910 8146 26962
rect 12574 26910 12626 26962
rect 15710 26910 15762 26962
rect 16494 26910 16546 26962
rect 16830 26910 16882 26962
rect 17166 26910 17218 26962
rect 17502 26910 17554 26962
rect 17838 26910 17890 26962
rect 18734 26910 18786 26962
rect 21422 26910 21474 26962
rect 21758 26910 21810 26962
rect 22094 26910 22146 26962
rect 22430 26910 22482 26962
rect 24558 26910 24610 26962
rect 30270 26910 30322 26962
rect 30606 26910 30658 26962
rect 31054 26910 31106 26962
rect 31614 26910 31666 26962
rect 32174 26910 32226 26962
rect 34414 26910 34466 26962
rect 39678 26910 39730 26962
rect 39902 26910 39954 26962
rect 43934 26910 43986 26962
rect 3614 26798 3666 26850
rect 4622 26798 4674 26850
rect 5630 26798 5682 26850
rect 6750 26798 6802 26850
rect 11566 26798 11618 26850
rect 11678 26798 11730 26850
rect 15486 26798 15538 26850
rect 18398 26798 18450 26850
rect 18622 26798 18674 26850
rect 19406 26798 19458 26850
rect 24222 26798 24274 26850
rect 44270 26798 44322 26850
rect 19838 26630 19890 26682
rect 19942 26630 19994 26682
rect 20046 26630 20098 26682
rect 2158 26462 2210 26514
rect 4174 26462 4226 26514
rect 4734 26462 4786 26514
rect 4958 26462 5010 26514
rect 5518 26462 5570 26514
rect 8990 26462 9042 26514
rect 10558 26462 10610 26514
rect 11790 26462 11842 26514
rect 12910 26462 12962 26514
rect 15822 26462 15874 26514
rect 16830 26462 16882 26514
rect 22430 26462 22482 26514
rect 26686 26462 26738 26514
rect 39678 26462 39730 26514
rect 5070 26350 5122 26402
rect 7870 26350 7922 26402
rect 11342 26350 11394 26402
rect 12350 26350 12402 26402
rect 16046 26350 16098 26402
rect 17614 26350 17666 26402
rect 18062 26350 18114 26402
rect 18286 26350 18338 26402
rect 18510 26350 18562 26402
rect 19966 26350 20018 26402
rect 24558 26350 24610 26402
rect 27806 26350 27858 26402
rect 2382 26238 2434 26290
rect 3390 26238 3442 26290
rect 4398 26238 4450 26290
rect 5854 26238 5906 26290
rect 6974 26238 7026 26290
rect 8094 26238 8146 26290
rect 8654 26238 8706 26290
rect 9550 26238 9602 26290
rect 9886 26238 9938 26290
rect 9998 26238 10050 26290
rect 10110 26238 10162 26290
rect 10782 26238 10834 26290
rect 11566 26238 11618 26290
rect 11902 26238 11954 26290
rect 12574 26238 12626 26290
rect 13806 26238 13858 26290
rect 14926 26238 14978 26290
rect 15150 26238 15202 26290
rect 15486 26238 15538 26290
rect 15598 26238 15650 26290
rect 16158 26238 16210 26290
rect 17502 26238 17554 26290
rect 17838 26238 17890 26290
rect 19294 26238 19346 26290
rect 22654 26238 22706 26290
rect 24446 26238 24498 26290
rect 27470 26238 27522 26290
rect 33070 26238 33122 26290
rect 39230 26238 39282 26290
rect 39454 26238 39506 26290
rect 39790 26238 39842 26290
rect 40014 26238 40066 26290
rect 44718 26238 44770 26290
rect 45614 26238 45666 26290
rect 2942 26126 2994 26178
rect 3838 26126 3890 26178
rect 7758 26126 7810 26178
rect 11790 26126 11842 26178
rect 13694 26126 13746 26178
rect 14254 26126 14306 26178
rect 15262 26126 15314 26178
rect 22094 26126 22146 26178
rect 33854 26126 33906 26178
rect 35982 26126 36034 26178
rect 36318 26126 36370 26178
rect 38446 26126 38498 26178
rect 40910 26126 40962 26178
rect 41918 26126 41970 26178
rect 44046 26126 44098 26178
rect 6078 26014 6130 26066
rect 6302 26014 6354 26066
rect 6750 26014 6802 26066
rect 10446 26014 10498 26066
rect 18398 26014 18450 26066
rect 23438 26014 23490 26066
rect 23774 26014 23826 26066
rect 27022 26014 27074 26066
rect 41134 26014 41186 26066
rect 41470 26014 41522 26066
rect 47966 26014 48018 26066
rect 4478 25846 4530 25898
rect 4582 25846 4634 25898
rect 4686 25846 4738 25898
rect 35198 25846 35250 25898
rect 35302 25846 35354 25898
rect 35406 25846 35458 25898
rect 8878 25678 8930 25730
rect 13470 25678 13522 25730
rect 2494 25566 2546 25618
rect 4622 25566 4674 25618
rect 5182 25566 5234 25618
rect 7310 25566 7362 25618
rect 12462 25566 12514 25618
rect 13582 25566 13634 25618
rect 14254 25566 14306 25618
rect 16382 25566 16434 25618
rect 18174 25566 18226 25618
rect 22318 25566 22370 25618
rect 23998 25566 24050 25618
rect 26126 25566 26178 25618
rect 32174 25566 32226 25618
rect 35198 25566 35250 25618
rect 37662 25566 37714 25618
rect 39454 25566 39506 25618
rect 40574 25566 40626 25618
rect 48190 25566 48242 25618
rect 1822 25454 1874 25506
rect 7198 25454 7250 25506
rect 7870 25454 7922 25506
rect 8094 25454 8146 25506
rect 10110 25454 10162 25506
rect 10446 25454 10498 25506
rect 10670 25454 10722 25506
rect 12014 25454 12066 25506
rect 12798 25454 12850 25506
rect 17054 25454 17106 25506
rect 17838 25454 17890 25506
rect 18734 25454 18786 25506
rect 19854 25454 19906 25506
rect 20638 25454 20690 25506
rect 21422 25454 21474 25506
rect 23214 25454 23266 25506
rect 29374 25454 29426 25506
rect 35646 25454 35698 25506
rect 38110 25454 38162 25506
rect 38334 25454 38386 25506
rect 38670 25454 38722 25506
rect 39566 25454 39618 25506
rect 39790 25454 39842 25506
rect 40014 25454 40066 25506
rect 40238 25454 40290 25506
rect 40798 25454 40850 25506
rect 41806 25454 41858 25506
rect 42366 25454 42418 25506
rect 43038 25454 43090 25506
rect 43598 25454 43650 25506
rect 45390 25454 45442 25506
rect 9774 25342 9826 25394
rect 11902 25342 11954 25394
rect 12462 25342 12514 25394
rect 19518 25342 19570 25394
rect 20414 25342 20466 25394
rect 26462 25342 26514 25394
rect 30046 25342 30098 25394
rect 33742 25342 33794 25394
rect 34078 25342 34130 25394
rect 37550 25342 37602 25394
rect 37774 25342 37826 25394
rect 39342 25342 39394 25394
rect 40686 25342 40738 25394
rect 41358 25342 41410 25394
rect 43486 25342 43538 25394
rect 46062 25342 46114 25394
rect 10110 25230 10162 25282
rect 17614 25230 17666 25282
rect 18174 25230 18226 25282
rect 18398 25230 18450 25282
rect 18846 25230 18898 25282
rect 19070 25230 19122 25282
rect 26798 25230 26850 25282
rect 38446 25230 38498 25282
rect 43374 25230 43426 25282
rect 19838 25062 19890 25114
rect 19942 25062 19994 25114
rect 20046 25062 20098 25114
rect 1710 24894 1762 24946
rect 3838 24894 3890 24946
rect 13246 24894 13298 24946
rect 15486 24894 15538 24946
rect 16718 24894 16770 24946
rect 17614 24894 17666 24946
rect 18174 24894 18226 24946
rect 19070 24894 19122 24946
rect 19406 24894 19458 24946
rect 30942 24894 30994 24946
rect 31278 24894 31330 24946
rect 34526 24894 34578 24946
rect 39230 24894 39282 24946
rect 43262 24894 43314 24946
rect 44606 24894 44658 24946
rect 45278 24894 45330 24946
rect 2046 24782 2098 24834
rect 7870 24782 7922 24834
rect 10782 24782 10834 24834
rect 11342 24782 11394 24834
rect 12238 24782 12290 24834
rect 13134 24782 13186 24834
rect 15038 24782 15090 24834
rect 16158 24782 16210 24834
rect 21310 24782 21362 24834
rect 22990 24782 23042 24834
rect 28702 24782 28754 24834
rect 35422 24782 35474 24834
rect 44942 24782 44994 24834
rect 2382 24670 2434 24722
rect 2942 24670 2994 24722
rect 5630 24670 5682 24722
rect 6974 24670 7026 24722
rect 7758 24670 7810 24722
rect 8318 24670 8370 24722
rect 8990 24670 9042 24722
rect 9550 24670 9602 24722
rect 10894 24670 10946 24722
rect 11454 24670 11506 24722
rect 12462 24670 12514 24722
rect 13022 24670 13074 24722
rect 13918 24670 13970 24722
rect 16046 24670 16098 24722
rect 16382 24670 16434 24722
rect 16606 24670 16658 24722
rect 16942 24670 16994 24722
rect 17838 24670 17890 24722
rect 20414 24670 20466 24722
rect 20750 24670 20802 24722
rect 23326 24670 23378 24722
rect 24670 24670 24722 24722
rect 25230 24670 25282 24722
rect 30830 24670 30882 24722
rect 31054 24670 31106 24722
rect 35646 24670 35698 24722
rect 38670 24670 38722 24722
rect 42478 24670 42530 24722
rect 42702 24670 42754 24722
rect 44382 24670 44434 24722
rect 48078 24670 48130 24722
rect 4174 24558 4226 24610
rect 4622 24558 4674 24610
rect 5070 24558 5122 24610
rect 6078 24558 6130 24610
rect 6302 24558 6354 24610
rect 6750 24558 6802 24610
rect 11678 24558 11730 24610
rect 21870 24558 21922 24610
rect 38446 24558 38498 24610
rect 39678 24558 39730 24610
rect 40238 24558 40290 24610
rect 41022 24558 41074 24610
rect 43374 24558 43426 24610
rect 46958 24558 47010 24610
rect 4174 24446 4226 24498
rect 5070 24446 5122 24498
rect 6526 24446 6578 24498
rect 7422 24446 7474 24498
rect 34862 24446 34914 24498
rect 38894 24446 38946 24498
rect 39678 24446 39730 24498
rect 40238 24446 40290 24498
rect 42142 24446 42194 24498
rect 43038 24446 43090 24498
rect 4478 24278 4530 24330
rect 4582 24278 4634 24330
rect 4686 24278 4738 24330
rect 35198 24278 35250 24330
rect 35302 24278 35354 24330
rect 35406 24278 35458 24330
rect 12798 24110 12850 24162
rect 13022 24110 13074 24162
rect 19854 24110 19906 24162
rect 2494 23998 2546 24050
rect 4622 23998 4674 24050
rect 5182 23998 5234 24050
rect 11230 23998 11282 24050
rect 12574 23998 12626 24050
rect 13022 23998 13074 24050
rect 23214 23998 23266 24050
rect 25342 23998 25394 24050
rect 25678 23998 25730 24050
rect 27806 23998 27858 24050
rect 29262 23998 29314 24050
rect 33742 23998 33794 24050
rect 43710 23998 43762 24050
rect 47966 23998 48018 24050
rect 1822 23886 1874 23938
rect 6750 23886 6802 23938
rect 8878 23886 8930 23938
rect 13694 23886 13746 23938
rect 14478 23886 14530 23938
rect 15262 23886 15314 23938
rect 16046 23886 16098 23938
rect 16830 23886 16882 23938
rect 17278 23886 17330 23938
rect 18062 23886 18114 23938
rect 20302 23886 20354 23938
rect 22430 23886 22482 23938
rect 28590 23886 28642 23938
rect 29038 23886 29090 23938
rect 29486 23886 29538 23938
rect 29598 23886 29650 23938
rect 30606 23886 30658 23938
rect 30830 23886 30882 23938
rect 37102 23886 37154 23938
rect 38894 23886 38946 23938
rect 39902 23886 39954 23938
rect 40462 23886 40514 23938
rect 41694 23886 41746 23938
rect 42590 23886 42642 23938
rect 42926 23886 42978 23938
rect 43262 23886 43314 23938
rect 45166 23886 45218 23938
rect 45614 23886 45666 23938
rect 6862 23774 6914 23826
rect 9998 23774 10050 23826
rect 13582 23774 13634 23826
rect 14254 23774 14306 23826
rect 16158 23774 16210 23826
rect 17838 23774 17890 23826
rect 18286 23774 18338 23826
rect 19070 23774 19122 23826
rect 19518 23774 19570 23826
rect 20638 23774 20690 23826
rect 30270 23774 30322 23826
rect 30382 23774 30434 23826
rect 31614 23774 31666 23826
rect 35982 23774 36034 23826
rect 37326 23774 37378 23826
rect 37998 23774 38050 23826
rect 40014 23774 40066 23826
rect 40686 23774 40738 23826
rect 43598 23774 43650 23826
rect 43822 23774 43874 23826
rect 44942 23774 44994 23826
rect 6078 23662 6130 23714
rect 6526 23662 6578 23714
rect 8430 23662 8482 23714
rect 11678 23662 11730 23714
rect 14366 23662 14418 23714
rect 17390 23662 17442 23714
rect 18398 23662 18450 23714
rect 18734 23662 18786 23714
rect 35646 23662 35698 23714
rect 37662 23662 37714 23714
rect 38334 23662 38386 23714
rect 40574 23662 40626 23714
rect 42926 23662 42978 23714
rect 19838 23494 19890 23546
rect 19942 23494 19994 23546
rect 20046 23494 20098 23546
rect 1710 23326 1762 23378
rect 2942 23326 2994 23378
rect 4510 23326 4562 23378
rect 7982 23326 8034 23378
rect 8206 23326 8258 23378
rect 8990 23326 9042 23378
rect 12574 23326 12626 23378
rect 13918 23326 13970 23378
rect 15710 23326 15762 23378
rect 16830 23326 16882 23378
rect 17614 23326 17666 23378
rect 23326 23326 23378 23378
rect 25678 23326 25730 23378
rect 26462 23326 26514 23378
rect 29374 23326 29426 23378
rect 30942 23326 30994 23378
rect 31166 23326 31218 23378
rect 35198 23326 35250 23378
rect 39006 23326 39058 23378
rect 39342 23326 39394 23378
rect 41806 23326 41858 23378
rect 46510 23326 46562 23378
rect 2046 23214 2098 23266
rect 8654 23214 8706 23266
rect 10894 23214 10946 23266
rect 13022 23214 13074 23266
rect 14142 23214 14194 23266
rect 18846 23214 18898 23266
rect 22878 23214 22930 23266
rect 24334 23214 24386 23266
rect 25454 23214 25506 23266
rect 27582 23214 27634 23266
rect 29486 23214 29538 23266
rect 31054 23214 31106 23266
rect 31726 23214 31778 23266
rect 31950 23214 32002 23266
rect 32062 23214 32114 23266
rect 36318 23214 36370 23266
rect 38670 23214 38722 23266
rect 39678 23214 39730 23266
rect 42030 23214 42082 23266
rect 42366 23214 42418 23266
rect 43598 23214 43650 23266
rect 47070 23214 47122 23266
rect 47406 23214 47458 23266
rect 4846 23102 4898 23154
rect 8318 23102 8370 23154
rect 9662 23102 9714 23154
rect 9886 23102 9938 23154
rect 10110 23102 10162 23154
rect 10558 23102 10610 23154
rect 11454 23102 11506 23154
rect 11790 23102 11842 23154
rect 12238 23102 12290 23154
rect 13246 23102 13298 23154
rect 14478 23102 14530 23154
rect 14926 23102 14978 23154
rect 16606 23102 16658 23154
rect 18062 23102 18114 23154
rect 22318 23102 22370 23154
rect 24222 23102 24274 23154
rect 25678 23102 25730 23154
rect 26014 23102 26066 23154
rect 26798 23102 26850 23154
rect 27470 23102 27522 23154
rect 29038 23102 29090 23154
rect 29710 23102 29762 23154
rect 31614 23102 31666 23154
rect 35534 23102 35586 23154
rect 35982 23102 36034 23154
rect 38446 23102 38498 23154
rect 40014 23102 40066 23154
rect 41246 23102 41298 23154
rect 42926 23102 42978 23154
rect 46846 23102 46898 23154
rect 2606 22990 2658 23042
rect 3502 22990 3554 23042
rect 3950 22990 4002 23042
rect 5518 22990 5570 23042
rect 7646 22990 7698 23042
rect 9774 22990 9826 23042
rect 16158 22990 16210 23042
rect 20974 22990 21026 23042
rect 37998 22990 38050 23042
rect 39790 22990 39842 23042
rect 45726 22990 45778 23042
rect 48190 22990 48242 23042
rect 2606 22878 2658 22930
rect 3166 22878 3218 22930
rect 3502 22878 3554 22930
rect 4510 22878 4562 22930
rect 10334 22878 10386 22930
rect 15598 22878 15650 22930
rect 16158 22878 16210 22930
rect 23662 22878 23714 22930
rect 40910 22878 40962 22930
rect 41246 22878 41298 22930
rect 4478 22710 4530 22762
rect 4582 22710 4634 22762
rect 4686 22710 4738 22762
rect 35198 22710 35250 22762
rect 35302 22710 35354 22762
rect 35406 22710 35458 22762
rect 7422 22542 7474 22594
rect 10670 22542 10722 22594
rect 10894 22542 10946 22594
rect 12014 22542 12066 22594
rect 12238 22542 12290 22594
rect 22318 22542 22370 22594
rect 35198 22542 35250 22594
rect 2494 22430 2546 22482
rect 4622 22430 4674 22482
rect 5854 22430 5906 22482
rect 6414 22430 6466 22482
rect 7310 22430 7362 22482
rect 10222 22430 10274 22482
rect 10894 22430 10946 22482
rect 11342 22430 11394 22482
rect 11902 22430 11954 22482
rect 12350 22430 12402 22482
rect 12798 22430 12850 22482
rect 14478 22430 14530 22482
rect 17838 22430 17890 22482
rect 19070 22430 19122 22482
rect 1822 22318 1874 22370
rect 6526 22318 6578 22370
rect 6750 22318 6802 22370
rect 7982 22318 8034 22370
rect 9214 22318 9266 22370
rect 10446 22318 10498 22370
rect 14030 22318 14082 22370
rect 14814 22318 14866 22370
rect 22094 22318 22146 22370
rect 6078 22206 6130 22258
rect 8766 22206 8818 22258
rect 8878 22206 8930 22258
rect 9326 22206 9378 22258
rect 9774 22206 9826 22258
rect 9998 22206 10050 22258
rect 13470 22206 13522 22258
rect 13694 22206 13746 22258
rect 15598 22206 15650 22258
rect 21758 22206 21810 22258
rect 5070 22094 5122 22146
rect 6302 22094 6354 22146
rect 7758 22094 7810 22146
rect 9550 22094 9602 22146
rect 12910 22094 12962 22146
rect 13806 22094 13858 22146
rect 22766 22430 22818 22482
rect 28142 22430 28194 22482
rect 32062 22430 32114 22482
rect 32734 22430 32786 22482
rect 44382 22430 44434 22482
rect 45054 22430 45106 22482
rect 48190 22430 48242 22482
rect 25230 22318 25282 22370
rect 29262 22318 29314 22370
rect 34078 22318 34130 22370
rect 35982 22318 36034 22370
rect 38782 22318 38834 22370
rect 39342 22318 39394 22370
rect 39902 22318 39954 22370
rect 40574 22318 40626 22370
rect 41806 22318 41858 22370
rect 42590 22318 42642 22370
rect 42814 22318 42866 22370
rect 43150 22318 43202 22370
rect 43486 22318 43538 22370
rect 45390 22318 45442 22370
rect 22542 22206 22594 22258
rect 23662 22206 23714 22258
rect 26014 22206 26066 22258
rect 29934 22206 29986 22258
rect 35758 22206 35810 22258
rect 39118 22206 39170 22258
rect 39790 22206 39842 22258
rect 40798 22206 40850 22258
rect 42254 22206 42306 22258
rect 43710 22206 43762 22258
rect 46062 22206 46114 22258
rect 21982 22094 22034 22146
rect 22318 22094 22370 22146
rect 22766 22094 22818 22146
rect 22990 22094 23042 22146
rect 23326 22094 23378 22146
rect 24222 22094 24274 22146
rect 34302 22094 34354 22146
rect 34862 22094 34914 22146
rect 37102 22094 37154 22146
rect 37550 22094 37602 22146
rect 38110 22094 38162 22146
rect 38446 22094 38498 22146
rect 39006 22094 39058 22146
rect 42030 22094 42082 22146
rect 43598 22094 43650 22146
rect 19838 21926 19890 21978
rect 19942 21926 19994 21978
rect 20046 21926 20098 21978
rect 5630 21758 5682 21810
rect 6302 21758 6354 21810
rect 6974 21758 7026 21810
rect 7982 21758 8034 21810
rect 8654 21758 8706 21810
rect 10110 21758 10162 21810
rect 15934 21758 15986 21810
rect 20638 21758 20690 21810
rect 22206 21758 22258 21810
rect 22878 21758 22930 21810
rect 26126 21758 26178 21810
rect 26238 21758 26290 21810
rect 27918 21758 27970 21810
rect 29150 21758 29202 21810
rect 29598 21758 29650 21810
rect 29710 21758 29762 21810
rect 30718 21758 30770 21810
rect 31390 21758 31442 21810
rect 39230 21758 39282 21810
rect 41806 21758 41858 21810
rect 42142 21758 42194 21810
rect 7422 21646 7474 21698
rect 7646 21646 7698 21698
rect 7758 21646 7810 21698
rect 8318 21646 8370 21698
rect 12910 21646 12962 21698
rect 21758 21646 21810 21698
rect 32062 21646 32114 21698
rect 32174 21646 32226 21698
rect 37550 21646 37602 21698
rect 39006 21646 39058 21698
rect 40014 21646 40066 21698
rect 42478 21646 42530 21698
rect 45390 21646 45442 21698
rect 47518 21646 47570 21698
rect 48078 21646 48130 21698
rect 1822 21534 1874 21586
rect 5742 21534 5794 21586
rect 6190 21534 6242 21586
rect 6414 21534 6466 21586
rect 10334 21534 10386 21586
rect 10894 21534 10946 21586
rect 11342 21534 11394 21586
rect 12238 21534 12290 21586
rect 15486 21534 15538 21586
rect 17502 21534 17554 21586
rect 20862 21534 20914 21586
rect 21422 21534 21474 21586
rect 21646 21534 21698 21586
rect 23102 21534 23154 21586
rect 23438 21534 23490 21586
rect 26350 21534 26402 21586
rect 26798 21534 26850 21586
rect 27694 21534 27746 21586
rect 28030 21534 28082 21586
rect 28926 21534 28978 21586
rect 29486 21534 29538 21586
rect 30158 21534 30210 21586
rect 30494 21534 30546 21586
rect 30830 21534 30882 21586
rect 31166 21534 31218 21586
rect 31838 21534 31890 21586
rect 33070 21534 33122 21586
rect 37886 21534 37938 21586
rect 39230 21534 39282 21586
rect 39902 21534 39954 21586
rect 40910 21534 40962 21586
rect 41358 21534 41410 21586
rect 42814 21534 42866 21586
rect 46062 21534 46114 21586
rect 47294 21534 47346 21586
rect 2494 21422 2546 21474
rect 4622 21422 4674 21474
rect 5182 21422 5234 21474
rect 7646 21422 7698 21474
rect 11790 21422 11842 21474
rect 15038 21422 15090 21474
rect 16494 21422 16546 21474
rect 18174 21422 18226 21474
rect 20302 21422 20354 21474
rect 22990 21422 23042 21474
rect 31278 21422 31330 21474
rect 35198 21422 35250 21474
rect 36990 21422 37042 21474
rect 43262 21422 43314 21474
rect 16158 21310 16210 21362
rect 16382 21310 16434 21362
rect 32174 21310 32226 21362
rect 37214 21310 37266 21362
rect 46958 21310 47010 21362
rect 4478 21142 4530 21194
rect 4582 21142 4634 21194
rect 4686 21142 4738 21194
rect 35198 21142 35250 21194
rect 35302 21142 35354 21194
rect 35406 21142 35458 21194
rect 7310 20974 7362 21026
rect 1710 20862 1762 20914
rect 5070 20862 5122 20914
rect 6078 20862 6130 20914
rect 7982 20862 8034 20914
rect 4510 20750 4562 20802
rect 6526 20750 6578 20802
rect 6750 20750 6802 20802
rect 7870 20750 7922 20802
rect 8878 20750 8930 20802
rect 9998 20974 10050 21026
rect 13582 20974 13634 21026
rect 15038 20974 15090 21026
rect 23662 20974 23714 21026
rect 34750 20974 34802 21026
rect 35086 20974 35138 21026
rect 47966 20974 48018 21026
rect 9886 20862 9938 20914
rect 10334 20862 10386 20914
rect 11006 20862 11058 20914
rect 11342 20862 11394 20914
rect 12798 20862 12850 20914
rect 22430 20862 22482 20914
rect 23998 20862 24050 20914
rect 32174 20862 32226 20914
rect 34302 20862 34354 20914
rect 36430 20862 36482 20914
rect 37662 20862 37714 20914
rect 39118 20862 39170 20914
rect 41246 20862 41298 20914
rect 43598 20862 43650 20914
rect 9214 20750 9266 20802
rect 9438 20750 9490 20802
rect 11566 20750 11618 20802
rect 11790 20750 11842 20802
rect 12126 20750 12178 20802
rect 12350 20750 12402 20802
rect 13470 20750 13522 20802
rect 13918 20750 13970 20802
rect 14478 20750 14530 20802
rect 14702 20750 14754 20802
rect 16158 20750 16210 20802
rect 16270 20750 16322 20802
rect 21422 20750 21474 20802
rect 21982 20750 22034 20802
rect 22990 20750 23042 20802
rect 23102 20750 23154 20802
rect 23214 20750 23266 20802
rect 25902 20750 25954 20802
rect 26350 20750 26402 20802
rect 31502 20750 31554 20802
rect 35870 20750 35922 20802
rect 38334 20750 38386 20802
rect 42030 20750 42082 20802
rect 42814 20750 42866 20802
rect 43710 20750 43762 20802
rect 45054 20750 45106 20802
rect 45614 20750 45666 20802
rect 3838 20638 3890 20690
rect 10558 20638 10610 20690
rect 10670 20638 10722 20690
rect 14142 20638 14194 20690
rect 15374 20638 15426 20690
rect 15486 20638 15538 20690
rect 15934 20638 15986 20690
rect 16718 20638 16770 20690
rect 24110 20638 24162 20690
rect 25454 20638 25506 20690
rect 26574 20638 26626 20690
rect 28366 20638 28418 20690
rect 30718 20638 30770 20690
rect 35758 20638 35810 20690
rect 37214 20638 37266 20690
rect 42926 20638 42978 20690
rect 43822 20638 43874 20690
rect 45278 20638 45330 20690
rect 8766 20526 8818 20578
rect 9102 20526 9154 20578
rect 10894 20526 10946 20578
rect 11566 20526 11618 20578
rect 13694 20526 13746 20578
rect 14926 20526 14978 20578
rect 15262 20526 15314 20578
rect 16382 20526 16434 20578
rect 16494 20526 16546 20578
rect 17278 20526 17330 20578
rect 24782 20526 24834 20578
rect 25118 20526 25170 20578
rect 26126 20526 26178 20578
rect 28030 20526 28082 20578
rect 31054 20526 31106 20578
rect 19838 20358 19890 20410
rect 19942 20358 19994 20410
rect 20046 20358 20098 20410
rect 15710 20190 15762 20242
rect 16046 20190 16098 20242
rect 31950 20190 32002 20242
rect 33182 20190 33234 20242
rect 42142 20190 42194 20242
rect 2158 20078 2210 20130
rect 2830 20078 2882 20130
rect 3278 20078 3330 20130
rect 3614 20078 3666 20130
rect 4174 20078 4226 20130
rect 4734 20078 4786 20130
rect 7982 20078 8034 20130
rect 8990 20078 9042 20130
rect 16606 20078 16658 20130
rect 16830 20078 16882 20130
rect 18398 20078 18450 20130
rect 20974 20078 21026 20130
rect 21534 20078 21586 20130
rect 28814 20078 28866 20130
rect 30158 20078 30210 20130
rect 35310 20078 35362 20130
rect 41246 20078 41298 20130
rect 43710 20078 43762 20130
rect 44382 20078 44434 20130
rect 45054 20078 45106 20130
rect 4398 19966 4450 20018
rect 5406 19966 5458 20018
rect 5630 19966 5682 20018
rect 6862 19966 6914 20018
rect 8318 19966 8370 20018
rect 8542 19966 8594 20018
rect 8766 19966 8818 20018
rect 9550 19966 9602 20018
rect 11118 19966 11170 20018
rect 11342 19966 11394 20018
rect 11902 19966 11954 20018
rect 12686 19966 12738 20018
rect 12798 19966 12850 20018
rect 13694 19966 13746 20018
rect 13918 19966 13970 20018
rect 14030 19966 14082 20018
rect 15150 19966 15202 20018
rect 16046 19966 16098 20018
rect 18734 19966 18786 20018
rect 25566 19966 25618 20018
rect 28926 19966 28978 20018
rect 30046 19966 30098 20018
rect 30382 19966 30434 20018
rect 31614 19966 31666 20018
rect 31838 19966 31890 20018
rect 32174 19966 32226 20018
rect 34638 19966 34690 20018
rect 37774 19966 37826 20018
rect 40910 19966 40962 20018
rect 41582 19966 41634 20018
rect 41806 19966 41858 20018
rect 42478 19966 42530 20018
rect 43038 19966 43090 20018
rect 43486 19966 43538 20018
rect 44046 19966 44098 20018
rect 45390 19966 45442 20018
rect 4062 19854 4114 19906
rect 4958 19854 5010 19906
rect 5742 19854 5794 19906
rect 6414 19854 6466 19906
rect 7422 19854 7474 19906
rect 8654 19854 8706 19906
rect 10110 19854 10162 19906
rect 11790 19854 11842 19906
rect 15374 19854 15426 19906
rect 26238 19854 26290 19906
rect 28366 19854 28418 19906
rect 30830 19854 30882 19906
rect 37438 19854 37490 19906
rect 40126 19854 40178 19906
rect 46062 19854 46114 19906
rect 48190 19854 48242 19906
rect 3726 19742 3778 19794
rect 5070 19742 5122 19794
rect 9886 19742 9938 19794
rect 13358 19742 13410 19794
rect 14478 19742 14530 19794
rect 16270 19742 16322 19794
rect 20414 19742 20466 19794
rect 20750 19742 20802 19794
rect 28814 19742 28866 19794
rect 30606 19742 30658 19794
rect 30830 19742 30882 19794
rect 4478 19574 4530 19626
rect 4582 19574 4634 19626
rect 4686 19574 4738 19626
rect 35198 19574 35250 19626
rect 35302 19574 35354 19626
rect 35406 19574 35458 19626
rect 2046 19406 2098 19458
rect 2942 19406 2994 19458
rect 4846 19406 4898 19458
rect 11230 19406 11282 19458
rect 11790 19406 11842 19458
rect 12238 19406 12290 19458
rect 14254 19406 14306 19458
rect 15262 19406 15314 19458
rect 42366 19406 42418 19458
rect 47966 19406 48018 19458
rect 2158 19294 2210 19346
rect 2494 19294 2546 19346
rect 2942 19294 2994 19346
rect 3502 19294 3554 19346
rect 5854 19294 5906 19346
rect 6302 19294 6354 19346
rect 7086 19294 7138 19346
rect 8766 19294 8818 19346
rect 10110 19294 10162 19346
rect 10782 19294 10834 19346
rect 11790 19294 11842 19346
rect 13022 19294 13074 19346
rect 15822 19294 15874 19346
rect 16718 19294 16770 19346
rect 18622 19294 18674 19346
rect 20750 19294 20802 19346
rect 25566 19294 25618 19346
rect 26462 19294 26514 19346
rect 30158 19294 30210 19346
rect 32174 19294 32226 19346
rect 33966 19294 34018 19346
rect 35982 19294 36034 19346
rect 39902 19294 39954 19346
rect 41022 19294 41074 19346
rect 42926 19294 42978 19346
rect 43374 19294 43426 19346
rect 43822 19294 43874 19346
rect 44942 19294 44994 19346
rect 3726 19182 3778 19234
rect 3950 19182 4002 19234
rect 4398 19182 4450 19234
rect 4958 19182 5010 19234
rect 8094 19182 8146 19234
rect 8206 19182 8258 19234
rect 8430 19182 8482 19234
rect 8990 19182 9042 19234
rect 10446 19182 10498 19234
rect 12238 19182 12290 19234
rect 13918 19182 13970 19234
rect 14142 19182 14194 19234
rect 14366 19182 14418 19234
rect 14702 19182 14754 19234
rect 14926 19182 14978 19234
rect 16494 19182 16546 19234
rect 17278 19182 17330 19234
rect 17838 19182 17890 19234
rect 21310 19182 21362 19234
rect 22654 19182 22706 19234
rect 26350 19182 26402 19234
rect 26574 19182 26626 19234
rect 27022 19182 27074 19234
rect 29486 19182 29538 19234
rect 29934 19182 29986 19234
rect 30270 19182 30322 19234
rect 30830 19182 30882 19234
rect 31278 19182 31330 19234
rect 31838 19182 31890 19234
rect 32286 19182 32338 19234
rect 32398 19182 32450 19234
rect 33182 19182 33234 19234
rect 33294 19182 33346 19234
rect 33518 19182 33570 19234
rect 33854 19182 33906 19234
rect 34414 19182 34466 19234
rect 37550 19182 37602 19234
rect 41694 19182 41746 19234
rect 42030 19182 42082 19234
rect 44718 19182 44770 19234
rect 45614 19182 45666 19234
rect 8654 19070 8706 19122
rect 9326 19070 9378 19122
rect 11342 19070 11394 19122
rect 13694 19070 13746 19122
rect 16270 19070 16322 19122
rect 16830 19070 16882 19122
rect 17390 19070 17442 19122
rect 23438 19070 23490 19122
rect 29150 19070 29202 19122
rect 29262 19070 29314 19122
rect 29710 19070 29762 19122
rect 30606 19070 30658 19122
rect 32846 19070 32898 19122
rect 34862 19070 34914 19122
rect 35422 19070 35474 19122
rect 41358 19070 41410 19122
rect 42254 19070 42306 19122
rect 4174 18958 4226 19010
rect 4286 18958 4338 19010
rect 7422 18958 7474 19010
rect 9214 18958 9266 19010
rect 16718 18958 16770 19010
rect 17614 18958 17666 19010
rect 21646 18958 21698 19010
rect 26126 18958 26178 19010
rect 28590 18958 28642 19010
rect 30942 18958 30994 19010
rect 32062 18958 32114 19010
rect 33070 18958 33122 19010
rect 34078 18958 34130 19010
rect 34302 18958 34354 19010
rect 36430 18958 36482 19010
rect 37214 18958 37266 19010
rect 40462 18958 40514 19010
rect 41694 18958 41746 19010
rect 42366 18958 42418 19010
rect 44270 18958 44322 19010
rect 45054 18958 45106 19010
rect 45278 18958 45330 19010
rect 19838 18790 19890 18842
rect 19942 18790 19994 18842
rect 20046 18790 20098 18842
rect 5294 18622 5346 18674
rect 7422 18622 7474 18674
rect 10222 18622 10274 18674
rect 7758 18566 7810 18618
rect 12126 18622 12178 18674
rect 16046 18622 16098 18674
rect 18622 18622 18674 18674
rect 25454 18622 25506 18674
rect 29710 18622 29762 18674
rect 30382 18622 30434 18674
rect 31278 18622 31330 18674
rect 31950 18622 32002 18674
rect 32174 18622 32226 18674
rect 39006 18622 39058 18674
rect 40462 18622 40514 18674
rect 42702 18622 42754 18674
rect 43710 18622 43762 18674
rect 45614 18622 45666 18674
rect 46510 18622 46562 18674
rect 47182 18622 47234 18674
rect 5070 18510 5122 18562
rect 7086 18510 7138 18562
rect 10782 18510 10834 18562
rect 11118 18510 11170 18562
rect 11454 18510 11506 18562
rect 12910 18510 12962 18562
rect 13246 18510 13298 18562
rect 13470 18510 13522 18562
rect 14590 18510 14642 18562
rect 16606 18510 16658 18562
rect 19518 18510 19570 18562
rect 21758 18510 21810 18562
rect 25902 18510 25954 18562
rect 26574 18510 26626 18562
rect 27246 18510 27298 18562
rect 28366 18510 28418 18562
rect 28478 18510 28530 18562
rect 29934 18510 29986 18562
rect 30158 18510 30210 18562
rect 31166 18510 31218 18562
rect 36430 18510 36482 18562
rect 45838 18510 45890 18562
rect 47854 18510 47906 18562
rect 1822 18398 1874 18450
rect 5518 18398 5570 18450
rect 7982 18398 8034 18450
rect 9774 18398 9826 18450
rect 11902 18398 11954 18450
rect 12574 18398 12626 18450
rect 13694 18398 13746 18450
rect 16270 18398 16322 18450
rect 18958 18398 19010 18450
rect 19630 18398 19682 18450
rect 21086 18398 21138 18450
rect 24222 18398 24274 18450
rect 25342 18398 25394 18450
rect 25678 18398 25730 18450
rect 26350 18398 26402 18450
rect 27022 18398 27074 18450
rect 27582 18398 27634 18450
rect 28142 18398 28194 18450
rect 30606 18398 30658 18450
rect 31502 18398 31554 18450
rect 31838 18398 31890 18450
rect 32398 18398 32450 18450
rect 35310 18398 35362 18450
rect 36094 18398 36146 18450
rect 37102 18398 37154 18450
rect 37886 18398 37938 18450
rect 38446 18398 38498 18450
rect 39454 18398 39506 18450
rect 39678 18398 39730 18450
rect 39902 18398 39954 18450
rect 40350 18398 40402 18450
rect 41806 18398 41858 18450
rect 42142 18398 42194 18450
rect 42590 18398 42642 18450
rect 43262 18398 43314 18450
rect 43486 18398 43538 18450
rect 43934 18398 43986 18450
rect 44830 18398 44882 18450
rect 46062 18398 46114 18450
rect 46734 18398 46786 18450
rect 47518 18398 47570 18450
rect 48190 18398 48242 18450
rect 2494 18286 2546 18338
rect 4622 18286 4674 18338
rect 5182 18286 5234 18338
rect 6190 18286 6242 18338
rect 6750 18286 6802 18338
rect 9102 18286 9154 18338
rect 11566 18286 11618 18338
rect 13582 18286 13634 18338
rect 14702 18286 14754 18338
rect 17502 18286 17554 18338
rect 23886 18286 23938 18338
rect 24334 18286 24386 18338
rect 25566 18286 25618 18338
rect 26798 18286 26850 18338
rect 30270 18286 30322 18338
rect 32286 18286 32338 18338
rect 34078 18286 34130 18338
rect 37550 18286 37602 18338
rect 40126 18286 40178 18338
rect 42254 18286 42306 18338
rect 44046 18286 44098 18338
rect 44382 18286 44434 18338
rect 45278 18286 45330 18338
rect 45726 18286 45778 18338
rect 46398 18286 46450 18338
rect 5742 18174 5794 18226
rect 9886 18174 9938 18226
rect 10334 18174 10386 18226
rect 12238 18174 12290 18226
rect 14814 18174 14866 18226
rect 16270 18174 16322 18226
rect 37102 18174 37154 18226
rect 42702 18174 42754 18226
rect 4478 18006 4530 18058
rect 4582 18006 4634 18058
rect 4686 18006 4738 18058
rect 35198 18006 35250 18058
rect 35302 18006 35354 18058
rect 35406 18006 35458 18058
rect 7198 17838 7250 17890
rect 8990 17838 9042 17890
rect 38670 17838 38722 17890
rect 1934 17726 1986 17778
rect 7086 17726 7138 17778
rect 9550 17726 9602 17778
rect 13582 17726 13634 17778
rect 14702 17726 14754 17778
rect 16830 17726 16882 17778
rect 20078 17726 20130 17778
rect 28590 17726 28642 17778
rect 30830 17726 30882 17778
rect 31278 17726 31330 17778
rect 36430 17726 36482 17778
rect 40462 17726 40514 17778
rect 42702 17726 42754 17778
rect 43486 17726 43538 17778
rect 44158 17726 44210 17778
rect 44942 17726 44994 17778
rect 48190 17726 48242 17778
rect 3838 17614 3890 17666
rect 5630 17614 5682 17666
rect 6414 17614 6466 17666
rect 8654 17614 8706 17666
rect 9774 17614 9826 17666
rect 9886 17614 9938 17666
rect 11454 17614 11506 17666
rect 11678 17614 11730 17666
rect 12238 17614 12290 17666
rect 12686 17614 12738 17666
rect 14030 17614 14082 17666
rect 19742 17614 19794 17666
rect 21870 17614 21922 17666
rect 25790 17614 25842 17666
rect 29598 17614 29650 17666
rect 29822 17614 29874 17666
rect 30046 17614 30098 17666
rect 30158 17614 30210 17666
rect 31838 17614 31890 17666
rect 32174 17614 32226 17666
rect 32286 17614 32338 17666
rect 32510 17614 32562 17666
rect 35198 17614 35250 17666
rect 35982 17614 36034 17666
rect 37102 17614 37154 17666
rect 38222 17614 38274 17666
rect 39230 17614 39282 17666
rect 40350 17614 40402 17666
rect 41918 17614 41970 17666
rect 42030 17614 42082 17666
rect 43598 17614 43650 17666
rect 45390 17614 45442 17666
rect 4734 17502 4786 17554
rect 5854 17502 5906 17554
rect 5966 17502 6018 17554
rect 6750 17502 6802 17554
rect 8206 17502 8258 17554
rect 8878 17502 8930 17554
rect 12910 17502 12962 17554
rect 17838 17502 17890 17554
rect 18958 17502 19010 17554
rect 26462 17502 26514 17554
rect 32958 17502 33010 17554
rect 33518 17502 33570 17554
rect 34302 17502 34354 17554
rect 35646 17502 35698 17554
rect 42366 17502 42418 17554
rect 42814 17502 42866 17554
rect 46062 17502 46114 17554
rect 5070 17390 5122 17442
rect 5742 17390 5794 17442
rect 10110 17390 10162 17442
rect 11566 17390 11618 17442
rect 12574 17390 12626 17442
rect 17502 17390 17554 17442
rect 18286 17390 18338 17442
rect 19294 17390 19346 17442
rect 22094 17390 22146 17442
rect 22542 17390 22594 17442
rect 29934 17390 29986 17442
rect 32622 17390 32674 17442
rect 32846 17390 32898 17442
rect 33854 17390 33906 17442
rect 34638 17390 34690 17442
rect 34974 17390 35026 17442
rect 42142 17390 42194 17442
rect 44046 17390 44098 17442
rect 44270 17390 44322 17442
rect 19838 17222 19890 17274
rect 19942 17222 19994 17274
rect 20046 17222 20098 17274
rect 3278 17054 3330 17106
rect 4286 17054 4338 17106
rect 5070 17054 5122 17106
rect 5742 17054 5794 17106
rect 6638 17054 6690 17106
rect 7422 17054 7474 17106
rect 7646 17054 7698 17106
rect 8542 17054 8594 17106
rect 9886 17054 9938 17106
rect 14478 17054 14530 17106
rect 15822 17054 15874 17106
rect 16606 17054 16658 17106
rect 23774 17054 23826 17106
rect 24222 17054 24274 17106
rect 25230 17054 25282 17106
rect 25566 17054 25618 17106
rect 29486 17054 29538 17106
rect 31390 17054 31442 17106
rect 31726 17054 31778 17106
rect 33294 17054 33346 17106
rect 35422 17054 35474 17106
rect 38670 17054 38722 17106
rect 40238 17054 40290 17106
rect 41358 17054 41410 17106
rect 43710 17054 43762 17106
rect 46062 17054 46114 17106
rect 4958 16942 5010 16994
rect 5294 16942 5346 16994
rect 6078 16942 6130 16994
rect 9550 16942 9602 16994
rect 11230 16942 11282 16994
rect 13806 16942 13858 16994
rect 14926 16942 14978 16994
rect 19518 16942 19570 16994
rect 26574 16942 26626 16994
rect 26910 16942 26962 16994
rect 28926 16942 28978 16994
rect 29262 16942 29314 16994
rect 30270 16942 30322 16994
rect 30494 16942 30546 16994
rect 31502 16942 31554 16994
rect 31950 16942 32002 16994
rect 33070 16942 33122 16994
rect 34974 16942 35026 16994
rect 36542 16942 36594 16994
rect 36878 16942 36930 16994
rect 39006 16942 39058 16994
rect 39902 16942 39954 16994
rect 42814 16942 42866 16994
rect 43262 16942 43314 16994
rect 44270 16942 44322 16994
rect 46958 16942 47010 16994
rect 47518 16942 47570 16994
rect 47630 16942 47682 16994
rect 48078 16942 48130 16994
rect 2830 16830 2882 16882
rect 4174 16830 4226 16882
rect 4510 16830 4562 16882
rect 8094 16830 8146 16882
rect 10334 16830 10386 16882
rect 12126 16830 12178 16882
rect 14142 16830 14194 16882
rect 16270 16830 16322 16882
rect 17502 16830 17554 16882
rect 17950 16830 18002 16882
rect 18734 16830 18786 16882
rect 22318 16830 22370 16882
rect 22542 16830 22594 16882
rect 23214 16830 23266 16882
rect 26350 16830 26402 16882
rect 26798 16830 26850 16882
rect 29486 16830 29538 16882
rect 29822 16830 29874 16882
rect 33518 16830 33570 16882
rect 34190 16830 34242 16882
rect 34414 16830 34466 16882
rect 36206 16830 36258 16882
rect 37214 16830 37266 16882
rect 37774 16830 37826 16882
rect 39230 16830 39282 16882
rect 39566 16830 39618 16882
rect 40910 16830 40962 16882
rect 41134 16830 41186 16882
rect 42702 16830 42754 16882
rect 43822 16830 43874 16882
rect 44830 16830 44882 16882
rect 45726 16830 45778 16882
rect 46174 16830 46226 16882
rect 46286 16830 46338 16882
rect 47294 16830 47346 16882
rect 3166 16718 3218 16770
rect 4398 16718 4450 16770
rect 7534 16718 7586 16770
rect 7870 16718 7922 16770
rect 16046 16718 16098 16770
rect 21646 16718 21698 16770
rect 30158 16718 30210 16770
rect 31614 16718 31666 16770
rect 38110 16718 38162 16770
rect 38222 16718 38274 16770
rect 39118 16718 39170 16770
rect 41022 16718 41074 16770
rect 41806 16718 41858 16770
rect 44718 16718 44770 16770
rect 45502 16718 45554 16770
rect 46846 16718 46898 16770
rect 3614 16606 3666 16658
rect 3838 16606 3890 16658
rect 22878 16606 22930 16658
rect 26126 16606 26178 16658
rect 41918 16606 41970 16658
rect 42142 16606 42194 16658
rect 42254 16606 42306 16658
rect 42814 16606 42866 16658
rect 46734 16606 46786 16658
rect 4478 16438 4530 16490
rect 4582 16438 4634 16490
rect 4686 16438 4738 16490
rect 35198 16438 35250 16490
rect 35302 16438 35354 16490
rect 35406 16438 35458 16490
rect 7198 16270 7250 16322
rect 11902 16270 11954 16322
rect 18958 16270 19010 16322
rect 19294 16270 19346 16322
rect 34862 16270 34914 16322
rect 37662 16270 37714 16322
rect 38670 16270 38722 16322
rect 39230 16270 39282 16322
rect 40686 16270 40738 16322
rect 43374 16270 43426 16322
rect 44942 16270 44994 16322
rect 1710 16158 1762 16210
rect 3838 16158 3890 16210
rect 5070 16158 5122 16210
rect 5854 16158 5906 16210
rect 6190 16158 6242 16210
rect 7646 16158 7698 16210
rect 14590 16158 14642 16210
rect 20750 16158 20802 16210
rect 21758 16158 21810 16210
rect 25902 16158 25954 16210
rect 27918 16158 27970 16210
rect 29262 16158 29314 16210
rect 30158 16158 30210 16210
rect 33854 16158 33906 16210
rect 35646 16158 35698 16210
rect 43038 16158 43090 16210
rect 44382 16158 44434 16210
rect 46398 16158 46450 16210
rect 46958 16158 47010 16210
rect 4622 16046 4674 16098
rect 7422 16046 7474 16098
rect 8094 16046 8146 16098
rect 9998 16046 10050 16098
rect 12238 16046 12290 16098
rect 12686 16046 12738 16098
rect 14030 16046 14082 16098
rect 16942 16046 16994 16098
rect 20078 16046 20130 16098
rect 22430 16046 22482 16098
rect 23662 16046 23714 16098
rect 23886 16046 23938 16098
rect 24670 16046 24722 16098
rect 25678 16046 25730 16098
rect 28254 16046 28306 16098
rect 29038 16046 29090 16098
rect 29710 16046 29762 16098
rect 31726 16046 31778 16098
rect 31950 16046 32002 16098
rect 34302 16046 34354 16098
rect 35198 16046 35250 16098
rect 35534 16046 35586 16098
rect 36206 16046 36258 16098
rect 37214 16046 37266 16098
rect 37662 16046 37714 16098
rect 37998 16046 38050 16098
rect 39454 16046 39506 16098
rect 40350 16046 40402 16098
rect 40798 16046 40850 16098
rect 41358 16046 41410 16098
rect 41582 16046 41634 16098
rect 45166 16046 45218 16098
rect 45614 16046 45666 16098
rect 45950 16046 46002 16098
rect 9886 15934 9938 15986
rect 12014 15934 12066 15986
rect 12910 15934 12962 15986
rect 17278 15934 17330 15986
rect 19966 15934 20018 15986
rect 22206 15934 22258 15986
rect 23214 15934 23266 15986
rect 24334 15934 24386 15986
rect 26014 15934 26066 15986
rect 28590 15934 28642 15986
rect 29486 15934 29538 15986
rect 30046 15934 30098 15986
rect 30270 15934 30322 15986
rect 31614 15934 31666 15986
rect 34526 15934 34578 15986
rect 38334 15934 38386 15986
rect 38894 15934 38946 15986
rect 40014 15934 40066 15986
rect 41470 15934 41522 15986
rect 42142 15934 42194 15986
rect 42478 15934 42530 15986
rect 43710 15934 43762 15986
rect 47294 15934 47346 15986
rect 7870 15822 7922 15874
rect 7982 15822 8034 15874
rect 11902 15822 11954 15874
rect 12574 15822 12626 15874
rect 16494 15822 16546 15874
rect 21310 15822 21362 15874
rect 22878 15822 22930 15874
rect 23998 15822 24050 15874
rect 24110 15822 24162 15874
rect 25006 15822 25058 15874
rect 31166 15822 31218 15874
rect 34974 15822 35026 15874
rect 35758 15822 35810 15874
rect 38222 15822 38274 15874
rect 39566 15822 39618 15874
rect 40238 15822 40290 15874
rect 41134 15822 41186 15874
rect 42030 15822 42082 15874
rect 42254 15822 42306 15874
rect 43486 15822 43538 15874
rect 47854 15822 47906 15874
rect 19838 15654 19890 15706
rect 19942 15654 19994 15706
rect 20046 15654 20098 15706
rect 4734 15486 4786 15538
rect 4958 15486 5010 15538
rect 11006 15486 11058 15538
rect 12238 15486 12290 15538
rect 24446 15486 24498 15538
rect 27918 15486 27970 15538
rect 28814 15486 28866 15538
rect 33070 15486 33122 15538
rect 34526 15486 34578 15538
rect 34862 15486 34914 15538
rect 35870 15486 35922 15538
rect 36654 15486 36706 15538
rect 37774 15486 37826 15538
rect 37998 15486 38050 15538
rect 40014 15486 40066 15538
rect 41470 15486 41522 15538
rect 41694 15486 41746 15538
rect 43486 15486 43538 15538
rect 5630 15374 5682 15426
rect 7086 15374 7138 15426
rect 9550 15374 9602 15426
rect 13246 15374 13298 15426
rect 16382 15374 16434 15426
rect 16606 15374 16658 15426
rect 17726 15374 17778 15426
rect 19406 15374 19458 15426
rect 25342 15374 25394 15426
rect 27694 15374 27746 15426
rect 31614 15374 31666 15426
rect 31726 15374 31778 15426
rect 36318 15374 36370 15426
rect 37550 15374 37602 15426
rect 39678 15374 39730 15426
rect 39790 15374 39842 15426
rect 40238 15374 40290 15426
rect 40350 15374 40402 15426
rect 41246 15374 41298 15426
rect 44830 15374 44882 15426
rect 47406 15374 47458 15426
rect 5406 15262 5458 15314
rect 6862 15262 6914 15314
rect 7198 15262 7250 15314
rect 7534 15262 7586 15314
rect 10782 15262 10834 15314
rect 11342 15262 11394 15314
rect 11790 15262 11842 15314
rect 12574 15250 12626 15302
rect 17390 15262 17442 15314
rect 19294 15262 19346 15314
rect 21310 15262 21362 15314
rect 24110 15262 24162 15314
rect 24222 15262 24274 15314
rect 24670 15262 24722 15314
rect 26126 15262 26178 15314
rect 26574 15262 26626 15314
rect 27582 15262 27634 15314
rect 31950 15262 32002 15314
rect 33294 15262 33346 15314
rect 34302 15262 34354 15314
rect 35086 15262 35138 15314
rect 35534 15262 35586 15314
rect 36542 15262 36594 15314
rect 36878 15262 36930 15314
rect 39118 15262 39170 15314
rect 41582 15262 41634 15314
rect 41918 15262 41970 15314
rect 43822 15262 43874 15314
rect 45950 15262 46002 15314
rect 46398 15262 46450 15314
rect 4846 15150 4898 15202
rect 5966 15150 6018 15202
rect 6974 15150 7026 15202
rect 9662 15150 9714 15202
rect 10222 15150 10274 15202
rect 11566 15150 11618 15202
rect 15374 15150 15426 15202
rect 15822 15150 15874 15202
rect 16270 15150 16322 15202
rect 18622 15150 18674 15202
rect 21870 15150 21922 15202
rect 24446 15150 24498 15202
rect 26686 15150 26738 15202
rect 29822 15150 29874 15202
rect 38782 15150 38834 15202
rect 42366 15150 42418 15202
rect 42814 15150 42866 15202
rect 44606 15150 44658 15202
rect 18286 15038 18338 15090
rect 31166 15038 31218 15090
rect 38110 15038 38162 15090
rect 39678 15038 39730 15090
rect 4478 14870 4530 14922
rect 4582 14870 4634 14922
rect 4686 14870 4738 14922
rect 35198 14870 35250 14922
rect 35302 14870 35354 14922
rect 35406 14870 35458 14922
rect 21758 14702 21810 14754
rect 26574 14702 26626 14754
rect 34414 14702 34466 14754
rect 38110 14702 38162 14754
rect 41582 14702 41634 14754
rect 2494 14590 2546 14642
rect 4622 14590 4674 14642
rect 7870 14590 7922 14642
rect 9998 14590 10050 14642
rect 10782 14590 10834 14642
rect 12014 14590 12066 14642
rect 13918 14590 13970 14642
rect 20078 14590 20130 14642
rect 21982 14590 22034 14642
rect 23662 14590 23714 14642
rect 26238 14590 26290 14642
rect 28590 14590 28642 14642
rect 35310 14590 35362 14642
rect 40574 14590 40626 14642
rect 43486 14590 43538 14642
rect 44942 14590 44994 14642
rect 46062 14590 46114 14642
rect 48190 14590 48242 14642
rect 1822 14478 1874 14530
rect 7198 14478 7250 14530
rect 10446 14478 10498 14530
rect 10670 14478 10722 14530
rect 12238 14478 12290 14530
rect 12910 14478 12962 14530
rect 16270 14478 16322 14530
rect 16606 14478 16658 14530
rect 16942 14478 16994 14530
rect 17278 14478 17330 14530
rect 20638 14478 20690 14530
rect 21870 14478 21922 14530
rect 22206 14478 22258 14530
rect 23550 14478 23602 14530
rect 24334 14478 24386 14530
rect 25006 14478 25058 14530
rect 26014 14478 26066 14530
rect 29486 14478 29538 14530
rect 30158 14478 30210 14530
rect 35646 14478 35698 14530
rect 35982 14478 36034 14530
rect 37886 14478 37938 14530
rect 39006 14478 39058 14530
rect 40014 14478 40066 14530
rect 40686 14478 40738 14530
rect 41022 14478 41074 14530
rect 41470 14478 41522 14530
rect 41694 14478 41746 14530
rect 43038 14478 43090 14530
rect 44270 14478 44322 14530
rect 45278 14478 45330 14530
rect 10334 14366 10386 14418
rect 17950 14366 18002 14418
rect 20414 14366 20466 14418
rect 23998 14366 24050 14418
rect 25678 14366 25730 14418
rect 27246 14366 27298 14418
rect 30382 14366 30434 14418
rect 31166 14366 31218 14418
rect 31278 14366 31330 14418
rect 34302 14366 34354 14418
rect 37214 14366 37266 14418
rect 37550 14366 37602 14418
rect 43486 14366 43538 14418
rect 43822 14366 43874 14418
rect 5070 14254 5122 14306
rect 12686 14254 12738 14306
rect 12798 14254 12850 14306
rect 16718 14254 16770 14306
rect 24558 14254 24610 14306
rect 24670 14254 24722 14306
rect 24782 14254 24834 14306
rect 25790 14254 25842 14306
rect 26350 14254 26402 14306
rect 27022 14254 27074 14306
rect 27358 14254 27410 14306
rect 27470 14254 27522 14306
rect 28030 14254 28082 14306
rect 29710 14254 29762 14306
rect 30718 14254 30770 14306
rect 35870 14254 35922 14306
rect 38446 14254 38498 14306
rect 38782 14254 38834 14306
rect 39454 14254 39506 14306
rect 39790 14254 39842 14306
rect 40462 14254 40514 14306
rect 41246 14254 41298 14306
rect 42030 14254 42082 14306
rect 42366 14254 42418 14306
rect 19838 14086 19890 14138
rect 19942 14086 19994 14138
rect 20046 14086 20098 14138
rect 4622 13918 4674 13970
rect 9662 13918 9714 13970
rect 10782 13918 10834 13970
rect 11454 13918 11506 13970
rect 12798 13918 12850 13970
rect 12910 13918 12962 13970
rect 13470 13918 13522 13970
rect 17502 13918 17554 13970
rect 17950 13918 18002 13970
rect 18734 13918 18786 13970
rect 23550 13918 23602 13970
rect 25342 13918 25394 13970
rect 26126 13918 26178 13970
rect 27918 13918 27970 13970
rect 30942 13918 30994 13970
rect 31054 13918 31106 13970
rect 37886 13918 37938 13970
rect 47070 13918 47122 13970
rect 6526 13806 6578 13858
rect 14478 13806 14530 13858
rect 18286 13806 18338 13858
rect 23326 13806 23378 13858
rect 24446 13806 24498 13858
rect 24670 13806 24722 13858
rect 27022 13806 27074 13858
rect 29262 13806 29314 13858
rect 31166 13806 31218 13858
rect 31278 13806 31330 13858
rect 37214 13806 37266 13858
rect 42254 13806 42306 13858
rect 43710 13806 43762 13858
rect 4846 13694 4898 13746
rect 5070 13694 5122 13746
rect 5854 13694 5906 13746
rect 9998 13694 10050 13746
rect 10222 13694 10274 13746
rect 10446 13694 10498 13746
rect 12238 13694 12290 13746
rect 12686 13694 12738 13746
rect 13806 13694 13858 13746
rect 22542 13694 22594 13746
rect 23774 13694 23826 13746
rect 23998 13694 24050 13746
rect 26910 13694 26962 13746
rect 27470 13694 27522 13746
rect 29598 13694 29650 13746
rect 30718 13694 30770 13746
rect 31726 13694 31778 13746
rect 33406 13694 33458 13746
rect 33966 13694 34018 13746
rect 34414 13694 34466 13746
rect 34862 13694 34914 13746
rect 35422 13694 35474 13746
rect 35870 13694 35922 13746
rect 36878 13694 36930 13746
rect 38558 13694 38610 13746
rect 40014 13694 40066 13746
rect 40798 13694 40850 13746
rect 41582 13694 41634 13746
rect 42142 13694 42194 13746
rect 43374 13694 43426 13746
rect 46286 13694 46338 13746
rect 46734 13694 46786 13746
rect 47742 13694 47794 13746
rect 4734 13582 4786 13634
rect 8654 13582 8706 13634
rect 12014 13582 12066 13634
rect 16606 13582 16658 13634
rect 19182 13582 19234 13634
rect 19630 13582 19682 13634
rect 21422 13582 21474 13634
rect 22990 13582 23042 13634
rect 23662 13582 23714 13634
rect 24446 13582 24498 13634
rect 28478 13582 28530 13634
rect 28926 13582 28978 13634
rect 30046 13582 30098 13634
rect 42702 13582 42754 13634
rect 43934 13582 43986 13634
rect 47966 13582 48018 13634
rect 5294 13470 5346 13522
rect 19406 13470 19458 13522
rect 22766 13470 22818 13522
rect 22990 13470 23042 13522
rect 26686 13470 26738 13522
rect 27246 13470 27298 13522
rect 28254 13470 28306 13522
rect 35870 13470 35922 13522
rect 47518 13470 47570 13522
rect 4478 13302 4530 13354
rect 4582 13302 4634 13354
rect 4686 13302 4738 13354
rect 35198 13302 35250 13354
rect 35302 13302 35354 13354
rect 35406 13302 35458 13354
rect 13694 13134 13746 13186
rect 20078 13134 20130 13186
rect 24782 13134 24834 13186
rect 27022 13134 27074 13186
rect 27246 13134 27298 13186
rect 35422 13134 35474 13186
rect 40350 13134 40402 13186
rect 40686 13134 40738 13186
rect 42702 13134 42754 13186
rect 44158 13134 44210 13186
rect 2494 13022 2546 13074
rect 4622 13022 4674 13074
rect 6638 13022 6690 13074
rect 10446 13022 10498 13074
rect 11454 13022 11506 13074
rect 13022 13022 13074 13074
rect 13470 13022 13522 13074
rect 17726 13022 17778 13074
rect 19630 13022 19682 13074
rect 24334 13022 24386 13074
rect 28702 13022 28754 13074
rect 29486 13022 29538 13074
rect 31614 13022 31666 13074
rect 33742 13022 33794 13074
rect 34190 13022 34242 13074
rect 34526 13022 34578 13074
rect 36430 13022 36482 13074
rect 39678 13022 39730 13074
rect 41470 13022 41522 13074
rect 48190 13022 48242 13074
rect 1822 12910 1874 12962
rect 4958 12910 5010 12962
rect 5630 12910 5682 12962
rect 5854 12910 5906 12962
rect 6078 12910 6130 12962
rect 8878 12910 8930 12962
rect 9214 12910 9266 12962
rect 9998 12910 10050 12962
rect 10110 12910 10162 12962
rect 10334 12910 10386 12962
rect 11006 12910 11058 12962
rect 14814 12910 14866 12962
rect 21310 12910 21362 12962
rect 26798 12910 26850 12962
rect 27470 12910 27522 12962
rect 30046 12910 30098 12962
rect 30606 12910 30658 12962
rect 30830 12910 30882 12962
rect 34750 12910 34802 12962
rect 34974 12910 35026 12962
rect 35646 12910 35698 12962
rect 36094 12910 36146 12962
rect 37662 12910 37714 12962
rect 38894 12910 38946 12962
rect 40014 12910 40066 12962
rect 40910 12910 40962 12962
rect 41246 12910 41298 12962
rect 43598 12910 43650 12962
rect 44382 12910 44434 12962
rect 44830 12910 44882 12962
rect 45278 12910 45330 12962
rect 5070 12798 5122 12850
rect 9438 12798 9490 12850
rect 10558 12798 10610 12850
rect 14366 12798 14418 12850
rect 14478 12798 14530 12850
rect 15598 12798 15650 12850
rect 20078 12798 20130 12850
rect 20190 12798 20242 12850
rect 22094 12798 22146 12850
rect 25006 12798 25058 12850
rect 26462 12798 26514 12850
rect 29598 12798 29650 12850
rect 30270 12798 30322 12850
rect 30382 12798 30434 12850
rect 41582 12798 41634 12850
rect 41694 12798 41746 12850
rect 42590 12798 42642 12850
rect 44942 12798 44994 12850
rect 46062 12798 46114 12850
rect 5742 12686 5794 12738
rect 9550 12686 9602 12738
rect 14030 12686 14082 12738
rect 18174 12686 18226 12738
rect 19182 12686 19234 12738
rect 20638 12686 20690 12738
rect 24894 12686 24946 12738
rect 26126 12686 26178 12738
rect 27918 12686 27970 12738
rect 29374 12686 29426 12738
rect 41470 12686 41522 12738
rect 19838 12518 19890 12570
rect 19942 12518 19994 12570
rect 20046 12518 20098 12570
rect 3166 12350 3218 12402
rect 4286 12350 4338 12402
rect 11118 12350 11170 12402
rect 13134 12350 13186 12402
rect 14478 12350 14530 12402
rect 15598 12350 15650 12402
rect 16718 12350 16770 12402
rect 18622 12350 18674 12402
rect 20078 12350 20130 12402
rect 22766 12350 22818 12402
rect 23998 12350 24050 12402
rect 29374 12350 29426 12402
rect 34638 12350 34690 12402
rect 47966 12350 48018 12402
rect 5406 12238 5458 12290
rect 6862 12238 6914 12290
rect 9662 12238 9714 12290
rect 11230 12238 11282 12290
rect 15150 12238 15202 12290
rect 15374 12238 15426 12290
rect 19518 12238 19570 12290
rect 22990 12238 23042 12290
rect 23438 12238 23490 12290
rect 24222 12238 24274 12290
rect 27246 12238 27298 12290
rect 29262 12238 29314 12290
rect 31838 12238 31890 12290
rect 31950 12238 32002 12290
rect 35982 12238 36034 12290
rect 37102 12238 37154 12290
rect 39902 12238 39954 12290
rect 40350 12238 40402 12290
rect 41918 12238 41970 12290
rect 43262 12238 43314 12290
rect 47406 12238 47458 12290
rect 3390 12126 3442 12178
rect 3614 12126 3666 12178
rect 3838 12126 3890 12178
rect 4510 12126 4562 12178
rect 4734 12126 4786 12178
rect 4958 12126 5010 12178
rect 5294 12126 5346 12178
rect 6190 12126 6242 12178
rect 10334 12126 10386 12178
rect 15934 12126 15986 12178
rect 18174 12126 18226 12178
rect 18734 12126 18786 12178
rect 18958 12126 19010 12178
rect 19294 12126 19346 12178
rect 26686 12126 26738 12178
rect 28702 12126 28754 12178
rect 30942 12126 30994 12178
rect 31166 12126 31218 12178
rect 31502 12126 31554 12178
rect 35534 12126 35586 12178
rect 37326 12126 37378 12178
rect 37774 12126 37826 12178
rect 37998 12126 38050 12178
rect 38782 12126 38834 12178
rect 39342 12126 39394 12178
rect 41470 12126 41522 12178
rect 42814 12126 42866 12178
rect 43150 12126 43202 12178
rect 44046 12126 44098 12178
rect 44494 12126 44546 12178
rect 46846 12126 46898 12178
rect 3278 12014 3330 12066
rect 4398 12014 4450 12066
rect 8990 12014 9042 12066
rect 10670 12014 10722 12066
rect 12126 12014 12178 12066
rect 14030 12014 14082 12066
rect 16606 12014 16658 12066
rect 18510 12014 18562 12066
rect 19518 12014 19570 12066
rect 22654 12014 22706 12066
rect 24110 12014 24162 12066
rect 31054 12014 31106 12066
rect 32622 12014 32674 12066
rect 33294 12014 33346 12066
rect 33742 12014 33794 12066
rect 34302 12014 34354 12066
rect 35086 12014 35138 12066
rect 36654 12014 36706 12066
rect 38446 12014 38498 12066
rect 39454 12014 39506 12066
rect 41022 12014 41074 12066
rect 42254 12014 42306 12066
rect 45950 12014 46002 12066
rect 46286 12014 46338 12066
rect 9438 11902 9490 11954
rect 9774 11902 9826 11954
rect 15710 11902 15762 11954
rect 16494 11902 16546 11954
rect 31950 11902 32002 11954
rect 34190 11902 34242 11954
rect 34974 11902 35026 11954
rect 38222 11902 38274 11954
rect 40238 11902 40290 11954
rect 45838 11902 45890 11954
rect 4478 11734 4530 11786
rect 4582 11734 4634 11786
rect 4686 11734 4738 11786
rect 35198 11734 35250 11786
rect 35302 11734 35354 11786
rect 35406 11734 35458 11786
rect 9998 11566 10050 11618
rect 11006 11566 11058 11618
rect 30046 11566 30098 11618
rect 37102 11566 37154 11618
rect 39902 11566 39954 11618
rect 2494 11454 2546 11506
rect 4622 11454 4674 11506
rect 6414 11454 6466 11506
rect 9326 11454 9378 11506
rect 12798 11454 12850 11506
rect 13806 11454 13858 11506
rect 18622 11454 18674 11506
rect 20750 11454 20802 11506
rect 24110 11454 24162 11506
rect 26238 11454 26290 11506
rect 28142 11454 28194 11506
rect 32510 11454 32562 11506
rect 34638 11454 34690 11506
rect 35086 11454 35138 11506
rect 36206 11454 36258 11506
rect 36990 11454 37042 11506
rect 37998 11454 38050 11506
rect 40686 11454 40738 11506
rect 47742 11454 47794 11506
rect 1822 11342 1874 11394
rect 4958 11342 5010 11394
rect 5630 11342 5682 11394
rect 7758 11342 7810 11394
rect 7982 11342 8034 11394
rect 8766 11342 8818 11394
rect 9774 11342 9826 11394
rect 10222 11342 10274 11394
rect 11230 11342 11282 11394
rect 11678 11342 11730 11394
rect 12238 11342 12290 11394
rect 12910 11342 12962 11394
rect 13470 11342 13522 11394
rect 17950 11342 18002 11394
rect 23326 11342 23378 11394
rect 28478 11342 28530 11394
rect 29038 11342 29090 11394
rect 29374 11342 29426 11394
rect 30606 11342 30658 11394
rect 31054 11342 31106 11394
rect 31838 11342 31890 11394
rect 39678 11342 39730 11394
rect 43598 11342 43650 11394
rect 44830 11342 44882 11394
rect 5070 11230 5122 11282
rect 5966 11230 6018 11282
rect 8990 11230 9042 11282
rect 10334 11230 10386 11282
rect 12686 11230 12738 11282
rect 13694 11230 13746 11282
rect 29598 11230 29650 11282
rect 29710 11230 29762 11282
rect 7870 11118 7922 11170
rect 8206 11118 8258 11170
rect 9438 11118 9490 11170
rect 10670 11118 10722 11170
rect 11790 11118 11842 11170
rect 12014 11118 12066 11170
rect 12462 11118 12514 11170
rect 14366 11118 14418 11170
rect 21422 11118 21474 11170
rect 22990 11118 23042 11170
rect 28590 11118 28642 11170
rect 29934 11174 29986 11226
rect 30046 11230 30098 11282
rect 31278 11230 31330 11282
rect 37550 11230 37602 11282
rect 39006 11230 39058 11282
rect 40238 11230 40290 11282
rect 42814 11230 42866 11282
rect 45614 11230 45666 11282
rect 30830 11118 30882 11170
rect 35870 11118 35922 11170
rect 40014 11118 40066 11170
rect 44270 11118 44322 11170
rect 48190 11118 48242 11170
rect 19838 10950 19890 11002
rect 19942 10950 19994 11002
rect 20046 10950 20098 11002
rect 8206 10782 8258 10834
rect 8430 10782 8482 10834
rect 9662 10782 9714 10834
rect 15038 10782 15090 10834
rect 16382 10782 16434 10834
rect 16942 10782 16994 10834
rect 17502 10782 17554 10834
rect 31726 10782 31778 10834
rect 40238 10782 40290 10834
rect 41134 10782 41186 10834
rect 41358 10782 41410 10834
rect 41470 10782 41522 10834
rect 41582 10782 41634 10834
rect 41918 10782 41970 10834
rect 42702 10782 42754 10834
rect 45054 10782 45106 10834
rect 45838 10782 45890 10834
rect 46174 10782 46226 10834
rect 6302 10670 6354 10722
rect 6638 10670 6690 10722
rect 9886 10670 9938 10722
rect 10110 10670 10162 10722
rect 13806 10670 13858 10722
rect 26014 10670 26066 10722
rect 29038 10670 29090 10722
rect 29374 10670 29426 10722
rect 30606 10670 30658 10722
rect 33854 10670 33906 10722
rect 37102 10670 37154 10722
rect 39678 10670 39730 10722
rect 43374 10670 43426 10722
rect 43934 10670 43986 10722
rect 44270 10670 44322 10722
rect 46510 10670 46562 10722
rect 46846 10670 46898 10722
rect 47182 10670 47234 10722
rect 4958 10558 5010 10610
rect 5182 10558 5234 10610
rect 8878 10558 8930 10610
rect 9438 10558 9490 10610
rect 10558 10558 10610 10610
rect 10894 10558 10946 10610
rect 14590 10558 14642 10610
rect 20526 10558 20578 10610
rect 25230 10558 25282 10610
rect 28478 10558 28530 10610
rect 28702 10558 28754 10610
rect 29598 10558 29650 10610
rect 30830 10558 30882 10610
rect 31166 10558 31218 10610
rect 31502 10558 31554 10610
rect 33182 10558 33234 10610
rect 36318 10558 36370 10610
rect 42142 10558 42194 10610
rect 43486 10558 43538 10610
rect 43710 10558 43762 10610
rect 44606 10558 44658 10610
rect 44830 10558 44882 10610
rect 47406 10558 47458 10610
rect 7534 10446 7586 10498
rect 8318 10446 8370 10498
rect 10782 10446 10834 10498
rect 11678 10446 11730 10498
rect 15486 10446 15538 10498
rect 15934 10446 15986 10498
rect 21198 10446 21250 10498
rect 23326 10446 23378 10498
rect 24670 10446 24722 10498
rect 28142 10446 28194 10498
rect 28590 10446 28642 10498
rect 30158 10446 30210 10498
rect 31054 10446 31106 10498
rect 32510 10446 32562 10498
rect 35982 10446 36034 10498
rect 39230 10446 39282 10498
rect 40350 10446 40402 10498
rect 45390 10446 45442 10498
rect 47966 10446 48018 10498
rect 4846 10334 4898 10386
rect 5294 10334 5346 10386
rect 10446 10334 10498 10386
rect 31838 10334 31890 10386
rect 39566 10334 39618 10386
rect 44830 10334 44882 10386
rect 45502 10334 45554 10386
rect 47854 10334 47906 10386
rect 4478 10166 4530 10218
rect 4582 10166 4634 10218
rect 4686 10166 4738 10218
rect 35198 10166 35250 10218
rect 35302 10166 35354 10218
rect 35406 10166 35458 10218
rect 10334 9998 10386 10050
rect 10446 9998 10498 10050
rect 30382 9998 30434 10050
rect 35534 9998 35586 10050
rect 1710 9886 1762 9938
rect 3838 9886 3890 9938
rect 9214 9886 9266 9938
rect 16494 9886 16546 9938
rect 19742 9886 19794 9938
rect 23214 9886 23266 9938
rect 25342 9886 25394 9938
rect 25678 9886 25730 9938
rect 27806 9886 27858 9938
rect 30046 9886 30098 9938
rect 31502 9886 31554 9938
rect 33630 9886 33682 9938
rect 34078 9886 34130 9938
rect 37438 9886 37490 9938
rect 37886 9886 37938 9938
rect 41022 9886 41074 9938
rect 44270 9886 44322 9938
rect 4622 9774 4674 9826
rect 5070 9774 5122 9826
rect 6190 9774 6242 9826
rect 6414 9774 6466 9826
rect 6638 9774 6690 9826
rect 6974 9774 7026 9826
rect 7870 9774 7922 9826
rect 7982 9774 8034 9826
rect 9998 9774 10050 9826
rect 10670 9774 10722 9826
rect 10894 9774 10946 9826
rect 12910 9774 12962 9826
rect 13582 9774 13634 9826
rect 16942 9774 16994 9826
rect 22430 9774 22482 9826
rect 28590 9774 28642 9826
rect 29038 9774 29090 9826
rect 29374 9774 29426 9826
rect 30718 9774 30770 9826
rect 36318 9774 36370 9826
rect 38110 9774 38162 9826
rect 41358 9774 41410 9826
rect 47854 9774 47906 9826
rect 7310 9662 7362 9714
rect 7534 9662 7586 9714
rect 11006 9662 11058 9714
rect 11342 9662 11394 9714
rect 11678 9662 11730 9714
rect 12574 9662 12626 9714
rect 14366 9662 14418 9714
rect 17614 9662 17666 9714
rect 30158 9662 30210 9714
rect 36094 9662 36146 9714
rect 38894 9662 38946 9714
rect 42142 9662 42194 9714
rect 44942 9662 44994 9714
rect 6526 9550 6578 9602
rect 7086 9550 7138 9602
rect 7646 9550 7698 9602
rect 12238 9550 12290 9602
rect 12686 9550 12738 9602
rect 20190 9550 20242 9602
rect 22094 9550 22146 9602
rect 29262 9550 29314 9602
rect 34862 9550 34914 9602
rect 35198 9550 35250 9602
rect 45054 9550 45106 9602
rect 45278 9550 45330 9602
rect 47182 9550 47234 9602
rect 19838 9382 19890 9434
rect 19942 9382 19994 9434
rect 20046 9382 20098 9434
rect 3838 9214 3890 9266
rect 4958 9214 5010 9266
rect 15038 9214 15090 9266
rect 17502 9214 17554 9266
rect 17950 9214 18002 9266
rect 18846 9214 18898 9266
rect 29150 9214 29202 9266
rect 33294 9214 33346 9266
rect 34302 9214 34354 9266
rect 34638 9214 34690 9266
rect 38222 9214 38274 9266
rect 38558 9214 38610 9266
rect 38782 9214 38834 9266
rect 41582 9214 41634 9266
rect 41918 9214 41970 9266
rect 4622 9102 4674 9154
rect 5742 9102 5794 9154
rect 6862 9102 6914 9154
rect 10670 9102 10722 9154
rect 18398 9102 18450 9154
rect 27582 9102 27634 9154
rect 28030 9102 28082 9154
rect 28142 9102 28194 9154
rect 33518 9102 33570 9154
rect 37326 9102 37378 9154
rect 42478 9102 42530 9154
rect 43822 9102 43874 9154
rect 44270 9102 44322 9154
rect 3950 8990 4002 9042
rect 4174 8990 4226 9042
rect 4398 8990 4450 9042
rect 4958 8990 5010 9042
rect 5294 8990 5346 9042
rect 5518 8990 5570 9042
rect 6190 8990 6242 9042
rect 10446 8990 10498 9042
rect 14590 8990 14642 9042
rect 14926 8990 14978 9042
rect 15150 8990 15202 9042
rect 15710 8990 15762 9042
rect 16382 8990 16434 9042
rect 16606 8990 16658 9042
rect 19630 8990 19682 9042
rect 20190 8990 20242 9042
rect 35198 8990 35250 9042
rect 36430 8990 36482 9042
rect 36878 8990 36930 9042
rect 39118 8990 39170 9042
rect 41470 8990 41522 9042
rect 41694 8990 41746 9042
rect 44158 8990 44210 9042
rect 44494 8990 44546 9042
rect 44718 8990 44770 9042
rect 44942 8990 44994 9042
rect 45838 8990 45890 9042
rect 8990 8878 9042 8930
rect 9998 8878 10050 8930
rect 11454 8878 11506 8930
rect 11678 8878 11730 8930
rect 13806 8878 13858 8930
rect 22542 8878 22594 8930
rect 22990 8878 23042 8930
rect 26238 8878 26290 8930
rect 28702 8878 28754 8930
rect 29934 8878 29986 8930
rect 30382 8878 30434 8930
rect 30830 8878 30882 8930
rect 31278 8878 31330 8930
rect 31726 8878 31778 8930
rect 32510 8878 32562 8930
rect 35758 8878 35810 8930
rect 36206 8878 36258 8930
rect 37886 8878 37938 8930
rect 38894 8878 38946 8930
rect 39454 8878 39506 8930
rect 40014 8878 40066 8930
rect 40350 8878 40402 8930
rect 41134 8878 41186 8930
rect 42814 8878 42866 8930
rect 43262 8878 43314 8930
rect 15486 8766 15538 8818
rect 16270 8766 16322 8818
rect 28142 8766 28194 8818
rect 30382 8766 30434 8818
rect 30830 8766 30882 8818
rect 33182 8766 33234 8818
rect 36654 8766 36706 8818
rect 39454 8766 39506 8818
rect 40350 8766 40402 8818
rect 42926 8766 42978 8818
rect 43374 8766 43426 8818
rect 43710 8766 43762 8818
rect 45278 8766 45330 8818
rect 47966 8766 48018 8818
rect 4478 8598 4530 8650
rect 4582 8598 4634 8650
rect 4686 8598 4738 8650
rect 35198 8598 35250 8650
rect 35302 8598 35354 8650
rect 35406 8598 35458 8650
rect 10782 8430 10834 8482
rect 13694 8430 13746 8482
rect 2494 8318 2546 8370
rect 4622 8318 4674 8370
rect 4958 8318 5010 8370
rect 5742 8318 5794 8370
rect 11454 8318 11506 8370
rect 13022 8318 13074 8370
rect 15150 8318 15202 8370
rect 17950 8318 18002 8370
rect 19966 8318 20018 8370
rect 20302 8318 20354 8370
rect 22430 8318 22482 8370
rect 25678 8318 25730 8370
rect 28702 8318 28754 8370
rect 33966 8318 34018 8370
rect 34414 8318 34466 8370
rect 35310 8318 35362 8370
rect 38334 8318 38386 8370
rect 44158 8318 44210 8370
rect 47966 8318 48018 8370
rect 1822 8206 1874 8258
rect 9438 8206 9490 8258
rect 10334 8206 10386 8258
rect 10782 8206 10834 8258
rect 13470 8206 13522 8258
rect 16830 8206 16882 8258
rect 19406 8206 19458 8258
rect 19742 8206 19794 8258
rect 21982 8206 22034 8258
rect 22766 8206 22818 8258
rect 30942 8206 30994 8258
rect 31614 8206 31666 8258
rect 33182 8206 33234 8258
rect 35646 8206 35698 8258
rect 35870 8206 35922 8258
rect 36542 8206 36594 8258
rect 38782 8206 38834 8258
rect 40014 8206 40066 8258
rect 40462 8206 40514 8258
rect 41358 8206 41410 8258
rect 45054 8206 45106 8258
rect 45950 8206 46002 8258
rect 12238 8094 12290 8146
rect 14030 8094 14082 8146
rect 14254 8094 14306 8146
rect 15598 8094 15650 8146
rect 19294 8094 19346 8146
rect 21646 8094 21698 8146
rect 23550 8094 23602 8146
rect 27134 8094 27186 8146
rect 27582 8094 27634 8146
rect 27806 8094 27858 8146
rect 29822 8094 29874 8146
rect 37326 8094 37378 8146
rect 39342 8094 39394 8146
rect 39678 8094 39730 8146
rect 40686 8094 40738 8146
rect 41918 8094 41970 8146
rect 42366 8094 42418 8146
rect 42478 8094 42530 8146
rect 42926 8094 42978 8146
rect 43822 8094 43874 8146
rect 43934 8094 43986 8146
rect 45278 8094 45330 8146
rect 5070 7982 5122 8034
rect 8878 7982 8930 8034
rect 9774 7982 9826 8034
rect 12014 7982 12066 8034
rect 12350 7982 12402 8034
rect 13918 7982 13970 8034
rect 14702 7982 14754 8034
rect 15486 7982 15538 8034
rect 16270 7982 16322 8034
rect 17054 7982 17106 8034
rect 17502 7982 17554 8034
rect 18398 7982 18450 8034
rect 18846 7982 18898 8034
rect 20862 7982 20914 8034
rect 27694 7982 27746 8034
rect 29486 7982 29538 8034
rect 29934 7982 29986 8034
rect 30046 7982 30098 8034
rect 30718 7982 30770 8034
rect 31390 7982 31442 8034
rect 32174 7982 32226 8034
rect 32622 7982 32674 8034
rect 33406 7982 33458 8034
rect 34974 7982 35026 8034
rect 36990 7982 37042 8034
rect 37774 7982 37826 8034
rect 39006 7982 39058 8034
rect 40126 7982 40178 8034
rect 40798 7982 40850 8034
rect 42142 7982 42194 8034
rect 42814 7982 42866 8034
rect 44046 7982 44098 8034
rect 44270 7982 44322 8034
rect 19838 7814 19890 7866
rect 19942 7814 19994 7866
rect 20046 7814 20098 7866
rect 6638 7646 6690 7698
rect 7086 7646 7138 7698
rect 19406 7646 19458 7698
rect 20078 7646 20130 7698
rect 26014 7646 26066 7698
rect 27918 7646 27970 7698
rect 32174 7646 32226 7698
rect 37214 7646 37266 7698
rect 38222 7646 38274 7698
rect 45278 7646 45330 7698
rect 4062 7534 4114 7586
rect 13246 7534 13298 7586
rect 19070 7534 19122 7586
rect 19742 7534 19794 7586
rect 21422 7534 21474 7586
rect 21982 7534 22034 7586
rect 26350 7534 26402 7586
rect 27134 7534 27186 7586
rect 36766 7534 36818 7586
rect 39902 7534 39954 7586
rect 40910 7534 40962 7586
rect 42142 7534 42194 7586
rect 3278 7422 3330 7474
rect 6526 7422 6578 7474
rect 9886 7422 9938 7474
rect 13134 7422 13186 7474
rect 13694 7422 13746 7474
rect 17950 7422 18002 7474
rect 21198 7422 21250 7474
rect 26574 7422 26626 7474
rect 27470 7422 27522 7474
rect 28366 7422 28418 7474
rect 28926 7422 28978 7474
rect 35422 7422 35474 7474
rect 35982 7422 36034 7474
rect 36430 7422 36482 7474
rect 38446 7422 38498 7474
rect 39566 7422 39618 7474
rect 41470 7422 41522 7474
rect 44718 7422 44770 7474
rect 44942 7422 44994 7474
rect 45726 7422 45778 7474
rect 6190 7310 6242 7362
rect 7534 7310 7586 7362
rect 8654 7310 8706 7362
rect 9102 7310 9154 7362
rect 10670 7310 10722 7362
rect 12798 7310 12850 7362
rect 14478 7310 14530 7362
rect 16606 7310 16658 7362
rect 17502 7310 17554 7362
rect 18398 7310 18450 7362
rect 18958 7310 19010 7362
rect 20190 7310 20242 7362
rect 22766 7310 22818 7362
rect 23550 7310 23602 7362
rect 24446 7310 24498 7362
rect 31278 7310 31330 7362
rect 31614 7310 31666 7362
rect 33070 7310 33122 7362
rect 37662 7310 37714 7362
rect 39342 7310 39394 7362
rect 40350 7310 40402 7362
rect 44270 7310 44322 7362
rect 47966 7310 48018 7362
rect 7422 7198 7474 7250
rect 13246 7198 13298 7250
rect 20862 7198 20914 7250
rect 22654 7198 22706 7250
rect 27470 7198 27522 7250
rect 31726 7198 31778 7250
rect 40238 7198 40290 7250
rect 41022 7198 41074 7250
rect 4478 7030 4530 7082
rect 4582 7030 4634 7082
rect 4686 7030 4738 7082
rect 35198 7030 35250 7082
rect 35302 7030 35354 7082
rect 35406 7030 35458 7082
rect 11566 6862 11618 6914
rect 31054 6862 31106 6914
rect 35310 6862 35362 6914
rect 7198 6750 7250 6802
rect 9326 6750 9378 6802
rect 11678 6750 11730 6802
rect 12126 6750 12178 6802
rect 19854 6750 19906 6802
rect 23214 6750 23266 6802
rect 27806 6750 27858 6802
rect 30718 6750 30770 6802
rect 32174 6750 32226 6802
rect 32958 6750 33010 6802
rect 38782 6750 38834 6802
rect 39342 6750 39394 6802
rect 43486 6750 43538 6802
rect 48190 6750 48242 6802
rect 6526 6638 6578 6690
rect 9774 6638 9826 6690
rect 10222 6638 10274 6690
rect 10670 6638 10722 6690
rect 12910 6638 12962 6690
rect 13694 6638 13746 6690
rect 17054 6638 17106 6690
rect 21982 6638 22034 6690
rect 23662 6638 23714 6690
rect 24782 6638 24834 6690
rect 25454 6638 25506 6690
rect 29486 6638 29538 6690
rect 29710 6638 29762 6690
rect 30382 6638 30434 6690
rect 32286 6638 32338 6690
rect 33294 6638 33346 6690
rect 34078 6638 34130 6690
rect 34302 6638 34354 6690
rect 34638 6638 34690 6690
rect 37886 6638 37938 6690
rect 38222 6638 38274 6690
rect 38446 6638 38498 6690
rect 39118 6638 39170 6690
rect 40574 6638 40626 6690
rect 45390 6638 45442 6690
rect 46062 6638 46114 6690
rect 11006 6526 11058 6578
rect 12462 6526 12514 6578
rect 12574 6526 12626 6578
rect 17726 6526 17778 6578
rect 23102 6526 23154 6578
rect 23214 6526 23266 6578
rect 23998 6526 24050 6578
rect 24334 6526 24386 6578
rect 33070 6526 33122 6578
rect 35198 6526 35250 6578
rect 36318 6526 36370 6578
rect 37326 6526 37378 6578
rect 40126 6526 40178 6578
rect 43710 6526 43762 6578
rect 43934 6526 43986 6578
rect 44270 6526 44322 6578
rect 44942 6526 44994 6578
rect 11118 6414 11170 6466
rect 11342 6414 11394 6466
rect 12686 6414 12738 6466
rect 14702 6414 14754 6466
rect 20302 6414 20354 6466
rect 20750 6414 20802 6466
rect 21422 6414 21474 6466
rect 22206 6414 22258 6466
rect 22542 6414 22594 6466
rect 22878 6414 22930 6466
rect 24110 6414 24162 6466
rect 28702 6414 28754 6466
rect 30158 6414 30210 6466
rect 30270 6414 30322 6466
rect 30830 6414 30882 6466
rect 31838 6414 31890 6466
rect 32062 6414 32114 6466
rect 34526 6414 34578 6466
rect 35758 6414 35810 6466
rect 36430 6414 36482 6466
rect 37438 6414 37490 6466
rect 37662 6414 37714 6466
rect 37998 6414 38050 6466
rect 40238 6414 40290 6466
rect 41582 6414 41634 6466
rect 44046 6414 44098 6466
rect 44830 6414 44882 6466
rect 19838 6246 19890 6298
rect 19942 6246 19994 6298
rect 20046 6246 20098 6298
rect 6302 6078 6354 6130
rect 6638 6078 6690 6130
rect 7422 6078 7474 6130
rect 7534 6078 7586 6130
rect 7646 6078 7698 6130
rect 8654 6078 8706 6130
rect 9774 6078 9826 6130
rect 11454 6078 11506 6130
rect 12350 6078 12402 6130
rect 12910 6078 12962 6130
rect 22542 6078 22594 6130
rect 22766 6078 22818 6130
rect 26350 6078 26402 6130
rect 27470 6078 27522 6130
rect 27694 6078 27746 6130
rect 29486 6078 29538 6130
rect 33182 6078 33234 6130
rect 33294 6078 33346 6130
rect 39454 6078 39506 6130
rect 46958 6078 47010 6130
rect 1710 5966 1762 6018
rect 7758 5966 7810 6018
rect 10782 5966 10834 6018
rect 11902 5966 11954 6018
rect 13134 5966 13186 6018
rect 13582 5966 13634 6018
rect 17502 5966 17554 6018
rect 19294 5966 19346 6018
rect 20078 5966 20130 6018
rect 21646 5966 21698 6018
rect 23102 5966 23154 6018
rect 23886 5966 23938 6018
rect 25790 5966 25842 6018
rect 28926 5966 28978 6018
rect 30382 5966 30434 6018
rect 31166 5966 31218 6018
rect 31502 5966 31554 6018
rect 32062 5966 32114 6018
rect 32398 5966 32450 6018
rect 33406 5966 33458 6018
rect 33742 5966 33794 6018
rect 33854 5966 33906 6018
rect 34414 5966 34466 6018
rect 36542 5966 36594 6018
rect 39790 5966 39842 6018
rect 40350 5966 40402 6018
rect 47294 5966 47346 6018
rect 48190 5966 48242 6018
rect 7086 5854 7138 5906
rect 8206 5854 8258 5906
rect 8542 5854 8594 5906
rect 9998 5854 10050 5906
rect 10446 5854 10498 5906
rect 11118 5854 11170 5906
rect 11790 5854 11842 5906
rect 12686 5854 12738 5906
rect 13246 5854 13298 5906
rect 13918 5854 13970 5906
rect 16718 5854 16770 5906
rect 17614 5854 17666 5906
rect 17950 5854 18002 5906
rect 19070 5854 19122 5906
rect 19854 5854 19906 5906
rect 20526 5854 20578 5906
rect 20862 5854 20914 5906
rect 21310 5854 21362 5906
rect 22206 5854 22258 5906
rect 22318 5854 22370 5906
rect 22766 5854 22818 5906
rect 23438 5854 23490 5906
rect 23774 5854 23826 5906
rect 26238 5854 26290 5906
rect 26462 5854 26514 5906
rect 26798 5854 26850 5906
rect 27022 5854 27074 5906
rect 27582 5854 27634 5906
rect 28590 5854 28642 5906
rect 29374 5854 29426 5906
rect 29598 5854 29650 5906
rect 30046 5854 30098 5906
rect 30494 5854 30546 5906
rect 34190 5854 34242 5906
rect 34526 5854 34578 5906
rect 35310 5854 35362 5906
rect 35870 5854 35922 5906
rect 39118 5854 39170 5906
rect 39902 5854 39954 5906
rect 40126 5854 40178 5906
rect 40910 5854 40962 5906
rect 43822 5854 43874 5906
rect 46734 5854 46786 5906
rect 47182 5854 47234 5906
rect 47854 5854 47906 5906
rect 5854 5742 5906 5794
rect 6974 5742 7026 5794
rect 14702 5742 14754 5794
rect 18062 5742 18114 5794
rect 18510 5742 18562 5794
rect 24446 5742 24498 5794
rect 25342 5742 25394 5794
rect 28142 5742 28194 5794
rect 34974 5742 35026 5794
rect 35422 5742 35474 5794
rect 38670 5742 38722 5794
rect 42030 5742 42082 5794
rect 47070 5742 47122 5794
rect 8654 5630 8706 5682
rect 11902 5630 11954 5682
rect 17502 5630 17554 5682
rect 18398 5630 18450 5682
rect 23886 5630 23938 5682
rect 25230 5630 25282 5682
rect 25902 5630 25954 5682
rect 29038 5630 29090 5682
rect 30382 5630 30434 5682
rect 33854 5630 33906 5682
rect 34862 5630 34914 5682
rect 44830 5630 44882 5682
rect 4478 5462 4530 5514
rect 4582 5462 4634 5514
rect 4686 5462 4738 5514
rect 35198 5462 35250 5514
rect 35302 5462 35354 5514
rect 35406 5462 35458 5514
rect 21534 5294 21586 5346
rect 21982 5294 22034 5346
rect 22094 5294 22146 5346
rect 22430 5294 22482 5346
rect 35198 5294 35250 5346
rect 37662 5294 37714 5346
rect 38894 5294 38946 5346
rect 10334 5182 10386 5234
rect 15150 5182 15202 5234
rect 16942 5182 16994 5234
rect 19070 5182 19122 5234
rect 20078 5182 20130 5234
rect 20750 5182 20802 5234
rect 21422 5182 21474 5234
rect 24222 5182 24274 5234
rect 26350 5182 26402 5234
rect 26798 5182 26850 5234
rect 28590 5182 28642 5234
rect 29150 5182 29202 5234
rect 32622 5182 32674 5234
rect 34750 5182 34802 5234
rect 36318 5182 36370 5234
rect 40126 5182 40178 5234
rect 42254 5182 42306 5234
rect 42702 5182 42754 5234
rect 5630 5070 5682 5122
rect 6414 5070 6466 5122
rect 6974 5070 7026 5122
rect 7422 5070 7474 5122
rect 8206 5070 8258 5122
rect 10670 5070 10722 5122
rect 11118 5070 11170 5122
rect 11342 5070 11394 5122
rect 12014 5070 12066 5122
rect 12798 5070 12850 5122
rect 13470 5070 13522 5122
rect 13806 5070 13858 5122
rect 14814 5070 14866 5122
rect 15038 5070 15090 5122
rect 16158 5070 16210 5122
rect 20190 5070 20242 5122
rect 22318 5070 22370 5122
rect 22878 5070 22930 5122
rect 23550 5070 23602 5122
rect 26686 5070 26738 5122
rect 27246 5070 27298 5122
rect 28030 5070 28082 5122
rect 29262 5070 29314 5122
rect 29486 5070 29538 5122
rect 30606 5070 30658 5122
rect 31054 5070 31106 5122
rect 31950 5070 32002 5122
rect 35646 5070 35698 5122
rect 36430 5070 36482 5122
rect 37102 5070 37154 5122
rect 37774 5070 37826 5122
rect 38110 5070 38162 5122
rect 39454 5070 39506 5122
rect 42590 5070 42642 5122
rect 43262 5070 43314 5122
rect 43710 5070 43762 5122
rect 44270 5070 44322 5122
rect 45054 5070 45106 5122
rect 47966 5070 48018 5122
rect 5070 4958 5122 5010
rect 6526 4958 6578 5010
rect 6638 4958 6690 5010
rect 10894 4958 10946 5010
rect 11790 4958 11842 5010
rect 12574 4958 12626 5010
rect 15262 4958 15314 5010
rect 19406 4958 19458 5010
rect 19742 4958 19794 5010
rect 23102 4958 23154 5010
rect 27806 4958 27858 5010
rect 29710 4958 29762 5010
rect 35310 4958 35362 5010
rect 36094 4958 36146 5010
rect 37326 4958 37378 5010
rect 38782 4958 38834 5010
rect 42926 4958 42978 5010
rect 47742 4958 47794 5010
rect 1710 4846 1762 4898
rect 5742 4846 5794 4898
rect 6302 4846 6354 4898
rect 10782 4846 10834 4898
rect 14030 4846 14082 4898
rect 14142 4846 14194 4898
rect 14254 4846 14306 4898
rect 15486 4846 15538 4898
rect 28478 4846 28530 4898
rect 29934 4846 29986 4898
rect 30270 4846 30322 4898
rect 31278 4846 31330 4898
rect 35198 4846 35250 4898
rect 36206 4846 36258 4898
rect 38222 4846 38274 4898
rect 38894 4846 38946 4898
rect 42814 4846 42866 4898
rect 45838 4846 45890 4898
rect 19838 4678 19890 4730
rect 19942 4678 19994 4730
rect 20046 4678 20098 4730
rect 4062 4510 4114 4562
rect 7534 4510 7586 4562
rect 8094 4510 8146 4562
rect 8542 4510 8594 4562
rect 17950 4510 18002 4562
rect 18062 4510 18114 4562
rect 21982 4510 22034 4562
rect 22094 4510 22146 4562
rect 22206 4510 22258 4562
rect 23438 4510 23490 4562
rect 24110 4510 24162 4562
rect 24558 4510 24610 4562
rect 25790 4510 25842 4562
rect 26014 4510 26066 4562
rect 33070 4510 33122 4562
rect 34078 4510 34130 4562
rect 34302 4510 34354 4562
rect 34638 4510 34690 4562
rect 36094 4510 36146 4562
rect 36318 4510 36370 4562
rect 40238 4510 40290 4562
rect 40462 4510 40514 4562
rect 43934 4510 43986 4562
rect 44158 4510 44210 4562
rect 47630 4510 47682 4562
rect 1710 4398 1762 4450
rect 6302 4398 6354 4450
rect 8430 4398 8482 4450
rect 8878 4398 8930 4450
rect 17838 4398 17890 4450
rect 19406 4398 19458 4450
rect 22318 4398 22370 4450
rect 23774 4398 23826 4450
rect 24670 4398 24722 4450
rect 25678 4398 25730 4450
rect 27470 4398 27522 4450
rect 33854 4398 33906 4450
rect 33966 4398 34018 4450
rect 34974 4398 35026 4450
rect 35982 4398 36034 4450
rect 38782 4398 38834 4450
rect 40126 4398 40178 4450
rect 43822 4398 43874 4450
rect 45166 4398 45218 4450
rect 7086 4286 7138 4338
rect 7422 4286 7474 4338
rect 9662 4286 9714 4338
rect 12910 4286 12962 4338
rect 16606 4286 16658 4338
rect 17502 4286 17554 4338
rect 18174 4286 18226 4338
rect 18734 4286 18786 4338
rect 22766 4286 22818 4338
rect 23102 4286 23154 4338
rect 25230 4286 25282 4338
rect 26798 4286 26850 4338
rect 29934 4286 29986 4338
rect 35534 4286 35586 4338
rect 39566 4286 39618 4338
rect 41134 4286 41186 4338
rect 44494 4286 44546 4338
rect 47854 4286 47906 4338
rect 7982 4174 8034 4226
rect 8990 4174 9042 4226
rect 13694 4174 13746 4226
rect 15822 4174 15874 4226
rect 16270 4174 16322 4226
rect 21534 4174 21586 4226
rect 25678 4174 25730 4226
rect 29598 4174 29650 4226
rect 33182 4174 33234 4226
rect 34190 4174 34242 4226
rect 35982 4174 36034 4226
rect 36654 4174 36706 4226
rect 42030 4174 42082 4226
rect 47294 4174 47346 4226
rect 7534 4062 7586 4114
rect 10670 4062 10722 4114
rect 24558 4062 24610 4114
rect 30942 4062 30994 4114
rect 4478 3894 4530 3946
rect 4582 3894 4634 3946
rect 4686 3894 4738 3946
rect 35198 3894 35250 3946
rect 35302 3894 35354 3946
rect 35406 3894 35458 3946
rect 6190 3726 6242 3778
rect 6638 3726 6690 3778
rect 4622 3614 4674 3666
rect 5070 3614 5122 3666
rect 5854 3614 5906 3666
rect 6526 3614 6578 3666
rect 16158 3614 16210 3666
rect 18622 3614 18674 3666
rect 22094 3614 22146 3666
rect 29374 3614 29426 3666
rect 33854 3614 33906 3666
rect 36990 3614 37042 3666
rect 40798 3614 40850 3666
rect 44606 3614 44658 3666
rect 48190 3614 48242 3666
rect 4174 3502 4226 3554
rect 7198 3502 7250 3554
rect 7870 3502 7922 3554
rect 8430 3502 8482 3554
rect 9550 3502 9602 3554
rect 10446 3502 10498 3554
rect 13470 3502 13522 3554
rect 14254 3502 14306 3554
rect 17054 3502 17106 3554
rect 17726 3502 17778 3554
rect 21086 3502 21138 3554
rect 24670 3502 24722 3554
rect 25454 3502 25506 3554
rect 28590 3502 28642 3554
rect 31278 3502 31330 3554
rect 32286 3502 32338 3554
rect 33294 3502 33346 3554
rect 36206 3502 36258 3554
rect 39118 3502 39170 3554
rect 40014 3502 40066 3554
rect 42702 3502 42754 3554
rect 43710 3502 43762 3554
rect 46734 3502 46786 3554
rect 47630 3502 47682 3554
rect 6078 3390 6130 3442
rect 6974 3390 7026 3442
rect 7646 3390 7698 3442
rect 8766 3390 8818 3442
rect 9326 3390 9378 3442
rect 11566 3390 11618 3442
rect 13134 3390 13186 3442
rect 17278 3390 17330 3442
rect 24894 3390 24946 3442
rect 26910 3390 26962 3442
rect 31614 3390 31666 3442
rect 32510 3390 32562 3442
rect 35982 3390 36034 3442
rect 43038 3390 43090 3442
rect 46510 3390 46562 3442
rect 47406 3390 47458 3442
rect 48078 3390 48130 3442
rect 1710 3278 1762 3330
rect 2158 3278 2210 3330
rect 19838 3110 19890 3162
rect 19942 3110 19994 3162
rect 20046 3110 20098 3162
<< metal2 >>
rect 13440 49200 13552 50000
rect 14784 49200 14896 50000
rect 18144 49200 18256 50000
rect 20160 49200 20272 50000
rect 22848 49200 22960 50000
rect 23520 49200 23632 50000
rect 25536 49200 25648 50000
rect 26208 49200 26320 50000
rect 26880 49200 26992 50000
rect 30240 49200 30352 50000
rect 30912 49200 31024 50000
rect 31584 49200 31696 50000
rect 32256 49200 32368 50000
rect 32928 49200 33040 50000
rect 33600 49200 33712 50000
rect 34944 49200 35056 50000
rect 36288 49200 36400 50000
rect 37632 49200 37744 50000
rect 38304 49200 38416 50000
rect 39648 49200 39760 50000
rect 44352 49200 44464 50000
rect 13468 47012 13524 49200
rect 13468 46956 13972 47012
rect 4476 46284 4740 46294
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4476 46218 4740 46228
rect 10668 46004 10724 46014
rect 10668 45910 10724 45948
rect 13916 46004 13972 46956
rect 14812 46116 14868 49200
rect 14812 46060 15316 46116
rect 13916 45890 13972 45948
rect 13916 45838 13918 45890
rect 13970 45838 13972 45890
rect 13916 45826 13972 45838
rect 15260 45892 15316 46060
rect 17724 46004 17780 46014
rect 18172 46004 18228 49200
rect 17724 46002 18228 46004
rect 17724 45950 17726 46002
rect 17778 45950 18228 46002
rect 17724 45948 18228 45950
rect 17724 45938 17780 45948
rect 15260 45798 15316 45836
rect 16268 45892 16324 45902
rect 18172 45892 18228 45948
rect 18396 45892 18452 45902
rect 18172 45890 18452 45892
rect 18172 45838 18398 45890
rect 18450 45838 18452 45890
rect 18172 45836 18452 45838
rect 16268 45798 16324 45836
rect 18396 45826 18452 45836
rect 19628 45890 19684 45902
rect 19628 45838 19630 45890
rect 19682 45838 19684 45890
rect 19404 45780 19460 45790
rect 19292 45778 19460 45780
rect 19292 45726 19406 45778
rect 19458 45726 19460 45778
rect 19292 45724 19460 45726
rect 1708 45666 1764 45678
rect 7420 45668 7476 45678
rect 1708 45614 1710 45666
rect 1762 45614 1764 45666
rect 1708 45444 1764 45614
rect 1708 45378 1764 45388
rect 7308 45612 7420 45668
rect 6188 44996 6244 45006
rect 4476 44716 4740 44726
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4476 44650 4740 44660
rect 1484 44100 1540 44110
rect 1372 39172 1428 39182
rect 1372 38668 1428 39116
rect 1260 38612 1428 38668
rect 1260 27972 1316 38612
rect 1484 36596 1540 44044
rect 4844 44098 4900 44110
rect 5852 44100 5908 44110
rect 4844 44046 4846 44098
rect 4898 44046 4900 44098
rect 3948 43652 4004 43662
rect 1820 43428 1876 43438
rect 1708 43426 1876 43428
rect 1708 43374 1822 43426
rect 1874 43374 1876 43426
rect 1708 43372 1876 43374
rect 1708 42196 1764 43372
rect 1820 43362 1876 43372
rect 2268 43426 2324 43438
rect 2268 43374 2270 43426
rect 2322 43374 2324 43426
rect 1820 42532 1876 42542
rect 2156 42532 2212 42542
rect 1820 42530 1988 42532
rect 1820 42478 1822 42530
rect 1874 42478 1988 42530
rect 1820 42476 1988 42478
rect 1820 42466 1876 42476
rect 1708 42140 1876 42196
rect 1708 41972 1764 41982
rect 1708 41524 1764 41916
rect 1596 41468 1764 41524
rect 1596 40404 1652 41468
rect 1820 41412 1876 42140
rect 1596 40338 1652 40348
rect 1708 41356 1876 41412
rect 1708 39618 1764 41356
rect 1708 39566 1710 39618
rect 1762 39566 1764 39618
rect 1708 38388 1764 39566
rect 1708 38322 1764 38332
rect 1820 40964 1876 40974
rect 1820 40402 1876 40908
rect 1820 40350 1822 40402
rect 1874 40350 1876 40402
rect 1820 38834 1876 40350
rect 1820 38782 1822 38834
rect 1874 38782 1876 38834
rect 1708 38052 1764 38062
rect 1708 37958 1764 37996
rect 1372 36540 1540 36596
rect 1708 37266 1764 37278
rect 1708 37214 1710 37266
rect 1762 37214 1764 37266
rect 1708 36932 1764 37214
rect 1372 33236 1428 36540
rect 1708 35700 1764 36876
rect 1820 36482 1876 38782
rect 1932 36820 1988 42476
rect 2156 41186 2212 42476
rect 2268 42084 2324 43374
rect 3948 43426 4004 43596
rect 4844 43652 4900 44046
rect 5740 44098 5908 44100
rect 5740 44046 5854 44098
rect 5906 44046 5908 44098
rect 5740 44044 5908 44046
rect 4844 43586 4900 43596
rect 5628 43652 5684 43662
rect 4396 43428 4452 43438
rect 3948 43374 3950 43426
rect 4002 43374 4004 43426
rect 3836 43314 3892 43326
rect 3836 43262 3838 43314
rect 3890 43262 3892 43314
rect 2268 42018 2324 42028
rect 2492 42530 2548 42542
rect 2940 42532 2996 42542
rect 2492 42478 2494 42530
rect 2546 42478 2548 42530
rect 2268 41858 2324 41870
rect 2268 41806 2270 41858
rect 2322 41806 2324 41858
rect 2268 41412 2324 41806
rect 2268 41346 2324 41356
rect 2156 41134 2158 41186
rect 2210 41134 2212 41186
rect 2156 40964 2212 41134
rect 2156 40898 2212 40908
rect 2492 40628 2548 42478
rect 2380 40572 2548 40628
rect 2828 42530 2996 42532
rect 2828 42478 2942 42530
rect 2994 42478 2996 42530
rect 2828 42476 2996 42478
rect 2268 39844 2324 39854
rect 2268 39730 2324 39788
rect 2268 39678 2270 39730
rect 2322 39678 2324 39730
rect 2268 39666 2324 39678
rect 2380 38668 2436 40572
rect 2492 40292 2548 40302
rect 2492 40198 2548 40236
rect 2604 39732 2660 39742
rect 2604 39618 2660 39676
rect 2604 39566 2606 39618
rect 2658 39566 2660 39618
rect 2604 39554 2660 39566
rect 2156 38612 2436 38668
rect 2492 38722 2548 38734
rect 2492 38670 2494 38722
rect 2546 38670 2548 38722
rect 2492 38668 2548 38670
rect 2828 38668 2884 42476
rect 2940 42466 2996 42476
rect 3388 42532 3444 42542
rect 3388 42530 3668 42532
rect 3388 42478 3390 42530
rect 3442 42478 3668 42530
rect 3388 42476 3668 42478
rect 3388 42466 3444 42476
rect 3164 41860 3220 41870
rect 3052 41858 3220 41860
rect 3052 41806 3166 41858
rect 3218 41806 3220 41858
rect 3052 41804 3220 41806
rect 2940 41074 2996 41086
rect 2940 41022 2942 41074
rect 2994 41022 2996 41074
rect 2940 40180 2996 41022
rect 2940 40114 2996 40124
rect 2940 39508 2996 39518
rect 2940 39414 2996 39452
rect 2492 38612 2772 38668
rect 2828 38612 2996 38668
rect 2044 37378 2100 37390
rect 2044 37326 2046 37378
rect 2098 37326 2100 37378
rect 2044 37044 2100 37326
rect 2044 36978 2100 36988
rect 1932 36764 2100 36820
rect 1820 36430 1822 36482
rect 1874 36430 1876 36482
rect 1820 36418 1876 36430
rect 1708 35634 1764 35644
rect 1932 35586 1988 35598
rect 1932 35534 1934 35586
rect 1986 35534 1988 35586
rect 1820 35252 1876 35262
rect 1708 34916 1764 34926
rect 1708 34132 1764 34860
rect 1820 34914 1876 35196
rect 1820 34862 1822 34914
rect 1874 34862 1876 34914
rect 1820 34850 1876 34862
rect 1596 34130 1764 34132
rect 1596 34078 1710 34130
rect 1762 34078 1764 34130
rect 1596 34076 1764 34078
rect 1596 34020 1652 34076
rect 1708 34066 1764 34076
rect 1820 34580 1876 34590
rect 1372 33170 1428 33180
rect 1484 33964 1652 34020
rect 1484 32340 1540 33964
rect 1708 33908 1764 33918
rect 1708 33234 1764 33852
rect 1708 33182 1710 33234
rect 1762 33182 1764 33234
rect 1708 33124 1764 33182
rect 1484 32274 1540 32284
rect 1596 33068 1764 33124
rect 1596 30772 1652 33068
rect 1820 33012 1876 34524
rect 1708 32956 1876 33012
rect 1708 31778 1764 32956
rect 1708 31726 1710 31778
rect 1762 31726 1764 31778
rect 1708 30996 1764 31726
rect 1820 32564 1876 32574
rect 1932 32564 1988 35534
rect 2044 33908 2100 36764
rect 2156 35252 2212 38612
rect 2268 38164 2324 38174
rect 2268 38070 2324 38108
rect 2716 38162 2772 38612
rect 2716 38110 2718 38162
rect 2770 38110 2772 38162
rect 2716 38098 2772 38110
rect 2828 38050 2884 38062
rect 2828 37998 2830 38050
rect 2882 37998 2884 38050
rect 2828 37940 2884 37998
rect 2828 37874 2884 37884
rect 2604 37828 2660 37838
rect 2268 37826 2660 37828
rect 2268 37774 2606 37826
rect 2658 37774 2660 37826
rect 2268 37772 2660 37774
rect 2268 36260 2324 37772
rect 2604 37762 2660 37772
rect 2828 37492 2884 37502
rect 2492 37156 2548 37166
rect 2492 37154 2660 37156
rect 2492 37102 2494 37154
rect 2546 37102 2660 37154
rect 2492 37100 2660 37102
rect 2492 37090 2548 37100
rect 2492 36372 2548 36382
rect 2268 35922 2324 36204
rect 2268 35870 2270 35922
rect 2322 35870 2324 35922
rect 2268 35858 2324 35870
rect 2380 36370 2548 36372
rect 2380 36318 2494 36370
rect 2546 36318 2548 36370
rect 2380 36316 2548 36318
rect 2380 35922 2436 36316
rect 2492 36306 2548 36316
rect 2380 35870 2382 35922
rect 2434 35870 2436 35922
rect 2380 35858 2436 35870
rect 2156 35186 2212 35196
rect 2492 35698 2548 35710
rect 2492 35646 2494 35698
rect 2546 35646 2548 35698
rect 2268 35140 2324 35150
rect 2268 35026 2324 35084
rect 2268 34974 2270 35026
rect 2322 34974 2324 35026
rect 2268 34962 2324 34974
rect 2492 34356 2548 35646
rect 2604 34580 2660 37100
rect 2604 34514 2660 34524
rect 2716 35252 2772 35262
rect 2716 34914 2772 35196
rect 2716 34862 2718 34914
rect 2770 34862 2772 34914
rect 2604 34356 2660 34366
rect 2492 34300 2604 34356
rect 2604 34262 2660 34300
rect 2044 33842 2100 33852
rect 2268 34018 2324 34030
rect 2268 33966 2270 34018
rect 2322 33966 2324 34018
rect 2156 33348 2212 33358
rect 1820 32562 1988 32564
rect 1820 32510 1822 32562
rect 1874 32510 1988 32562
rect 1820 32508 1988 32510
rect 2044 33122 2100 33134
rect 2044 33070 2046 33122
rect 2098 33070 2100 33122
rect 1820 31668 1876 32508
rect 1820 31602 1876 31612
rect 1708 30930 1764 30940
rect 1932 30884 1988 30894
rect 2044 30884 2100 33070
rect 2156 31890 2212 33292
rect 2268 32900 2324 33966
rect 2604 33684 2660 33694
rect 2716 33684 2772 34862
rect 2828 34244 2884 37436
rect 2940 36932 2996 38612
rect 3052 37604 3108 41804
rect 3164 41794 3220 41804
rect 3388 40180 3444 40190
rect 3164 39844 3220 39854
rect 3164 38948 3220 39788
rect 3164 38882 3220 38892
rect 3276 39732 3332 39742
rect 3276 39618 3332 39676
rect 3388 39730 3444 40124
rect 3388 39678 3390 39730
rect 3442 39678 3444 39730
rect 3388 39666 3444 39678
rect 3500 40068 3556 40078
rect 3276 39566 3278 39618
rect 3330 39566 3332 39618
rect 3276 38668 3332 39566
rect 3500 39620 3556 40012
rect 3500 39554 3556 39564
rect 3500 39396 3556 39406
rect 3500 39302 3556 39340
rect 3612 39172 3668 42476
rect 3836 42308 3892 43262
rect 3948 42532 4004 43374
rect 3948 42438 4004 42476
rect 4060 43426 4452 43428
rect 4060 43374 4398 43426
rect 4450 43374 4452 43426
rect 4060 43372 4452 43374
rect 3836 42252 4004 42308
rect 3836 41972 3892 41982
rect 3836 41878 3892 41916
rect 3052 37538 3108 37548
rect 3164 38612 3332 38668
rect 3388 39116 3668 39172
rect 3724 40292 3780 40302
rect 3052 37380 3108 37390
rect 3052 37286 3108 37324
rect 2940 36866 2996 36876
rect 3164 36260 3220 38612
rect 3164 36194 3220 36204
rect 3276 38050 3332 38062
rect 3276 37998 3278 38050
rect 3330 37998 3332 38050
rect 2940 35698 2996 35710
rect 2940 35646 2942 35698
rect 2994 35646 2996 35698
rect 2940 34916 2996 35646
rect 3276 35700 3332 37998
rect 3388 38052 3444 39116
rect 3724 39060 3780 40236
rect 3948 39844 4004 42252
rect 4060 40068 4116 43372
rect 4396 43362 4452 43372
rect 4844 43428 4900 43438
rect 4844 43314 4900 43372
rect 4844 43262 4846 43314
rect 4898 43262 4900 43314
rect 4844 43250 4900 43262
rect 5404 43426 5460 43438
rect 5404 43374 5406 43426
rect 5458 43374 5460 43426
rect 4476 43148 4740 43158
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4476 43082 4740 43092
rect 4396 42532 4452 42542
rect 4844 42532 4900 42542
rect 4060 40002 4116 40012
rect 4172 42530 4452 42532
rect 4172 42478 4398 42530
rect 4450 42478 4452 42530
rect 4172 42476 4452 42478
rect 3948 39778 4004 39788
rect 3836 39620 3892 39630
rect 4060 39620 4116 39630
rect 3836 39618 4116 39620
rect 3836 39566 3838 39618
rect 3890 39566 4062 39618
rect 4114 39566 4116 39618
rect 3836 39564 4116 39566
rect 3836 39554 3892 39564
rect 4060 39554 4116 39564
rect 3612 39004 3780 39060
rect 3388 37986 3444 37996
rect 3500 38164 3556 38174
rect 3500 37380 3556 38108
rect 3612 38162 3668 39004
rect 4172 38948 4228 42476
rect 4396 42466 4452 42476
rect 4508 42530 4900 42532
rect 4508 42478 4846 42530
rect 4898 42478 4900 42530
rect 4508 42476 4900 42478
rect 4284 42084 4340 42094
rect 4284 41970 4340 42028
rect 4284 41918 4286 41970
rect 4338 41918 4340 41970
rect 4284 41906 4340 41918
rect 4508 41748 4564 42476
rect 4844 42466 4900 42476
rect 4844 42082 4900 42094
rect 4844 42030 4846 42082
rect 4898 42030 4900 42082
rect 4284 41692 4564 41748
rect 4620 41970 4676 41982
rect 4620 41918 4622 41970
rect 4674 41918 4676 41970
rect 4620 41748 4676 41918
rect 4844 41860 4900 42030
rect 5404 41972 5460 43374
rect 5628 42754 5684 43596
rect 5740 43428 5796 44044
rect 5852 44034 5908 44044
rect 6076 43652 6132 43662
rect 6188 43652 6244 44940
rect 7308 44324 7364 45612
rect 7420 45602 7476 45612
rect 8092 45668 8148 45678
rect 8092 45574 8148 45612
rect 9548 45666 9604 45678
rect 9548 45614 9550 45666
rect 9602 45614 9604 45666
rect 7420 44996 7476 45006
rect 7980 44996 8036 45006
rect 7420 44994 7588 44996
rect 7420 44942 7422 44994
rect 7474 44942 7588 44994
rect 7420 44940 7588 44942
rect 7420 44930 7476 44940
rect 7532 44882 7588 44940
rect 7980 44902 8036 44940
rect 8428 44996 8484 45006
rect 7532 44830 7534 44882
rect 7586 44830 7588 44882
rect 7420 44324 7476 44334
rect 7308 44322 7476 44324
rect 7308 44270 7422 44322
rect 7474 44270 7476 44322
rect 7308 44268 7476 44270
rect 7420 44258 7476 44268
rect 6132 43596 6244 43652
rect 6076 43586 6132 43596
rect 6188 43538 6244 43596
rect 6188 43486 6190 43538
rect 6242 43486 6244 43538
rect 6188 43474 6244 43486
rect 6412 44098 6468 44110
rect 6860 44100 6916 44110
rect 6412 44046 6414 44098
rect 6466 44046 6468 44098
rect 5740 43362 5796 43372
rect 5852 43428 5908 43438
rect 5852 43426 6132 43428
rect 5852 43374 5854 43426
rect 5906 43374 6132 43426
rect 5852 43372 6132 43374
rect 5852 43362 5908 43372
rect 6076 42868 6132 43372
rect 6412 42980 6468 44046
rect 6748 44098 6916 44100
rect 6748 44046 6862 44098
rect 6914 44046 6916 44098
rect 6748 44044 6916 44046
rect 6636 42980 6692 42990
rect 6412 42924 6636 42980
rect 6076 42812 6580 42868
rect 5628 42702 5630 42754
rect 5682 42702 5684 42754
rect 5628 42690 5684 42702
rect 6412 42644 6468 42654
rect 6412 42550 6468 42588
rect 6300 42308 6356 42318
rect 5404 41906 5460 41916
rect 5852 42082 5908 42094
rect 5852 42030 5854 42082
rect 5906 42030 5908 42082
rect 4956 41860 5012 41870
rect 4844 41804 4956 41860
rect 4956 41794 5012 41804
rect 4620 41692 4900 41748
rect 4284 39732 4340 41692
rect 4476 41580 4740 41590
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4476 41514 4740 41524
rect 4844 41300 4900 41692
rect 5068 41300 5124 41310
rect 4844 41298 5124 41300
rect 4844 41246 5070 41298
rect 5122 41246 5124 41298
rect 4844 41244 5124 41246
rect 5068 41076 5124 41244
rect 5852 41300 5908 42030
rect 5852 41206 5908 41244
rect 5068 41010 5124 41020
rect 5628 41186 5684 41198
rect 5628 41134 5630 41186
rect 5682 41134 5684 41186
rect 5628 40740 5684 41134
rect 5068 40684 5684 40740
rect 5740 41188 5796 41198
rect 5068 40402 5124 40684
rect 5068 40350 5070 40402
rect 5122 40350 5124 40402
rect 4620 40292 4676 40302
rect 5068 40292 5124 40350
rect 4620 40290 5124 40292
rect 4620 40238 4622 40290
rect 4674 40238 5124 40290
rect 4620 40236 5124 40238
rect 5292 40514 5348 40526
rect 5292 40462 5294 40514
rect 5346 40462 5348 40514
rect 4620 40226 4676 40236
rect 4476 40012 4740 40022
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4476 39946 4740 39956
rect 4284 39676 4564 39732
rect 4396 39506 4452 39518
rect 4396 39454 4398 39506
rect 4450 39454 4452 39506
rect 4284 39394 4340 39406
rect 4284 39342 4286 39394
rect 4338 39342 4340 39394
rect 4284 39060 4340 39342
rect 4396 39172 4452 39454
rect 4396 39106 4452 39116
rect 4284 38994 4340 39004
rect 3612 38110 3614 38162
rect 3666 38110 3668 38162
rect 3612 38098 3668 38110
rect 4060 38892 4228 38948
rect 3612 37828 3668 37838
rect 3612 37734 3668 37772
rect 3724 37828 3780 37838
rect 3724 37826 3892 37828
rect 3724 37774 3726 37826
rect 3778 37774 3892 37826
rect 3724 37772 3892 37774
rect 3724 37762 3780 37772
rect 3836 37716 3892 37772
rect 3612 37492 3668 37502
rect 3612 37398 3668 37436
rect 3388 37324 3556 37380
rect 3836 37378 3892 37660
rect 3948 37826 4004 37838
rect 3948 37774 3950 37826
rect 4002 37774 4004 37826
rect 3948 37492 4004 37774
rect 3948 37426 4004 37436
rect 3836 37326 3838 37378
rect 3890 37326 3892 37378
rect 3388 35924 3444 37324
rect 3500 37156 3556 37166
rect 3500 37062 3556 37100
rect 3724 37044 3780 37054
rect 3388 35868 3556 35924
rect 3276 35634 3332 35644
rect 3388 35698 3444 35710
rect 3388 35646 3390 35698
rect 3442 35646 3444 35698
rect 3276 35476 3332 35486
rect 3164 35474 3332 35476
rect 3164 35422 3278 35474
rect 3330 35422 3332 35474
rect 3164 35420 3332 35422
rect 3164 35308 3220 35420
rect 3276 35410 3332 35420
rect 2940 34850 2996 34860
rect 3052 35252 3220 35308
rect 2940 34692 2996 34702
rect 2940 34598 2996 34636
rect 2940 34356 2996 34366
rect 2940 34262 2996 34300
rect 2828 34178 2884 34188
rect 2660 33628 2772 33684
rect 2604 33618 2660 33628
rect 2268 32834 2324 32844
rect 2828 33572 2884 33582
rect 2828 33346 2884 33516
rect 2828 33294 2830 33346
rect 2882 33294 2884 33346
rect 2828 32674 2884 33294
rect 3052 32788 3108 35252
rect 3276 34802 3332 34814
rect 3276 34750 3278 34802
rect 3330 34750 3332 34802
rect 3276 33572 3332 34750
rect 3388 34804 3444 35646
rect 3500 35140 3556 35868
rect 3724 35698 3780 36988
rect 3724 35646 3726 35698
rect 3778 35646 3780 35698
rect 3724 35634 3780 35646
rect 3500 35084 3668 35140
rect 3612 35028 3668 35084
rect 3612 34962 3668 34972
rect 3836 35028 3892 37326
rect 3948 37266 4004 37278
rect 3948 37214 3950 37266
rect 4002 37214 4004 37266
rect 3948 37156 4004 37214
rect 3948 37090 4004 37100
rect 4060 35252 4116 38892
rect 4508 38724 4564 39676
rect 4844 39396 4900 39406
rect 4172 38668 4564 38724
rect 4620 39394 4900 39396
rect 4620 39342 4846 39394
rect 4898 39342 4900 39394
rect 4620 39340 4900 39342
rect 4172 38164 4228 38668
rect 4620 38612 4676 39340
rect 4844 39330 4900 39340
rect 5292 39060 5348 40462
rect 5292 38946 5348 39004
rect 5292 38894 5294 38946
rect 5346 38894 5348 38946
rect 5292 38882 5348 38894
rect 5404 39508 5460 39518
rect 4732 38836 4788 38846
rect 4732 38724 4788 38780
rect 5180 38724 5236 38734
rect 4732 38722 4900 38724
rect 4732 38670 4734 38722
rect 4786 38670 4900 38722
rect 4732 38668 4900 38670
rect 4732 38658 4788 38668
rect 4620 38546 4676 38556
rect 4476 38444 4740 38454
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4476 38378 4740 38388
rect 4172 38098 4228 38108
rect 4844 38162 4900 38668
rect 4844 38110 4846 38162
rect 4898 38110 4900 38162
rect 4844 38098 4900 38110
rect 4956 38722 5236 38724
rect 4956 38670 5182 38722
rect 5234 38670 5236 38722
rect 4956 38668 5236 38670
rect 4396 38052 4452 38062
rect 4284 37996 4396 38052
rect 4172 37940 4228 37950
rect 4284 37940 4340 37996
rect 4396 37986 4452 37996
rect 4956 38052 5012 38668
rect 5180 38658 5236 38668
rect 4172 37938 4340 37940
rect 4172 37886 4174 37938
rect 4226 37886 4340 37938
rect 4172 37884 4340 37886
rect 4508 37940 4564 37950
rect 4172 37874 4228 37884
rect 4172 37716 4228 37726
rect 4172 37268 4228 37660
rect 4172 37202 4228 37212
rect 4508 37044 4564 37884
rect 4956 37716 5012 37996
rect 4844 37660 5012 37716
rect 5180 37940 5236 37950
rect 4620 37266 4676 37278
rect 4620 37214 4622 37266
rect 4674 37214 4676 37266
rect 4620 37044 4676 37214
rect 4284 36988 4676 37044
rect 4732 37268 4788 37278
rect 4732 37154 4788 37212
rect 4732 37102 4734 37154
rect 4786 37102 4788 37154
rect 4732 37044 4788 37102
rect 4060 35186 4116 35196
rect 4172 36596 4228 36606
rect 3836 34962 3892 34972
rect 3948 35028 4004 35038
rect 4172 35028 4228 36540
rect 3948 35026 4228 35028
rect 3948 34974 3950 35026
rect 4002 34974 4228 35026
rect 3948 34972 4228 34974
rect 4284 35476 4340 36988
rect 4732 36978 4788 36988
rect 4844 37266 4900 37660
rect 5068 37604 5124 37614
rect 4844 37214 4846 37266
rect 4898 37214 4900 37266
rect 4476 36876 4740 36886
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4476 36810 4740 36820
rect 4620 36620 4676 36632
rect 4620 36568 4622 36620
rect 4674 36596 4676 36620
rect 4732 36596 4788 36606
rect 4674 36568 4732 36596
rect 4620 36540 4732 36568
rect 4732 36530 4788 36540
rect 4844 35810 4900 37214
rect 4844 35758 4846 35810
rect 4898 35758 4900 35810
rect 4844 35746 4900 35758
rect 4956 37492 5012 37502
rect 4508 35586 4564 35598
rect 4508 35534 4510 35586
rect 4562 35534 4564 35586
rect 4508 35476 4564 35534
rect 4284 35420 4564 35476
rect 3948 34962 4004 34972
rect 3388 34710 3444 34748
rect 3500 34916 3556 34926
rect 3500 34242 3556 34860
rect 3724 34916 3780 34926
rect 4284 34916 4340 35420
rect 4476 35308 4740 35318
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4476 35242 4740 35252
rect 3612 34692 3668 34702
rect 3612 34598 3668 34636
rect 3612 34468 3668 34478
rect 3612 34354 3668 34412
rect 3612 34302 3614 34354
rect 3666 34302 3668 34354
rect 3612 34290 3668 34302
rect 3500 34190 3502 34242
rect 3554 34190 3556 34242
rect 3500 34178 3556 34190
rect 3724 34242 3780 34860
rect 4060 34860 4340 34916
rect 3836 34690 3892 34702
rect 3836 34638 3838 34690
rect 3890 34638 3892 34690
rect 3836 34356 3892 34638
rect 3836 34290 3892 34300
rect 3724 34190 3726 34242
rect 3778 34190 3780 34242
rect 3724 34178 3780 34190
rect 3276 33506 3332 33516
rect 3388 34130 3444 34142
rect 3388 34078 3390 34130
rect 3442 34078 3444 34130
rect 3388 33908 3444 34078
rect 3276 33348 3332 33358
rect 3388 33348 3444 33852
rect 3836 33572 3892 33582
rect 3612 33460 3668 33470
rect 3612 33366 3668 33404
rect 2828 32622 2830 32674
rect 2882 32622 2884 32674
rect 2828 32610 2884 32622
rect 2940 32676 2996 32686
rect 2940 32582 2996 32620
rect 3052 32674 3108 32732
rect 3052 32622 3054 32674
rect 3106 32622 3108 32674
rect 3052 32610 3108 32622
rect 3164 33346 3444 33348
rect 3164 33294 3278 33346
rect 3330 33294 3444 33346
rect 3164 33292 3444 33294
rect 2268 32452 2324 32462
rect 2268 32358 2324 32396
rect 2156 31838 2158 31890
rect 2210 31838 2212 31890
rect 2156 31826 2212 31838
rect 3164 31780 3220 33292
rect 3276 33254 3332 33292
rect 3836 33124 3892 33516
rect 3836 33058 3892 33068
rect 3612 32788 3668 32798
rect 3612 32564 3668 32732
rect 3948 32676 4004 32686
rect 3948 32582 4004 32620
rect 3836 32564 3892 32574
rect 3612 32562 3892 32564
rect 3612 32510 3838 32562
rect 3890 32510 3892 32562
rect 3612 32508 3892 32510
rect 3500 32338 3556 32350
rect 3500 32286 3502 32338
rect 3554 32286 3556 32338
rect 3164 31714 3220 31724
rect 3388 31890 3444 31902
rect 3388 31838 3390 31890
rect 3442 31838 3444 31890
rect 3276 31668 3332 31678
rect 3276 31574 3332 31612
rect 2828 31554 2884 31566
rect 2828 31502 2830 31554
rect 2882 31502 2884 31554
rect 2380 31106 2436 31118
rect 2380 31054 2382 31106
rect 2434 31054 2436 31106
rect 2380 30996 2436 31054
rect 2380 30930 2436 30940
rect 1932 30882 2100 30884
rect 1932 30830 1934 30882
rect 1986 30830 2100 30882
rect 1932 30828 2100 30830
rect 1596 30716 1876 30772
rect 1820 30324 1876 30716
rect 1820 30258 1876 30268
rect 1708 30212 1764 30222
rect 1708 29426 1764 30156
rect 1708 29374 1710 29426
rect 1762 29374 1764 29426
rect 1708 28308 1764 29374
rect 1820 29204 1876 29214
rect 1820 28420 1876 29148
rect 1932 28644 1988 30828
rect 2492 30098 2548 30110
rect 2492 30046 2494 30098
rect 2546 30046 2548 30098
rect 2492 29652 2548 30046
rect 2492 29586 2548 29596
rect 2044 29540 2100 29550
rect 2716 29540 2772 29550
rect 2044 29538 2324 29540
rect 2044 29486 2046 29538
rect 2098 29486 2324 29538
rect 2044 29484 2324 29486
rect 2044 29474 2100 29484
rect 2156 28644 2212 28654
rect 1932 28642 2212 28644
rect 1932 28590 2158 28642
rect 2210 28590 2212 28642
rect 1932 28588 2212 28590
rect 2156 28578 2212 28588
rect 1932 28420 1988 28430
rect 1820 28418 1988 28420
rect 1820 28366 1934 28418
rect 1986 28366 1988 28418
rect 1820 28364 1988 28366
rect 1932 28354 1988 28364
rect 1708 28242 1764 28252
rect 2268 28308 2324 29484
rect 2716 29446 2772 29484
rect 2492 29428 2548 29438
rect 2492 29334 2548 29372
rect 2604 29426 2660 29438
rect 2604 29374 2606 29426
rect 2658 29374 2660 29426
rect 2604 28756 2660 29374
rect 2828 29428 2884 31502
rect 2828 29362 2884 29372
rect 3164 29428 3220 29438
rect 3388 29428 3444 31838
rect 3500 31332 3556 32286
rect 3724 31778 3780 32508
rect 3836 32498 3892 32508
rect 4060 32452 4116 34860
rect 4396 34804 4452 34814
rect 4172 34132 4228 34142
rect 4396 34132 4452 34748
rect 4732 34692 4788 34702
rect 4732 34690 4900 34692
rect 4732 34638 4734 34690
rect 4786 34638 4900 34690
rect 4732 34636 4900 34638
rect 4732 34626 4788 34636
rect 4732 34356 4788 34366
rect 4732 34262 4788 34300
rect 4172 34130 4340 34132
rect 4172 34078 4174 34130
rect 4226 34078 4340 34130
rect 4172 34076 4340 34078
rect 4172 34066 4228 34076
rect 4172 33460 4228 33470
rect 4172 33366 4228 33404
rect 4284 33348 4340 34076
rect 4396 34066 4452 34076
rect 4476 33740 4740 33750
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4476 33674 4740 33684
rect 4844 33572 4900 34636
rect 4844 33506 4900 33516
rect 4844 33348 4900 33358
rect 4956 33348 5012 37436
rect 5068 36594 5124 37548
rect 5068 36542 5070 36594
rect 5122 36542 5124 36594
rect 5068 36530 5124 36542
rect 5068 35812 5124 35822
rect 5068 35028 5124 35756
rect 5068 34934 5124 34972
rect 5180 34356 5236 37884
rect 5180 34290 5236 34300
rect 5068 34132 5124 34142
rect 5404 34132 5460 39452
rect 5740 38836 5796 41132
rect 6300 40626 6356 42252
rect 6300 40574 6302 40626
rect 6354 40574 6356 40626
rect 5964 40514 6020 40526
rect 5964 40462 5966 40514
rect 6018 40462 6020 40514
rect 5964 39732 6020 40462
rect 6300 40516 6356 40574
rect 6300 40450 6356 40460
rect 6188 40404 6244 40414
rect 6188 39844 6244 40348
rect 6300 39844 6356 39854
rect 6188 39842 6356 39844
rect 6188 39790 6302 39842
rect 6354 39790 6356 39842
rect 6188 39788 6356 39790
rect 6300 39778 6356 39788
rect 5964 39666 6020 39676
rect 5852 39620 5908 39630
rect 5852 39508 5908 39564
rect 5964 39508 6020 39518
rect 5852 39506 6020 39508
rect 5852 39454 5966 39506
rect 6018 39454 6020 39506
rect 5852 39452 6020 39454
rect 5964 39442 6020 39452
rect 6188 39508 6244 39518
rect 6188 39414 6244 39452
rect 6524 39284 6580 42812
rect 6636 42308 6692 42924
rect 6636 42242 6692 42252
rect 6748 42084 6804 44044
rect 6860 44034 6916 44044
rect 7196 44100 7252 44110
rect 7196 44006 7252 44044
rect 7308 44098 7364 44110
rect 7308 44046 7310 44098
rect 7362 44046 7364 44098
rect 7308 43764 7364 44046
rect 6860 43708 7364 43764
rect 6860 43650 6916 43708
rect 6860 43598 6862 43650
rect 6914 43598 6916 43650
rect 6860 43586 6916 43598
rect 7532 42756 7588 44830
rect 8428 44882 8484 44940
rect 9100 44994 9156 45006
rect 9100 44942 9102 44994
rect 9154 44942 9156 44994
rect 8428 44830 8430 44882
rect 8482 44830 8484 44882
rect 8428 44818 8484 44830
rect 8764 44884 8820 44894
rect 7868 44324 7924 44334
rect 8092 44324 8148 44334
rect 7868 44322 8148 44324
rect 7868 44270 7870 44322
rect 7922 44270 8094 44322
rect 8146 44270 8148 44322
rect 7868 44268 8148 44270
rect 7868 44258 7924 44268
rect 8092 44258 8148 44268
rect 8764 44322 8820 44828
rect 8764 44270 8766 44322
rect 8818 44270 8820 44322
rect 8764 44258 8820 44270
rect 8428 44212 8484 44222
rect 8428 44118 8484 44156
rect 8316 44100 8372 44110
rect 8316 44006 8372 44044
rect 8988 44100 9044 44110
rect 6636 42028 6804 42084
rect 7308 42700 7588 42756
rect 8988 43426 9044 44044
rect 8988 43374 8990 43426
rect 9042 43374 9044 43426
rect 6636 41636 6692 42028
rect 6972 41970 7028 41982
rect 6972 41918 6974 41970
rect 7026 41918 7028 41970
rect 6748 41860 6804 41870
rect 6972 41860 7028 41918
rect 7308 41860 7364 42700
rect 8652 42532 8708 42542
rect 8428 42476 8652 42532
rect 7980 42196 8036 42206
rect 7980 42102 8036 42140
rect 7420 41972 7476 41982
rect 7420 41878 7476 41916
rect 6804 41804 6916 41860
rect 6972 41804 7364 41860
rect 6748 41794 6804 41804
rect 6636 41580 6804 41636
rect 6636 40290 6692 40302
rect 6636 40238 6638 40290
rect 6690 40238 6692 40290
rect 6636 40180 6692 40238
rect 6636 40114 6692 40124
rect 6748 39620 6804 41580
rect 6860 39620 6916 41804
rect 6972 41300 7028 41310
rect 6972 39732 7028 41244
rect 7084 41076 7140 41086
rect 7084 40982 7140 41020
rect 7196 41076 7252 41804
rect 7420 41076 7476 41086
rect 7196 41020 7420 41076
rect 7196 40626 7252 41020
rect 7196 40574 7198 40626
rect 7250 40574 7252 40626
rect 7196 40562 7252 40574
rect 7420 39842 7476 41020
rect 7980 41074 8036 41086
rect 7980 41022 7982 41074
rect 8034 41022 8036 41074
rect 7980 40628 8036 41022
rect 7980 40562 8036 40572
rect 8092 40740 8148 40750
rect 7420 39790 7422 39842
rect 7474 39790 7476 39842
rect 7420 39778 7476 39790
rect 7532 40292 7588 40302
rect 8092 40292 8148 40684
rect 7532 39844 7588 40236
rect 7868 40290 8148 40292
rect 7868 40238 8094 40290
rect 8146 40238 8148 40290
rect 7868 40236 8148 40238
rect 7644 40180 7700 40190
rect 7644 40178 7812 40180
rect 7644 40126 7646 40178
rect 7698 40126 7812 40178
rect 7644 40124 7812 40126
rect 7644 40114 7700 40124
rect 7644 39844 7700 39854
rect 7532 39842 7700 39844
rect 7532 39790 7646 39842
rect 7698 39790 7700 39842
rect 7532 39788 7700 39790
rect 7196 39732 7252 39742
rect 6972 39730 7252 39732
rect 6972 39678 7198 39730
rect 7250 39678 7252 39730
rect 6972 39676 7252 39678
rect 7196 39666 7252 39676
rect 6860 39564 7028 39620
rect 6748 39554 6804 39564
rect 5740 38742 5796 38780
rect 5852 39060 5908 39070
rect 5852 38834 5908 39004
rect 6524 39058 6580 39228
rect 6524 39006 6526 39058
rect 6578 39006 6580 39058
rect 6524 38994 6580 39006
rect 6636 39396 6692 39406
rect 5852 38782 5854 38834
rect 5906 38782 5908 38834
rect 5852 38770 5908 38782
rect 6300 38948 6356 38958
rect 6300 38834 6356 38892
rect 6636 38836 6692 39340
rect 6860 39394 6916 39406
rect 6860 39342 6862 39394
rect 6914 39342 6916 39394
rect 6860 39284 6916 39342
rect 6860 39218 6916 39228
rect 6300 38782 6302 38834
rect 6354 38782 6356 38834
rect 6300 38770 6356 38782
rect 6524 38780 6692 38836
rect 6748 39060 6804 39070
rect 6076 38722 6132 38734
rect 6076 38670 6078 38722
rect 6130 38670 6132 38722
rect 6076 38668 6132 38670
rect 5964 38612 6020 38622
rect 6076 38612 6356 38668
rect 5964 38164 6020 38556
rect 6188 38164 6244 38174
rect 5964 38162 6244 38164
rect 5964 38110 6190 38162
rect 6242 38110 6244 38162
rect 5964 38108 6244 38110
rect 5628 37268 5684 37278
rect 5628 37266 5908 37268
rect 5628 37214 5630 37266
rect 5682 37214 5908 37266
rect 5628 37212 5908 37214
rect 5628 37202 5684 37212
rect 5852 36484 5908 37212
rect 5964 37266 6020 38108
rect 6188 38098 6244 38108
rect 6188 37940 6244 37950
rect 6076 37828 6132 37838
rect 6076 37490 6132 37772
rect 6076 37438 6078 37490
rect 6130 37438 6132 37490
rect 6076 37426 6132 37438
rect 6188 37490 6244 37884
rect 6188 37438 6190 37490
rect 6242 37438 6244 37490
rect 6188 37426 6244 37438
rect 5964 37214 5966 37266
rect 6018 37214 6020 37266
rect 5964 37044 6020 37214
rect 5964 36978 6020 36988
rect 6300 36596 6356 38612
rect 6524 38500 6580 38780
rect 6748 38724 6804 39004
rect 6076 36594 6356 36596
rect 6076 36542 6302 36594
rect 6354 36542 6356 36594
rect 6076 36540 6356 36542
rect 5964 36484 6020 36494
rect 5852 36482 6020 36484
rect 5852 36430 5966 36482
rect 6018 36430 6020 36482
rect 5852 36428 6020 36430
rect 5852 36260 5908 36428
rect 5964 36418 6020 36428
rect 5516 36204 5908 36260
rect 5516 35028 5572 36204
rect 5852 36036 5908 36046
rect 5628 35924 5684 35934
rect 5628 35252 5684 35868
rect 5852 35922 5908 35980
rect 6076 35924 6132 36540
rect 6300 36530 6356 36540
rect 6412 38444 6580 38500
rect 6636 38668 6804 38724
rect 6972 38668 7028 39564
rect 7084 38948 7140 38958
rect 7084 38834 7140 38892
rect 7084 38782 7086 38834
rect 7138 38782 7140 38834
rect 7084 38770 7140 38782
rect 7532 38834 7588 39788
rect 7644 39778 7700 39788
rect 7532 38782 7534 38834
rect 7586 38782 7588 38834
rect 7532 38770 7588 38782
rect 7756 38668 7812 40124
rect 7868 39842 7924 40236
rect 8092 40226 8148 40236
rect 8316 40178 8372 40190
rect 8316 40126 8318 40178
rect 8370 40126 8372 40178
rect 8316 39844 8372 40126
rect 7868 39790 7870 39842
rect 7922 39790 7924 39842
rect 7868 39778 7924 39790
rect 7980 39788 8316 39844
rect 7980 38946 8036 39788
rect 8316 39778 8372 39788
rect 7980 38894 7982 38946
rect 8034 38894 8036 38946
rect 7980 38882 8036 38894
rect 8316 39394 8372 39406
rect 8316 39342 8318 39394
rect 8370 39342 8372 39394
rect 6188 36372 6244 36382
rect 6188 36278 6244 36316
rect 6412 35924 6468 38444
rect 6636 38388 6692 38668
rect 6860 38610 6916 38622
rect 6860 38558 6862 38610
rect 6914 38558 6916 38610
rect 6860 38388 6916 38558
rect 6524 38332 6692 38388
rect 6748 38332 6916 38388
rect 6972 38612 7588 38668
rect 7756 38612 7924 38668
rect 6524 38050 6580 38332
rect 6748 38276 6804 38332
rect 6524 37998 6526 38050
rect 6578 37998 6580 38050
rect 6524 37986 6580 37998
rect 6636 38220 6804 38276
rect 6636 37266 6692 38220
rect 6636 37214 6638 37266
rect 6690 37214 6692 37266
rect 6636 37202 6692 37214
rect 6860 38164 6916 38174
rect 6860 37716 6916 38108
rect 6748 37042 6804 37054
rect 6748 36990 6750 37042
rect 6802 36990 6804 37042
rect 5852 35870 5854 35922
rect 5906 35870 5908 35922
rect 5852 35858 5908 35870
rect 5964 35868 6132 35924
rect 6300 35868 6468 35924
rect 6636 36482 6692 36494
rect 6636 36430 6638 36482
rect 6690 36430 6692 36482
rect 6636 35924 6692 36430
rect 5740 35700 5796 35710
rect 5964 35700 6020 35868
rect 5740 35606 5796 35644
rect 5852 35644 6020 35700
rect 6076 35698 6132 35710
rect 6076 35646 6078 35698
rect 6130 35646 6132 35698
rect 5628 35196 5796 35252
rect 5628 35028 5684 35038
rect 5516 35026 5684 35028
rect 5516 34974 5630 35026
rect 5682 34974 5684 35026
rect 5516 34972 5684 34974
rect 5628 34962 5684 34972
rect 5068 34130 5460 34132
rect 5068 34078 5070 34130
rect 5122 34078 5460 34130
rect 5068 34076 5460 34078
rect 5068 34066 5124 34076
rect 4284 33292 4788 33348
rect 4508 33124 4564 33134
rect 4508 33030 4564 33068
rect 4508 32788 4564 32798
rect 4508 32694 4564 32732
rect 4732 32786 4788 33292
rect 4844 33346 5012 33348
rect 4844 33294 4846 33346
rect 4898 33294 5012 33346
rect 4844 33292 5012 33294
rect 5180 33572 5236 33582
rect 4844 33012 4900 33292
rect 4844 32946 4900 32956
rect 4732 32734 4734 32786
rect 4786 32734 4788 32786
rect 4732 32722 4788 32734
rect 4844 32788 4900 32798
rect 4172 32564 4228 32574
rect 4396 32564 4452 32574
rect 4172 32562 4452 32564
rect 4172 32510 4174 32562
rect 4226 32510 4398 32562
rect 4450 32510 4452 32562
rect 4172 32508 4452 32510
rect 4172 32498 4228 32508
rect 4396 32498 4452 32508
rect 3724 31726 3726 31778
rect 3778 31726 3780 31778
rect 3724 31714 3780 31726
rect 3948 32396 4116 32452
rect 3948 31556 4004 32396
rect 4284 32340 4340 32350
rect 4172 31892 4228 31902
rect 4060 31780 4116 31818
rect 4060 31714 4116 31724
rect 4060 31556 4116 31566
rect 3948 31500 4060 31556
rect 4060 31490 4116 31500
rect 3500 31276 3892 31332
rect 3724 31106 3780 31118
rect 3724 31054 3726 31106
rect 3778 31054 3780 31106
rect 3724 30996 3780 31054
rect 3724 30930 3780 30940
rect 3500 29428 3556 29438
rect 3388 29426 3556 29428
rect 3388 29374 3502 29426
rect 3554 29374 3556 29426
rect 3388 29372 3556 29374
rect 3164 29334 3220 29372
rect 3500 29362 3556 29372
rect 3836 29426 3892 31276
rect 3948 30884 4004 30894
rect 3948 30790 4004 30828
rect 4172 30212 4228 31836
rect 4284 30436 4340 32284
rect 4476 32172 4740 32182
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4476 32106 4740 32116
rect 4508 32004 4564 32014
rect 4844 32004 4900 32732
rect 4508 31778 4564 31948
rect 4508 31726 4510 31778
rect 4562 31726 4564 31778
rect 4508 31714 4564 31726
rect 4620 31948 4900 32004
rect 5068 32450 5124 32462
rect 5068 32398 5070 32450
rect 5122 32398 5124 32450
rect 4620 31668 4676 31948
rect 5068 31892 5124 32398
rect 5180 32340 5236 33516
rect 5404 32564 5460 34076
rect 5404 32498 5460 32508
rect 5516 34020 5572 34030
rect 5740 34020 5796 35196
rect 5852 35138 5908 35644
rect 6076 35308 6132 35646
rect 5964 35252 6132 35308
rect 5964 35186 6020 35196
rect 5852 35086 5854 35138
rect 5906 35086 5908 35138
rect 5852 35074 5908 35086
rect 5516 34018 5796 34020
rect 5516 33966 5518 34018
rect 5570 33966 5796 34018
rect 5516 33964 5796 33966
rect 5964 35028 6020 35038
rect 5964 34018 6020 34972
rect 6300 35028 6356 35868
rect 6636 35858 6692 35868
rect 6412 35700 6468 35710
rect 6636 35700 6692 35710
rect 6412 35698 6692 35700
rect 6412 35646 6414 35698
rect 6466 35646 6638 35698
rect 6690 35646 6692 35698
rect 6412 35644 6692 35646
rect 6412 35634 6468 35644
rect 6636 35634 6692 35644
rect 6748 35588 6804 36990
rect 6860 35922 6916 37660
rect 6972 37042 7028 38612
rect 7084 37940 7140 37950
rect 7084 37938 7364 37940
rect 7084 37886 7086 37938
rect 7138 37886 7364 37938
rect 7084 37884 7364 37886
rect 7084 37874 7140 37884
rect 7308 37378 7364 37884
rect 7532 37938 7588 38612
rect 7756 38388 7812 38398
rect 7756 38274 7812 38332
rect 7756 38222 7758 38274
rect 7810 38222 7812 38274
rect 7756 38210 7812 38222
rect 7644 38164 7700 38174
rect 7644 38070 7700 38108
rect 7532 37886 7534 37938
rect 7586 37886 7588 37938
rect 7532 37874 7588 37886
rect 7308 37326 7310 37378
rect 7362 37326 7364 37378
rect 7308 37314 7364 37326
rect 7868 37268 7924 38612
rect 8316 38612 8372 39342
rect 8316 38546 8372 38556
rect 8316 38164 8372 38174
rect 8316 38070 8372 38108
rect 8092 38050 8148 38062
rect 8092 37998 8094 38050
rect 8146 37998 8148 38050
rect 8092 37604 8148 37998
rect 8092 37548 8372 37604
rect 8204 37380 8260 37418
rect 8204 37314 8260 37324
rect 8092 37268 8148 37278
rect 7868 37212 8092 37268
rect 8092 37174 8148 37212
rect 7084 37156 7140 37166
rect 8204 37156 8260 37166
rect 8316 37156 8372 37548
rect 7084 37154 7252 37156
rect 7084 37102 7086 37154
rect 7138 37102 7252 37154
rect 7084 37100 7252 37102
rect 7084 37090 7140 37100
rect 6972 36990 6974 37042
rect 7026 36990 7028 37042
rect 6972 36978 7028 36990
rect 6860 35870 6862 35922
rect 6914 35870 6916 35922
rect 6860 35812 6916 35870
rect 6860 35746 6916 35756
rect 7084 36148 7140 36158
rect 6972 35698 7028 35710
rect 6972 35646 6974 35698
rect 7026 35646 7028 35698
rect 6748 35532 6916 35588
rect 6300 34962 6356 34972
rect 6636 35028 6692 35038
rect 6188 34692 6244 34702
rect 6188 34690 6356 34692
rect 6188 34638 6190 34690
rect 6242 34638 6356 34690
rect 6188 34636 6356 34638
rect 6188 34626 6244 34636
rect 5964 33966 5966 34018
rect 6018 33966 6020 34018
rect 5180 32274 5236 32284
rect 5068 31826 5124 31836
rect 4844 31780 4900 31790
rect 4844 31778 5012 31780
rect 4844 31726 4846 31778
rect 4898 31726 5012 31778
rect 4844 31724 5012 31726
rect 4844 31714 4900 31724
rect 4732 31668 4788 31678
rect 4620 31666 4788 31668
rect 4620 31614 4734 31666
rect 4786 31614 4788 31666
rect 4620 31612 4788 31614
rect 4732 31602 4788 31612
rect 4956 31332 5012 31724
rect 4956 31276 5348 31332
rect 4844 31108 4900 31118
rect 4844 30994 4900 31052
rect 5292 31106 5348 31276
rect 5292 31054 5294 31106
rect 5346 31054 5348 31106
rect 5292 31042 5348 31054
rect 4844 30942 4846 30994
rect 4898 30942 4900 30994
rect 4844 30930 4900 30942
rect 4956 30996 5012 31006
rect 4956 30882 5012 30940
rect 4956 30830 4958 30882
rect 5010 30830 5012 30882
rect 4476 30604 4740 30614
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4476 30538 4740 30548
rect 4284 30380 4452 30436
rect 4172 30146 4228 30156
rect 4284 30210 4340 30222
rect 4284 30158 4286 30210
rect 4338 30158 4340 30210
rect 4284 30100 4340 30158
rect 4284 30034 4340 30044
rect 3836 29374 3838 29426
rect 3890 29374 3892 29426
rect 3836 29362 3892 29374
rect 4284 29652 4340 29662
rect 2604 28690 2660 28700
rect 2716 29316 2772 29326
rect 2716 28754 2772 29260
rect 3500 29204 3556 29214
rect 2716 28702 2718 28754
rect 2770 28702 2772 28754
rect 2716 28690 2772 28702
rect 3052 28980 3108 28990
rect 2268 28242 2324 28252
rect 3052 28642 3108 28924
rect 3500 28868 3556 29148
rect 3388 28812 3556 28868
rect 3052 28590 3054 28642
rect 3106 28590 3108 28642
rect 2268 28084 2324 28094
rect 1372 27972 1428 27982
rect 1260 27916 1372 27972
rect 1372 27906 1428 27916
rect 1820 27858 1876 27870
rect 1820 27806 1822 27858
rect 1874 27806 1876 27858
rect 1708 26962 1764 26974
rect 1708 26910 1710 26962
rect 1762 26910 1764 26962
rect 1708 26292 1764 26910
rect 1708 25844 1764 26236
rect 1708 25778 1764 25788
rect 1708 25620 1764 25630
rect 1708 24946 1764 25564
rect 1708 24894 1710 24946
rect 1762 24894 1764 24946
rect 1708 24882 1764 24894
rect 1820 25506 1876 27806
rect 2268 27186 2324 28028
rect 2492 27748 2548 27758
rect 2492 27654 2548 27692
rect 2268 27134 2270 27186
rect 2322 27134 2324 27186
rect 2268 27122 2324 27134
rect 2940 27074 2996 27086
rect 2940 27022 2942 27074
rect 2994 27022 2996 27074
rect 2380 26852 2436 26862
rect 2716 26852 2772 26862
rect 2156 26628 2212 26638
rect 2156 26514 2212 26572
rect 2156 26462 2158 26514
rect 2210 26462 2212 26514
rect 2156 26450 2212 26462
rect 1820 25454 1822 25506
rect 1874 25454 1876 25506
rect 1820 23938 1876 25454
rect 2380 26290 2436 26796
rect 2604 26796 2716 26852
rect 2380 26238 2382 26290
rect 2434 26238 2436 26290
rect 2380 25284 2436 26238
rect 2492 26740 2548 26750
rect 2492 25618 2548 26684
rect 2492 25566 2494 25618
rect 2546 25566 2548 25618
rect 2492 25554 2548 25566
rect 2492 25284 2548 25294
rect 2380 25228 2492 25284
rect 2492 25218 2548 25228
rect 2044 24834 2100 24846
rect 2044 24782 2046 24834
rect 2098 24782 2100 24834
rect 2044 24164 2100 24782
rect 2380 24724 2436 24734
rect 2044 24098 2100 24108
rect 2156 24612 2212 24622
rect 1820 23886 1822 23938
rect 1874 23886 1876 23938
rect 1708 23604 1764 23614
rect 1708 23378 1764 23548
rect 1708 23326 1710 23378
rect 1762 23326 1764 23378
rect 1708 21364 1764 23326
rect 1820 23044 1876 23886
rect 1820 22370 1876 22988
rect 2044 23266 2100 23278
rect 2044 23214 2046 23266
rect 2098 23214 2100 23266
rect 2044 22932 2100 23214
rect 2044 22866 2100 22876
rect 1820 22318 1822 22370
rect 1874 22318 1876 22370
rect 1820 21586 1876 22318
rect 1820 21534 1822 21586
rect 1874 21534 1876 21586
rect 1820 21522 1876 21534
rect 1708 21308 1988 21364
rect 1708 20914 1764 20926
rect 1708 20862 1710 20914
rect 1762 20862 1764 20914
rect 1708 20132 1764 20862
rect 1932 20188 1988 21308
rect 1932 20132 2100 20188
rect 1708 20066 1764 20076
rect 2044 19458 2100 20132
rect 2156 20130 2212 24556
rect 2156 20078 2158 20130
rect 2210 20078 2212 20130
rect 2156 20066 2212 20078
rect 2044 19406 2046 19458
rect 2098 19406 2100 19458
rect 2044 19394 2100 19406
rect 2156 19348 2212 19358
rect 2380 19348 2436 24668
rect 2492 24052 2548 24062
rect 2604 24052 2660 26796
rect 2716 26786 2772 26796
rect 2940 26516 2996 27022
rect 3052 26628 3108 28590
rect 3164 28644 3220 28654
rect 3164 27188 3220 28588
rect 3388 28530 3444 28812
rect 4284 28642 4340 29596
rect 4396 29316 4452 30380
rect 4956 30324 5012 30830
rect 5404 30884 5460 30894
rect 4956 30258 5012 30268
rect 5068 30436 5124 30446
rect 5068 30322 5124 30380
rect 5068 30270 5070 30322
rect 5122 30270 5124 30322
rect 5068 30258 5124 30270
rect 5404 29426 5460 30828
rect 5404 29374 5406 29426
rect 5458 29374 5460 29426
rect 5404 29362 5460 29374
rect 4396 29250 4452 29260
rect 4956 29316 5012 29326
rect 4476 29036 4740 29046
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4476 28970 4740 28980
rect 4844 28980 4900 28990
rect 4284 28590 4286 28642
rect 4338 28590 4340 28642
rect 4284 28578 4340 28590
rect 4396 28756 4452 28766
rect 3388 28478 3390 28530
rect 3442 28478 3444 28530
rect 3388 28466 3444 28478
rect 4396 28530 4452 28700
rect 4396 28478 4398 28530
rect 4450 28478 4452 28530
rect 4396 28466 4452 28478
rect 4620 28644 4676 28654
rect 4620 27746 4676 28588
rect 4844 28642 4900 28924
rect 4844 28590 4846 28642
rect 4898 28590 4900 28642
rect 4844 28578 4900 28590
rect 4956 28418 5012 29260
rect 4956 28366 4958 28418
rect 5010 28366 5012 28418
rect 4956 28354 5012 28366
rect 5180 28868 5236 28878
rect 5180 28082 5236 28812
rect 5180 28030 5182 28082
rect 5234 28030 5236 28082
rect 5180 28018 5236 28030
rect 4956 27860 5012 27870
rect 4620 27694 4622 27746
rect 4674 27694 4676 27746
rect 4620 27682 4676 27694
rect 4844 27858 5012 27860
rect 4844 27806 4958 27858
rect 5010 27806 5012 27858
rect 4844 27804 5012 27806
rect 3164 26962 3220 27132
rect 3164 26910 3166 26962
rect 3218 26910 3220 26962
rect 3164 26898 3220 26910
rect 3388 27636 3444 27646
rect 3052 26572 3220 26628
rect 2940 26450 2996 26460
rect 2940 26180 2996 26190
rect 2940 26086 2996 26124
rect 3052 25844 3108 25854
rect 2716 25620 2772 25630
rect 2772 25564 2884 25620
rect 2716 25554 2772 25564
rect 2492 24050 2660 24052
rect 2492 23998 2494 24050
rect 2546 23998 2660 24050
rect 2492 23996 2660 23998
rect 2492 23986 2548 23996
rect 2828 23380 2884 25564
rect 2940 25172 2996 25182
rect 2940 24722 2996 25116
rect 2940 24670 2942 24722
rect 2994 24670 2996 24722
rect 2940 24658 2996 24670
rect 2940 23380 2996 23390
rect 2828 23378 2996 23380
rect 2828 23326 2942 23378
rect 2994 23326 2996 23378
rect 2828 23324 2996 23326
rect 2940 23314 2996 23324
rect 2604 23042 2660 23054
rect 2604 22990 2606 23042
rect 2658 22990 2660 23042
rect 2604 22930 2660 22990
rect 2604 22878 2606 22930
rect 2658 22878 2660 22930
rect 2604 22866 2660 22878
rect 2492 22596 2548 22606
rect 2492 22482 2548 22540
rect 2492 22430 2494 22482
rect 2546 22430 2548 22482
rect 2492 22418 2548 22430
rect 2492 21474 2548 21486
rect 2492 21422 2494 21474
rect 2546 21422 2548 21474
rect 2492 19908 2548 21422
rect 3052 20188 3108 25788
rect 3164 22930 3220 26572
rect 3388 26290 3444 27580
rect 3724 27636 3780 27646
rect 3500 26962 3556 26974
rect 3500 26910 3502 26962
rect 3554 26910 3556 26962
rect 3500 26628 3556 26910
rect 3724 26962 3780 27580
rect 4476 27468 4740 27478
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4476 27402 4740 27412
rect 3724 26910 3726 26962
rect 3778 26910 3780 26962
rect 3612 26852 3668 26862
rect 3612 26758 3668 26796
rect 3500 26562 3556 26572
rect 3388 26238 3390 26290
rect 3442 26238 3444 26290
rect 3164 22878 3166 22930
rect 3218 22878 3220 22930
rect 3164 22866 3220 22878
rect 3276 25284 3332 25294
rect 2828 20132 3108 20188
rect 2828 20130 2884 20132
rect 2828 20078 2830 20130
rect 2882 20078 2884 20130
rect 2828 20066 2884 20078
rect 3276 20130 3332 25228
rect 3388 24612 3444 26238
rect 3724 24948 3780 26910
rect 4060 27300 4116 27310
rect 4060 26516 4116 27244
rect 4844 27188 4900 27804
rect 4956 27794 5012 27804
rect 5068 27748 5124 27758
rect 5068 27654 5124 27692
rect 5516 27524 5572 33964
rect 5964 33124 6020 33966
rect 5964 33058 6020 33068
rect 6188 34356 6244 34366
rect 6188 32786 6244 34300
rect 6300 33684 6356 34636
rect 6636 34690 6692 34972
rect 6636 34638 6638 34690
rect 6690 34638 6692 34690
rect 6412 34356 6468 34366
rect 6468 34300 6580 34356
rect 6412 34262 6468 34300
rect 6412 33684 6468 33694
rect 6300 33628 6412 33684
rect 6412 33618 6468 33628
rect 6188 32734 6190 32786
rect 6242 32734 6244 32786
rect 6188 32722 6244 32734
rect 6300 33236 6356 33246
rect 6300 32786 6356 33180
rect 6524 33234 6580 34300
rect 6636 34020 6692 34638
rect 6748 34356 6804 34366
rect 6748 34262 6804 34300
rect 6860 34244 6916 35532
rect 6860 34178 6916 34188
rect 6636 33348 6692 33964
rect 6972 33684 7028 35646
rect 6972 33618 7028 33628
rect 6636 33254 6692 33292
rect 6524 33182 6526 33234
rect 6578 33182 6580 33234
rect 6524 33170 6580 33182
rect 6300 32734 6302 32786
rect 6354 32734 6356 32786
rect 6300 32722 6356 32734
rect 5740 32562 5796 32574
rect 5740 32510 5742 32562
rect 5794 32510 5796 32562
rect 5628 32452 5684 32462
rect 5628 31780 5684 32396
rect 5740 32004 5796 32510
rect 5740 31938 5796 31948
rect 6300 32564 6356 32574
rect 5852 31780 5908 31790
rect 5628 31724 5852 31780
rect 6300 31780 6356 32508
rect 6412 32562 6468 32574
rect 6412 32510 6414 32562
rect 6466 32510 6468 32562
rect 6412 32452 6468 32510
rect 6636 32452 6692 32462
rect 6412 32396 6636 32452
rect 6636 32386 6692 32396
rect 6972 32450 7028 32462
rect 6972 32398 6974 32450
rect 7026 32398 7028 32450
rect 6748 32116 6804 32126
rect 6636 31892 6692 31902
rect 6636 31798 6692 31836
rect 6412 31780 6468 31790
rect 6300 31778 6468 31780
rect 6300 31726 6414 31778
rect 6466 31726 6468 31778
rect 6300 31724 6468 31726
rect 5852 31686 5908 31724
rect 6412 31714 6468 31724
rect 6412 31556 6468 31566
rect 6636 31556 6692 31566
rect 6468 31554 6692 31556
rect 6468 31502 6638 31554
rect 6690 31502 6692 31554
rect 6468 31500 6692 31502
rect 6412 31490 6468 31500
rect 6636 31490 6692 31500
rect 6636 31332 6692 31342
rect 6076 31220 6132 31230
rect 6524 31220 6580 31230
rect 6076 31218 6580 31220
rect 6076 31166 6078 31218
rect 6130 31166 6526 31218
rect 6578 31166 6580 31218
rect 6076 31164 6580 31166
rect 6076 31154 6132 31164
rect 5852 30996 5908 31006
rect 5852 30994 6020 30996
rect 5852 30942 5854 30994
rect 5906 30942 6020 30994
rect 5852 30940 6020 30942
rect 5852 30930 5908 30940
rect 5964 30098 6020 30940
rect 6412 30994 6468 31006
rect 6412 30942 6414 30994
rect 6466 30942 6468 30994
rect 5964 30046 5966 30098
rect 6018 30046 6020 30098
rect 5740 28868 5796 28878
rect 5740 28774 5796 28812
rect 5628 28644 5684 28654
rect 5964 28644 6020 30046
rect 6188 30884 6244 30894
rect 5684 28588 6020 28644
rect 6076 29314 6132 29326
rect 6076 29262 6078 29314
rect 6130 29262 6132 29314
rect 5628 28550 5684 28588
rect 5852 28420 5908 28430
rect 5740 28084 5796 28094
rect 5628 28028 5740 28084
rect 5628 27858 5684 28028
rect 5740 28018 5796 28028
rect 5628 27806 5630 27858
rect 5682 27806 5684 27858
rect 5628 27794 5684 27806
rect 5068 27468 5572 27524
rect 4508 27132 4900 27188
rect 4172 27074 4228 27086
rect 4172 27022 4174 27074
rect 4226 27022 4228 27074
rect 4172 26908 4228 27022
rect 4508 27074 4564 27132
rect 4508 27022 4510 27074
rect 4562 27022 4564 27074
rect 4508 27010 4564 27022
rect 4732 26964 4788 26974
rect 4172 26852 4564 26908
rect 4732 26870 4788 26908
rect 4172 26516 4228 26526
rect 4060 26514 4228 26516
rect 4060 26462 4174 26514
rect 4226 26462 4228 26514
rect 4060 26460 4228 26462
rect 4172 26450 4228 26460
rect 4396 26516 4452 26526
rect 4508 26516 4564 26852
rect 4620 26850 4676 26862
rect 4620 26798 4622 26850
rect 4674 26798 4676 26850
rect 4620 26740 4676 26798
rect 4620 26674 4676 26684
rect 4844 26628 4900 27132
rect 4732 26516 4788 26526
rect 4508 26514 4788 26516
rect 4508 26462 4734 26514
rect 4786 26462 4788 26514
rect 4508 26460 4788 26462
rect 4396 26292 4452 26460
rect 4732 26450 4788 26460
rect 4284 26290 4452 26292
rect 4284 26238 4398 26290
rect 4450 26238 4452 26290
rect 4284 26236 4452 26238
rect 3836 26178 3892 26190
rect 3836 26126 3838 26178
rect 3890 26126 3892 26178
rect 3836 25844 3892 26126
rect 3836 25778 3892 25788
rect 3836 24948 3892 24958
rect 3724 24946 3892 24948
rect 3724 24894 3838 24946
rect 3890 24894 3892 24946
rect 3724 24892 3892 24894
rect 3836 24882 3892 24892
rect 3388 24546 3444 24556
rect 4172 24610 4228 24622
rect 4172 24558 4174 24610
rect 4226 24558 4228 24610
rect 4172 24498 4228 24558
rect 4172 24446 4174 24498
rect 4226 24446 4228 24498
rect 4172 24434 4228 24446
rect 4284 23548 4340 26236
rect 4396 26226 4452 26236
rect 4476 25900 4740 25910
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4476 25834 4740 25844
rect 4620 25620 4676 25630
rect 4620 25526 4676 25564
rect 4620 24610 4676 24622
rect 4620 24558 4622 24610
rect 4674 24558 4676 24610
rect 4620 24500 4676 24558
rect 4844 24612 4900 26572
rect 4956 27188 5012 27198
rect 4956 26514 5012 27132
rect 5068 26628 5124 27468
rect 5740 27188 5796 27198
rect 5180 27186 5796 27188
rect 5180 27134 5742 27186
rect 5794 27134 5796 27186
rect 5180 27132 5796 27134
rect 5180 27074 5236 27132
rect 5740 27122 5796 27132
rect 5180 27022 5182 27074
rect 5234 27022 5236 27074
rect 5180 27010 5236 27022
rect 5852 26962 5908 28364
rect 5852 26910 5854 26962
rect 5906 26910 5908 26962
rect 5628 26852 5684 26862
rect 5068 26562 5124 26572
rect 5180 26740 5236 26750
rect 4956 26462 4958 26514
rect 5010 26462 5012 26514
rect 4956 26450 5012 26462
rect 5068 26404 5124 26414
rect 5068 26310 5124 26348
rect 5180 25618 5236 26684
rect 5516 26516 5572 26526
rect 5516 26422 5572 26460
rect 5628 26292 5684 26796
rect 5740 26740 5796 26750
rect 5852 26740 5908 26910
rect 5964 27300 6020 27310
rect 5964 26962 6020 27244
rect 5964 26910 5966 26962
rect 6018 26910 6020 26962
rect 5964 26898 6020 26910
rect 5796 26684 5908 26740
rect 5964 26740 6020 26750
rect 5740 26674 5796 26684
rect 5852 26292 5908 26302
rect 5628 26290 5908 26292
rect 5628 26238 5854 26290
rect 5906 26238 5908 26290
rect 5628 26236 5908 26238
rect 5852 26226 5908 26236
rect 5180 25566 5182 25618
rect 5234 25566 5236 25618
rect 5180 25554 5236 25566
rect 5404 26180 5460 26190
rect 5180 25172 5236 25182
rect 5068 24612 5124 24622
rect 4844 24610 5124 24612
rect 4844 24558 5070 24610
rect 5122 24558 5124 24610
rect 4844 24556 5124 24558
rect 4620 24444 4900 24500
rect 4476 24332 4740 24342
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4476 24266 4740 24276
rect 4620 24052 4676 24062
rect 4620 23958 4676 23996
rect 4284 23492 4564 23548
rect 4508 23378 4564 23492
rect 4508 23326 4510 23378
rect 4562 23326 4564 23378
rect 3500 23042 3556 23054
rect 3500 22990 3502 23042
rect 3554 22990 3556 23042
rect 3500 22930 3556 22990
rect 3948 23044 4004 23054
rect 3948 22950 4004 22988
rect 3500 22878 3502 22930
rect 3554 22878 3556 22930
rect 3500 22866 3556 22878
rect 4508 22930 4564 23326
rect 4508 22878 4510 22930
rect 4562 22878 4564 22930
rect 4508 22866 4564 22878
rect 4844 23154 4900 24444
rect 5068 24498 5124 24556
rect 5068 24446 5070 24498
rect 5122 24446 5124 24498
rect 5068 24388 5124 24446
rect 5068 24322 5124 24332
rect 5180 24050 5236 25116
rect 5180 23998 5182 24050
rect 5234 23998 5236 24050
rect 5180 23986 5236 23998
rect 4844 23102 4846 23154
rect 4898 23102 4900 23154
rect 4844 23044 4900 23102
rect 4476 22764 4740 22774
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4476 22698 4740 22708
rect 4620 22484 4676 22494
rect 4620 22390 4676 22428
rect 4844 22148 4900 22988
rect 5068 22148 5124 22158
rect 4844 22146 5124 22148
rect 4844 22094 5070 22146
rect 5122 22094 5124 22146
rect 4844 22092 5124 22094
rect 5068 21588 5124 22092
rect 5404 21812 5460 26124
rect 5964 26068 6020 26684
rect 6076 26292 6132 29262
rect 6188 28530 6244 30828
rect 6412 30772 6468 30942
rect 6524 30996 6580 31164
rect 6524 30930 6580 30940
rect 6300 30436 6356 30446
rect 6300 29988 6356 30380
rect 6412 30210 6468 30716
rect 6412 30158 6414 30210
rect 6466 30158 6468 30210
rect 6412 30146 6468 30158
rect 6300 29932 6468 29988
rect 6188 28478 6190 28530
rect 6242 28478 6244 28530
rect 6188 26908 6244 28478
rect 6412 29764 6468 29932
rect 6412 28530 6468 29708
rect 6636 28644 6692 31276
rect 6748 31218 6804 32060
rect 6972 31780 7028 32398
rect 7084 31892 7140 36092
rect 7196 35028 7252 37100
rect 8260 37100 8372 37156
rect 7420 37044 7476 37054
rect 7420 36950 7476 36988
rect 8204 37042 8260 37100
rect 8204 36990 8206 37042
rect 8258 36990 8260 37042
rect 8204 36978 8260 36990
rect 7420 36596 7476 36606
rect 7420 36502 7476 36540
rect 7308 36484 7364 36494
rect 7308 36258 7364 36428
rect 7532 36484 7588 36494
rect 7532 36390 7588 36428
rect 7756 36484 7812 36494
rect 7812 36428 7924 36484
rect 7756 36418 7812 36428
rect 7308 36206 7310 36258
rect 7362 36206 7364 36258
rect 7308 36194 7364 36206
rect 7756 36258 7812 36270
rect 7756 36206 7758 36258
rect 7810 36206 7812 36258
rect 7644 36148 7700 36158
rect 7644 35700 7700 36092
rect 7196 34962 7252 34972
rect 7308 35698 7700 35700
rect 7308 35646 7646 35698
rect 7698 35646 7700 35698
rect 7308 35644 7700 35646
rect 7196 34802 7252 34814
rect 7196 34750 7198 34802
rect 7250 34750 7252 34802
rect 7196 33906 7252 34750
rect 7308 34580 7364 35644
rect 7644 35634 7700 35644
rect 7420 35252 7476 35262
rect 7420 34802 7476 35196
rect 7644 35028 7700 35038
rect 7756 35028 7812 36206
rect 7868 35700 7924 36428
rect 8428 35924 8484 42476
rect 8652 42438 8708 42476
rect 8876 42084 8932 42094
rect 8876 41990 8932 42028
rect 8764 41412 8820 41422
rect 8820 41356 8932 41412
rect 8764 41346 8820 41356
rect 8764 41188 8820 41198
rect 8764 41094 8820 41132
rect 8764 40402 8820 40414
rect 8764 40350 8766 40402
rect 8818 40350 8820 40402
rect 8540 40180 8596 40190
rect 8540 40086 8596 40124
rect 8540 39508 8596 39518
rect 8764 39508 8820 40350
rect 8540 39506 8820 39508
rect 8540 39454 8542 39506
rect 8594 39454 8820 39506
rect 8540 39452 8820 39454
rect 8540 39396 8596 39452
rect 8540 39330 8596 39340
rect 8652 39172 8708 39182
rect 8540 39060 8596 39070
rect 8540 38966 8596 39004
rect 8540 38500 8596 38510
rect 8540 38050 8596 38444
rect 8652 38162 8708 39116
rect 8876 39060 8932 41356
rect 8988 40964 9044 43374
rect 9100 42754 9156 44942
rect 9548 44884 9604 45614
rect 11116 45666 11172 45678
rect 11116 45614 11118 45666
rect 11170 45614 11172 45666
rect 11116 45444 11172 45614
rect 11116 45378 11172 45388
rect 11564 45668 11620 45678
rect 11676 45668 11732 45678
rect 11620 45666 11732 45668
rect 11620 45614 11678 45666
rect 11730 45614 11732 45666
rect 11620 45612 11732 45614
rect 10108 45108 10164 45118
rect 9660 44996 9716 45006
rect 9660 44902 9716 44940
rect 10108 44994 10164 45052
rect 10108 44942 10110 44994
rect 10162 44942 10164 44994
rect 9548 44818 9604 44828
rect 10108 44884 10164 44942
rect 10444 44996 10500 45006
rect 10444 44994 10612 44996
rect 10444 44942 10446 44994
rect 10498 44942 10612 44994
rect 10444 44940 10612 44942
rect 10444 44930 10500 44940
rect 10108 44818 10164 44828
rect 9548 44210 9604 44222
rect 9548 44158 9550 44210
rect 9602 44158 9604 44210
rect 9548 43652 9604 44158
rect 9548 43586 9604 43596
rect 9996 43538 10052 43550
rect 9996 43486 9998 43538
rect 10050 43486 10052 43538
rect 9548 43428 9604 43438
rect 9100 42702 9102 42754
rect 9154 42702 9156 42754
rect 9100 41860 9156 42702
rect 9324 43426 9604 43428
rect 9324 43374 9550 43426
rect 9602 43374 9604 43426
rect 9324 43372 9604 43374
rect 9212 42644 9268 42654
rect 9212 42550 9268 42588
rect 9100 41794 9156 41804
rect 9324 41188 9380 43372
rect 9548 43362 9604 43372
rect 9436 42530 9492 42542
rect 9436 42478 9438 42530
rect 9490 42478 9492 42530
rect 9436 41972 9492 42478
rect 9996 42196 10052 43486
rect 10444 43426 10500 43438
rect 10444 43374 10446 43426
rect 10498 43374 10500 43426
rect 9996 42130 10052 42140
rect 10108 42868 10164 42878
rect 10108 42084 10164 42812
rect 10220 42642 10276 42654
rect 10220 42590 10222 42642
rect 10274 42590 10276 42642
rect 10220 42532 10276 42590
rect 10220 42466 10276 42476
rect 10444 42196 10500 43374
rect 10556 42756 10612 44940
rect 11004 43764 11060 43774
rect 10892 43538 10948 43550
rect 10892 43486 10894 43538
rect 10946 43486 10948 43538
rect 10892 42868 10948 43486
rect 10892 42802 10948 42812
rect 10556 42690 10612 42700
rect 11004 42754 11060 43708
rect 11452 43652 11508 43662
rect 11452 43558 11508 43596
rect 11340 43538 11396 43550
rect 11340 43486 11342 43538
rect 11394 43486 11396 43538
rect 11340 42980 11396 43486
rect 11564 43540 11620 45612
rect 11676 45602 11732 45612
rect 12124 45666 12180 45678
rect 12124 45614 12126 45666
rect 12178 45614 12180 45666
rect 11788 44996 11844 45006
rect 12124 44996 12180 45614
rect 12572 45666 12628 45678
rect 12572 45614 12574 45666
rect 12626 45614 12628 45666
rect 11844 44940 12180 44996
rect 12236 45444 12292 45454
rect 12572 45444 12628 45614
rect 12292 45388 12628 45444
rect 13468 45666 13524 45678
rect 13468 45614 13470 45666
rect 13522 45614 13524 45666
rect 11788 44930 11844 44940
rect 11676 44434 11732 44446
rect 11676 44382 11678 44434
rect 11730 44382 11732 44434
rect 11676 44100 11732 44382
rect 12012 44100 12068 44110
rect 11676 44098 12068 44100
rect 11676 44046 12014 44098
rect 12066 44046 12068 44098
rect 11676 44044 12068 44046
rect 11676 43764 11732 44044
rect 12012 44034 12068 44044
rect 11676 43698 11732 43708
rect 11900 43764 11956 43774
rect 11620 43484 11732 43540
rect 11564 43446 11620 43484
rect 11676 43092 11732 43484
rect 11900 43538 11956 43708
rect 11900 43486 11902 43538
rect 11954 43486 11956 43538
rect 11900 43474 11956 43486
rect 11676 43026 11732 43036
rect 11340 42924 11620 42980
rect 11004 42702 11006 42754
rect 11058 42702 11060 42754
rect 11004 42690 11060 42702
rect 11340 42756 11396 42766
rect 11340 42662 11396 42700
rect 11452 42644 11508 42654
rect 11452 42550 11508 42588
rect 10108 42018 10164 42028
rect 10220 42140 10500 42196
rect 9436 41906 9492 41916
rect 9884 41972 9940 41982
rect 9772 41860 9828 41870
rect 9660 41858 9828 41860
rect 9660 41806 9774 41858
rect 9826 41806 9828 41858
rect 9660 41804 9828 41806
rect 9324 41186 9604 41188
rect 9324 41134 9326 41186
rect 9378 41134 9604 41186
rect 9324 41132 9604 41134
rect 9324 41122 9380 41132
rect 8988 40908 9268 40964
rect 8876 38994 8932 39004
rect 8988 38722 9044 38734
rect 8988 38670 8990 38722
rect 9042 38670 9044 38722
rect 8988 38668 9044 38670
rect 8988 38612 9156 38668
rect 8652 38110 8654 38162
rect 8706 38110 8708 38162
rect 8652 38098 8708 38110
rect 8988 38052 9044 38062
rect 8540 37998 8542 38050
rect 8594 37998 8596 38050
rect 8540 37986 8596 37998
rect 8876 37996 8988 38052
rect 8764 37828 8820 37838
rect 8652 37826 8820 37828
rect 8652 37774 8766 37826
rect 8818 37774 8820 37826
rect 8652 37772 8820 37774
rect 8540 36258 8596 36270
rect 8540 36206 8542 36258
rect 8594 36206 8596 36258
rect 8540 36148 8596 36206
rect 8540 36082 8596 36092
rect 8652 35924 8708 37772
rect 8764 37762 8820 37772
rect 8316 35868 8484 35924
rect 8540 35868 8708 35924
rect 8764 37268 8820 37278
rect 8876 37268 8932 37996
rect 8988 37986 9044 37996
rect 8764 37266 8932 37268
rect 8764 37214 8766 37266
rect 8818 37214 8932 37266
rect 8764 37212 8932 37214
rect 8988 37378 9044 37390
rect 8988 37326 8990 37378
rect 9042 37326 9044 37378
rect 8092 35812 8148 35822
rect 8092 35718 8148 35756
rect 7868 35606 7924 35644
rect 8204 35700 8260 35710
rect 7980 35586 8036 35598
rect 7980 35534 7982 35586
rect 8034 35534 8036 35586
rect 7980 35028 8036 35534
rect 8092 35140 8148 35150
rect 8204 35140 8260 35644
rect 8092 35138 8260 35140
rect 8092 35086 8094 35138
rect 8146 35086 8260 35138
rect 8092 35084 8260 35086
rect 8092 35074 8148 35084
rect 7644 35026 7812 35028
rect 7644 34974 7646 35026
rect 7698 34974 7812 35026
rect 7644 34972 7812 34974
rect 7868 34972 8036 35028
rect 7644 34962 7700 34972
rect 7420 34750 7422 34802
rect 7474 34750 7476 34802
rect 7420 34738 7476 34750
rect 7532 34804 7588 34814
rect 7868 34804 7924 34972
rect 8204 34916 8260 34926
rect 8316 34916 8372 35868
rect 8428 35700 8484 35710
rect 8428 35606 8484 35644
rect 8540 35252 8596 35868
rect 8652 35700 8708 35710
rect 8764 35700 8820 37212
rect 8652 35698 8820 35700
rect 8652 35646 8654 35698
rect 8706 35646 8820 35698
rect 8652 35644 8820 35646
rect 8876 36258 8932 36270
rect 8876 36206 8878 36258
rect 8930 36206 8932 36258
rect 8652 35634 8708 35644
rect 8540 35196 8820 35252
rect 8428 35140 8484 35150
rect 8484 35084 8708 35140
rect 8428 35074 8484 35084
rect 8652 35026 8708 35084
rect 8652 34974 8654 35026
rect 8706 34974 8708 35026
rect 8652 34962 8708 34974
rect 8204 34914 8484 34916
rect 8204 34862 8206 34914
rect 8258 34862 8484 34914
rect 8204 34860 8484 34862
rect 8204 34850 8260 34860
rect 7532 34710 7588 34748
rect 7756 34748 7924 34804
rect 7756 34692 7812 34748
rect 7644 34690 7812 34692
rect 7644 34638 7758 34690
rect 7810 34638 7812 34690
rect 7644 34636 7812 34638
rect 7308 34524 7588 34580
rect 7308 34020 7364 34030
rect 7308 33926 7364 33964
rect 7196 33854 7198 33906
rect 7250 33854 7252 33906
rect 7196 33842 7252 33854
rect 7420 33684 7476 33694
rect 7308 32452 7364 32462
rect 7308 32358 7364 32396
rect 7084 31836 7252 31892
rect 7028 31724 7140 31780
rect 6972 31686 7028 31724
rect 6748 31166 6750 31218
rect 6802 31166 6804 31218
rect 6748 31154 6804 31166
rect 6860 31554 6916 31566
rect 6860 31502 6862 31554
rect 6914 31502 6916 31554
rect 6748 29428 6804 29438
rect 6748 29334 6804 29372
rect 6860 28868 6916 31502
rect 7084 31106 7140 31724
rect 7084 31054 7086 31106
rect 7138 31054 7140 31106
rect 7084 30884 7140 31054
rect 7084 30818 7140 30828
rect 6972 30772 7028 30782
rect 6972 30678 7028 30716
rect 6972 29316 7028 29326
rect 6972 29222 7028 29260
rect 6860 28802 6916 28812
rect 7196 28866 7252 31836
rect 7196 28814 7198 28866
rect 7250 28814 7252 28866
rect 7196 28802 7252 28814
rect 7308 30770 7364 30782
rect 7308 30718 7310 30770
rect 7362 30718 7364 30770
rect 6412 28478 6414 28530
rect 6466 28478 6468 28530
rect 6300 28418 6356 28430
rect 6300 28366 6302 28418
rect 6354 28366 6356 28418
rect 6300 28084 6356 28366
rect 6412 28420 6468 28478
rect 6412 28354 6468 28364
rect 6524 28642 6692 28644
rect 6524 28590 6638 28642
rect 6690 28590 6692 28642
rect 6524 28588 6692 28590
rect 6300 28018 6356 28028
rect 6300 27748 6356 27758
rect 6524 27748 6580 28588
rect 6636 28578 6692 28588
rect 6972 28644 7028 28654
rect 7196 28644 7252 28654
rect 6972 28642 7196 28644
rect 6972 28590 6974 28642
rect 7026 28590 7196 28642
rect 6972 28588 7196 28590
rect 6972 28578 7028 28588
rect 7196 28578 7252 28588
rect 6300 27746 6580 27748
rect 6300 27694 6302 27746
rect 6354 27694 6580 27746
rect 6300 27692 6580 27694
rect 6636 27858 6692 27870
rect 6636 27806 6638 27858
rect 6690 27806 6692 27858
rect 6300 27682 6356 27692
rect 6412 27412 6468 27422
rect 6300 27356 6412 27412
rect 6300 27074 6356 27356
rect 6412 27346 6468 27356
rect 6300 27022 6302 27074
rect 6354 27022 6356 27074
rect 6300 27010 6356 27022
rect 6524 27300 6580 27310
rect 6524 26964 6580 27244
rect 6188 26852 6468 26908
rect 6524 26898 6580 26908
rect 6076 26236 6244 26292
rect 6076 26068 6132 26078
rect 5964 26066 6132 26068
rect 5964 26014 6078 26066
rect 6130 26014 6132 26066
rect 5964 26012 6132 26014
rect 6076 26002 6132 26012
rect 5628 24724 5684 24734
rect 5628 24630 5684 24668
rect 6076 24610 6132 24622
rect 6076 24558 6078 24610
rect 6130 24558 6132 24610
rect 6076 23940 6132 24558
rect 6188 24612 6244 26236
rect 6300 26068 6356 26078
rect 6300 25974 6356 26012
rect 6412 24724 6468 26852
rect 6636 26740 6692 27806
rect 7084 27858 7140 27870
rect 7084 27806 7086 27858
rect 7138 27806 7140 27858
rect 6860 27412 6916 27422
rect 6860 27186 6916 27356
rect 6860 27134 6862 27186
rect 6914 27134 6916 27186
rect 6860 27122 6916 27134
rect 6972 26964 7028 27002
rect 6972 26898 7028 26908
rect 6748 26852 6804 26862
rect 6748 26850 6916 26852
rect 6748 26798 6750 26850
rect 6802 26798 6916 26850
rect 6748 26796 6916 26798
rect 6748 26786 6804 26796
rect 6636 26516 6692 26684
rect 6636 26450 6692 26460
rect 6748 26628 6804 26638
rect 6748 26292 6804 26572
rect 6748 26226 6804 26236
rect 6748 26066 6804 26078
rect 6748 26014 6750 26066
rect 6802 26014 6804 26066
rect 6748 25508 6804 26014
rect 6860 26068 6916 26796
rect 7084 26740 7140 27806
rect 7196 27860 7252 27870
rect 7196 27766 7252 27804
rect 7196 27076 7252 27086
rect 7196 26962 7252 27020
rect 7196 26910 7198 26962
rect 7250 26910 7252 26962
rect 7196 26898 7252 26910
rect 6860 26002 6916 26012
rect 6972 26684 7140 26740
rect 6972 26290 7028 26684
rect 7308 26628 7364 30718
rect 7420 26908 7476 33628
rect 7532 33346 7588 34524
rect 7532 33294 7534 33346
rect 7586 33294 7588 33346
rect 7532 32004 7588 33294
rect 7644 32786 7700 34636
rect 7756 34626 7812 34636
rect 8204 34468 8260 34478
rect 8204 34242 8260 34412
rect 8204 34190 8206 34242
rect 8258 34190 8260 34242
rect 7980 34130 8036 34142
rect 7980 34078 7982 34130
rect 8034 34078 8036 34130
rect 7756 34018 7812 34030
rect 7756 33966 7758 34018
rect 7810 33966 7812 34018
rect 7756 33796 7812 33966
rect 7868 33908 7924 33918
rect 7980 33908 8036 34078
rect 7868 33906 8036 33908
rect 7868 33854 7870 33906
rect 7922 33854 8036 33906
rect 7868 33852 8036 33854
rect 7868 33842 7924 33852
rect 7756 33730 7812 33740
rect 7644 32734 7646 32786
rect 7698 32734 7700 32786
rect 7644 32722 7700 32734
rect 8092 33122 8148 33134
rect 8092 33070 8094 33122
rect 8146 33070 8148 33122
rect 8092 32786 8148 33070
rect 8092 32734 8094 32786
rect 8146 32734 8148 32786
rect 8092 32722 8148 32734
rect 7868 32564 7924 32574
rect 7868 32470 7924 32508
rect 7532 31938 7588 31948
rect 7756 32450 7812 32462
rect 7756 32398 7758 32450
rect 7810 32398 7812 32450
rect 7532 31668 7588 31678
rect 7532 31574 7588 31612
rect 7756 30996 7812 32398
rect 8204 32004 8260 34190
rect 8316 34130 8372 34142
rect 8316 34078 8318 34130
rect 8370 34078 8372 34130
rect 8316 32564 8372 34078
rect 8428 33236 8484 34860
rect 8540 34804 8596 34814
rect 8540 33684 8596 34748
rect 8764 34804 8820 35196
rect 8876 35028 8932 36206
rect 8988 35812 9044 37326
rect 9100 36260 9156 38612
rect 9212 37492 9268 40908
rect 9324 40962 9380 40974
rect 9324 40910 9326 40962
rect 9378 40910 9380 40962
rect 9324 38388 9380 40910
rect 9548 40292 9604 41132
rect 9548 40226 9604 40236
rect 9324 38322 9380 38332
rect 9436 40178 9492 40190
rect 9436 40126 9438 40178
rect 9490 40126 9492 40178
rect 9436 38052 9492 40126
rect 9660 38500 9716 41804
rect 9772 41794 9828 41804
rect 9772 41074 9828 41086
rect 9772 41022 9774 41074
rect 9826 41022 9828 41074
rect 9772 40740 9828 41022
rect 9772 40674 9828 40684
rect 9660 38434 9716 38444
rect 9772 40516 9828 40526
rect 9436 37986 9492 37996
rect 9660 38050 9716 38062
rect 9660 37998 9662 38050
rect 9714 37998 9716 38050
rect 9660 37492 9716 37998
rect 9212 37436 9604 37492
rect 9100 36194 9156 36204
rect 9324 37268 9380 37278
rect 8988 35746 9044 35756
rect 8988 35476 9044 35486
rect 8988 35474 9156 35476
rect 8988 35422 8990 35474
rect 9042 35422 9156 35474
rect 8988 35420 9156 35422
rect 8988 35410 9044 35420
rect 8876 34962 8932 34972
rect 8988 34804 9044 34814
rect 8764 34802 9044 34804
rect 8764 34750 8990 34802
rect 9042 34750 9044 34802
rect 8764 34748 9044 34750
rect 8764 34356 8820 34748
rect 8988 34738 9044 34748
rect 8764 34242 8820 34300
rect 8764 34190 8766 34242
rect 8818 34190 8820 34242
rect 8764 34178 8820 34190
rect 8876 34244 8932 34254
rect 8876 34150 8932 34188
rect 8540 33618 8596 33628
rect 8652 33908 8708 33918
rect 8652 33460 8708 33852
rect 8428 33170 8484 33180
rect 8540 33404 8708 33460
rect 8876 33906 8932 33918
rect 8876 33854 8878 33906
rect 8930 33854 8932 33906
rect 8540 33346 8596 33404
rect 8876 33348 8932 33854
rect 9100 33572 9156 35420
rect 9324 35140 9380 37212
rect 9436 36258 9492 36270
rect 9436 36206 9438 36258
rect 9490 36206 9492 36258
rect 9436 36148 9492 36206
rect 9436 36082 9492 36092
rect 9548 35252 9604 37436
rect 9660 37044 9716 37436
rect 9660 36978 9716 36988
rect 9772 36596 9828 40460
rect 9884 40290 9940 41916
rect 10108 41860 10164 41870
rect 10108 40516 10164 41804
rect 10220 40740 10276 42140
rect 11116 42084 11172 42094
rect 11564 42084 11620 42924
rect 11900 42084 11956 42094
rect 10444 41970 10500 41982
rect 10444 41918 10446 41970
rect 10498 41918 10500 41970
rect 10220 40674 10276 40684
rect 10332 41746 10388 41758
rect 10332 41694 10334 41746
rect 10386 41694 10388 41746
rect 10108 40460 10276 40516
rect 9884 40238 9886 40290
rect 9938 40238 9940 40290
rect 9884 40226 9940 40238
rect 10108 40292 10164 40302
rect 10108 40198 10164 40236
rect 9996 39620 10052 39630
rect 9884 39394 9940 39406
rect 9884 39342 9886 39394
rect 9938 39342 9940 39394
rect 9884 38948 9940 39342
rect 9884 38162 9940 38892
rect 9884 38110 9886 38162
rect 9938 38110 9940 38162
rect 9884 38098 9940 38110
rect 9996 39058 10052 39564
rect 9996 39006 9998 39058
rect 10050 39006 10052 39058
rect 9996 37380 10052 39006
rect 10220 38668 10276 40460
rect 10332 40404 10388 41694
rect 10444 40516 10500 41918
rect 10668 41972 10724 41982
rect 10668 41878 10724 41916
rect 11004 41186 11060 41198
rect 11004 41134 11006 41186
rect 11058 41134 11060 41186
rect 11004 41076 11060 41134
rect 11004 41010 11060 41020
rect 10556 40516 10612 40526
rect 10444 40514 10836 40516
rect 10444 40462 10558 40514
rect 10610 40462 10836 40514
rect 10444 40460 10836 40462
rect 10556 40450 10612 40460
rect 10332 40348 10500 40404
rect 10332 40178 10388 40190
rect 10332 40126 10334 40178
rect 10386 40126 10388 40178
rect 10332 39618 10388 40126
rect 10332 39566 10334 39618
rect 10386 39566 10388 39618
rect 10332 39508 10388 39566
rect 10332 39442 10388 39452
rect 10444 39060 10500 40348
rect 10780 40292 10836 40460
rect 11004 40404 11060 40414
rect 11116 40404 11172 42028
rect 11452 42028 11620 42084
rect 11676 42082 11956 42084
rect 11676 42030 11902 42082
rect 11954 42030 11956 42082
rect 11676 42028 11956 42030
rect 11004 40402 11172 40404
rect 11004 40350 11006 40402
rect 11058 40350 11172 40402
rect 11004 40348 11172 40350
rect 11228 40740 11284 40750
rect 10892 40292 10948 40302
rect 10780 40290 10948 40292
rect 10780 40238 10894 40290
rect 10946 40238 10948 40290
rect 10780 40236 10948 40238
rect 10444 39004 10612 39060
rect 10444 38834 10500 38846
rect 10444 38782 10446 38834
rect 10498 38782 10500 38834
rect 10444 38668 10500 38782
rect 10220 38612 10500 38668
rect 10220 37604 10276 38612
rect 9996 37314 10052 37324
rect 10108 37378 10164 37390
rect 10108 37326 10110 37378
rect 10162 37326 10164 37378
rect 9884 37268 9940 37278
rect 9884 37174 9940 37212
rect 10108 37156 10164 37326
rect 10108 37044 10164 37100
rect 9660 36540 9828 36596
rect 9884 36988 10164 37044
rect 9660 35924 9716 36540
rect 9772 36370 9828 36382
rect 9772 36318 9774 36370
rect 9826 36318 9828 36370
rect 9772 36260 9828 36318
rect 9772 36194 9828 36204
rect 9884 36370 9940 36988
rect 10220 36932 10276 37548
rect 10332 37938 10388 37950
rect 10332 37886 10334 37938
rect 10386 37886 10388 37938
rect 10332 37380 10388 37886
rect 10332 37314 10388 37324
rect 10556 37268 10612 39004
rect 10108 36876 10276 36932
rect 10444 37266 10612 37268
rect 10444 37214 10558 37266
rect 10610 37214 10612 37266
rect 10444 37212 10612 37214
rect 9996 36820 10052 36830
rect 9996 36482 10052 36764
rect 9996 36430 9998 36482
rect 10050 36430 10052 36482
rect 9996 36418 10052 36430
rect 9884 36318 9886 36370
rect 9938 36318 9940 36370
rect 9772 35924 9828 35934
rect 9660 35922 9828 35924
rect 9660 35870 9774 35922
rect 9826 35870 9828 35922
rect 9660 35868 9828 35870
rect 9772 35858 9828 35868
rect 9884 35812 9940 36318
rect 9884 35746 9940 35756
rect 9660 35700 9716 35710
rect 9716 35644 9828 35700
rect 9660 35606 9716 35644
rect 9772 35308 9828 35644
rect 9548 35186 9604 35196
rect 9660 35252 9828 35308
rect 9996 35698 10052 35710
rect 9996 35646 9998 35698
rect 10050 35646 10052 35698
rect 9436 35140 9492 35150
rect 9324 35084 9436 35140
rect 9436 35074 9492 35084
rect 9436 34916 9492 34926
rect 9436 34822 9492 34860
rect 9660 34914 9716 35252
rect 9660 34862 9662 34914
rect 9714 34862 9716 34914
rect 9660 34850 9716 34862
rect 9884 34804 9940 34814
rect 9996 34804 10052 35646
rect 10108 35588 10164 36876
rect 10444 36820 10500 37212
rect 10556 37202 10612 37212
rect 10668 37826 10724 37838
rect 10668 37774 10670 37826
rect 10722 37774 10724 37826
rect 10668 37268 10724 37774
rect 10668 37202 10724 37212
rect 10780 37044 10836 40236
rect 10892 40226 10948 40236
rect 10892 39732 10948 39742
rect 10892 39058 10948 39676
rect 10892 39006 10894 39058
rect 10946 39006 10948 39058
rect 10892 37828 10948 39006
rect 10892 37762 10948 37772
rect 11004 37716 11060 40348
rect 11228 39506 11284 40684
rect 11452 40516 11508 42028
rect 11452 40450 11508 40460
rect 11564 41858 11620 41870
rect 11564 41806 11566 41858
rect 11618 41806 11620 41858
rect 11340 40404 11396 40414
rect 11340 40310 11396 40348
rect 11564 39844 11620 41806
rect 11676 40180 11732 42028
rect 11900 42018 11956 42028
rect 11900 41188 11956 41198
rect 11900 40514 11956 41132
rect 11900 40462 11902 40514
rect 11954 40462 11956 40514
rect 11900 40450 11956 40462
rect 12124 41076 12180 41086
rect 12236 41076 12292 45388
rect 13244 45108 13300 45118
rect 13468 45108 13524 45614
rect 13692 45668 13748 45678
rect 14588 45668 14644 45678
rect 15036 45668 15092 45678
rect 15820 45668 15876 45678
rect 13692 45666 13860 45668
rect 13692 45614 13694 45666
rect 13746 45614 13860 45666
rect 13692 45612 13860 45614
rect 13692 45602 13748 45612
rect 13692 45108 13748 45118
rect 13244 45106 13692 45108
rect 13244 45054 13246 45106
rect 13298 45054 13692 45106
rect 13244 45052 13692 45054
rect 12572 44996 12628 45006
rect 12572 44994 12740 44996
rect 12572 44942 12574 44994
rect 12626 44942 12740 44994
rect 12572 44940 12740 44942
rect 12572 44930 12628 44940
rect 12348 44098 12404 44110
rect 12348 44046 12350 44098
rect 12402 44046 12404 44098
rect 12348 43652 12404 44046
rect 12572 44098 12628 44110
rect 12572 44046 12574 44098
rect 12626 44046 12628 44098
rect 12572 43764 12628 44046
rect 12572 43698 12628 43708
rect 12348 42084 12404 43596
rect 12460 43538 12516 43550
rect 12460 43486 12462 43538
rect 12514 43486 12516 43538
rect 12460 43204 12516 43486
rect 12684 43540 12740 44940
rect 12908 44212 12964 44222
rect 12796 44098 12852 44110
rect 12796 44046 12798 44098
rect 12850 44046 12852 44098
rect 12796 43652 12852 44046
rect 12908 43764 12964 44156
rect 12908 43698 12964 43708
rect 12796 43586 12852 43596
rect 12684 43474 12740 43484
rect 13132 43428 13188 43438
rect 13132 43334 13188 43372
rect 13244 43204 13300 45052
rect 13692 45014 13748 45052
rect 13692 44098 13748 44110
rect 13692 44046 13694 44098
rect 13746 44046 13748 44098
rect 13692 43876 13748 44046
rect 13692 43810 13748 43820
rect 13804 43652 13860 45612
rect 14252 45666 14644 45668
rect 14252 45614 14590 45666
rect 14642 45614 14644 45666
rect 14252 45612 14644 45614
rect 14140 44100 14196 44110
rect 12460 43148 13300 43204
rect 13468 43596 13860 43652
rect 14028 44098 14196 44100
rect 14028 44046 14142 44098
rect 14194 44046 14196 44098
rect 14028 44044 14196 44046
rect 12460 42756 12516 42766
rect 12460 42194 12516 42700
rect 12460 42142 12462 42194
rect 12514 42142 12516 42194
rect 12460 42130 12516 42142
rect 12348 42018 12404 42028
rect 12908 41860 12964 41870
rect 12572 41748 12628 41758
rect 12460 41692 12572 41748
rect 12124 41074 12292 41076
rect 12124 41022 12126 41074
rect 12178 41022 12292 41074
rect 12124 41020 12292 41022
rect 12348 41074 12404 41086
rect 12348 41022 12350 41074
rect 12402 41022 12404 41074
rect 11788 40180 11844 40190
rect 11676 40124 11788 40180
rect 11788 40114 11844 40124
rect 11564 39778 11620 39788
rect 11228 39454 11230 39506
rect 11282 39454 11284 39506
rect 11228 39442 11284 39454
rect 11788 39060 11844 39070
rect 11788 38946 11844 39004
rect 12124 39060 12180 41020
rect 12348 40740 12404 41022
rect 12460 40962 12516 41692
rect 12572 41682 12628 41692
rect 12684 41636 12740 41646
rect 12684 41410 12740 41580
rect 12908 41524 12964 41804
rect 12908 41458 12964 41468
rect 12684 41358 12686 41410
rect 12738 41358 12740 41410
rect 12684 41346 12740 41358
rect 12460 40910 12462 40962
rect 12514 40910 12516 40962
rect 12460 40898 12516 40910
rect 12908 41186 12964 41198
rect 12908 41134 12910 41186
rect 12962 41134 12964 41186
rect 12572 40852 12628 40862
rect 12572 40740 12628 40796
rect 12348 40684 12628 40740
rect 12348 39844 12404 39854
rect 12348 39618 12404 39788
rect 12348 39566 12350 39618
rect 12402 39566 12404 39618
rect 12124 38994 12180 39004
rect 12236 39396 12292 39406
rect 11788 38894 11790 38946
rect 11842 38894 11844 38946
rect 11788 38882 11844 38894
rect 12236 38946 12292 39340
rect 12236 38894 12238 38946
rect 12290 38894 12292 38946
rect 12236 38882 12292 38894
rect 11340 38836 11396 38846
rect 11340 38722 11396 38780
rect 11340 38670 11342 38722
rect 11394 38670 11396 38722
rect 11340 38388 11396 38670
rect 11340 38322 11396 38332
rect 11676 38610 11732 38622
rect 11676 38558 11678 38610
rect 11730 38558 11732 38610
rect 11116 38052 11172 38062
rect 11116 37958 11172 37996
rect 11452 38052 11508 38062
rect 11676 38052 11732 38558
rect 12348 38610 12404 39566
rect 12348 38558 12350 38610
rect 12402 38558 12404 38610
rect 12348 38546 12404 38558
rect 12012 38052 12068 38062
rect 12348 38052 12404 38062
rect 11452 38050 12180 38052
rect 11452 37998 11454 38050
rect 11506 37998 12014 38050
rect 12066 37998 12180 38050
rect 11452 37996 12180 37998
rect 11452 37986 11508 37996
rect 12012 37986 12068 37996
rect 11228 37940 11284 37950
rect 11228 37846 11284 37884
rect 11004 37660 11284 37716
rect 11116 37490 11172 37502
rect 11116 37438 11118 37490
rect 11170 37438 11172 37490
rect 11004 37268 11060 37278
rect 10444 36754 10500 36764
rect 10556 36988 10836 37044
rect 10892 37266 11060 37268
rect 10892 37214 11006 37266
rect 11058 37214 11060 37266
rect 10892 37212 11060 37214
rect 10444 36260 10500 36270
rect 10220 36258 10500 36260
rect 10220 36206 10446 36258
rect 10498 36206 10500 36258
rect 10220 36204 10500 36206
rect 10220 35810 10276 36204
rect 10444 36194 10500 36204
rect 10220 35758 10222 35810
rect 10274 35758 10276 35810
rect 10220 35746 10276 35758
rect 10108 35532 10388 35588
rect 9940 34748 10052 34804
rect 10108 35028 10164 35038
rect 10108 34914 10164 34972
rect 10108 34862 10110 34914
rect 10162 34862 10164 34914
rect 10108 34804 10164 34862
rect 9884 34738 9940 34748
rect 10108 34738 10164 34748
rect 10220 34802 10276 34814
rect 10220 34750 10222 34802
rect 10274 34750 10276 34802
rect 9212 34690 9268 34702
rect 9212 34638 9214 34690
rect 9266 34638 9268 34690
rect 9212 34244 9268 34638
rect 9212 34178 9268 34188
rect 9324 34690 9380 34702
rect 9324 34638 9326 34690
rect 9378 34638 9380 34690
rect 9324 34020 9380 34638
rect 9436 34356 9492 34366
rect 10220 34356 10276 34750
rect 9492 34300 9604 34356
rect 9436 34290 9492 34300
rect 9548 34242 9604 34300
rect 9548 34190 9550 34242
rect 9602 34190 9604 34242
rect 9548 34178 9604 34190
rect 10108 34300 10276 34356
rect 9996 34130 10052 34142
rect 9996 34078 9998 34130
rect 10050 34078 10052 34130
rect 9324 33954 9380 33964
rect 9660 34018 9716 34030
rect 9660 33966 9662 34018
rect 9714 33966 9716 34018
rect 9660 33908 9716 33966
rect 9660 33842 9716 33852
rect 9100 33506 9156 33516
rect 9212 33684 9268 33694
rect 8540 33294 8542 33346
rect 8594 33294 8596 33346
rect 8540 32788 8596 33294
rect 8652 33292 8932 33348
rect 8652 32900 8708 33292
rect 8764 33124 8820 33134
rect 8764 33030 8820 33068
rect 8876 33012 8932 33022
rect 8652 32844 8820 32900
rect 8540 32732 8708 32788
rect 8316 32498 8372 32508
rect 8092 31948 8260 32004
rect 7980 30996 8036 31006
rect 7756 30994 8036 30996
rect 7756 30942 7982 30994
rect 8034 30942 8036 30994
rect 7756 30940 8036 30942
rect 7980 30930 8036 30940
rect 7756 30772 7812 30782
rect 7756 30678 7812 30716
rect 7868 30212 7924 30222
rect 7868 30118 7924 30156
rect 7644 30098 7700 30110
rect 7644 30046 7646 30098
rect 7698 30046 7700 30098
rect 7644 29652 7700 30046
rect 8092 29988 8148 31948
rect 8204 31780 8260 31790
rect 8260 31724 8484 31780
rect 8204 31686 8260 31724
rect 8428 31332 8484 31724
rect 8540 31668 8596 31678
rect 8540 31574 8596 31612
rect 8652 31444 8708 32732
rect 8764 31780 8820 32844
rect 8876 32002 8932 32956
rect 8988 32452 9044 32462
rect 8988 32358 9044 32396
rect 8876 31950 8878 32002
rect 8930 31950 8932 32002
rect 8876 31938 8932 31950
rect 9100 32004 9156 32014
rect 9100 31890 9156 31948
rect 9100 31838 9102 31890
rect 9154 31838 9156 31890
rect 9100 31826 9156 31838
rect 8764 31714 8820 31724
rect 8764 31444 8820 31454
rect 8652 31388 8764 31444
rect 8764 31378 8820 31388
rect 8428 31276 8708 31332
rect 8204 30884 8260 30894
rect 8204 30790 8260 30828
rect 8428 30882 8484 30894
rect 8428 30830 8430 30882
rect 8482 30830 8484 30882
rect 7644 29586 7700 29596
rect 7868 29932 8148 29988
rect 8204 30324 8260 30334
rect 8204 29986 8260 30268
rect 8428 30212 8484 30830
rect 8428 30146 8484 30156
rect 8652 30210 8708 31276
rect 8764 31220 8820 31230
rect 8820 31164 8932 31220
rect 8764 31154 8820 31164
rect 8876 31106 8932 31164
rect 8876 31054 8878 31106
rect 8930 31054 8932 31106
rect 8876 31042 8932 31054
rect 8988 30996 9044 31006
rect 8988 30212 9044 30940
rect 8652 30158 8654 30210
rect 8706 30158 8708 30210
rect 8652 30146 8708 30158
rect 8876 30210 9044 30212
rect 8876 30158 8990 30210
rect 9042 30158 9044 30210
rect 8876 30156 9044 30158
rect 8204 29934 8206 29986
rect 8258 29934 8260 29986
rect 7532 28754 7588 28766
rect 7532 28702 7534 28754
rect 7586 28702 7588 28754
rect 7532 28644 7588 28702
rect 7532 28642 7812 28644
rect 7532 28590 7534 28642
rect 7586 28590 7812 28642
rect 7532 28588 7812 28590
rect 7532 28578 7588 28588
rect 7756 28082 7812 28588
rect 7756 28030 7758 28082
rect 7810 28030 7812 28082
rect 7756 26908 7812 28030
rect 7868 27972 7924 29932
rect 8204 29876 8260 29934
rect 7980 29820 8260 29876
rect 8764 30098 8820 30110
rect 8764 30046 8766 30098
rect 8818 30046 8820 30098
rect 7980 28642 8036 29820
rect 8316 29540 8372 29550
rect 8316 29446 8372 29484
rect 8652 29428 8708 29438
rect 8764 29428 8820 30046
rect 8876 29538 8932 30156
rect 8988 30146 9044 30156
rect 8876 29486 8878 29538
rect 8930 29486 8932 29538
rect 8876 29474 8932 29486
rect 8652 29426 8820 29428
rect 8652 29374 8654 29426
rect 8706 29374 8820 29426
rect 8652 29372 8820 29374
rect 8428 29316 8484 29326
rect 8204 29314 8484 29316
rect 8204 29262 8430 29314
rect 8482 29262 8484 29314
rect 8204 29260 8484 29262
rect 7980 28590 7982 28642
rect 8034 28590 8036 28642
rect 7980 28578 8036 28590
rect 8092 28644 8148 28654
rect 8092 28550 8148 28588
rect 8204 28530 8260 29260
rect 8428 29250 8484 29260
rect 8652 28868 8708 29372
rect 9212 29316 9268 33628
rect 9996 33684 10052 34078
rect 9996 33618 10052 33628
rect 9884 33458 9940 33470
rect 9884 33406 9886 33458
rect 9938 33406 9940 33458
rect 9884 33348 9940 33406
rect 10108 33460 10164 34300
rect 10332 34244 10388 35532
rect 10556 34916 10612 36988
rect 10780 36484 10836 36494
rect 10892 36484 10948 37212
rect 11004 37202 11060 37212
rect 11116 37156 11172 37438
rect 11116 37090 11172 37100
rect 10780 36482 10948 36484
rect 10780 36430 10782 36482
rect 10834 36430 10948 36482
rect 10780 36428 10948 36430
rect 11004 37044 11060 37054
rect 11004 36482 11060 36988
rect 11004 36430 11006 36482
rect 11058 36430 11060 36482
rect 10780 35476 10836 36428
rect 11004 36418 11060 36430
rect 11116 36820 11172 36830
rect 11116 36482 11172 36764
rect 11116 36430 11118 36482
rect 11170 36430 11172 36482
rect 11116 36418 11172 36430
rect 10892 35812 10948 35822
rect 10892 35718 10948 35756
rect 10556 34850 10612 34860
rect 10668 35474 10836 35476
rect 10668 35422 10782 35474
rect 10834 35422 10836 35474
rect 10668 35420 10836 35422
rect 10444 34804 10500 34814
rect 10444 34354 10500 34748
rect 10444 34302 10446 34354
rect 10498 34302 10500 34354
rect 10444 34290 10500 34302
rect 10556 34356 10612 34366
rect 10332 34178 10388 34188
rect 10220 34132 10276 34142
rect 10220 34038 10276 34076
rect 10444 34020 10500 34030
rect 9884 33282 9940 33292
rect 9996 33346 10052 33358
rect 9996 33294 9998 33346
rect 10050 33294 10052 33346
rect 9548 33236 9604 33246
rect 9548 33142 9604 33180
rect 9324 32900 9380 32910
rect 9324 31890 9380 32844
rect 9548 32676 9604 32686
rect 9324 31838 9326 31890
rect 9378 31838 9380 31890
rect 9324 31826 9380 31838
rect 9436 32620 9548 32676
rect 8876 29260 9268 29316
rect 9324 31444 9380 31454
rect 8764 28868 8820 28878
rect 8652 28812 8764 28868
rect 8764 28802 8820 28812
rect 8540 28644 8596 28654
rect 8204 28478 8206 28530
rect 8258 28478 8260 28530
rect 8204 28466 8260 28478
rect 8428 28532 8484 28542
rect 8428 28082 8484 28476
rect 8428 28030 8430 28082
rect 8482 28030 8484 28082
rect 8428 28018 8484 28030
rect 8092 27972 8148 27982
rect 8204 27972 8260 27982
rect 7868 27970 8204 27972
rect 7868 27918 8094 27970
rect 8146 27918 8204 27970
rect 7868 27916 8204 27918
rect 8092 27906 8148 27916
rect 7420 26852 7588 26908
rect 6972 26238 6974 26290
rect 7026 26238 7028 26290
rect 6972 25620 7028 26238
rect 6972 25554 7028 25564
rect 7084 26572 7364 26628
rect 6748 25442 6804 25452
rect 6972 25172 7028 25182
rect 6412 24668 6692 24724
rect 6300 24612 6356 24622
rect 6188 24610 6356 24612
rect 6188 24558 6302 24610
rect 6354 24558 6356 24610
rect 6188 24556 6356 24558
rect 6076 23884 6244 23940
rect 6076 23716 6132 23726
rect 6076 23622 6132 23660
rect 6188 23604 6244 23884
rect 6300 23828 6356 24556
rect 6300 23762 6356 23772
rect 6412 24500 6468 24510
rect 6412 23716 6468 24444
rect 6524 24498 6580 24510
rect 6524 24446 6526 24498
rect 6578 24446 6580 24498
rect 6524 23940 6580 24446
rect 6524 23874 6580 23884
rect 6524 23716 6580 23726
rect 6412 23714 6580 23716
rect 6412 23662 6526 23714
rect 6578 23662 6580 23714
rect 6412 23660 6580 23662
rect 6524 23650 6580 23660
rect 6300 23604 6356 23614
rect 6188 23548 6300 23604
rect 6300 23538 6356 23548
rect 6636 23380 6692 24668
rect 6972 24722 7028 25116
rect 6972 24670 6974 24722
rect 7026 24670 7028 24722
rect 6972 24658 7028 24670
rect 6748 24612 6804 24622
rect 6748 24518 6804 24556
rect 7084 24388 7140 26572
rect 7532 26516 7588 26852
rect 7308 26460 7588 26516
rect 7644 26852 7812 26908
rect 7868 27748 7924 27758
rect 7868 27074 7924 27692
rect 7868 27022 7870 27074
rect 7922 27022 7924 27074
rect 7868 26908 7924 27022
rect 8092 27076 8148 27086
rect 8092 26962 8148 27020
rect 8092 26910 8094 26962
rect 8146 26910 8148 26962
rect 7868 26852 8036 26908
rect 8092 26898 8148 26910
rect 6748 24332 7140 24388
rect 7196 26292 7252 26302
rect 7196 25506 7252 26236
rect 7308 25618 7364 26460
rect 7644 26180 7700 26852
rect 7868 26402 7924 26414
rect 7868 26350 7870 26402
rect 7922 26350 7924 26402
rect 7644 26114 7700 26124
rect 7756 26178 7812 26190
rect 7756 26126 7758 26178
rect 7810 26126 7812 26178
rect 7308 25566 7310 25618
rect 7362 25566 7364 25618
rect 7308 25554 7364 25566
rect 7756 26068 7812 26126
rect 7196 25454 7198 25506
rect 7250 25454 7252 25506
rect 6748 23940 6804 24332
rect 6748 23846 6804 23884
rect 7196 23940 7252 25454
rect 7756 24722 7812 26012
rect 7868 25956 7924 26350
rect 7868 25890 7924 25900
rect 7868 25506 7924 25518
rect 7868 25454 7870 25506
rect 7922 25454 7924 25506
rect 7868 24834 7924 25454
rect 7980 24948 8036 26852
rect 8092 26292 8148 26302
rect 8092 26198 8148 26236
rect 8204 25844 8260 27916
rect 8204 25778 8260 25788
rect 8316 27074 8372 27086
rect 8316 27022 8318 27074
rect 8370 27022 8372 27074
rect 8316 26852 8372 27022
rect 8540 27076 8596 28588
rect 8764 28530 8820 28542
rect 8764 28478 8766 28530
rect 8818 28478 8820 28530
rect 8764 27188 8820 28478
rect 8764 27122 8820 27132
rect 8652 27076 8708 27086
rect 8540 27020 8652 27076
rect 8652 26982 8708 27020
rect 8876 26908 8932 29260
rect 9324 29204 9380 31388
rect 9436 31108 9492 32620
rect 9548 32610 9604 32620
rect 9996 32564 10052 33294
rect 10108 33236 10164 33404
rect 10332 33908 10388 33918
rect 10332 33346 10388 33852
rect 10332 33294 10334 33346
rect 10386 33294 10388 33346
rect 10332 33282 10388 33294
rect 10108 33180 10276 33236
rect 9996 32470 10052 32508
rect 9660 32452 9716 32462
rect 9660 32358 9716 32396
rect 9772 32228 9828 32238
rect 9660 32004 9716 32014
rect 9548 31780 9604 31790
rect 9660 31780 9716 31948
rect 9548 31778 9716 31780
rect 9548 31726 9550 31778
rect 9602 31726 9716 31778
rect 9548 31724 9716 31726
rect 9772 31778 9828 32172
rect 9772 31726 9774 31778
rect 9826 31726 9828 31778
rect 9548 31714 9604 31724
rect 9660 31554 9716 31566
rect 9660 31502 9662 31554
rect 9714 31502 9716 31554
rect 9548 31220 9604 31258
rect 9548 31154 9604 31164
rect 9436 30322 9492 31052
rect 9548 30996 9604 31006
rect 9548 30902 9604 30940
rect 9660 30772 9716 31502
rect 9772 31444 9828 31726
rect 10220 31778 10276 33180
rect 10220 31726 10222 31778
rect 10274 31726 10276 31778
rect 10220 31714 10276 31726
rect 10332 32900 10388 32910
rect 10332 32674 10388 32844
rect 10332 32622 10334 32674
rect 10386 32622 10388 32674
rect 9772 31378 9828 31388
rect 10108 31668 10164 31678
rect 9660 30706 9716 30716
rect 9772 31108 9828 31118
rect 9436 30270 9438 30322
rect 9490 30270 9492 30322
rect 9436 30258 9492 30270
rect 9660 30324 9716 30334
rect 9772 30324 9828 31052
rect 9660 30322 9828 30324
rect 9660 30270 9662 30322
rect 9714 30270 9828 30322
rect 9660 30268 9828 30270
rect 9996 30994 10052 31006
rect 9996 30942 9998 30994
rect 10050 30942 10052 30994
rect 9660 30258 9716 30268
rect 9660 29652 9716 29662
rect 9660 29558 9716 29596
rect 9996 29428 10052 30942
rect 10108 30996 10164 31612
rect 10108 30902 10164 30940
rect 10332 30212 10388 32622
rect 9212 29148 9380 29204
rect 9660 29372 10052 29428
rect 10220 30156 10388 30212
rect 8988 27746 9044 27758
rect 8988 27694 8990 27746
rect 9042 27694 9044 27746
rect 8988 27636 9044 27694
rect 8988 27570 9044 27580
rect 8092 25508 8148 25518
rect 8092 25414 8148 25452
rect 7980 24892 8148 24948
rect 7868 24782 7870 24834
rect 7922 24782 7924 24834
rect 7868 24770 7924 24782
rect 7756 24670 7758 24722
rect 7810 24670 7812 24722
rect 7756 24658 7812 24670
rect 7420 24500 7476 24510
rect 7420 24498 7588 24500
rect 7420 24446 7422 24498
rect 7474 24446 7588 24498
rect 7420 24444 7588 24446
rect 7420 24434 7476 24444
rect 6860 23828 6916 23838
rect 6860 23734 6916 23772
rect 6636 23314 6692 23324
rect 6524 23268 6580 23278
rect 5516 23044 5572 23054
rect 5516 23042 6468 23044
rect 5516 22990 5518 23042
rect 5570 22990 6468 23042
rect 5516 22988 6468 22990
rect 5516 22978 5572 22988
rect 5852 22820 5908 22830
rect 5852 22482 5908 22764
rect 5852 22430 5854 22482
rect 5906 22430 5908 22482
rect 5852 22418 5908 22430
rect 6412 22482 6468 22988
rect 6412 22430 6414 22482
rect 6466 22430 6468 22482
rect 6412 22418 6468 22430
rect 6524 22370 6580 23212
rect 7196 22820 7252 23884
rect 7196 22754 7252 22764
rect 7420 23156 7476 23166
rect 7420 22594 7476 23100
rect 7420 22542 7422 22594
rect 7474 22542 7476 22594
rect 7420 22530 7476 22542
rect 7308 22484 7364 22494
rect 7308 22390 7364 22428
rect 6524 22318 6526 22370
rect 6578 22318 6580 22370
rect 6524 22306 6580 22318
rect 6748 22370 6804 22382
rect 6748 22318 6750 22370
rect 6802 22318 6804 22370
rect 6076 22258 6132 22270
rect 6076 22206 6078 22258
rect 6130 22206 6132 22258
rect 6076 22148 6132 22206
rect 6748 22260 6804 22318
rect 6804 22204 6916 22260
rect 6748 22194 6804 22204
rect 5628 21812 5684 21822
rect 5404 21756 5628 21812
rect 5628 21718 5684 21756
rect 4620 21474 4676 21486
rect 4620 21422 4622 21474
rect 4674 21422 4676 21474
rect 4620 21364 4676 21422
rect 4620 21298 4676 21308
rect 4476 21196 4740 21206
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4476 21130 4740 21140
rect 5068 20914 5124 21532
rect 5740 21586 5796 21598
rect 5740 21534 5742 21586
rect 5794 21534 5796 21586
rect 5180 21476 5236 21486
rect 5180 21382 5236 21420
rect 5068 20862 5070 20914
rect 5122 20862 5124 20914
rect 5068 20850 5124 20862
rect 4508 20804 4564 20814
rect 4284 20802 4564 20804
rect 4284 20750 4510 20802
rect 4562 20750 4564 20802
rect 4284 20748 4564 20750
rect 3836 20690 3892 20702
rect 3836 20638 3838 20690
rect 3890 20638 3892 20690
rect 3276 20078 3278 20130
rect 3330 20078 3332 20130
rect 3276 20066 3332 20078
rect 3612 20132 3668 20142
rect 3612 20038 3668 20076
rect 3500 20020 3556 20030
rect 2492 19842 2548 19852
rect 3388 19964 3500 20020
rect 2940 19458 2996 19470
rect 2940 19406 2942 19458
rect 2994 19406 2996 19458
rect 2492 19348 2548 19358
rect 2380 19346 2548 19348
rect 2380 19294 2494 19346
rect 2546 19294 2548 19346
rect 2380 19292 2548 19294
rect 2156 19254 2212 19292
rect 2492 19282 2548 19292
rect 2940 19346 2996 19406
rect 2940 19294 2942 19346
rect 2994 19294 2996 19346
rect 2940 19282 2996 19294
rect 1820 18452 1876 18462
rect 1708 16772 1764 16782
rect 1708 16210 1764 16716
rect 1708 16158 1710 16210
rect 1762 16158 1764 16210
rect 1708 16146 1764 16158
rect 1820 14530 1876 18396
rect 2492 18340 2548 18350
rect 2492 18246 2548 18284
rect 1932 17780 1988 17790
rect 1932 17686 1988 17724
rect 3276 17108 3332 17118
rect 3276 17014 3332 17052
rect 2828 16884 2884 16894
rect 2828 16790 2884 16828
rect 3164 16772 3220 16782
rect 3164 16678 3220 16716
rect 3388 16772 3444 19964
rect 3500 19954 3556 19964
rect 3724 19796 3780 19806
rect 3612 19794 3780 19796
rect 3612 19742 3726 19794
rect 3778 19742 3780 19794
rect 3612 19740 3780 19742
rect 3500 19348 3556 19358
rect 3500 19254 3556 19292
rect 3612 19236 3668 19740
rect 3724 19730 3780 19740
rect 3612 19170 3668 19180
rect 3724 19234 3780 19246
rect 3724 19182 3726 19234
rect 3778 19182 3780 19234
rect 3724 18676 3780 19182
rect 3836 19012 3892 20638
rect 4172 20132 4228 20142
rect 4172 20038 4228 20076
rect 4060 19908 4116 19918
rect 4060 19814 4116 19852
rect 3948 19236 4004 19246
rect 4284 19236 4340 20748
rect 4508 20738 4564 20748
rect 5740 20244 5796 21534
rect 5740 20178 5796 20188
rect 5852 21588 5908 21598
rect 4732 20130 4788 20142
rect 4732 20078 4734 20130
rect 4786 20078 4788 20130
rect 4396 20020 4452 20030
rect 4396 19926 4452 19964
rect 4732 19796 4788 20078
rect 5628 20132 5684 20142
rect 5404 20020 5460 20030
rect 5292 20018 5460 20020
rect 5292 19966 5406 20018
rect 5458 19966 5460 20018
rect 5292 19964 5460 19966
rect 4956 19908 5012 19918
rect 4956 19814 5012 19852
rect 4732 19730 4788 19740
rect 5068 19794 5124 19806
rect 5068 19742 5070 19794
rect 5122 19742 5124 19794
rect 4476 19628 4740 19638
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4476 19562 4740 19572
rect 4844 19460 4900 19470
rect 3948 19142 4004 19180
rect 4060 19180 4340 19236
rect 4396 19404 4844 19460
rect 4396 19234 4452 19404
rect 4844 19366 4900 19404
rect 4956 19236 5012 19246
rect 4396 19182 4398 19234
rect 4450 19182 4452 19234
rect 3836 18946 3892 18956
rect 3724 18620 4004 18676
rect 3948 17892 4004 18620
rect 4060 18452 4116 19180
rect 4396 19170 4452 19182
rect 4732 19234 5012 19236
rect 4732 19182 4958 19234
rect 5010 19182 5012 19234
rect 4732 19180 5012 19182
rect 4060 18386 4116 18396
rect 4172 19010 4228 19022
rect 4172 18958 4174 19010
rect 4226 18958 4228 19010
rect 3836 17666 3892 17678
rect 3836 17614 3838 17666
rect 3890 17614 3892 17666
rect 3836 17332 3892 17614
rect 3388 16706 3444 16716
rect 3500 16884 3556 16894
rect 3836 16884 3892 17276
rect 3556 16828 3892 16884
rect 2492 15204 2548 15214
rect 2492 14642 2548 15148
rect 3500 15148 3556 16828
rect 3612 16658 3668 16670
rect 3612 16606 3614 16658
rect 3666 16606 3668 16658
rect 3612 16324 3668 16606
rect 3836 16660 3892 16670
rect 3948 16660 4004 17836
rect 4172 18228 4228 18958
rect 4284 19012 4340 19022
rect 4284 18918 4340 18956
rect 4620 18452 4676 18462
rect 4732 18452 4788 19180
rect 4956 19170 5012 19180
rect 5068 19236 5124 19742
rect 5068 18900 5124 19180
rect 4956 18844 5124 18900
rect 5180 19460 5236 19470
rect 4676 18396 4788 18452
rect 4844 18564 4900 18574
rect 4620 18338 4676 18396
rect 4620 18286 4622 18338
rect 4674 18286 4676 18338
rect 4620 18274 4676 18286
rect 4172 17332 4228 18172
rect 4476 18060 4740 18070
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4476 17994 4740 18004
rect 4732 17556 4788 17566
rect 4844 17556 4900 18508
rect 4732 17554 4900 17556
rect 4732 17502 4734 17554
rect 4786 17502 4900 17554
rect 4732 17500 4900 17502
rect 4732 17490 4788 17500
rect 4172 17276 4340 17332
rect 4172 17108 4228 17118
rect 4172 16882 4228 17052
rect 4284 17106 4340 17276
rect 4284 17054 4286 17106
rect 4338 17054 4340 17106
rect 4284 17042 4340 17054
rect 4172 16830 4174 16882
rect 4226 16830 4228 16882
rect 4172 16818 4228 16830
rect 4508 16882 4564 16894
rect 4508 16830 4510 16882
rect 4562 16830 4564 16882
rect 4396 16770 4452 16782
rect 4396 16718 4398 16770
rect 4450 16718 4452 16770
rect 4396 16660 4452 16718
rect 3836 16658 4004 16660
rect 3836 16606 3838 16658
rect 3890 16606 4004 16658
rect 3836 16604 4004 16606
rect 4172 16604 4452 16660
rect 4508 16660 4564 16830
rect 3836 16594 3892 16604
rect 4172 16324 4228 16604
rect 4508 16594 4564 16604
rect 4476 16492 4740 16502
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4476 16426 4740 16436
rect 3612 16258 3668 16268
rect 3836 16268 4228 16324
rect 3836 16210 3892 16268
rect 3836 16158 3838 16210
rect 3890 16158 3892 16210
rect 3836 16146 3892 16158
rect 4620 16212 4676 16222
rect 4620 16098 4676 16156
rect 4620 16046 4622 16098
rect 4674 16046 4676 16098
rect 4620 16034 4676 16046
rect 4732 15540 4788 15550
rect 4844 15540 4900 17500
rect 4956 16994 5012 18844
rect 5180 18676 5236 19404
rect 5292 19348 5348 19964
rect 5404 19954 5460 19964
rect 5628 20018 5684 20076
rect 5628 19966 5630 20018
rect 5682 19966 5684 20018
rect 5628 19796 5684 19966
rect 5292 19012 5348 19292
rect 5292 18946 5348 18956
rect 5404 19740 5684 19796
rect 5740 19908 5796 19918
rect 5404 19236 5460 19740
rect 5740 19348 5796 19852
rect 5292 18676 5348 18686
rect 5180 18674 5348 18676
rect 5180 18622 5294 18674
rect 5346 18622 5348 18674
rect 5180 18620 5348 18622
rect 5292 18610 5348 18620
rect 5068 18564 5124 18574
rect 5068 18470 5124 18508
rect 5180 18340 5236 18350
rect 5180 18246 5236 18284
rect 5180 18004 5236 18014
rect 5068 17444 5124 17454
rect 5068 17350 5124 17388
rect 5068 17108 5124 17118
rect 5180 17108 5236 17948
rect 5124 17052 5236 17108
rect 5068 17014 5124 17052
rect 4956 16942 4958 16994
rect 5010 16942 5012 16994
rect 4956 16930 5012 16942
rect 5292 16996 5348 17006
rect 5292 16902 5348 16940
rect 5292 16772 5348 16782
rect 4732 15538 4900 15540
rect 4732 15486 4734 15538
rect 4786 15486 4900 15538
rect 4732 15484 4900 15486
rect 4956 16660 5012 16670
rect 4956 15538 5012 16604
rect 5180 16548 5236 16558
rect 4956 15486 4958 15538
rect 5010 15486 5012 15538
rect 4732 15148 4788 15484
rect 4956 15474 5012 15486
rect 5068 16212 5124 16222
rect 4956 15316 5012 15326
rect 3500 15092 3780 15148
rect 2492 14590 2494 14642
rect 2546 14590 2548 14642
rect 2492 14578 2548 14590
rect 1820 14478 1822 14530
rect 1874 14478 1876 14530
rect 1820 12962 1876 14478
rect 2492 13636 2548 13646
rect 2492 13074 2548 13580
rect 2492 13022 2494 13074
rect 2546 13022 2548 13074
rect 2492 13010 2548 13022
rect 1820 12910 1822 12962
rect 1874 12910 1876 12962
rect 1820 11394 1876 12910
rect 3164 12404 3220 12414
rect 3164 12310 3220 12348
rect 3612 12292 3668 12302
rect 3388 12178 3444 12190
rect 3388 12126 3390 12178
rect 3442 12126 3444 12178
rect 2492 12068 2548 12078
rect 2492 11506 2548 12012
rect 3276 12068 3332 12078
rect 3276 11974 3332 12012
rect 3388 11620 3444 12126
rect 3612 12178 3668 12236
rect 3612 12126 3614 12178
rect 3666 12126 3668 12178
rect 3612 12114 3668 12126
rect 3388 11554 3444 11564
rect 2492 11454 2494 11506
rect 2546 11454 2548 11506
rect 2492 11442 2548 11454
rect 1820 11342 1822 11394
rect 1874 11342 1876 11394
rect 1708 9940 1764 9950
rect 1708 9846 1764 9884
rect 1820 8260 1876 11342
rect 2492 9268 2548 9278
rect 2492 8370 2548 9212
rect 2492 8318 2494 8370
rect 2546 8318 2548 8370
rect 2492 8306 2548 8318
rect 1820 8166 1876 8204
rect 3276 8260 3332 8270
rect 3276 7474 3332 8204
rect 3276 7422 3278 7474
rect 3330 7422 3332 7474
rect 3276 7410 3332 7422
rect 3724 7252 3780 15092
rect 4284 15092 4788 15148
rect 4844 15204 4900 15242
rect 4844 15138 4900 15148
rect 4284 12404 4340 15092
rect 4476 14924 4740 14934
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4476 14858 4740 14868
rect 4620 14644 4676 14654
rect 4620 14550 4676 14588
rect 4620 13972 4676 13982
rect 4956 13972 5012 15260
rect 5068 14306 5124 16156
rect 5068 14254 5070 14306
rect 5122 14254 5124 14306
rect 5068 14084 5124 14254
rect 5068 14018 5124 14028
rect 4620 13970 5012 13972
rect 4620 13918 4622 13970
rect 4674 13918 5012 13970
rect 4620 13916 5012 13918
rect 4620 13906 4676 13916
rect 4844 13746 4900 13758
rect 4844 13694 4846 13746
rect 4898 13694 4900 13746
rect 4732 13636 4788 13646
rect 4732 13542 4788 13580
rect 4476 13356 4740 13366
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4476 13290 4740 13300
rect 4844 13300 4900 13694
rect 5068 13748 5124 13758
rect 5180 13748 5236 16492
rect 5292 15316 5348 16716
rect 5292 15250 5348 15260
rect 5404 15314 5460 19180
rect 5516 19292 5796 19348
rect 5852 19348 5908 21532
rect 6076 21140 6132 22092
rect 6300 22146 6356 22158
rect 6300 22094 6302 22146
rect 6354 22094 6356 22146
rect 6300 21810 6356 22094
rect 6300 21758 6302 21810
rect 6354 21758 6356 21810
rect 6300 21746 6356 21758
rect 6748 21700 6804 21710
rect 5964 21084 6132 21140
rect 6188 21586 6244 21598
rect 6188 21534 6190 21586
rect 6242 21534 6244 21586
rect 5964 20132 6020 21084
rect 5964 20066 6020 20076
rect 6076 20916 6132 20926
rect 6188 20916 6244 21534
rect 6076 20914 6244 20916
rect 6076 20862 6078 20914
rect 6130 20862 6244 20914
rect 6076 20860 6244 20862
rect 6412 21586 6468 21598
rect 6412 21534 6414 21586
rect 6466 21534 6468 21586
rect 6076 20020 6132 20860
rect 6076 19954 6132 19964
rect 6412 19908 6468 21534
rect 6524 20804 6580 20814
rect 6524 20710 6580 20748
rect 6748 20802 6804 21644
rect 6748 20750 6750 20802
rect 6802 20750 6804 20802
rect 6300 19348 6356 19358
rect 5852 19346 6356 19348
rect 5852 19294 5854 19346
rect 5906 19294 6302 19346
rect 6354 19294 6356 19346
rect 5852 19292 6356 19294
rect 5516 18450 5572 19292
rect 5852 19282 5908 19292
rect 6300 19282 6356 19292
rect 6412 19124 6468 19852
rect 6300 19068 6468 19124
rect 6524 20244 6580 20254
rect 5516 18398 5518 18450
rect 5570 18398 5572 18450
rect 5516 18386 5572 18398
rect 6076 19012 6132 19022
rect 5740 18226 5796 18238
rect 5740 18174 5742 18226
rect 5794 18174 5796 18226
rect 5740 18004 5796 18174
rect 5740 17938 5796 17948
rect 5852 17780 5908 17790
rect 5628 17668 5684 17678
rect 5628 17574 5684 17612
rect 5852 17554 5908 17724
rect 5852 17502 5854 17554
rect 5906 17502 5908 17554
rect 5852 17490 5908 17502
rect 5964 17556 6020 17566
rect 5964 17462 6020 17500
rect 5740 17444 5796 17454
rect 5740 17106 5796 17388
rect 6076 17332 6132 18956
rect 5740 17054 5742 17106
rect 5794 17054 5796 17106
rect 5740 17042 5796 17054
rect 5852 17276 6132 17332
rect 6188 18338 6244 18350
rect 6188 18286 6190 18338
rect 6242 18286 6244 18338
rect 5628 16660 5684 16670
rect 5628 15426 5684 16604
rect 5852 16324 5908 17276
rect 6076 16994 6132 17006
rect 6076 16942 6078 16994
rect 6130 16942 6132 16994
rect 6076 16772 6132 16942
rect 6076 16706 6132 16716
rect 5852 16210 5908 16268
rect 5852 16158 5854 16210
rect 5906 16158 5908 16210
rect 5852 16146 5908 16158
rect 6188 16212 6244 18286
rect 6300 17668 6356 19068
rect 6524 18116 6580 20188
rect 6748 18564 6804 20750
rect 6860 20244 6916 22204
rect 6972 21812 7028 21822
rect 6972 21718 7028 21756
rect 7420 21698 7476 21710
rect 7420 21646 7422 21698
rect 7474 21646 7476 21698
rect 7420 21476 7476 21646
rect 7308 21026 7364 21038
rect 7308 20974 7310 21026
rect 7362 20974 7364 21026
rect 6860 20188 7028 20244
rect 6524 18050 6580 18060
rect 6636 18508 6804 18564
rect 6860 20020 6916 20030
rect 6300 17602 6356 17612
rect 6412 17668 6468 17678
rect 6412 17666 6580 17668
rect 6412 17614 6414 17666
rect 6466 17614 6580 17666
rect 6412 17612 6580 17614
rect 6412 17602 6468 17612
rect 6524 17108 6580 17612
rect 6636 17556 6692 18508
rect 6636 17490 6692 17500
rect 6748 18338 6804 18350
rect 6748 18286 6750 18338
rect 6802 18286 6804 18338
rect 6748 17554 6804 18286
rect 6860 17780 6916 19964
rect 6972 19348 7028 20188
rect 7084 19348 7140 19358
rect 6972 19346 7140 19348
rect 6972 19294 7086 19346
rect 7138 19294 7140 19346
rect 6972 19292 7140 19294
rect 7084 19282 7140 19292
rect 7308 18788 7364 20974
rect 7420 20356 7476 21420
rect 7420 20290 7476 20300
rect 7532 20244 7588 24444
rect 7980 23380 8036 23390
rect 8092 23380 8148 24892
rect 8316 24722 8372 26796
rect 8764 26852 8932 26908
rect 8988 27300 9044 27310
rect 8988 26908 9044 27244
rect 9100 27188 9156 27198
rect 9100 27074 9156 27132
rect 9100 27022 9102 27074
rect 9154 27022 9156 27074
rect 9100 27010 9156 27022
rect 8988 26852 9156 26908
rect 8652 26292 8708 26302
rect 8316 24670 8318 24722
rect 8370 24670 8372 24722
rect 8316 24658 8372 24670
rect 8428 26290 8708 26292
rect 8428 26238 8654 26290
rect 8706 26238 8708 26290
rect 8428 26236 8708 26238
rect 7980 23378 8148 23380
rect 7980 23326 7982 23378
rect 8034 23326 8148 23378
rect 7980 23324 8148 23326
rect 8204 24052 8260 24062
rect 8428 24052 8484 26236
rect 8652 26226 8708 26236
rect 8260 23996 8484 24052
rect 8652 25844 8708 25854
rect 8204 23378 8260 23996
rect 8204 23326 8206 23378
rect 8258 23326 8260 23378
rect 7980 23314 8036 23324
rect 8204 23314 8260 23326
rect 8428 23714 8484 23726
rect 8428 23662 8430 23714
rect 8482 23662 8484 23714
rect 8316 23154 8372 23166
rect 8316 23102 8318 23154
rect 8370 23102 8372 23154
rect 7644 23044 7700 23054
rect 7644 22950 7700 22988
rect 8092 22708 8148 22718
rect 7980 22372 8036 22382
rect 7868 22370 8036 22372
rect 7868 22318 7982 22370
rect 8034 22318 8036 22370
rect 7868 22316 8036 22318
rect 7756 22148 7812 22158
rect 7756 22054 7812 22092
rect 7868 21812 7924 22316
rect 7980 22306 8036 22316
rect 8092 21924 8148 22652
rect 7868 21746 7924 21756
rect 7980 21868 8148 21924
rect 8316 21924 8372 23102
rect 8428 22708 8484 23662
rect 8652 23716 8708 25788
rect 8652 23650 8708 23660
rect 8652 23268 8708 23278
rect 8764 23268 8820 26852
rect 8988 26516 9044 26526
rect 8988 26422 9044 26460
rect 8876 25730 8932 25742
rect 8876 25678 8878 25730
rect 8930 25678 8932 25730
rect 8876 24612 8932 25678
rect 8988 24724 9044 24734
rect 9100 24724 9156 26852
rect 8988 24722 9156 24724
rect 8988 24670 8990 24722
rect 9042 24670 9156 24722
rect 8988 24668 9156 24670
rect 8988 24658 9044 24668
rect 8876 23938 8932 24556
rect 8876 23886 8878 23938
rect 8930 23886 8932 23938
rect 8876 23874 8932 23886
rect 9212 23828 9268 29148
rect 9436 28868 9492 28878
rect 9660 28868 9716 29372
rect 9492 28812 9716 28868
rect 9772 29204 9828 29214
rect 9436 28082 9492 28812
rect 9772 28644 9828 29148
rect 10108 29202 10164 29214
rect 10108 29150 10110 29202
rect 10162 29150 10164 29202
rect 10108 29092 10164 29150
rect 10108 29026 10164 29036
rect 9772 28550 9828 28588
rect 9996 28642 10052 28654
rect 9996 28590 9998 28642
rect 10050 28590 10052 28642
rect 9436 28030 9438 28082
rect 9490 28030 9492 28082
rect 9436 28018 9492 28030
rect 9772 27748 9828 27758
rect 9772 27654 9828 27692
rect 9548 27636 9604 27646
rect 9548 27186 9604 27580
rect 9996 27636 10052 28590
rect 10108 27860 10164 27870
rect 10108 27766 10164 27804
rect 9996 27570 10052 27580
rect 9548 27134 9550 27186
rect 9602 27134 9604 27186
rect 9548 27122 9604 27134
rect 10108 27524 10164 27534
rect 10220 27524 10276 30156
rect 10332 29988 10388 29998
rect 10444 29988 10500 33964
rect 10556 34018 10612 34300
rect 10668 34130 10724 35420
rect 10780 35410 10836 35420
rect 11228 35308 11284 37660
rect 11788 37492 11844 37502
rect 11788 37490 12068 37492
rect 11788 37438 11790 37490
rect 11842 37438 12068 37490
rect 11788 37436 12068 37438
rect 11788 37426 11844 37436
rect 11676 37380 11732 37390
rect 11676 37286 11732 37324
rect 11564 37268 11620 37278
rect 11564 37174 11620 37212
rect 11452 36820 11508 36830
rect 11116 35252 11284 35308
rect 11340 35812 11396 35822
rect 10668 34078 10670 34130
rect 10722 34078 10724 34130
rect 10668 34066 10724 34078
rect 10892 35140 10948 35150
rect 10892 34914 10948 35084
rect 10892 34862 10894 34914
rect 10946 34862 10948 34914
rect 10556 33966 10558 34018
rect 10610 33966 10612 34018
rect 10556 33954 10612 33966
rect 10556 33684 10612 33694
rect 10556 30548 10612 33628
rect 10668 33236 10724 33246
rect 10668 32674 10724 33180
rect 10668 32622 10670 32674
rect 10722 32622 10724 32674
rect 10668 32610 10724 32622
rect 10668 32004 10724 32014
rect 10668 31556 10724 31948
rect 10668 31490 10724 31500
rect 10780 31668 10836 31678
rect 10780 31220 10836 31612
rect 10556 30482 10612 30492
rect 10668 31218 10836 31220
rect 10668 31166 10782 31218
rect 10834 31166 10836 31218
rect 10668 31164 10836 31166
rect 10668 30436 10724 31164
rect 10780 31154 10836 31164
rect 10892 30996 10948 34862
rect 11116 34804 11172 35196
rect 11340 35140 11396 35756
rect 11340 35074 11396 35084
rect 11116 34738 11172 34748
rect 11340 34914 11396 34926
rect 11340 34862 11342 34914
rect 11394 34862 11396 34914
rect 11340 34356 11396 34862
rect 11452 34916 11508 36764
rect 11564 36708 11620 36718
rect 11564 36614 11620 36652
rect 11676 36596 11732 36606
rect 11676 35924 11732 36540
rect 11676 35922 11956 35924
rect 11676 35870 11678 35922
rect 11730 35870 11956 35922
rect 11676 35868 11956 35870
rect 11676 35858 11732 35868
rect 11900 35028 11956 35868
rect 12012 35698 12068 37436
rect 12012 35646 12014 35698
rect 12066 35646 12068 35698
rect 12012 35634 12068 35646
rect 12012 35028 12068 35038
rect 11900 35026 12068 35028
rect 11900 34974 12014 35026
rect 12066 34974 12068 35026
rect 11900 34972 12068 34974
rect 12012 34962 12068 34972
rect 11452 34860 11620 34916
rect 11340 34290 11396 34300
rect 11452 34692 11508 34702
rect 11452 34130 11508 34636
rect 11452 34078 11454 34130
rect 11506 34078 11508 34130
rect 11452 34066 11508 34078
rect 11452 33796 11508 33806
rect 11116 33460 11172 33470
rect 11116 33346 11172 33404
rect 11116 33294 11118 33346
rect 11170 33294 11172 33346
rect 11116 32116 11172 33294
rect 11116 32050 11172 32060
rect 11340 32004 11396 32014
rect 11004 31780 11060 31790
rect 11004 31686 11060 31724
rect 10668 30370 10724 30380
rect 10780 30940 10948 30996
rect 11116 31444 11172 31454
rect 11116 31218 11172 31388
rect 11116 31166 11118 31218
rect 11170 31166 11172 31218
rect 10332 29986 10444 29988
rect 10332 29934 10334 29986
rect 10386 29934 10444 29986
rect 10332 29932 10444 29934
rect 10332 29922 10388 29932
rect 10444 29894 10500 29932
rect 10556 30210 10612 30222
rect 10556 30158 10558 30210
rect 10610 30158 10612 30210
rect 10556 29652 10612 30158
rect 10780 29764 10836 30940
rect 11116 30660 11172 31166
rect 11116 30594 11172 30604
rect 11228 30436 11284 30446
rect 10892 30212 10948 30222
rect 10892 29986 10948 30156
rect 11228 30210 11284 30380
rect 11228 30158 11230 30210
rect 11282 30158 11284 30210
rect 11228 30146 11284 30158
rect 10892 29934 10894 29986
rect 10946 29934 10948 29986
rect 10892 29922 10948 29934
rect 11004 30098 11060 30110
rect 11004 30046 11006 30098
rect 11058 30046 11060 30098
rect 10780 29708 10948 29764
rect 10556 29586 10612 29596
rect 10668 29540 10724 29550
rect 10332 29204 10388 29214
rect 10332 29110 10388 29148
rect 10556 29204 10612 29214
rect 10444 29092 10500 29102
rect 10444 28866 10500 29036
rect 10444 28814 10446 28866
rect 10498 28814 10500 28866
rect 10444 28756 10500 28814
rect 10444 28690 10500 28700
rect 10556 28642 10612 29148
rect 10556 28590 10558 28642
rect 10610 28590 10612 28642
rect 10332 27860 10388 27870
rect 10332 27636 10388 27804
rect 10444 27860 10500 27870
rect 10556 27860 10612 28590
rect 10444 27858 10612 27860
rect 10444 27806 10446 27858
rect 10498 27806 10612 27858
rect 10444 27804 10612 27806
rect 10444 27794 10500 27804
rect 10332 27580 10612 27636
rect 10220 27468 10500 27524
rect 10108 27188 10164 27468
rect 10220 27188 10276 27198
rect 10108 27186 10276 27188
rect 10108 27134 10222 27186
rect 10274 27134 10276 27186
rect 10108 27132 10276 27134
rect 10220 27122 10276 27132
rect 9324 27076 9380 27086
rect 9324 25620 9380 27020
rect 10332 26852 10388 26862
rect 9548 26290 9604 26302
rect 9548 26238 9550 26290
rect 9602 26238 9604 26290
rect 9548 25844 9604 26238
rect 9884 26290 9940 26302
rect 9884 26238 9886 26290
rect 9938 26238 9940 26290
rect 9884 25956 9940 26238
rect 9996 26292 10052 26302
rect 9996 26198 10052 26236
rect 10108 26290 10164 26302
rect 10108 26238 10110 26290
rect 10162 26238 10164 26290
rect 10108 26180 10164 26238
rect 10332 26180 10388 26796
rect 10444 26292 10500 27468
rect 10556 27074 10612 27580
rect 10556 27022 10558 27074
rect 10610 27022 10612 27074
rect 10556 26964 10612 27022
rect 10556 26898 10612 26908
rect 10668 26852 10724 29484
rect 10780 29426 10836 29438
rect 10780 29374 10782 29426
rect 10834 29374 10836 29426
rect 10780 27860 10836 29374
rect 10892 28868 10948 29708
rect 11004 29092 11060 30046
rect 11116 29540 11172 29550
rect 11116 29446 11172 29484
rect 11004 29026 11060 29036
rect 10892 28812 11060 28868
rect 10780 27794 10836 27804
rect 10892 28644 10948 28654
rect 10668 26786 10724 26796
rect 10780 27076 10836 27086
rect 10780 26628 10836 27020
rect 10892 26740 10948 28588
rect 11004 26908 11060 28812
rect 11228 28644 11284 28654
rect 11228 28550 11284 28588
rect 11228 27970 11284 27982
rect 11228 27918 11230 27970
rect 11282 27918 11284 27970
rect 11228 27748 11284 27918
rect 11228 27682 11284 27692
rect 11340 27412 11396 31948
rect 11452 32002 11508 33740
rect 11564 33234 11620 34860
rect 11676 34804 11732 34814
rect 11676 34710 11732 34748
rect 12012 34130 12068 34142
rect 12012 34078 12014 34130
rect 12066 34078 12068 34130
rect 12012 33460 12068 34078
rect 12124 33572 12180 37996
rect 12348 37958 12404 37996
rect 12460 37940 12516 37950
rect 12460 37846 12516 37884
rect 12460 37716 12516 37726
rect 12348 36260 12404 36270
rect 12348 36166 12404 36204
rect 12348 35476 12404 35486
rect 12236 35252 12292 35262
rect 12236 34914 12292 35196
rect 12236 34862 12238 34914
rect 12290 34862 12292 34914
rect 12236 34850 12292 34862
rect 12124 33506 12180 33516
rect 12012 33394 12068 33404
rect 12348 33460 12404 35420
rect 12460 34244 12516 37660
rect 12572 34468 12628 40684
rect 12908 39844 12964 41134
rect 13020 40516 13076 40526
rect 13020 40422 13076 40460
rect 12908 39778 12964 39788
rect 12684 39396 12740 39406
rect 12684 36372 12740 39340
rect 13020 39394 13076 39406
rect 13020 39342 13022 39394
rect 13074 39342 13076 39394
rect 12796 38162 12852 38174
rect 12796 38110 12798 38162
rect 12850 38110 12852 38162
rect 12796 37268 12852 38110
rect 12796 37202 12852 37212
rect 12796 36820 12852 36830
rect 12796 36706 12852 36764
rect 12796 36654 12798 36706
rect 12850 36654 12852 36706
rect 12796 36642 12852 36654
rect 12908 36596 12964 36606
rect 12908 36482 12964 36540
rect 12908 36430 12910 36482
rect 12962 36430 12964 36482
rect 12908 36418 12964 36430
rect 12796 36372 12852 36382
rect 12684 36370 12852 36372
rect 12684 36318 12798 36370
rect 12850 36318 12852 36370
rect 12684 36316 12852 36318
rect 12796 36306 12852 36316
rect 13020 36260 13076 39342
rect 12908 34916 12964 34926
rect 12908 34822 12964 34860
rect 12572 34402 12628 34412
rect 13020 34356 13076 36204
rect 12908 34300 13076 34356
rect 12460 34150 12516 34188
rect 12684 34244 12740 34254
rect 11788 33348 11844 33358
rect 11788 33346 11956 33348
rect 11788 33294 11790 33346
rect 11842 33294 11956 33346
rect 11788 33292 11956 33294
rect 11788 33282 11844 33292
rect 11564 33182 11566 33234
rect 11618 33182 11620 33234
rect 11564 33170 11620 33182
rect 11676 33124 11732 33134
rect 11676 33030 11732 33068
rect 11788 32564 11844 32574
rect 11788 32470 11844 32508
rect 11452 31950 11454 32002
rect 11506 31950 11508 32002
rect 11452 31938 11508 31950
rect 11900 31890 11956 33292
rect 12348 33346 12404 33404
rect 12572 34130 12628 34142
rect 12572 34078 12574 34130
rect 12626 34078 12628 34130
rect 12572 33348 12628 34078
rect 12348 33294 12350 33346
rect 12402 33294 12404 33346
rect 12348 33282 12404 33294
rect 12460 33292 12628 33348
rect 12236 33178 12292 33190
rect 12012 33124 12068 33134
rect 12236 33126 12238 33178
rect 12290 33126 12292 33178
rect 12012 33122 12180 33124
rect 12012 33070 12014 33122
rect 12066 33070 12180 33122
rect 12012 33068 12180 33070
rect 12012 33058 12068 33068
rect 11900 31838 11902 31890
rect 11954 31838 11956 31890
rect 11900 31826 11956 31838
rect 12012 32452 12068 32462
rect 11564 31780 11620 31818
rect 11564 31714 11620 31724
rect 11452 31668 11508 31678
rect 11452 31574 11508 31612
rect 11564 30996 11620 31006
rect 11452 30940 11564 30996
rect 11452 29650 11508 30940
rect 11564 30902 11620 30940
rect 11900 30994 11956 31006
rect 11900 30942 11902 30994
rect 11954 30942 11956 30994
rect 11452 29598 11454 29650
rect 11506 29598 11508 29650
rect 11452 29586 11508 29598
rect 11900 30210 11956 30942
rect 11900 30158 11902 30210
rect 11954 30158 11956 30210
rect 11900 29650 11956 30158
rect 11900 29598 11902 29650
rect 11954 29598 11956 29650
rect 11900 29586 11956 29598
rect 12012 29988 12068 32396
rect 12124 31780 12180 33068
rect 12236 32452 12292 33126
rect 12236 32386 12292 32396
rect 12348 33012 12404 33022
rect 12124 31686 12180 31724
rect 12124 29988 12180 29998
rect 12012 29986 12180 29988
rect 12012 29934 12126 29986
rect 12178 29934 12180 29986
rect 12012 29932 12180 29934
rect 11788 29316 11844 29326
rect 11788 29092 11844 29260
rect 11564 29036 11844 29092
rect 11564 28420 11620 29036
rect 11788 28642 11844 28654
rect 11788 28590 11790 28642
rect 11842 28590 11844 28642
rect 11340 27346 11396 27356
rect 11452 28364 11620 28420
rect 11676 28418 11732 28430
rect 11676 28366 11678 28418
rect 11730 28366 11732 28418
rect 11116 27188 11172 27226
rect 11116 27122 11172 27132
rect 11004 26852 11172 26908
rect 10892 26684 11060 26740
rect 10556 26572 10836 26628
rect 10556 26514 10612 26572
rect 10892 26516 10948 26526
rect 10556 26462 10558 26514
rect 10610 26462 10612 26514
rect 10556 26450 10612 26462
rect 10780 26460 10892 26516
rect 10444 26236 10612 26292
rect 10164 26124 10500 26180
rect 10108 26114 10164 26124
rect 10444 26066 10500 26124
rect 10444 26014 10446 26066
rect 10498 26014 10500 26066
rect 10444 26002 10500 26014
rect 9884 25890 9940 25900
rect 9548 25778 9604 25788
rect 10108 25844 10164 25854
rect 9324 25554 9380 25564
rect 10108 25506 10164 25788
rect 10108 25454 10110 25506
rect 10162 25454 10164 25506
rect 10108 25442 10164 25454
rect 10444 25508 10500 25518
rect 10556 25508 10612 26236
rect 10780 26290 10836 26460
rect 10892 26450 10948 26460
rect 10780 26238 10782 26290
rect 10834 26238 10836 26290
rect 10780 26226 10836 26238
rect 10668 25508 10724 25518
rect 10556 25506 10724 25508
rect 10556 25454 10670 25506
rect 10722 25454 10724 25506
rect 10556 25452 10724 25454
rect 10444 25414 10500 25452
rect 10668 25442 10724 25452
rect 9772 25396 9828 25406
rect 9212 23762 9268 23772
rect 9324 25394 9828 25396
rect 9324 25342 9774 25394
rect 9826 25342 9828 25394
rect 9324 25340 9828 25342
rect 8988 23716 9044 23726
rect 8988 23378 9044 23660
rect 9212 23604 9268 23614
rect 8988 23326 8990 23378
rect 9042 23326 9044 23378
rect 8988 23314 9044 23326
rect 9100 23548 9212 23604
rect 8708 23212 8820 23268
rect 8652 23174 8708 23212
rect 8428 22642 8484 22652
rect 8764 22820 8820 22830
rect 8764 22258 8820 22764
rect 8764 22206 8766 22258
rect 8818 22206 8820 22258
rect 8764 21924 8820 22206
rect 8876 22260 8932 22270
rect 8876 22166 8932 22204
rect 8316 21868 8484 21924
rect 7980 21810 8036 21868
rect 7980 21758 7982 21810
rect 8034 21758 8036 21810
rect 7644 21700 7700 21710
rect 7644 21606 7700 21644
rect 7756 21698 7812 21710
rect 7756 21646 7758 21698
rect 7810 21646 7812 21698
rect 7532 20178 7588 20188
rect 7644 21474 7700 21486
rect 7644 21422 7646 21474
rect 7698 21422 7700 21474
rect 7420 19908 7476 19918
rect 7420 19814 7476 19852
rect 7420 19012 7476 19022
rect 7420 18918 7476 18956
rect 7644 18788 7700 21422
rect 7756 20804 7812 21646
rect 7980 20914 8036 21758
rect 8092 21700 8148 21710
rect 8316 21700 8372 21710
rect 8148 21698 8372 21700
rect 8148 21646 8318 21698
rect 8370 21646 8372 21698
rect 8148 21644 8372 21646
rect 8092 21634 8148 21644
rect 8316 21634 8372 21644
rect 8428 21252 8484 21868
rect 8764 21858 8820 21868
rect 8652 21812 8708 21822
rect 8652 21718 8708 21756
rect 8428 21186 8484 21196
rect 8988 21476 9044 21486
rect 7980 20862 7982 20914
rect 8034 20862 8036 20914
rect 7868 20804 7924 20814
rect 7756 20748 7868 20804
rect 7868 20710 7924 20748
rect 7980 20580 8036 20862
rect 8876 20804 8932 20814
rect 8876 20710 8932 20748
rect 8764 20580 8820 20590
rect 7756 20524 8036 20580
rect 8652 20578 8820 20580
rect 8652 20526 8766 20578
rect 8818 20526 8820 20578
rect 8652 20524 8820 20526
rect 7756 20132 7812 20524
rect 8204 20244 8260 20254
rect 8092 20188 8204 20244
rect 8260 20188 8372 20244
rect 7980 20132 8036 20142
rect 7756 20130 8036 20132
rect 7756 20078 7982 20130
rect 8034 20078 8036 20130
rect 7756 20076 8036 20078
rect 7980 20066 8036 20076
rect 8092 19234 8148 20188
rect 8204 20178 8260 20188
rect 8316 20018 8372 20188
rect 8652 20132 8708 20524
rect 8764 20514 8820 20524
rect 8652 20066 8708 20076
rect 8988 20130 9044 21420
rect 9100 20804 9156 23548
rect 9212 23538 9268 23548
rect 9212 22484 9268 22494
rect 9212 22370 9268 22428
rect 9212 22318 9214 22370
rect 9266 22318 9268 22370
rect 9212 22306 9268 22318
rect 9324 22260 9380 25340
rect 9772 25330 9828 25340
rect 10108 25282 10164 25294
rect 10108 25230 10110 25282
rect 10162 25230 10164 25282
rect 9996 25172 10052 25182
rect 9548 24724 9604 24734
rect 9548 24630 9604 24668
rect 9996 23826 10052 25116
rect 9996 23774 9998 23826
rect 10050 23774 10052 23826
rect 9996 23716 10052 23774
rect 9996 23650 10052 23660
rect 10108 23604 10164 25230
rect 10780 24836 10836 24846
rect 10556 23716 10612 23726
rect 10612 23660 10724 23716
rect 10556 23650 10612 23660
rect 10108 23538 10164 23548
rect 9436 23380 9492 23390
rect 9436 22932 9492 23324
rect 10108 23268 10164 23278
rect 9660 23156 9716 23166
rect 9660 23062 9716 23100
rect 9884 23156 9940 23166
rect 9884 23154 10052 23156
rect 9884 23102 9886 23154
rect 9938 23102 10052 23154
rect 9884 23100 10052 23102
rect 9884 23090 9940 23100
rect 9436 22866 9492 22876
rect 9772 23042 9828 23054
rect 9772 22990 9774 23042
rect 9826 22990 9828 23042
rect 9772 22484 9828 22990
rect 9772 22418 9828 22428
rect 9884 22932 9940 22942
rect 9324 22166 9380 22204
rect 9772 22258 9828 22270
rect 9772 22206 9774 22258
rect 9826 22206 9828 22258
rect 9548 22148 9604 22158
rect 9548 22146 9716 22148
rect 9548 22094 9550 22146
rect 9602 22094 9716 22146
rect 9548 22092 9716 22094
rect 9548 22082 9604 22092
rect 9212 20804 9268 20814
rect 9436 20804 9492 20814
rect 9100 20802 9492 20804
rect 9100 20750 9214 20802
rect 9266 20750 9438 20802
rect 9490 20750 9492 20802
rect 9100 20748 9492 20750
rect 9212 20738 9268 20748
rect 9436 20738 9492 20748
rect 9100 20580 9156 20590
rect 9100 20578 9268 20580
rect 9100 20526 9102 20578
rect 9154 20526 9268 20578
rect 9100 20524 9268 20526
rect 9100 20514 9156 20524
rect 8988 20078 8990 20130
rect 9042 20078 9044 20130
rect 8988 20066 9044 20078
rect 9100 20356 9156 20366
rect 8316 19966 8318 20018
rect 8370 19966 8372 20018
rect 8316 19954 8372 19966
rect 8540 20020 8596 20030
rect 8540 19460 8596 19964
rect 8764 20020 8820 20030
rect 8764 20018 8932 20020
rect 8764 19966 8766 20018
rect 8818 19966 8932 20018
rect 8764 19964 8932 19966
rect 8764 19954 8820 19964
rect 8092 19182 8094 19234
rect 8146 19182 8148 19234
rect 8092 19170 8148 19182
rect 8204 19404 8596 19460
rect 8652 19906 8708 19918
rect 8652 19854 8654 19906
rect 8706 19854 8708 19906
rect 8204 19234 8260 19404
rect 8652 19348 8708 19854
rect 8540 19292 8708 19348
rect 8764 19796 8820 19806
rect 8764 19346 8820 19740
rect 8764 19294 8766 19346
rect 8818 19294 8820 19346
rect 8204 19182 8206 19234
rect 8258 19182 8260 19234
rect 8204 19170 8260 19182
rect 8428 19236 8484 19246
rect 8428 19142 8484 19180
rect 8204 19012 8260 19022
rect 6972 18732 7364 18788
rect 7420 18732 8036 18788
rect 6972 18004 7028 18732
rect 7420 18674 7476 18732
rect 7420 18622 7422 18674
rect 7474 18622 7476 18674
rect 7420 18610 7476 18622
rect 7532 18620 7812 18676
rect 7084 18562 7140 18574
rect 7084 18510 7086 18562
rect 7138 18510 7140 18562
rect 7084 18228 7140 18510
rect 7084 18162 7140 18172
rect 7308 18228 7364 18238
rect 6972 17938 7028 17948
rect 7196 17890 7252 17902
rect 7196 17838 7198 17890
rect 7250 17838 7252 17890
rect 7084 17780 7140 17790
rect 6860 17724 7084 17780
rect 7084 17686 7140 17724
rect 7196 17668 7252 17838
rect 7196 17602 7252 17612
rect 6748 17502 6750 17554
rect 6802 17502 6804 17554
rect 6748 17332 6804 17502
rect 6748 17266 6804 17276
rect 7308 17220 7364 18172
rect 7196 17164 7364 17220
rect 6636 17108 6692 17118
rect 6524 17106 6692 17108
rect 6524 17054 6638 17106
rect 6690 17054 6692 17106
rect 6524 17052 6692 17054
rect 6636 16436 6692 17052
rect 6636 16370 6692 16380
rect 6188 16118 6244 16156
rect 7196 16322 7252 17164
rect 7420 17108 7476 17118
rect 7532 17108 7588 18620
rect 7756 18618 7812 18620
rect 7756 18566 7758 18618
rect 7810 18566 7812 18618
rect 7756 18554 7812 18566
rect 7980 18450 8036 18732
rect 7980 18398 7982 18450
rect 8034 18398 8036 18450
rect 7980 18386 8036 18398
rect 7868 18116 7924 18126
rect 7868 17780 7924 18060
rect 8204 18004 8260 18956
rect 8204 17938 8260 17948
rect 7420 17106 7588 17108
rect 7420 17054 7422 17106
rect 7474 17054 7588 17106
rect 7420 17052 7588 17054
rect 7644 17724 7924 17780
rect 7644 17106 7700 17724
rect 8204 17556 8260 17566
rect 8092 17554 8260 17556
rect 8092 17502 8206 17554
rect 8258 17502 8260 17554
rect 8092 17500 8260 17502
rect 7644 17054 7646 17106
rect 7698 17054 7700 17106
rect 7420 16548 7476 17052
rect 7644 17042 7700 17054
rect 7980 17444 8036 17454
rect 7420 16482 7476 16492
rect 7532 16770 7588 16782
rect 7532 16718 7534 16770
rect 7586 16718 7588 16770
rect 7196 16270 7198 16322
rect 7250 16270 7252 16322
rect 5628 15374 5630 15426
rect 5682 15374 5684 15426
rect 5628 15362 5684 15374
rect 7084 15428 7140 15438
rect 5404 15262 5406 15314
rect 5458 15262 5460 15314
rect 5404 15250 5460 15262
rect 6860 15316 6916 15354
rect 7084 15334 7140 15372
rect 6860 15250 6916 15260
rect 7196 15314 7252 16270
rect 7420 16100 7476 16110
rect 7420 16006 7476 16044
rect 7532 15876 7588 16718
rect 7868 16772 7924 16782
rect 7980 16772 8036 17388
rect 8092 16884 8148 17500
rect 8204 17490 8260 17500
rect 8540 17444 8596 19292
rect 8764 19282 8820 19294
rect 8876 19236 8932 19964
rect 8988 19236 9044 19246
rect 8876 19234 9044 19236
rect 8876 19182 8990 19234
rect 9042 19182 9044 19234
rect 8876 19180 9044 19182
rect 8988 19170 9044 19180
rect 8652 19122 8708 19134
rect 8652 19070 8654 19122
rect 8706 19070 8708 19122
rect 8652 18564 8708 19070
rect 9100 18788 9156 20300
rect 9212 19908 9268 20524
rect 9548 20020 9604 20030
rect 9548 19926 9604 19964
rect 9436 19908 9492 19918
rect 9212 19852 9436 19908
rect 9436 19842 9492 19852
rect 9660 19236 9716 22092
rect 9772 20132 9828 22206
rect 9884 20914 9940 22876
rect 9996 22484 10052 23100
rect 10108 23154 10164 23212
rect 10108 23102 10110 23154
rect 10162 23102 10164 23154
rect 10108 23090 10164 23102
rect 10556 23156 10612 23166
rect 10332 22930 10388 22942
rect 10332 22878 10334 22930
rect 10386 22878 10388 22930
rect 10332 22820 10388 22878
rect 10332 22754 10388 22764
rect 10220 22484 10276 22494
rect 9996 22482 10276 22484
rect 9996 22430 10222 22482
rect 10274 22430 10276 22482
rect 9996 22428 10276 22430
rect 10220 22418 10276 22428
rect 10444 22372 10500 22382
rect 10444 22278 10500 22316
rect 9996 22260 10052 22270
rect 9996 22166 10052 22204
rect 10556 22148 10612 23100
rect 10668 22594 10724 23660
rect 10780 23604 10836 24780
rect 10892 24724 10948 24734
rect 10892 24630 10948 24668
rect 10780 23538 10836 23548
rect 10892 23828 10948 23838
rect 10892 23268 10948 23772
rect 10668 22542 10670 22594
rect 10722 22542 10724 22594
rect 10668 22530 10724 22542
rect 10780 23266 10948 23268
rect 10780 23214 10894 23266
rect 10946 23214 10948 23266
rect 10780 23212 10948 23214
rect 10108 22092 10612 22148
rect 10108 21810 10164 22092
rect 10780 22036 10836 23212
rect 10892 23202 10948 23212
rect 10892 22594 10948 22606
rect 10892 22542 10894 22594
rect 10946 22542 10948 22594
rect 10892 22482 10948 22542
rect 10892 22430 10894 22482
rect 10946 22430 10948 22482
rect 10892 22418 10948 22430
rect 10108 21758 10110 21810
rect 10162 21758 10164 21810
rect 10108 21746 10164 21758
rect 10444 21980 10836 22036
rect 10332 21586 10388 21598
rect 10332 21534 10334 21586
rect 10386 21534 10388 21586
rect 10332 21364 10388 21534
rect 10108 21308 10332 21364
rect 9884 20862 9886 20914
rect 9938 20862 9940 20914
rect 9884 20850 9940 20862
rect 9996 21026 10052 21038
rect 9996 20974 9998 21026
rect 10050 20974 10052 21026
rect 9772 20066 9828 20076
rect 9436 19180 9716 19236
rect 9772 19908 9828 19918
rect 9324 19124 9380 19134
rect 9100 18722 9156 18732
rect 9212 19010 9268 19022
rect 9212 18958 9214 19010
rect 9266 18958 9268 19010
rect 8988 18564 9044 18574
rect 8652 18508 8988 18564
rect 8988 17890 9044 18508
rect 8988 17838 8990 17890
rect 9042 17838 9044 17890
rect 8988 17826 9044 17838
rect 9100 18340 9156 18350
rect 9212 18340 9268 18958
rect 9100 18338 9268 18340
rect 9100 18286 9102 18338
rect 9154 18286 9268 18338
rect 9100 18284 9268 18286
rect 8652 17666 8708 17678
rect 8652 17614 8654 17666
rect 8706 17614 8708 17666
rect 8652 17556 8708 17614
rect 8652 17490 8708 17500
rect 8876 17554 8932 17566
rect 8876 17502 8878 17554
rect 8930 17502 8932 17554
rect 8540 17378 8596 17388
rect 8428 17332 8484 17342
rect 8428 17108 8484 17276
rect 8540 17108 8596 17118
rect 8876 17108 8932 17502
rect 9100 17556 9156 18284
rect 9324 18004 9380 19068
rect 9100 17490 9156 17500
rect 9212 17948 9380 18004
rect 8428 17106 8932 17108
rect 8428 17054 8542 17106
rect 8594 17054 8932 17106
rect 8428 17052 8932 17054
rect 8540 17042 8596 17052
rect 8092 16790 8148 16828
rect 8540 16884 8596 16894
rect 7868 16770 8036 16772
rect 7868 16718 7870 16770
rect 7922 16718 8036 16770
rect 7868 16716 8036 16718
rect 7868 16706 7924 16716
rect 7644 16212 7700 16222
rect 7644 16118 7700 16156
rect 8428 16212 8484 16222
rect 8092 16100 8148 16110
rect 7196 15262 7198 15314
rect 7250 15262 7252 15314
rect 7196 15250 7252 15262
rect 7420 15820 7588 15876
rect 7756 16044 8092 16100
rect 5964 15202 6020 15214
rect 5964 15150 5966 15202
rect 6018 15150 6020 15202
rect 5964 15148 6020 15150
rect 6972 15202 7028 15214
rect 6972 15150 6974 15202
rect 7026 15150 7028 15202
rect 6972 15148 7028 15150
rect 5964 15092 6132 15148
rect 6076 14644 6132 15092
rect 5852 14084 5908 14094
rect 5068 13746 5236 13748
rect 5068 13694 5070 13746
rect 5122 13694 5236 13746
rect 5068 13692 5236 13694
rect 5068 13682 5124 13692
rect 4844 13244 5124 13300
rect 4732 13188 4788 13198
rect 4620 13074 4676 13086
rect 4620 13022 4622 13074
rect 4674 13022 4676 13074
rect 4620 12852 4676 13022
rect 4620 12786 4676 12796
rect 4284 12310 4340 12348
rect 4732 12292 4788 13132
rect 5068 13076 5124 13244
rect 5180 13188 5236 13692
rect 5404 13972 5460 13982
rect 5180 13122 5236 13132
rect 5292 13522 5348 13534
rect 5292 13470 5294 13522
rect 5346 13470 5348 13522
rect 3836 12180 3892 12190
rect 3836 12086 3892 12124
rect 4508 12180 4564 12190
rect 4508 12086 4564 12124
rect 4732 12178 4788 12236
rect 4732 12126 4734 12178
rect 4786 12126 4788 12178
rect 4732 12114 4788 12126
rect 4956 13020 5124 13076
rect 5292 13076 5348 13470
rect 4956 12962 5012 13020
rect 5292 13010 5348 13020
rect 4956 12910 4958 12962
rect 5010 12910 5012 12962
rect 4956 12178 5012 12910
rect 4956 12126 4958 12178
rect 5010 12126 5012 12178
rect 4956 12114 5012 12126
rect 5068 12852 5124 12862
rect 4396 12066 4452 12078
rect 4396 12014 4398 12066
rect 4450 12014 4452 12066
rect 4396 11956 4452 12014
rect 3948 11900 4452 11956
rect 3836 9940 3892 9950
rect 3948 9940 4004 11900
rect 4476 11788 4740 11798
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 5068 11788 5124 12796
rect 5404 12290 5460 13916
rect 5852 13746 5908 14028
rect 5852 13694 5854 13746
rect 5906 13694 5908 13746
rect 5852 13682 5908 13694
rect 5404 12238 5406 12290
rect 5458 12238 5460 12290
rect 5292 12180 5348 12190
rect 5292 12086 5348 12124
rect 5068 11732 5348 11788
rect 4476 11722 4740 11732
rect 4732 11620 4788 11630
rect 4788 11564 4900 11620
rect 4732 11554 4788 11564
rect 4620 11508 4676 11518
rect 4620 11414 4676 11452
rect 4844 11396 4900 11564
rect 4956 11396 5012 11406
rect 4844 11394 5012 11396
rect 4844 11342 4958 11394
rect 5010 11342 5012 11394
rect 4844 11340 5012 11342
rect 4956 11330 5012 11340
rect 5068 11284 5124 11294
rect 5124 11228 5236 11284
rect 5068 11190 5124 11228
rect 4956 10612 5012 10622
rect 4956 10518 5012 10556
rect 5180 10610 5236 11228
rect 5180 10558 5182 10610
rect 5234 10558 5236 10610
rect 5180 10546 5236 10558
rect 5292 10612 5348 11732
rect 5292 10546 5348 10556
rect 4844 10388 4900 10398
rect 3836 9938 4004 9940
rect 3836 9886 3838 9938
rect 3890 9886 4004 9938
rect 3836 9884 4004 9886
rect 4172 10386 4900 10388
rect 4172 10334 4846 10386
rect 4898 10334 4900 10386
rect 4172 10332 4900 10334
rect 3836 9874 3892 9884
rect 3836 9268 3892 9306
rect 3836 9202 3892 9212
rect 4060 9268 4116 9278
rect 3948 9044 4004 9054
rect 3948 8950 4004 8988
rect 4060 7586 4116 9212
rect 4172 9042 4228 10332
rect 4844 10322 4900 10332
rect 5292 10386 5348 10398
rect 5292 10334 5294 10386
rect 5346 10334 5348 10386
rect 4476 10220 4740 10230
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4476 10154 4740 10164
rect 5292 10052 5348 10334
rect 4620 9828 4676 9838
rect 5068 9828 5124 9838
rect 5292 9828 5348 9996
rect 5404 9940 5460 12238
rect 5628 12962 5684 12974
rect 5628 12910 5630 12962
rect 5682 12910 5684 12962
rect 5628 11508 5684 12910
rect 5852 12962 5908 12974
rect 5852 12910 5854 12962
rect 5906 12910 5908 12962
rect 5852 12852 5908 12910
rect 6076 12962 6132 14588
rect 6524 15092 7028 15148
rect 6524 13858 6580 15092
rect 7196 14530 7252 14542
rect 7196 14478 7198 14530
rect 7250 14478 7252 14530
rect 6524 13806 6526 13858
rect 6578 13806 6580 13858
rect 6524 13794 6580 13806
rect 6636 14084 6692 14094
rect 6636 13076 6692 14028
rect 7196 14084 7252 14478
rect 7196 14018 7252 14028
rect 7420 13636 7476 15820
rect 7532 15316 7588 15326
rect 7756 15316 7812 16044
rect 8092 16006 8148 16044
rect 8428 15988 8484 16156
rect 8316 15932 8484 15988
rect 7532 15314 7812 15316
rect 7532 15262 7534 15314
rect 7586 15262 7812 15314
rect 7532 15260 7812 15262
rect 7868 15874 7924 15886
rect 7868 15822 7870 15874
rect 7922 15822 7924 15874
rect 7868 15316 7924 15822
rect 7532 15250 7588 15260
rect 7868 15250 7924 15260
rect 7980 15874 8036 15886
rect 7980 15822 7982 15874
rect 8034 15822 8036 15874
rect 7980 15148 8036 15822
rect 7868 15092 8036 15148
rect 7868 14642 7924 15092
rect 7868 14590 7870 14642
rect 7922 14590 7924 14642
rect 7868 14578 7924 14590
rect 6076 12910 6078 12962
rect 6130 12910 6132 12962
rect 6076 12898 6132 12910
rect 6188 13074 6692 13076
rect 6188 13022 6638 13074
rect 6690 13022 6692 13074
rect 6188 13020 6692 13022
rect 5852 12786 5908 12796
rect 5740 12740 5796 12750
rect 5740 12646 5796 12684
rect 6188 12180 6244 13020
rect 6636 13010 6692 13020
rect 6860 13580 7476 13636
rect 6860 12290 6916 13580
rect 6860 12238 6862 12290
rect 6914 12238 6916 12290
rect 6860 12226 6916 12238
rect 6188 12178 6468 12180
rect 6188 12126 6190 12178
rect 6242 12126 6468 12178
rect 6188 12124 6468 12126
rect 6188 12114 6244 12124
rect 5628 11394 5684 11452
rect 5628 11342 5630 11394
rect 5682 11342 5684 11394
rect 5628 11330 5684 11342
rect 6412 11506 6468 12124
rect 8316 11956 8372 15932
rect 8540 12180 8596 16828
rect 9212 15148 9268 17948
rect 9436 15148 9492 19180
rect 9548 18452 9604 18462
rect 9548 17778 9604 18396
rect 9772 18450 9828 19852
rect 9884 19794 9940 19806
rect 9884 19742 9886 19794
rect 9938 19742 9940 19794
rect 9884 19124 9940 19742
rect 9884 19058 9940 19068
rect 9772 18398 9774 18450
rect 9826 18398 9828 18450
rect 9772 18386 9828 18398
rect 9548 17726 9550 17778
rect 9602 17726 9604 17778
rect 9548 17714 9604 17726
rect 9884 18226 9940 18238
rect 9884 18174 9886 18226
rect 9938 18174 9940 18226
rect 9772 17666 9828 17678
rect 9772 17614 9774 17666
rect 9826 17614 9828 17666
rect 9548 16994 9604 17006
rect 9548 16942 9550 16994
rect 9602 16942 9604 16994
rect 9548 16212 9604 16942
rect 9772 16772 9828 17614
rect 9884 17666 9940 18174
rect 9884 17614 9886 17666
rect 9938 17614 9940 17666
rect 9884 17602 9940 17614
rect 9884 17108 9940 17118
rect 9996 17108 10052 20974
rect 10108 20132 10164 21308
rect 10332 21298 10388 21308
rect 10332 20916 10388 20926
rect 10444 20916 10500 21980
rect 10892 21924 10948 21934
rect 10892 21586 10948 21868
rect 10892 21534 10894 21586
rect 10946 21534 10948 21586
rect 10332 20914 10500 20916
rect 10332 20862 10334 20914
rect 10386 20862 10500 20914
rect 10332 20860 10500 20862
rect 10668 20916 10724 20926
rect 10332 20850 10388 20860
rect 10556 20692 10612 20702
rect 10556 20598 10612 20636
rect 10668 20690 10724 20860
rect 10892 20804 10948 21534
rect 10892 20738 10948 20748
rect 11004 20914 11060 26684
rect 11116 25172 11172 26852
rect 11340 26852 11396 26862
rect 11340 26402 11396 26796
rect 11452 26516 11508 28364
rect 11564 28084 11620 28094
rect 11564 27990 11620 28028
rect 11564 27188 11620 27198
rect 11676 27188 11732 28366
rect 11788 28308 11844 28590
rect 11788 28084 11844 28252
rect 11788 28018 11844 28028
rect 11900 27748 11956 27758
rect 11900 27300 11956 27692
rect 12012 27524 12068 29932
rect 12124 29922 12180 29932
rect 12012 27458 12068 27468
rect 12124 28868 12180 28878
rect 11956 27244 12068 27300
rect 11900 27234 11956 27244
rect 11620 27132 11732 27188
rect 11788 27188 11844 27198
rect 11564 27122 11620 27132
rect 11788 27074 11844 27132
rect 11788 27022 11790 27074
rect 11842 27022 11844 27074
rect 11788 27010 11844 27022
rect 11900 27076 11956 27086
rect 11900 26982 11956 27020
rect 12012 26908 12068 27244
rect 11564 26852 11620 26862
rect 11564 26758 11620 26796
rect 11676 26850 11732 26862
rect 11676 26798 11678 26850
rect 11730 26798 11732 26850
rect 11452 26450 11508 26460
rect 11340 26350 11342 26402
rect 11394 26350 11396 26402
rect 11340 26338 11396 26350
rect 11676 26404 11732 26798
rect 11788 26852 12068 26908
rect 12124 26852 12180 28812
rect 12236 28644 12292 28654
rect 12236 27860 12292 28588
rect 12348 28642 12404 32956
rect 12460 32564 12516 33292
rect 12460 31666 12516 32508
rect 12460 31614 12462 31666
rect 12514 31614 12516 31666
rect 12460 31602 12516 31614
rect 12572 33122 12628 33134
rect 12572 33070 12574 33122
rect 12626 33070 12628 33122
rect 12572 31668 12628 33070
rect 12684 31778 12740 34188
rect 12796 34132 12852 34142
rect 12796 34038 12852 34076
rect 12908 33460 12964 34300
rect 13020 34132 13076 34170
rect 13020 34066 13076 34076
rect 13132 33684 13188 43148
rect 13356 41970 13412 41982
rect 13356 41918 13358 41970
rect 13410 41918 13412 41970
rect 13356 41748 13412 41918
rect 13356 41682 13412 41692
rect 13244 40180 13300 40190
rect 13244 38834 13300 40124
rect 13468 40068 13524 43596
rect 13916 43540 13972 43550
rect 13692 43428 13748 43438
rect 13692 42866 13748 43372
rect 13692 42814 13694 42866
rect 13746 42814 13748 42866
rect 13692 42802 13748 42814
rect 13804 43316 13860 43326
rect 13804 42754 13860 43260
rect 13804 42702 13806 42754
rect 13858 42702 13860 42754
rect 13580 42532 13636 42542
rect 13580 42530 13748 42532
rect 13580 42478 13582 42530
rect 13634 42478 13748 42530
rect 13580 42476 13748 42478
rect 13580 42466 13636 42476
rect 13580 41970 13636 41982
rect 13580 41918 13582 41970
rect 13634 41918 13636 41970
rect 13580 41860 13636 41918
rect 13580 41188 13636 41804
rect 13580 41122 13636 41132
rect 13580 40964 13636 40974
rect 13580 40870 13636 40908
rect 13692 40628 13748 42476
rect 13804 42420 13860 42702
rect 13804 42354 13860 42364
rect 13804 41972 13860 41982
rect 13916 41972 13972 43484
rect 14028 43092 14084 44044
rect 14140 44034 14196 44044
rect 14028 42868 14084 43036
rect 14028 42532 14084 42812
rect 14028 42466 14084 42476
rect 14140 43876 14196 43886
rect 13804 41970 13972 41972
rect 13804 41918 13806 41970
rect 13858 41918 13972 41970
rect 13804 41916 13972 41918
rect 14028 41972 14084 41982
rect 13804 41906 13860 41916
rect 14028 41878 14084 41916
rect 13804 41300 13860 41310
rect 13804 41186 13860 41244
rect 13804 41134 13806 41186
rect 13858 41134 13860 41186
rect 13804 41122 13860 41134
rect 13916 41188 13972 41198
rect 13916 40964 13972 41132
rect 13356 40012 13524 40068
rect 13580 40572 13748 40628
rect 13804 40908 13972 40964
rect 13356 39620 13412 40012
rect 13468 39844 13524 39854
rect 13468 39750 13524 39788
rect 13356 39564 13524 39620
rect 13244 38782 13246 38834
rect 13298 38782 13300 38834
rect 13244 38770 13300 38782
rect 13468 37940 13524 39564
rect 13580 38164 13636 40572
rect 13692 40404 13748 40414
rect 13692 40310 13748 40348
rect 13804 38834 13860 40908
rect 14028 40852 14084 40862
rect 14140 40852 14196 43820
rect 14252 43316 14308 45612
rect 14588 45602 14644 45612
rect 14924 45666 15092 45668
rect 14924 45614 15038 45666
rect 15090 45614 15092 45666
rect 14924 45612 15092 45614
rect 14476 44994 14532 45006
rect 14476 44942 14478 44994
rect 14530 44942 14532 44994
rect 14252 43250 14308 43260
rect 14364 44098 14420 44110
rect 14364 44046 14366 44098
rect 14418 44046 14420 44098
rect 14252 42756 14308 42766
rect 14364 42756 14420 44046
rect 14476 43652 14532 44942
rect 14700 44210 14756 44222
rect 14700 44158 14702 44210
rect 14754 44158 14756 44210
rect 14476 43586 14532 43596
rect 14588 44098 14644 44110
rect 14588 44046 14590 44098
rect 14642 44046 14644 44098
rect 14588 42868 14644 44046
rect 14700 43764 14756 44158
rect 14700 43698 14756 43708
rect 14588 42866 14868 42868
rect 14588 42814 14590 42866
rect 14642 42814 14868 42866
rect 14588 42812 14868 42814
rect 14588 42802 14644 42812
rect 14252 42754 14420 42756
rect 14252 42702 14254 42754
rect 14306 42702 14420 42754
rect 14252 42700 14420 42702
rect 14252 42690 14308 42700
rect 14364 42532 14420 42542
rect 14364 41970 14420 42476
rect 14364 41918 14366 41970
rect 14418 41918 14420 41970
rect 14364 41906 14420 41918
rect 14700 42532 14756 42542
rect 14700 42308 14756 42476
rect 14084 40796 14196 40852
rect 14252 41074 14308 41086
rect 14252 41022 14254 41074
rect 14306 41022 14308 41074
rect 14028 40786 14084 40796
rect 14252 40404 14308 41022
rect 14252 40338 14308 40348
rect 14252 39620 14308 39630
rect 14252 39526 14308 39564
rect 13804 38782 13806 38834
rect 13858 38782 13860 38834
rect 13804 38770 13860 38782
rect 13916 39506 13972 39518
rect 13916 39454 13918 39506
rect 13970 39454 13972 39506
rect 13916 38668 13972 39454
rect 13804 38612 13972 38668
rect 14028 39506 14084 39518
rect 14028 39454 14030 39506
rect 14082 39454 14084 39506
rect 14028 38668 14084 39454
rect 14700 39506 14756 42252
rect 14812 40964 14868 42812
rect 14924 42196 14980 45612
rect 15036 45602 15092 45612
rect 15708 45666 15876 45668
rect 15708 45614 15822 45666
rect 15874 45614 15876 45666
rect 15708 45612 15876 45614
rect 15484 44100 15540 44110
rect 15372 44098 15540 44100
rect 15372 44046 15486 44098
rect 15538 44046 15540 44098
rect 15372 44044 15540 44046
rect 15260 43426 15316 43438
rect 15260 43374 15262 43426
rect 15314 43374 15316 43426
rect 15260 42644 15316 43374
rect 15036 42532 15092 42542
rect 15036 42438 15092 42476
rect 14924 42140 15092 42196
rect 14924 41970 14980 41982
rect 14924 41918 14926 41970
rect 14978 41918 14980 41970
rect 14924 41636 14980 41918
rect 14924 41570 14980 41580
rect 14924 41412 14980 41422
rect 14924 41186 14980 41356
rect 15036 41300 15092 42140
rect 15260 42194 15316 42588
rect 15260 42142 15262 42194
rect 15314 42142 15316 42194
rect 15260 42130 15316 42142
rect 15372 41860 15428 44044
rect 15484 44034 15540 44044
rect 15596 43762 15652 43774
rect 15596 43710 15598 43762
rect 15650 43710 15652 43762
rect 15596 43652 15652 43710
rect 15596 43586 15652 43596
rect 15708 43540 15764 45612
rect 15820 45602 15876 45612
rect 17164 45666 17220 45678
rect 17164 45614 17166 45666
rect 17218 45614 17220 45666
rect 17164 45108 17220 45614
rect 18172 45668 18228 45678
rect 18172 45574 18228 45612
rect 18732 45666 18788 45678
rect 18732 45614 18734 45666
rect 18786 45614 18788 45666
rect 17612 45444 17668 45454
rect 17220 45052 17444 45108
rect 17164 45042 17220 45052
rect 16604 44996 16660 45006
rect 16380 44994 16660 44996
rect 16380 44942 16606 44994
rect 16658 44942 16660 44994
rect 16380 44940 16660 44942
rect 16380 44324 16436 44940
rect 16604 44930 16660 44940
rect 17388 44434 17444 45052
rect 17388 44382 17390 44434
rect 17442 44382 17444 44434
rect 17388 44370 17444 44382
rect 17612 45106 17668 45388
rect 17612 45054 17614 45106
rect 17666 45054 17668 45106
rect 16044 44268 16436 44324
rect 17612 44324 17668 45054
rect 18284 44996 18340 45006
rect 18284 44994 18452 44996
rect 18284 44942 18286 44994
rect 18338 44942 18452 44994
rect 18284 44940 18452 44942
rect 18284 44930 18340 44940
rect 17836 44324 17892 44334
rect 17612 44322 18004 44324
rect 17612 44270 17838 44322
rect 17890 44270 18004 44322
rect 17612 44268 18004 44270
rect 15708 43446 15764 43484
rect 15820 44098 15876 44110
rect 15820 44046 15822 44098
rect 15874 44046 15876 44098
rect 15708 42866 15764 42878
rect 15708 42814 15710 42866
rect 15762 42814 15764 42866
rect 15596 42196 15652 42206
rect 15596 42102 15652 42140
rect 15372 41804 15652 41860
rect 15036 41206 15092 41244
rect 15260 41748 15316 41758
rect 15260 41300 15316 41692
rect 15260 41234 15316 41244
rect 15372 41636 15428 41646
rect 14924 41134 14926 41186
rect 14978 41134 14980 41186
rect 14924 41122 14980 41134
rect 14812 40908 14980 40964
rect 14700 39454 14702 39506
rect 14754 39454 14756 39506
rect 14588 39396 14644 39406
rect 14588 39302 14644 39340
rect 14700 39172 14756 39454
rect 14700 39106 14756 39116
rect 14812 40402 14868 40414
rect 14812 40350 14814 40402
rect 14866 40350 14868 40402
rect 14476 39060 14532 39070
rect 14476 38948 14532 39004
rect 14812 38948 14868 40350
rect 14476 38892 14868 38948
rect 14924 39060 14980 40908
rect 15260 39396 15316 39406
rect 15260 39302 15316 39340
rect 14028 38612 14420 38668
rect 13804 38610 13860 38612
rect 13804 38558 13806 38610
rect 13858 38558 13860 38610
rect 13692 38164 13748 38174
rect 13580 38162 13748 38164
rect 13580 38110 13694 38162
rect 13746 38110 13748 38162
rect 13580 38108 13748 38110
rect 13692 38098 13748 38108
rect 13804 38052 13860 38558
rect 13804 37986 13860 37996
rect 13916 38164 13972 38174
rect 13580 37940 13636 37950
rect 13468 37938 13748 37940
rect 13468 37886 13582 37938
rect 13634 37886 13748 37938
rect 13468 37884 13748 37886
rect 13580 37874 13636 37884
rect 13244 37492 13300 37502
rect 13244 35700 13300 37436
rect 13580 37268 13636 37278
rect 13580 37174 13636 37212
rect 13692 36596 13748 37884
rect 13804 37828 13860 37838
rect 13916 37828 13972 38108
rect 14364 37940 14420 38612
rect 14364 37846 14420 37884
rect 13860 37772 13972 37828
rect 14028 37828 14084 37838
rect 13804 37734 13860 37772
rect 14028 37734 14084 37772
rect 14140 37378 14196 37390
rect 14140 37326 14142 37378
rect 14194 37326 14196 37378
rect 14140 36708 14196 37326
rect 14140 36642 14196 36652
rect 13692 36502 13748 36540
rect 13356 36372 13412 36382
rect 13356 35812 13412 36316
rect 13804 36260 13860 36270
rect 13804 36166 13860 36204
rect 13580 36036 13636 36046
rect 13468 35812 13524 35822
rect 13356 35810 13524 35812
rect 13356 35758 13470 35810
rect 13522 35758 13524 35810
rect 13356 35756 13524 35758
rect 13468 35746 13524 35756
rect 13244 35644 13412 35700
rect 13244 35364 13300 35374
rect 13244 34354 13300 35308
rect 13356 34804 13412 35644
rect 13580 35252 13636 35980
rect 13580 35186 13636 35196
rect 13692 35586 13748 35598
rect 13692 35534 13694 35586
rect 13746 35534 13748 35586
rect 13580 34804 13636 34814
rect 13356 34802 13636 34804
rect 13356 34750 13582 34802
rect 13634 34750 13636 34802
rect 13356 34748 13636 34750
rect 13580 34468 13636 34748
rect 13580 34402 13636 34412
rect 13244 34302 13246 34354
rect 13298 34302 13300 34354
rect 13244 34290 13300 34302
rect 13580 34242 13636 34254
rect 13580 34190 13582 34242
rect 13634 34190 13636 34242
rect 13468 33796 13524 33806
rect 13580 33796 13636 34190
rect 13524 33740 13636 33796
rect 13468 33730 13524 33740
rect 13132 33618 13188 33628
rect 12908 33404 13188 33460
rect 12908 33236 12964 33246
rect 12908 33142 12964 33180
rect 12796 33122 12852 33134
rect 12796 33070 12798 33122
rect 12850 33070 12852 33122
rect 12796 32676 12852 33070
rect 12796 32610 12852 32620
rect 12684 31726 12686 31778
rect 12738 31726 12740 31778
rect 12684 31714 12740 31726
rect 12796 31778 12852 31790
rect 12796 31726 12798 31778
rect 12850 31726 12852 31778
rect 12572 31602 12628 31612
rect 12796 31668 12852 31726
rect 12796 31602 12852 31612
rect 13020 31556 13076 31566
rect 13020 31106 13076 31500
rect 13020 31054 13022 31106
rect 13074 31054 13076 31106
rect 13020 31042 13076 31054
rect 12460 30548 12516 30558
rect 12460 30100 12516 30492
rect 12572 30436 12628 30446
rect 12572 30342 12628 30380
rect 12908 30324 12964 30334
rect 12908 30230 12964 30268
rect 12460 30044 12740 30100
rect 12572 29876 12628 29886
rect 12460 29426 12516 29438
rect 12460 29374 12462 29426
rect 12514 29374 12516 29426
rect 12460 28754 12516 29374
rect 12460 28702 12462 28754
rect 12514 28702 12516 28754
rect 12460 28690 12516 28702
rect 12348 28590 12350 28642
rect 12402 28590 12404 28642
rect 12348 28578 12404 28590
rect 12572 28530 12628 29820
rect 12684 28980 12740 30044
rect 12684 28644 12740 28924
rect 12796 29988 12852 29998
rect 12796 28756 12852 29932
rect 13020 29540 13076 29550
rect 13020 29446 13076 29484
rect 12908 28756 12964 28766
rect 12796 28700 12908 28756
rect 12908 28690 12964 28700
rect 13020 28644 13076 28654
rect 12684 28588 12852 28644
rect 12572 28478 12574 28530
rect 12626 28478 12628 28530
rect 12572 28466 12628 28478
rect 12684 28084 12740 28094
rect 12460 27860 12516 27870
rect 12236 27804 12460 27860
rect 12460 27766 12516 27804
rect 12572 27524 12628 27534
rect 12236 27300 12292 27310
rect 12236 27206 12292 27244
rect 11788 26514 11844 26852
rect 11788 26462 11790 26514
rect 11842 26462 11844 26514
rect 11788 26450 11844 26462
rect 11676 26338 11732 26348
rect 11564 26290 11620 26302
rect 11564 26238 11566 26290
rect 11618 26238 11620 26290
rect 11116 25106 11172 25116
rect 11340 26180 11396 26190
rect 11340 25396 11396 26124
rect 11340 24948 11396 25340
rect 11116 24892 11396 24948
rect 11116 21476 11172 24892
rect 11340 24834 11396 24892
rect 11340 24782 11342 24834
rect 11394 24782 11396 24834
rect 11340 24770 11396 24782
rect 11452 25172 11508 25182
rect 11228 24724 11284 24734
rect 11228 24050 11284 24668
rect 11452 24722 11508 25116
rect 11452 24670 11454 24722
rect 11506 24670 11508 24722
rect 11340 24500 11396 24510
rect 11452 24500 11508 24670
rect 11564 24724 11620 26238
rect 11900 26290 11956 26302
rect 11900 26238 11902 26290
rect 11954 26238 11956 26290
rect 11788 26178 11844 26190
rect 11788 26126 11790 26178
rect 11842 26126 11844 26178
rect 11564 24658 11620 24668
rect 11676 25060 11732 25070
rect 11676 24610 11732 25004
rect 11676 24558 11678 24610
rect 11730 24558 11732 24610
rect 11676 24546 11732 24558
rect 11396 24444 11508 24500
rect 11340 24434 11396 24444
rect 11228 23998 11230 24050
rect 11282 23998 11284 24050
rect 11228 23986 11284 23998
rect 11340 24276 11396 24286
rect 11340 22708 11396 24220
rect 11788 24052 11844 26126
rect 11900 26180 11956 26238
rect 11900 26114 11956 26124
rect 12012 25506 12068 25518
rect 12012 25454 12014 25506
rect 12066 25454 12068 25506
rect 11900 25394 11956 25406
rect 11900 25342 11902 25394
rect 11954 25342 11956 25394
rect 11900 24836 11956 25342
rect 11900 24770 11956 24780
rect 12012 24724 12068 25454
rect 12012 24658 12068 24668
rect 11788 23986 11844 23996
rect 11900 23940 11956 23950
rect 11676 23716 11732 23726
rect 11340 22482 11396 22652
rect 11340 22430 11342 22482
rect 11394 22430 11396 22482
rect 11340 22418 11396 22430
rect 11452 23660 11676 23716
rect 11452 23154 11508 23660
rect 11676 23622 11732 23660
rect 11452 23102 11454 23154
rect 11506 23102 11508 23154
rect 11452 21700 11508 23102
rect 11564 23492 11620 23502
rect 11564 21812 11620 23436
rect 11788 23380 11844 23390
rect 11788 23154 11844 23324
rect 11788 23102 11790 23154
rect 11842 23102 11844 23154
rect 11788 23090 11844 23102
rect 11900 22482 11956 23884
rect 11900 22430 11902 22482
rect 11954 22430 11956 22482
rect 11900 22418 11956 22430
rect 12012 22594 12068 22606
rect 12012 22542 12014 22594
rect 12066 22542 12068 22594
rect 11564 21756 11732 21812
rect 11452 21634 11508 21644
rect 11340 21586 11396 21598
rect 11340 21534 11342 21586
rect 11394 21534 11396 21586
rect 11228 21476 11284 21486
rect 11116 21420 11228 21476
rect 11228 21410 11284 21420
rect 11004 20862 11006 20914
rect 11058 20862 11060 20914
rect 10668 20638 10670 20690
rect 10722 20638 10724 20690
rect 10556 20132 10612 20142
rect 10108 20076 10388 20132
rect 10108 19908 10164 19918
rect 10108 19814 10164 19852
rect 10220 19796 10276 19806
rect 10108 19348 10164 19358
rect 10220 19348 10276 19740
rect 10108 19346 10276 19348
rect 10108 19294 10110 19346
rect 10162 19294 10276 19346
rect 10108 19292 10276 19294
rect 10108 19282 10164 19292
rect 10220 19124 10276 19134
rect 10220 18674 10276 19068
rect 10220 18622 10222 18674
rect 10274 18622 10276 18674
rect 10220 18610 10276 18622
rect 10332 18340 10388 20076
rect 10332 18226 10388 18284
rect 10332 18174 10334 18226
rect 10386 18174 10388 18226
rect 10332 18162 10388 18174
rect 10444 19234 10500 19246
rect 10444 19182 10446 19234
rect 10498 19182 10500 19234
rect 10444 19124 10500 19182
rect 9884 17106 10052 17108
rect 9884 17054 9886 17106
rect 9938 17054 10052 17106
rect 9884 17052 10052 17054
rect 10108 17442 10164 17454
rect 10108 17390 10110 17442
rect 10162 17390 10164 17442
rect 9884 17042 9940 17052
rect 9772 16706 9828 16716
rect 9548 16156 10052 16212
rect 9548 15428 9604 15438
rect 9548 15334 9604 15372
rect 9100 15092 9268 15148
rect 9324 15092 9492 15148
rect 9660 15202 9716 15214
rect 9660 15150 9662 15202
rect 9714 15150 9716 15202
rect 8652 14532 8708 14542
rect 8652 13634 8708 14476
rect 8652 13582 8654 13634
rect 8706 13582 8708 13634
rect 8652 13570 8708 13582
rect 8876 12962 8932 12974
rect 8876 12910 8878 12962
rect 8930 12910 8932 12962
rect 8876 12740 8932 12910
rect 8876 12674 8932 12684
rect 8540 12114 8596 12124
rect 8876 12516 8932 12526
rect 7980 11900 8372 11956
rect 6412 11454 6414 11506
rect 6466 11454 6468 11506
rect 5964 11284 6020 11294
rect 5964 11190 6020 11228
rect 6300 10724 6356 10734
rect 6188 10722 6356 10724
rect 6188 10670 6302 10722
rect 6354 10670 6356 10722
rect 6188 10668 6356 10670
rect 6188 10052 6244 10668
rect 6300 10658 6356 10668
rect 6412 10052 6468 11454
rect 7756 11732 7812 11742
rect 7756 11394 7812 11676
rect 7756 11342 7758 11394
rect 7810 11342 7812 11394
rect 7756 11330 7812 11342
rect 7980 11394 8036 11900
rect 7980 11342 7982 11394
rect 8034 11342 8036 11394
rect 7980 11330 8036 11342
rect 8316 11508 8372 11900
rect 6188 9986 6244 9996
rect 6300 9996 6468 10052
rect 6524 11284 6580 11294
rect 5404 9874 5460 9884
rect 6076 9940 6132 9950
rect 4620 9826 5124 9828
rect 4620 9774 4622 9826
rect 4674 9774 5070 9826
rect 5122 9774 5124 9826
rect 4620 9772 5124 9774
rect 4620 9762 4676 9772
rect 4956 9268 5012 9306
rect 4956 9202 5012 9212
rect 4620 9156 4676 9166
rect 4620 9062 4676 9100
rect 4172 8990 4174 9042
rect 4226 8990 4228 9042
rect 4172 8978 4228 8990
rect 4396 9042 4452 9054
rect 4396 8990 4398 9042
rect 4450 8990 4452 9042
rect 4396 8820 4452 8990
rect 4956 9044 5012 9054
rect 4956 8950 5012 8988
rect 5068 8820 5124 9772
rect 5180 9772 5348 9828
rect 6076 9828 6132 9884
rect 6188 9828 6244 9838
rect 6076 9826 6244 9828
rect 6076 9774 6190 9826
rect 6242 9774 6244 9826
rect 6076 9772 6244 9774
rect 5180 9156 5236 9772
rect 6188 9762 6244 9772
rect 5516 9604 5572 9614
rect 5180 9090 5236 9100
rect 5292 9548 5516 9604
rect 5292 9042 5348 9548
rect 5516 9538 5572 9548
rect 5740 9156 5796 9166
rect 5740 9062 5796 9100
rect 5292 8990 5294 9042
rect 5346 8990 5348 9042
rect 5292 8978 5348 8990
rect 5516 9042 5572 9054
rect 6188 9044 6244 9054
rect 6300 9044 6356 9996
rect 6412 9828 6468 9838
rect 6524 9828 6580 11228
rect 6412 9826 6580 9828
rect 6412 9774 6414 9826
rect 6466 9774 6580 9826
rect 6412 9772 6580 9774
rect 6636 11172 6692 11182
rect 6636 10722 6692 11116
rect 7868 11172 7924 11182
rect 7868 11078 7924 11116
rect 8204 11172 8260 11182
rect 8204 11078 8260 11116
rect 8204 10836 8260 10846
rect 8316 10836 8372 11452
rect 8764 11732 8820 11742
rect 8764 11394 8820 11676
rect 8764 11342 8766 11394
rect 8818 11342 8820 11394
rect 8764 11330 8820 11342
rect 8428 10836 8484 10846
rect 8316 10834 8484 10836
rect 8316 10782 8430 10834
rect 8482 10782 8484 10834
rect 8316 10780 8484 10782
rect 8204 10742 8260 10780
rect 8428 10770 8484 10780
rect 6636 10670 6638 10722
rect 6690 10670 6692 10722
rect 6636 9826 6692 10670
rect 8876 10610 8932 12460
rect 8988 12292 9044 12302
rect 8988 12066 9044 12236
rect 8988 12014 8990 12066
rect 9042 12014 9044 12066
rect 8988 12002 9044 12014
rect 8988 11284 9044 11294
rect 9100 11284 9156 15092
rect 9212 13636 9268 13646
rect 9212 12962 9268 13580
rect 9212 12910 9214 12962
rect 9266 12910 9268 12962
rect 9212 12898 9268 12910
rect 9324 11620 9380 15092
rect 9660 14532 9716 15150
rect 9660 14466 9716 14476
rect 9660 14084 9716 14094
rect 9660 13970 9716 14028
rect 9660 13918 9662 13970
rect 9714 13918 9716 13970
rect 9436 13524 9492 13534
rect 9436 12850 9492 13468
rect 9436 12798 9438 12850
rect 9490 12798 9492 12850
rect 9436 12786 9492 12798
rect 9548 12738 9604 12750
rect 9548 12686 9550 12738
rect 9602 12686 9604 12738
rect 9548 12628 9604 12686
rect 9436 12572 9604 12628
rect 9436 11954 9492 12572
rect 9660 12292 9716 13918
rect 9772 12628 9828 16156
rect 9996 16098 10052 16156
rect 9996 16046 9998 16098
rect 10050 16046 10052 16098
rect 9996 16034 10052 16046
rect 9884 15988 9940 15998
rect 9884 15894 9940 15932
rect 9884 15540 9940 15550
rect 9884 13860 9940 15484
rect 9996 14644 10052 14654
rect 9996 14550 10052 14588
rect 9884 12964 9940 13804
rect 9996 13746 10052 13758
rect 9996 13694 9998 13746
rect 10050 13694 10052 13746
rect 9996 13188 10052 13694
rect 10108 13748 10164 17390
rect 10332 16882 10388 16894
rect 10332 16830 10334 16882
rect 10386 16830 10388 16882
rect 10332 15988 10388 16830
rect 10332 15922 10388 15932
rect 10220 15204 10276 15242
rect 10332 15204 10388 15214
rect 10220 15202 10332 15204
rect 10220 15150 10222 15202
rect 10274 15150 10332 15202
rect 10220 15148 10332 15150
rect 10220 14084 10276 15148
rect 10332 15138 10388 15148
rect 10444 15148 10500 19068
rect 10556 18900 10612 20076
rect 10668 19236 10724 20638
rect 10892 20580 10948 20590
rect 10892 20486 10948 20524
rect 10892 20356 10948 20366
rect 10780 20300 10892 20356
rect 10780 19346 10836 20300
rect 10892 20290 10948 20300
rect 11004 19796 11060 20862
rect 11340 20916 11396 21534
rect 11340 20822 11396 20860
rect 11564 20804 11620 20842
rect 11564 20738 11620 20748
rect 11564 20578 11620 20590
rect 11564 20526 11566 20578
rect 11618 20526 11620 20578
rect 11116 20132 11172 20142
rect 11116 20018 11172 20076
rect 11340 20020 11396 20030
rect 11116 19966 11118 20018
rect 11170 19966 11172 20018
rect 11116 19954 11172 19966
rect 11228 20018 11396 20020
rect 11228 19966 11342 20018
rect 11394 19966 11396 20018
rect 11228 19964 11396 19966
rect 11004 19730 11060 19740
rect 11228 19460 11284 19964
rect 11340 19954 11396 19964
rect 11564 20020 11620 20526
rect 11564 19954 11620 19964
rect 10780 19294 10782 19346
rect 10834 19294 10836 19346
rect 10780 19282 10836 19294
rect 11004 19458 11284 19460
rect 11004 19406 11230 19458
rect 11282 19406 11284 19458
rect 11004 19404 11284 19406
rect 10668 19170 10724 19180
rect 10556 18844 10724 18900
rect 10556 18676 10612 18686
rect 10556 16212 10612 18620
rect 10668 16884 10724 18844
rect 10780 18562 10836 18574
rect 10780 18510 10782 18562
rect 10834 18510 10836 18562
rect 10780 18116 10836 18510
rect 10780 18050 10836 18060
rect 10892 18228 10948 18238
rect 10668 16818 10724 16828
rect 10556 16146 10612 16156
rect 10780 16772 10836 16782
rect 10780 15314 10836 16716
rect 10780 15262 10782 15314
rect 10834 15262 10836 15314
rect 10780 15250 10836 15262
rect 10444 15092 10836 15148
rect 10780 14644 10836 15092
rect 10780 14550 10836 14588
rect 10444 14530 10500 14542
rect 10444 14478 10446 14530
rect 10498 14478 10500 14530
rect 10220 14018 10276 14028
rect 10332 14418 10388 14430
rect 10332 14366 10334 14418
rect 10386 14366 10388 14418
rect 10220 13748 10276 13758
rect 10108 13746 10276 13748
rect 10108 13694 10222 13746
rect 10274 13694 10276 13746
rect 10108 13692 10276 13694
rect 10332 13748 10388 14366
rect 10444 13972 10500 14478
rect 10444 13906 10500 13916
rect 10668 14532 10724 14542
rect 10444 13748 10500 13758
rect 10332 13746 10500 13748
rect 10332 13694 10446 13746
rect 10498 13694 10500 13746
rect 10332 13692 10500 13694
rect 10220 13524 10276 13692
rect 10444 13636 10500 13692
rect 10444 13570 10500 13580
rect 10220 13458 10276 13468
rect 10668 13412 10724 14476
rect 10780 13972 10836 13982
rect 10892 13972 10948 18172
rect 11004 16100 11060 19404
rect 11228 19394 11284 19404
rect 11116 19124 11172 19134
rect 11340 19124 11396 19134
rect 11172 19122 11396 19124
rect 11172 19070 11342 19122
rect 11394 19070 11396 19122
rect 11172 19068 11396 19070
rect 11116 19058 11172 19068
rect 11340 19058 11396 19068
rect 11116 18564 11172 18574
rect 11452 18564 11508 18574
rect 11116 18562 11508 18564
rect 11116 18510 11118 18562
rect 11170 18510 11454 18562
rect 11506 18510 11508 18562
rect 11116 18508 11508 18510
rect 11116 17780 11172 18508
rect 11452 18498 11508 18508
rect 11564 18340 11620 18350
rect 11564 18246 11620 18284
rect 11676 18116 11732 21756
rect 11788 21476 11844 21486
rect 11788 21382 11844 21420
rect 11788 20802 11844 20814
rect 11788 20750 11790 20802
rect 11842 20750 11844 20802
rect 11788 20580 11844 20750
rect 11788 19906 11844 20524
rect 11788 19854 11790 19906
rect 11842 19854 11844 19906
rect 11788 19842 11844 19854
rect 11900 20018 11956 20030
rect 11900 19966 11902 20018
rect 11954 19966 11956 20018
rect 11788 19458 11844 19470
rect 11788 19406 11790 19458
rect 11842 19406 11844 19458
rect 11788 19346 11844 19406
rect 11788 19294 11790 19346
rect 11842 19294 11844 19346
rect 11788 19282 11844 19294
rect 11900 18676 11956 19966
rect 11564 18060 11732 18116
rect 11788 18620 11956 18676
rect 11788 18116 11844 18620
rect 11900 18452 11956 18462
rect 11900 18358 11956 18396
rect 11116 17714 11172 17724
rect 11452 17780 11508 17790
rect 11452 17666 11508 17724
rect 11452 17614 11454 17666
rect 11506 17614 11508 17666
rect 11452 17602 11508 17614
rect 11564 17442 11620 18060
rect 11788 18050 11844 18060
rect 11564 17390 11566 17442
rect 11618 17390 11620 17442
rect 11564 17378 11620 17390
rect 11676 17666 11732 17678
rect 11676 17614 11678 17666
rect 11730 17614 11732 17666
rect 11340 17220 11396 17230
rect 11228 17164 11340 17220
rect 11396 17164 11508 17220
rect 11228 16994 11284 17164
rect 11340 17154 11396 17164
rect 11228 16942 11230 16994
rect 11282 16942 11284 16994
rect 11228 16930 11284 16942
rect 11004 16034 11060 16044
rect 11004 15540 11060 15550
rect 11004 15446 11060 15484
rect 11340 15428 11396 15438
rect 10780 13970 10948 13972
rect 10780 13918 10782 13970
rect 10834 13918 10948 13970
rect 10780 13916 10948 13918
rect 11116 15316 11172 15326
rect 10780 13906 10836 13916
rect 10332 13356 10724 13412
rect 9996 13132 10276 13188
rect 9996 12964 10052 12974
rect 9884 12962 10052 12964
rect 9884 12910 9998 12962
rect 10050 12910 10052 12962
rect 9884 12908 10052 12910
rect 9996 12898 10052 12908
rect 10108 12962 10164 12974
rect 10108 12910 10110 12962
rect 10162 12910 10164 12962
rect 10108 12740 10164 12910
rect 9996 12684 10164 12740
rect 9772 12572 9940 12628
rect 9436 11902 9438 11954
rect 9490 11902 9492 11954
rect 9436 11890 9492 11902
rect 9548 12290 9716 12292
rect 9548 12238 9662 12290
rect 9714 12238 9716 12290
rect 9548 12236 9716 12238
rect 9324 11506 9380 11564
rect 9324 11454 9326 11506
rect 9378 11454 9380 11506
rect 9324 11442 9380 11454
rect 8988 11282 9156 11284
rect 8988 11230 8990 11282
rect 9042 11230 9156 11282
rect 8988 11228 9156 11230
rect 8988 10836 9044 11228
rect 8988 10770 9044 10780
rect 9436 11170 9492 11182
rect 9436 11118 9438 11170
rect 9490 11118 9492 11170
rect 8876 10558 8878 10610
rect 8930 10558 8932 10610
rect 7532 10498 7588 10510
rect 7532 10446 7534 10498
rect 7586 10446 7588 10498
rect 6636 9774 6638 9826
rect 6690 9774 6692 9826
rect 6412 9762 6468 9772
rect 6636 9762 6692 9774
rect 6972 10052 7028 10062
rect 6972 9826 7028 9996
rect 7532 9940 7588 10446
rect 8316 10498 8372 10510
rect 8316 10446 8318 10498
rect 8370 10446 8372 10498
rect 8316 10052 8372 10446
rect 8876 10500 8932 10558
rect 9436 10610 9492 11118
rect 9436 10558 9438 10610
rect 9490 10558 9492 10610
rect 9436 10546 9492 10558
rect 8876 10434 8932 10444
rect 9548 10276 9604 12236
rect 9660 12226 9716 12236
rect 9772 11954 9828 11966
rect 9772 11902 9774 11954
rect 9826 11902 9828 11954
rect 9772 11394 9828 11902
rect 9884 11732 9940 12572
rect 9996 12516 10052 12684
rect 10220 12516 10276 13132
rect 10332 12962 10388 13356
rect 11116 13188 11172 15260
rect 11340 15314 11396 15372
rect 11340 15262 11342 15314
rect 11394 15262 11396 15314
rect 11340 15250 11396 15262
rect 11452 13970 11508 17164
rect 11676 16100 11732 17614
rect 11900 17332 11956 17342
rect 11900 16322 11956 17276
rect 12012 16660 12068 22542
rect 12124 22036 12180 26796
rect 12348 26964 12404 26974
rect 12348 26402 12404 26908
rect 12572 26962 12628 27468
rect 12572 26910 12574 26962
rect 12626 26910 12628 26962
rect 12572 26898 12628 26910
rect 12348 26350 12350 26402
rect 12402 26350 12404 26402
rect 12348 26338 12404 26350
rect 12460 26404 12516 26414
rect 12460 25618 12516 26348
rect 12572 26292 12628 26302
rect 12684 26292 12740 28028
rect 12572 26290 12740 26292
rect 12572 26238 12574 26290
rect 12626 26238 12740 26290
rect 12572 26236 12740 26238
rect 12572 26226 12628 26236
rect 12460 25566 12462 25618
rect 12514 25566 12516 25618
rect 12460 25554 12516 25566
rect 12684 25508 12740 25518
rect 12572 25452 12684 25508
rect 12460 25396 12516 25406
rect 12460 25302 12516 25340
rect 12236 24834 12292 24846
rect 12236 24782 12238 24834
rect 12290 24782 12292 24834
rect 12236 23828 12292 24782
rect 12460 24722 12516 24734
rect 12460 24670 12462 24722
rect 12514 24670 12516 24722
rect 12236 23154 12292 23772
rect 12236 23102 12238 23154
rect 12290 23102 12292 23154
rect 12236 22594 12292 23102
rect 12236 22542 12238 22594
rect 12290 22542 12292 22594
rect 12236 22530 12292 22542
rect 12348 24500 12404 24510
rect 12348 22482 12404 24444
rect 12460 23940 12516 24670
rect 12572 24050 12628 25452
rect 12684 25442 12740 25452
rect 12796 25506 12852 28588
rect 12908 27636 12964 27646
rect 12908 27074 12964 27580
rect 12908 27022 12910 27074
rect 12962 27022 12964 27074
rect 12908 27010 12964 27022
rect 12908 26516 12964 26526
rect 13020 26516 13076 28588
rect 12908 26514 13076 26516
rect 12908 26462 12910 26514
rect 12962 26462 13076 26514
rect 12908 26460 13076 26462
rect 12908 26450 12964 26460
rect 13132 26292 13188 33404
rect 13692 33348 13748 35534
rect 14252 35028 14308 35038
rect 14252 34934 14308 34972
rect 13580 33292 13748 33348
rect 13804 34914 13860 34926
rect 13804 34862 13806 34914
rect 13858 34862 13860 34914
rect 13804 33572 13860 34862
rect 14028 34916 14084 34926
rect 14028 34822 14084 34860
rect 14476 34916 14532 38892
rect 14924 38834 14980 39004
rect 14924 38782 14926 38834
rect 14978 38782 14980 38834
rect 14924 38770 14980 38782
rect 15148 39284 15204 39294
rect 14700 38050 14756 38062
rect 14700 37998 14702 38050
rect 14754 37998 14756 38050
rect 14700 37380 14756 37998
rect 15036 38050 15092 38062
rect 15036 37998 15038 38050
rect 15090 37998 15092 38050
rect 15036 37604 15092 37998
rect 15036 37538 15092 37548
rect 15148 37492 15204 39228
rect 15260 39172 15316 39182
rect 15260 38388 15316 39116
rect 15372 38612 15428 41580
rect 15596 41188 15652 41804
rect 15708 41412 15764 42814
rect 15820 41972 15876 44046
rect 16044 43764 16100 44268
rect 16380 44210 16436 44268
rect 17836 44258 17892 44268
rect 16380 44158 16382 44210
rect 16434 44158 16436 44210
rect 16380 44146 16436 44158
rect 16492 44212 16548 44222
rect 16492 44210 16660 44212
rect 16492 44158 16494 44210
rect 16546 44158 16660 44210
rect 16492 44156 16660 44158
rect 16492 44146 16548 44156
rect 16156 44098 16212 44110
rect 16156 44046 16158 44098
rect 16210 44046 16212 44098
rect 16156 43988 16212 44046
rect 16156 43932 16548 43988
rect 16044 43708 16212 43764
rect 15932 43316 15988 43326
rect 15932 43314 16100 43316
rect 15932 43262 15934 43314
rect 15986 43262 16100 43314
rect 15932 43260 16100 43262
rect 15932 43250 15988 43260
rect 15932 41972 15988 41982
rect 15820 41970 15988 41972
rect 15820 41918 15934 41970
rect 15986 41918 15988 41970
rect 15820 41916 15988 41918
rect 15820 41524 15876 41916
rect 15932 41906 15988 41916
rect 15820 41458 15876 41468
rect 15708 41346 15764 41356
rect 15708 41188 15764 41198
rect 15596 41186 15764 41188
rect 15596 41134 15710 41186
rect 15762 41134 15764 41186
rect 15596 41132 15764 41134
rect 15596 40964 15652 41132
rect 15708 41122 15764 41132
rect 15932 41076 15988 41086
rect 15932 40982 15988 41020
rect 15484 40628 15540 40638
rect 15484 40514 15540 40572
rect 15484 40462 15486 40514
rect 15538 40462 15540 40514
rect 15484 40450 15540 40462
rect 15596 39396 15652 40908
rect 16044 40740 16100 43260
rect 16156 43092 16212 43708
rect 16492 43650 16548 43932
rect 16492 43598 16494 43650
rect 16546 43598 16548 43650
rect 16492 43586 16548 43598
rect 16268 43538 16324 43550
rect 16268 43486 16270 43538
rect 16322 43486 16324 43538
rect 16268 43316 16324 43486
rect 16268 43250 16324 43260
rect 16156 43036 16324 43092
rect 16044 40674 16100 40684
rect 16156 41860 16212 41870
rect 15932 40626 15988 40638
rect 15932 40574 15934 40626
rect 15986 40574 15988 40626
rect 15932 39732 15988 40574
rect 16156 40628 16212 41804
rect 16268 41636 16324 43036
rect 16604 42420 16660 44156
rect 17052 44100 17108 44110
rect 17052 44006 17108 44044
rect 17500 43428 17556 43438
rect 16492 42364 16660 42420
rect 17164 43426 17556 43428
rect 17164 43374 17502 43426
rect 17554 43374 17556 43426
rect 17164 43372 17556 43374
rect 16492 41860 16548 42364
rect 16492 41794 16548 41804
rect 16604 42196 16660 42206
rect 16604 42082 16660 42140
rect 16604 42030 16606 42082
rect 16658 42030 16660 42082
rect 16268 41570 16324 41580
rect 16156 40562 16212 40572
rect 16268 41410 16324 41422
rect 16268 41358 16270 41410
rect 16322 41358 16324 41410
rect 16268 41300 16324 41358
rect 16604 41412 16660 42030
rect 16716 41748 16772 41758
rect 16716 41746 17108 41748
rect 16716 41694 16718 41746
rect 16770 41694 17108 41746
rect 16716 41692 17108 41694
rect 16716 41682 16772 41692
rect 16604 41346 16660 41356
rect 16268 40516 16324 41244
rect 16268 40450 16324 40460
rect 16380 41186 16436 41198
rect 17052 41188 17108 41692
rect 16380 41134 16382 41186
rect 16434 41134 16436 41186
rect 16044 40292 16100 40302
rect 16044 40198 16100 40236
rect 16268 40180 16324 40190
rect 16268 40086 16324 40124
rect 16380 39844 16436 41134
rect 16940 41186 17108 41188
rect 16940 41134 17054 41186
rect 17106 41134 17108 41186
rect 16940 41132 17108 41134
rect 16828 41076 16884 41086
rect 16492 41074 16884 41076
rect 16492 41022 16830 41074
rect 16882 41022 16884 41074
rect 16492 41020 16884 41022
rect 16492 40962 16548 41020
rect 16828 41010 16884 41020
rect 16492 40910 16494 40962
rect 16546 40910 16548 40962
rect 16492 40898 16548 40910
rect 16828 40516 16884 40526
rect 16940 40516 16996 41132
rect 17052 41122 17108 41132
rect 16828 40514 16996 40516
rect 16828 40462 16830 40514
rect 16882 40462 16996 40514
rect 16828 40460 16996 40462
rect 16828 40450 16884 40460
rect 16716 40404 16772 40414
rect 16492 39844 16548 39854
rect 16380 39842 16548 39844
rect 16380 39790 16494 39842
rect 16546 39790 16548 39842
rect 16380 39788 16548 39790
rect 16492 39778 16548 39788
rect 16044 39732 16100 39742
rect 15932 39676 16044 39732
rect 15596 39330 15652 39340
rect 15820 39620 15876 39630
rect 15820 39172 15876 39564
rect 16044 39618 16100 39676
rect 16044 39566 16046 39618
rect 16098 39566 16100 39618
rect 16044 39554 16100 39566
rect 15820 39106 15876 39116
rect 15932 39506 15988 39518
rect 15932 39454 15934 39506
rect 15986 39454 15988 39506
rect 15708 39060 15764 39070
rect 15484 38834 15540 38846
rect 15484 38782 15486 38834
rect 15538 38782 15540 38834
rect 15484 38724 15540 38782
rect 15484 38658 15540 38668
rect 15596 38722 15652 38734
rect 15596 38670 15598 38722
rect 15650 38670 15652 38722
rect 15372 38546 15428 38556
rect 15260 38332 15540 38388
rect 15148 37426 15204 37436
rect 15372 38052 15428 38062
rect 14812 37380 14868 37390
rect 14700 37324 14812 37380
rect 14812 37314 14868 37324
rect 14588 36596 14644 36606
rect 14588 36260 14644 36540
rect 14588 35476 14644 36204
rect 14924 36372 14980 36382
rect 14700 35924 14756 35934
rect 14700 35810 14756 35868
rect 14700 35758 14702 35810
rect 14754 35758 14756 35810
rect 14700 35746 14756 35758
rect 14588 35410 14644 35420
rect 14924 35308 14980 36316
rect 15036 36260 15092 36270
rect 15036 35698 15092 36204
rect 15036 35646 15038 35698
rect 15090 35646 15092 35698
rect 15036 35634 15092 35646
rect 14924 35252 15092 35308
rect 14924 35028 14980 35038
rect 14924 34934 14980 34972
rect 14476 34850 14532 34860
rect 15036 34916 15092 35252
rect 15036 34850 15092 34860
rect 15260 35028 15316 35038
rect 15260 34914 15316 34972
rect 15260 34862 15262 34914
rect 15314 34862 15316 34914
rect 15260 34850 15316 34862
rect 13804 33348 13860 33516
rect 14140 34804 14196 34814
rect 14028 33348 14084 33358
rect 13804 33346 14084 33348
rect 13804 33294 14030 33346
rect 14082 33294 14084 33346
rect 13804 33292 14084 33294
rect 13244 33236 13300 33246
rect 13244 32562 13300 33180
rect 13244 32510 13246 32562
rect 13298 32510 13300 32562
rect 13244 32498 13300 32510
rect 13580 32004 13636 33292
rect 14028 33282 14084 33292
rect 14140 33234 14196 34748
rect 15148 34802 15204 34814
rect 15148 34750 15150 34802
rect 15202 34750 15204 34802
rect 14588 34692 14644 34702
rect 14476 34636 14588 34692
rect 14140 33182 14142 33234
rect 14194 33182 14196 33234
rect 14140 33170 14196 33182
rect 14364 34468 14420 34478
rect 13692 33122 13748 33134
rect 13692 33070 13694 33122
rect 13746 33070 13748 33122
rect 13692 33012 13748 33070
rect 13804 33012 13860 33022
rect 13692 32956 13804 33012
rect 13580 31938 13636 31948
rect 13804 31444 13860 32956
rect 13916 32562 13972 32574
rect 13916 32510 13918 32562
rect 13970 32510 13972 32562
rect 13916 32340 13972 32510
rect 13916 32274 13972 32284
rect 13916 31668 13972 31678
rect 13916 31666 14196 31668
rect 13916 31614 13918 31666
rect 13970 31614 14196 31666
rect 13916 31612 14196 31614
rect 13916 31602 13972 31612
rect 13804 31388 13972 31444
rect 13244 31332 13300 31342
rect 13244 27524 13300 31276
rect 13356 30996 13412 31006
rect 13356 30436 13412 30940
rect 13916 30884 13972 31388
rect 14028 31220 14084 31230
rect 14028 31106 14084 31164
rect 14028 31054 14030 31106
rect 14082 31054 14084 31106
rect 14028 31042 14084 31054
rect 13916 30828 14084 30884
rect 13692 30772 13748 30782
rect 13692 30678 13748 30716
rect 13804 30770 13860 30782
rect 13804 30718 13806 30770
rect 13858 30718 13860 30770
rect 13356 30380 13524 30436
rect 13468 30210 13524 30380
rect 13580 30324 13636 30334
rect 13804 30324 13860 30718
rect 13580 30322 13860 30324
rect 13580 30270 13582 30322
rect 13634 30270 13860 30322
rect 13580 30268 13860 30270
rect 13580 30258 13636 30268
rect 13468 30158 13470 30210
rect 13522 30158 13524 30210
rect 13468 30146 13524 30158
rect 13916 30210 13972 30222
rect 13916 30158 13918 30210
rect 13970 30158 13972 30210
rect 13804 30098 13860 30110
rect 13804 30046 13806 30098
rect 13858 30046 13860 30098
rect 13804 29876 13860 30046
rect 13916 29988 13972 30158
rect 13916 29922 13972 29932
rect 13804 29316 13860 29820
rect 14028 29764 14084 30828
rect 13804 29250 13860 29260
rect 13916 29708 14084 29764
rect 13468 28756 13524 28766
rect 13244 27458 13300 27468
rect 13356 28420 13412 28430
rect 12796 25454 12798 25506
rect 12850 25454 12852 25506
rect 12572 23998 12574 24050
rect 12626 23998 12628 24050
rect 12572 23986 12628 23998
rect 12684 25284 12740 25294
rect 12460 23874 12516 23884
rect 12572 23380 12628 23390
rect 12572 23286 12628 23324
rect 12348 22430 12350 22482
rect 12402 22430 12404 22482
rect 12348 22418 12404 22430
rect 12124 21970 12180 21980
rect 12124 21700 12180 21710
rect 12124 20802 12180 21644
rect 12236 21588 12292 21598
rect 12236 21494 12292 21532
rect 12684 20916 12740 25228
rect 12796 24162 12852 25454
rect 12796 24110 12798 24162
rect 12850 24110 12852 24162
rect 12796 24098 12852 24110
rect 12908 26236 13188 26292
rect 13356 27188 13412 28364
rect 12796 22708 12852 22718
rect 12796 22482 12852 22652
rect 12796 22430 12798 22482
rect 12850 22430 12852 22482
rect 12796 21140 12852 22430
rect 12908 22372 12964 26236
rect 13356 25508 13412 27132
rect 13468 27186 13524 28700
rect 13692 28756 13748 28766
rect 13692 28662 13748 28700
rect 13916 28308 13972 29708
rect 14028 29426 14084 29438
rect 14028 29374 14030 29426
rect 14082 29374 14084 29426
rect 14028 28644 14084 29374
rect 14028 28578 14084 28588
rect 14140 28420 14196 31612
rect 14252 31666 14308 31678
rect 14252 31614 14254 31666
rect 14306 31614 14308 31666
rect 14252 30436 14308 31614
rect 14364 31106 14420 34412
rect 14476 31332 14532 34636
rect 14588 34626 14644 34636
rect 14700 34690 14756 34702
rect 14700 34638 14702 34690
rect 14754 34638 14756 34690
rect 14588 34132 14644 34142
rect 14700 34132 14756 34638
rect 15148 34468 15204 34750
rect 15148 34412 15316 34468
rect 15036 34132 15092 34142
rect 14700 34130 15092 34132
rect 14700 34078 15038 34130
rect 15090 34078 15092 34130
rect 14700 34076 15092 34078
rect 14588 31554 14644 34076
rect 15036 34066 15092 34076
rect 15260 33908 15316 34412
rect 15260 33842 15316 33852
rect 14812 33234 14868 33246
rect 14812 33182 14814 33234
rect 14866 33182 14868 33234
rect 14700 32340 14756 32350
rect 14700 31778 14756 32284
rect 14700 31726 14702 31778
rect 14754 31726 14756 31778
rect 14700 31714 14756 31726
rect 14588 31502 14590 31554
rect 14642 31502 14644 31554
rect 14588 31490 14644 31502
rect 14476 31276 14644 31332
rect 14364 31054 14366 31106
rect 14418 31054 14420 31106
rect 14364 31042 14420 31054
rect 14588 31106 14644 31276
rect 14588 31054 14590 31106
rect 14642 31054 14644 31106
rect 14588 31042 14644 31054
rect 14476 30994 14532 31006
rect 14476 30942 14478 30994
rect 14530 30942 14532 30994
rect 14476 30884 14532 30942
rect 14476 30818 14532 30828
rect 14812 30772 14868 33182
rect 15372 32788 15428 37996
rect 15484 35700 15540 38332
rect 15596 37380 15652 38670
rect 15708 38668 15764 39004
rect 15932 38724 15988 39454
rect 16044 39396 16100 39406
rect 16044 39060 16100 39340
rect 16492 39060 16548 39070
rect 16044 39058 16212 39060
rect 16044 39006 16046 39058
rect 16098 39006 16212 39058
rect 16044 39004 16212 39006
rect 16044 38994 16100 39004
rect 15708 38612 15876 38668
rect 15932 38658 15988 38668
rect 15820 38050 15876 38612
rect 15820 37998 15822 38050
rect 15874 37998 15876 38050
rect 15820 37986 15876 37998
rect 15932 38052 15988 38062
rect 15708 37938 15764 37950
rect 15708 37886 15710 37938
rect 15762 37886 15764 37938
rect 15708 37604 15764 37886
rect 15708 37538 15764 37548
rect 15820 37492 15876 37502
rect 15820 37398 15876 37436
rect 15708 37380 15764 37390
rect 15596 37378 15764 37380
rect 15596 37326 15710 37378
rect 15762 37326 15764 37378
rect 15596 37324 15764 37326
rect 15708 37314 15764 37324
rect 15932 36708 15988 37996
rect 16044 37828 16100 37838
rect 16156 37828 16212 39004
rect 16380 38724 16436 38734
rect 16268 38052 16324 38090
rect 16268 37986 16324 37996
rect 16156 37772 16324 37828
rect 16044 37490 16100 37772
rect 16044 37438 16046 37490
rect 16098 37438 16100 37490
rect 16044 37426 16100 37438
rect 15932 36642 15988 36652
rect 16268 36148 16324 37772
rect 16380 37378 16436 38668
rect 16492 38050 16548 39004
rect 16492 37998 16494 38050
rect 16546 37998 16548 38050
rect 16492 37986 16548 37998
rect 16716 38050 16772 40348
rect 17164 40292 17220 43372
rect 17500 43362 17556 43372
rect 17948 43426 18004 44268
rect 18284 43652 18340 43662
rect 17948 43374 17950 43426
rect 18002 43374 18004 43426
rect 17836 42644 17892 42654
rect 17276 42642 17892 42644
rect 17276 42590 17838 42642
rect 17890 42590 17892 42642
rect 17276 42588 17892 42590
rect 17276 41298 17332 42588
rect 17836 42578 17892 42588
rect 17948 42644 18004 43374
rect 17948 42578 18004 42588
rect 18172 43650 18340 43652
rect 18172 43598 18286 43650
rect 18338 43598 18340 43650
rect 18172 43596 18340 43598
rect 17500 42084 17556 42094
rect 17276 41246 17278 41298
rect 17330 41246 17332 41298
rect 17276 41234 17332 41246
rect 17388 41972 17444 41982
rect 17388 41186 17444 41916
rect 17500 41858 17556 42028
rect 17500 41806 17502 41858
rect 17554 41806 17556 41858
rect 17500 41794 17556 41806
rect 18060 41860 18116 41870
rect 17388 41134 17390 41186
rect 17442 41134 17444 41186
rect 17388 41076 17444 41134
rect 17388 41010 17444 41020
rect 17948 40964 18004 40974
rect 17724 40962 18004 40964
rect 17724 40910 17950 40962
rect 18002 40910 18004 40962
rect 17724 40908 18004 40910
rect 16828 40236 17220 40292
rect 17276 40740 17332 40750
rect 16828 39842 16884 40236
rect 16828 39790 16830 39842
rect 16882 39790 16884 39842
rect 16828 39172 16884 39790
rect 17164 39844 17220 39854
rect 17276 39844 17332 40684
rect 17164 39842 17332 39844
rect 17164 39790 17166 39842
rect 17218 39790 17332 39842
rect 17164 39788 17332 39790
rect 17612 40290 17668 40302
rect 17612 40238 17614 40290
rect 17666 40238 17668 40290
rect 17164 39778 17220 39788
rect 17164 39618 17220 39630
rect 17164 39566 17166 39618
rect 17218 39566 17220 39618
rect 17164 39508 17220 39566
rect 16828 39116 16996 39172
rect 16716 37998 16718 38050
rect 16770 37998 16772 38050
rect 16716 37986 16772 37998
rect 16828 38724 16884 38762
rect 16828 38050 16884 38668
rect 16828 37998 16830 38050
rect 16882 37998 16884 38050
rect 16828 37986 16884 37998
rect 16604 37828 16660 37838
rect 16604 37826 16772 37828
rect 16604 37774 16606 37826
rect 16658 37774 16772 37826
rect 16604 37772 16772 37774
rect 16604 37762 16660 37772
rect 16380 37326 16382 37378
rect 16434 37326 16436 37378
rect 16380 37268 16436 37326
rect 16604 37268 16660 37278
rect 16380 37202 16436 37212
rect 16492 37212 16604 37268
rect 16380 36372 16436 36382
rect 16492 36372 16548 37212
rect 16604 37174 16660 37212
rect 16380 36370 16548 36372
rect 16380 36318 16382 36370
rect 16434 36318 16548 36370
rect 16380 36316 16548 36318
rect 16604 36372 16660 36382
rect 16380 36306 16436 36316
rect 16604 36278 16660 36316
rect 16324 36092 16436 36148
rect 16268 36054 16324 36092
rect 16044 35812 16100 35850
rect 16044 35746 16100 35756
rect 15484 35644 15988 35700
rect 16380 35698 16436 36092
rect 16716 36036 16772 37772
rect 15596 35474 15652 35486
rect 15596 35422 15598 35474
rect 15650 35422 15652 35474
rect 15484 34916 15540 34926
rect 15484 34802 15540 34860
rect 15484 34750 15486 34802
rect 15538 34750 15540 34802
rect 15484 34738 15540 34750
rect 15596 34468 15652 35422
rect 15708 35476 15764 35486
rect 15708 34914 15764 35420
rect 15708 34862 15710 34914
rect 15762 34862 15764 34914
rect 15708 34850 15764 34862
rect 15596 34402 15652 34412
rect 15596 34244 15652 34254
rect 15596 34150 15652 34188
rect 15708 33796 15764 33806
rect 15708 33346 15764 33740
rect 15708 33294 15710 33346
rect 15762 33294 15764 33346
rect 15708 33282 15764 33294
rect 15596 33236 15652 33246
rect 15596 33142 15652 33180
rect 15820 33236 15876 33246
rect 15372 32722 15428 32732
rect 15708 32788 15764 32798
rect 15708 32694 15764 32732
rect 15036 32676 15092 32686
rect 15036 32562 15092 32620
rect 15820 32674 15876 33180
rect 15820 32622 15822 32674
rect 15874 32622 15876 32674
rect 15820 32610 15876 32622
rect 15932 32676 15988 35644
rect 16156 35642 16212 35654
rect 16156 35590 16158 35642
rect 16210 35590 16212 35642
rect 16380 35646 16382 35698
rect 16434 35646 16436 35698
rect 16380 35634 16436 35646
rect 16492 35980 16772 36036
rect 16828 36596 16884 36606
rect 16156 35588 16212 35590
rect 16156 35522 16212 35532
rect 16380 35476 16436 35486
rect 16268 35364 16324 35374
rect 16044 34804 16100 34814
rect 16268 34804 16324 35308
rect 16380 34914 16436 35420
rect 16380 34862 16382 34914
rect 16434 34862 16436 34914
rect 16380 34850 16436 34862
rect 16044 34802 16324 34804
rect 16044 34750 16046 34802
rect 16098 34750 16324 34802
rect 16044 34748 16324 34750
rect 16044 33012 16100 34748
rect 16380 34692 16436 34702
rect 16380 34598 16436 34636
rect 16268 34356 16324 34366
rect 16044 32946 16100 32956
rect 16156 34300 16268 34356
rect 15932 32610 15988 32620
rect 15036 32510 15038 32562
rect 15090 32510 15092 32562
rect 15036 32498 15092 32510
rect 15484 32564 15540 32574
rect 15484 32470 15540 32508
rect 16156 32562 16212 34300
rect 16268 34290 16324 34300
rect 16268 33346 16324 33358
rect 16268 33294 16270 33346
rect 16322 33294 16324 33346
rect 16268 32788 16324 33294
rect 16268 32722 16324 32732
rect 16156 32510 16158 32562
rect 16210 32510 16212 32562
rect 15148 32452 15204 32462
rect 15148 32358 15204 32396
rect 14700 30716 14868 30772
rect 15036 32116 15092 32126
rect 14700 30548 14756 30716
rect 15036 30548 15092 32060
rect 16156 32116 16212 32510
rect 16156 32050 16212 32060
rect 14700 30492 14868 30548
rect 14252 30324 14308 30380
rect 14364 30324 14420 30334
rect 14252 30322 14420 30324
rect 14252 30270 14366 30322
rect 14418 30270 14420 30322
rect 14252 30268 14420 30270
rect 14364 30258 14420 30268
rect 14476 30324 14532 30334
rect 14476 30098 14532 30268
rect 14476 30046 14478 30098
rect 14530 30046 14532 30098
rect 14476 30034 14532 30046
rect 14588 30212 14644 30222
rect 14588 29876 14644 30156
rect 14812 30098 14868 30492
rect 15036 30482 15092 30492
rect 15148 31666 15204 31678
rect 15148 31614 15150 31666
rect 15202 31614 15204 31666
rect 15036 30324 15092 30334
rect 15036 30210 15092 30268
rect 15036 30158 15038 30210
rect 15090 30158 15092 30210
rect 15036 30146 15092 30158
rect 14812 30046 14814 30098
rect 14866 30046 14868 30098
rect 14812 30034 14868 30046
rect 14588 29810 14644 29820
rect 14252 29538 14308 29550
rect 14252 29486 14254 29538
rect 14306 29486 14308 29538
rect 14252 28756 14308 29486
rect 15036 29316 15092 29326
rect 15148 29316 15204 31614
rect 15484 31668 15540 31678
rect 15260 31554 15316 31566
rect 15260 31502 15262 31554
rect 15314 31502 15316 31554
rect 15260 30324 15316 31502
rect 15484 30994 15540 31612
rect 16156 31556 16212 31566
rect 15596 31108 15652 31118
rect 15596 31106 16100 31108
rect 15596 31054 15598 31106
rect 15650 31054 16100 31106
rect 15596 31052 16100 31054
rect 15596 31042 15652 31052
rect 15484 30942 15486 30994
rect 15538 30942 15540 30994
rect 15484 30930 15540 30942
rect 15372 30772 15428 30782
rect 15428 30716 15540 30772
rect 15372 30706 15428 30716
rect 15260 30258 15316 30268
rect 15372 29988 15428 29998
rect 15372 29894 15428 29932
rect 15036 29314 15204 29316
rect 15036 29262 15038 29314
rect 15090 29262 15204 29314
rect 15036 29260 15204 29262
rect 15372 29540 15428 29550
rect 15036 29250 15092 29260
rect 14252 28690 14308 28700
rect 15260 28532 15316 28542
rect 14140 28364 14308 28420
rect 13916 28242 13972 28252
rect 13468 27134 13470 27186
rect 13522 27134 13524 27186
rect 13468 27122 13524 27134
rect 13804 27746 13860 27758
rect 13804 27694 13806 27746
rect 13858 27694 13860 27746
rect 13692 27074 13748 27086
rect 13692 27022 13694 27074
rect 13746 27022 13748 27074
rect 13692 26180 13748 27022
rect 13804 26740 13860 27694
rect 14252 27748 14308 28364
rect 13804 26674 13860 26684
rect 13916 27074 13972 27086
rect 13916 27022 13918 27074
rect 13970 27022 13972 27074
rect 13916 26964 13972 27022
rect 13916 26740 13972 26908
rect 13916 26684 14196 26740
rect 13468 25956 13524 25966
rect 13468 25730 13524 25900
rect 13468 25678 13470 25730
rect 13522 25678 13524 25730
rect 13468 25666 13524 25678
rect 13580 25620 13636 25630
rect 13580 25526 13636 25564
rect 13356 25442 13412 25452
rect 13244 24948 13300 24958
rect 13692 24948 13748 26124
rect 13244 24946 13412 24948
rect 13244 24894 13246 24946
rect 13298 24894 13412 24946
rect 13244 24892 13412 24894
rect 13244 24882 13300 24892
rect 13132 24834 13188 24846
rect 13132 24782 13134 24834
rect 13186 24782 13188 24834
rect 13020 24724 13076 24734
rect 13020 24630 13076 24668
rect 13020 24162 13076 24174
rect 13020 24110 13022 24162
rect 13074 24110 13076 24162
rect 13020 24050 13076 24110
rect 13020 23998 13022 24050
rect 13074 23998 13076 24050
rect 13020 23986 13076 23998
rect 13020 23268 13076 23278
rect 13132 23268 13188 24782
rect 13020 23266 13188 23268
rect 13020 23214 13022 23266
rect 13074 23214 13188 23266
rect 13020 23212 13188 23214
rect 13020 22596 13076 23212
rect 13244 23156 13300 23166
rect 13244 23062 13300 23100
rect 13020 22540 13300 22596
rect 12908 22316 13076 22372
rect 12908 22148 12964 22158
rect 12908 22054 12964 22092
rect 12908 21700 12964 21710
rect 12908 21606 12964 21644
rect 12796 21084 12964 21140
rect 12796 20916 12852 20926
rect 12124 20750 12126 20802
rect 12178 20750 12180 20802
rect 12124 20356 12180 20750
rect 12348 20914 12852 20916
rect 12348 20862 12798 20914
rect 12850 20862 12852 20914
rect 12348 20860 12852 20862
rect 12348 20802 12404 20860
rect 12796 20850 12852 20860
rect 12348 20750 12350 20802
rect 12402 20750 12404 20802
rect 12348 20738 12404 20750
rect 12684 20580 12740 20590
rect 12124 20290 12180 20300
rect 12236 20468 12292 20478
rect 12236 19460 12292 20412
rect 12684 20018 12740 20524
rect 12684 19966 12686 20018
rect 12738 19966 12740 20018
rect 12684 19954 12740 19966
rect 12796 20018 12852 20030
rect 12796 19966 12798 20018
rect 12850 19966 12852 20018
rect 12236 19458 12404 19460
rect 12236 19406 12238 19458
rect 12290 19406 12404 19458
rect 12236 19404 12404 19406
rect 12236 19394 12292 19404
rect 12236 19236 12292 19246
rect 12236 19142 12292 19180
rect 12124 19012 12180 19022
rect 12124 18674 12180 18956
rect 12124 18622 12126 18674
rect 12178 18622 12180 18674
rect 12124 18610 12180 18622
rect 12236 18228 12292 18238
rect 12236 18134 12292 18172
rect 12236 17666 12292 17678
rect 12236 17614 12238 17666
rect 12290 17614 12292 17666
rect 12236 16996 12292 17614
rect 12236 16930 12292 16940
rect 12124 16884 12180 16894
rect 12124 16790 12180 16828
rect 12012 16604 12180 16660
rect 11900 16270 11902 16322
rect 11954 16270 11956 16322
rect 11900 16258 11956 16270
rect 11676 16044 11844 16100
rect 11788 15316 11844 16044
rect 12012 15988 12068 15998
rect 12012 15894 12068 15932
rect 11900 15874 11956 15886
rect 11900 15822 11902 15874
rect 11954 15822 11956 15874
rect 11900 15540 11956 15822
rect 11900 15474 11956 15484
rect 11788 15222 11844 15260
rect 11564 15202 11620 15214
rect 11564 15150 11566 15202
rect 11618 15150 11620 15202
rect 11564 14644 11620 15150
rect 11564 14578 11620 14588
rect 12012 14644 12068 14654
rect 12012 14550 12068 14588
rect 11452 13918 11454 13970
rect 11506 13918 11508 13970
rect 10892 13132 11172 13188
rect 11340 13748 11396 13758
rect 10444 13076 10500 13086
rect 10444 12982 10500 13020
rect 10332 12910 10334 12962
rect 10386 12910 10388 12962
rect 10332 12898 10388 12910
rect 10556 12850 10612 12862
rect 10556 12798 10558 12850
rect 10610 12798 10612 12850
rect 10220 12460 10500 12516
rect 9996 12450 10052 12460
rect 10444 12404 10500 12460
rect 9884 11666 9940 11676
rect 9996 12292 10052 12302
rect 9996 11618 10052 12236
rect 10332 12180 10388 12190
rect 10444 12180 10500 12348
rect 10556 12292 10612 12798
rect 10892 12292 10948 13132
rect 11004 12964 11060 12974
rect 11004 12962 11284 12964
rect 11004 12910 11006 12962
rect 11058 12910 11284 12962
rect 11004 12908 11284 12910
rect 11004 12898 11060 12908
rect 11116 12404 11172 12414
rect 11116 12310 11172 12348
rect 10556 12236 10948 12292
rect 11228 12292 11284 12908
rect 10332 12178 10500 12180
rect 10332 12126 10334 12178
rect 10386 12126 10500 12178
rect 10332 12124 10500 12126
rect 10332 12114 10388 12124
rect 9996 11566 9998 11618
rect 10050 11566 10052 11618
rect 9996 11554 10052 11566
rect 10108 12068 10164 12078
rect 9772 11342 9774 11394
rect 9826 11342 9828 11394
rect 9660 11172 9716 11182
rect 9660 10834 9716 11116
rect 9660 10782 9662 10834
rect 9714 10782 9716 10834
rect 9660 10770 9716 10782
rect 9772 10612 9828 11342
rect 9884 11396 9940 11406
rect 9884 10722 9940 11340
rect 10108 10948 10164 12012
rect 10668 12066 10724 12078
rect 10668 12014 10670 12066
rect 10722 12014 10724 12066
rect 10668 11508 10724 12014
rect 10668 11442 10724 11452
rect 10220 11396 10276 11406
rect 10220 11302 10276 11340
rect 9884 10670 9886 10722
rect 9938 10670 9940 10722
rect 9884 10658 9940 10670
rect 9996 10892 10164 10948
rect 10332 11282 10388 11294
rect 10332 11230 10334 11282
rect 10386 11230 10388 11282
rect 9772 10546 9828 10556
rect 9996 10500 10052 10892
rect 10108 10724 10164 10734
rect 10332 10724 10388 11230
rect 10668 11170 10724 11182
rect 10668 11118 10670 11170
rect 10722 11118 10724 11170
rect 10108 10722 10388 10724
rect 10108 10670 10110 10722
rect 10162 10670 10388 10722
rect 10108 10668 10388 10670
rect 10108 10658 10164 10668
rect 9996 10444 10164 10500
rect 7868 9996 8372 10052
rect 9212 10220 9604 10276
rect 7532 9884 7812 9940
rect 6972 9774 6974 9826
rect 7026 9774 7028 9826
rect 6972 9762 7028 9774
rect 7308 9716 7364 9726
rect 7532 9716 7588 9726
rect 7308 9714 7588 9716
rect 7308 9662 7310 9714
rect 7362 9662 7534 9714
rect 7586 9662 7588 9714
rect 7308 9660 7588 9662
rect 7308 9650 7364 9660
rect 7532 9650 7588 9660
rect 6524 9604 6580 9614
rect 6524 9510 6580 9548
rect 7084 9604 7140 9614
rect 7084 9510 7140 9548
rect 7644 9602 7700 9614
rect 7644 9550 7646 9602
rect 7698 9550 7700 9602
rect 7644 9268 7700 9550
rect 7756 9604 7812 9884
rect 7868 9826 7924 9996
rect 9212 9938 9268 10220
rect 9212 9886 9214 9938
rect 9266 9886 9268 9938
rect 9212 9874 9268 9886
rect 7868 9774 7870 9826
rect 7922 9774 7924 9826
rect 7868 9762 7924 9774
rect 7980 9826 8036 9838
rect 7980 9774 7982 9826
rect 8034 9774 8036 9826
rect 7756 9538 7812 9548
rect 6860 9212 7700 9268
rect 6860 9154 6916 9212
rect 6860 9102 6862 9154
rect 6914 9102 6916 9154
rect 6860 9090 6916 9102
rect 5516 8990 5518 9042
rect 5570 8990 5572 9042
rect 5068 8764 5348 8820
rect 4396 8754 4452 8764
rect 4476 8652 4740 8662
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4476 8586 4740 8596
rect 5180 8596 5236 8606
rect 4620 8372 4676 8382
rect 4956 8372 5012 8382
rect 4620 8370 5012 8372
rect 4620 8318 4622 8370
rect 4674 8318 4958 8370
rect 5010 8318 5012 8370
rect 4620 8316 5012 8318
rect 4620 8306 4676 8316
rect 4956 8306 5012 8316
rect 5068 8036 5124 8046
rect 5180 8036 5236 8540
rect 5068 8034 5236 8036
rect 5068 7982 5070 8034
rect 5122 7982 5236 8034
rect 5068 7980 5236 7982
rect 5068 7970 5124 7980
rect 4060 7534 4062 7586
rect 4114 7534 4116 7586
rect 4060 7522 4116 7534
rect 3724 7196 4116 7252
rect 1708 6018 1764 6030
rect 1708 5966 1710 6018
rect 1762 5966 1764 6018
rect 1708 5460 1764 5966
rect 1708 5394 1764 5404
rect 4060 5012 4116 7196
rect 5292 7140 5348 8764
rect 5516 8148 5572 8990
rect 5852 9042 6356 9044
rect 5852 8990 6190 9042
rect 6242 8990 6356 9042
rect 5852 8988 6356 8990
rect 7980 9044 8036 9774
rect 9996 9828 10052 9838
rect 9996 9734 10052 9772
rect 5740 8372 5796 8382
rect 5852 8372 5908 8988
rect 6188 8978 6244 8988
rect 7980 8978 8036 8988
rect 8988 9604 9044 9614
rect 8988 8930 9044 9548
rect 8988 8878 8990 8930
rect 9042 8878 9044 8930
rect 8988 8708 9044 8878
rect 9996 8932 10052 8942
rect 9996 8838 10052 8876
rect 8988 8642 9044 8652
rect 5740 8370 5852 8372
rect 5740 8318 5742 8370
rect 5794 8318 5852 8370
rect 5740 8316 5852 8318
rect 5740 8306 5796 8316
rect 5852 8278 5908 8316
rect 7084 8372 7140 8382
rect 5516 8082 5572 8092
rect 6636 8148 6692 8158
rect 6636 7698 6692 8092
rect 7084 7700 7140 8316
rect 9436 8260 9492 8270
rect 9436 8166 9492 8204
rect 8876 8036 8932 8046
rect 8988 8036 9044 8046
rect 8876 8034 8988 8036
rect 8876 7982 8878 8034
rect 8930 7982 8988 8034
rect 8876 7980 8988 7982
rect 8876 7970 8932 7980
rect 6636 7646 6638 7698
rect 6690 7646 6692 7698
rect 6636 7634 6692 7646
rect 6748 7698 7140 7700
rect 6748 7646 7086 7698
rect 7138 7646 7140 7698
rect 6748 7644 7140 7646
rect 6524 7476 6580 7486
rect 6188 7474 6580 7476
rect 6188 7422 6526 7474
rect 6578 7422 6580 7474
rect 6188 7420 6580 7422
rect 6188 7362 6244 7420
rect 6524 7410 6580 7420
rect 6188 7310 6190 7362
rect 6242 7310 6244 7362
rect 6188 7298 6244 7310
rect 4476 7084 4740 7094
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 5292 7074 5348 7084
rect 6524 7140 6580 7150
rect 4476 7018 4740 7028
rect 6524 6690 6580 7084
rect 6524 6638 6526 6690
rect 6578 6638 6580 6690
rect 6524 6626 6580 6638
rect 6524 6244 6580 6254
rect 6300 6132 6356 6142
rect 6300 6038 6356 6076
rect 5852 5796 5908 5806
rect 5516 5794 5908 5796
rect 5516 5742 5854 5794
rect 5906 5742 5908 5794
rect 5516 5740 5908 5742
rect 4476 5516 4740 5526
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4476 5450 4740 5460
rect 1708 4900 1764 4910
rect 1708 4806 1764 4844
rect 4060 4562 4116 4956
rect 5068 5012 5124 5022
rect 5068 4918 5124 4956
rect 4060 4510 4062 4562
rect 4114 4510 4116 4562
rect 4060 4498 4116 4510
rect 1708 4450 1764 4462
rect 1708 4398 1710 4450
rect 1762 4398 1764 4450
rect 1708 4116 1764 4398
rect 1708 4050 1764 4060
rect 5516 4116 5572 5740
rect 5852 5730 5908 5740
rect 5628 5124 5684 5134
rect 6412 5124 6468 5134
rect 5628 5122 6468 5124
rect 5628 5070 5630 5122
rect 5682 5070 6414 5122
rect 6466 5070 6468 5122
rect 5628 5068 6468 5070
rect 5628 5058 5684 5068
rect 6412 5058 6468 5068
rect 6524 5010 6580 6188
rect 6636 6132 6692 6142
rect 6748 6132 6804 7644
rect 7084 7634 7140 7644
rect 7532 7362 7588 7374
rect 7532 7310 7534 7362
rect 7586 7310 7588 7362
rect 7420 7252 7476 7262
rect 7196 7250 7476 7252
rect 7196 7198 7422 7250
rect 7474 7198 7476 7250
rect 7196 7196 7476 7198
rect 7196 6802 7252 7196
rect 7420 7186 7476 7196
rect 7196 6750 7198 6802
rect 7250 6750 7252 6802
rect 7196 6738 7252 6750
rect 6636 6130 6804 6132
rect 6636 6078 6638 6130
rect 6690 6078 6804 6130
rect 6636 6076 6804 6078
rect 6636 6066 6692 6076
rect 6748 5796 6804 6076
rect 7420 6132 7476 6142
rect 7420 6038 7476 6076
rect 7532 6130 7588 7310
rect 8652 7364 8708 7374
rect 8652 7362 8932 7364
rect 8652 7310 8654 7362
rect 8706 7310 8932 7362
rect 8652 7308 8932 7310
rect 8652 7298 8708 7308
rect 8092 6580 8148 6590
rect 7532 6078 7534 6130
rect 7586 6078 7588 6130
rect 7532 6066 7588 6078
rect 7644 6244 7700 6254
rect 7644 6130 7700 6188
rect 7644 6078 7646 6130
rect 7698 6078 7700 6130
rect 7644 6066 7700 6078
rect 7756 6018 7812 6030
rect 7756 5966 7758 6018
rect 7810 5966 7812 6018
rect 7084 5908 7140 5918
rect 7084 5814 7140 5852
rect 6972 5796 7028 5806
rect 6748 5730 6804 5740
rect 6860 5794 7028 5796
rect 6860 5742 6974 5794
rect 7026 5742 7028 5794
rect 6860 5740 7028 5742
rect 6748 5348 6804 5358
rect 6524 4958 6526 5010
rect 6578 4958 6580 5010
rect 6524 4946 6580 4958
rect 6636 5292 6748 5348
rect 6636 5010 6692 5292
rect 6748 5282 6804 5292
rect 6636 4958 6638 5010
rect 6690 4958 6692 5010
rect 6636 4946 6692 4958
rect 6748 5124 6804 5134
rect 5740 4900 5796 4910
rect 6300 4900 6356 4910
rect 5740 4898 6244 4900
rect 5740 4846 5742 4898
rect 5794 4846 6244 4898
rect 5740 4844 6244 4846
rect 5740 4834 5796 4844
rect 6188 4452 6244 4844
rect 6300 4806 6356 4844
rect 6748 4788 6804 5068
rect 6636 4732 6804 4788
rect 6300 4452 6356 4462
rect 6188 4450 6356 4452
rect 6188 4398 6302 4450
rect 6354 4398 6356 4450
rect 6188 4396 6356 4398
rect 6300 4386 6356 4396
rect 6524 4452 6580 4462
rect 5516 4050 5572 4060
rect 5852 4340 5908 4350
rect 4476 3948 4740 3958
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4476 3882 4740 3892
rect 5068 3892 5124 3902
rect 4620 3668 4676 3678
rect 4620 3574 4676 3612
rect 5068 3666 5124 3836
rect 5068 3614 5070 3666
rect 5122 3614 5124 3666
rect 5068 3602 5124 3614
rect 5852 3666 5908 4284
rect 6188 4228 6244 4238
rect 6188 3778 6244 4172
rect 6188 3726 6190 3778
rect 6242 3726 6244 3778
rect 6188 3714 6244 3726
rect 5852 3614 5854 3666
rect 5906 3614 5908 3666
rect 5852 3602 5908 3614
rect 6524 3666 6580 4396
rect 6636 3778 6692 4732
rect 6636 3726 6638 3778
rect 6690 3726 6692 3778
rect 6636 3714 6692 3726
rect 6748 4116 6804 4126
rect 6524 3614 6526 3666
rect 6578 3614 6580 3666
rect 6524 3602 6580 3614
rect 6748 3668 6804 4060
rect 6860 4004 6916 5740
rect 6972 5730 7028 5740
rect 7420 5796 7476 5806
rect 6972 5122 7028 5134
rect 7420 5124 7476 5740
rect 7756 5348 7812 5966
rect 7756 5282 7812 5292
rect 6972 5070 6974 5122
rect 7026 5070 7028 5122
rect 6972 4116 7028 5070
rect 7084 5122 7476 5124
rect 7084 5070 7422 5122
rect 7474 5070 7476 5122
rect 7084 5068 7476 5070
rect 7084 4340 7140 5068
rect 7420 5058 7476 5068
rect 7532 4564 7588 4574
rect 7532 4470 7588 4508
rect 8092 4562 8148 6524
rect 8652 6356 8708 6366
rect 8652 6130 8708 6300
rect 8652 6078 8654 6130
rect 8706 6078 8708 6130
rect 8652 6066 8708 6078
rect 8204 5906 8260 5918
rect 8204 5854 8206 5906
rect 8258 5854 8260 5906
rect 8204 5684 8260 5854
rect 8540 5908 8596 5918
rect 8540 5814 8596 5852
rect 8764 5908 8820 5918
rect 8652 5684 8708 5694
rect 8204 5682 8708 5684
rect 8204 5630 8654 5682
rect 8706 5630 8708 5682
rect 8204 5628 8708 5630
rect 8652 5618 8708 5628
rect 8540 5236 8596 5246
rect 8204 5124 8260 5134
rect 8204 5030 8260 5068
rect 8428 5124 8484 5134
rect 8092 4510 8094 4562
rect 8146 4510 8148 4562
rect 8092 4498 8148 4510
rect 8428 4450 8484 5068
rect 8540 4562 8596 5180
rect 8540 4510 8542 4562
rect 8594 4510 8596 4562
rect 8540 4498 8596 4510
rect 8428 4398 8430 4450
rect 8482 4398 8484 4450
rect 8428 4386 8484 4398
rect 7084 4246 7140 4284
rect 7420 4340 7476 4350
rect 7420 4246 7476 4284
rect 7980 4226 8036 4238
rect 7980 4174 7982 4226
rect 8034 4174 8036 4226
rect 7532 4116 7588 4126
rect 6972 4114 7588 4116
rect 6972 4062 7534 4114
rect 7586 4062 7588 4114
rect 6972 4060 7588 4062
rect 7532 4050 7588 4060
rect 6860 3948 7476 4004
rect 7420 3892 7476 3948
rect 7420 3836 7700 3892
rect 6748 3612 7252 3668
rect 4172 3556 4228 3566
rect 4172 3462 4228 3500
rect 1708 3444 1764 3454
rect 1708 3330 1764 3388
rect 6076 3444 6132 3482
rect 6076 3378 6132 3388
rect 1708 3278 1710 3330
rect 1762 3278 1764 3330
rect 1708 3266 1764 3278
rect 2156 3330 2212 3342
rect 2156 3278 2158 3330
rect 2210 3278 2212 3330
rect 2156 2772 2212 3278
rect 2156 2706 2212 2716
rect 6748 800 6804 3612
rect 7196 3554 7252 3612
rect 7196 3502 7198 3554
rect 7250 3502 7252 3554
rect 7196 3490 7252 3502
rect 7420 3556 7476 3566
rect 6972 3444 7028 3482
rect 6972 3378 7028 3388
rect 7420 800 7476 3500
rect 7644 3442 7700 3836
rect 7980 3780 8036 4174
rect 7980 3714 8036 3724
rect 8428 3668 8484 3678
rect 7868 3556 7924 3566
rect 7868 3462 7924 3500
rect 8428 3554 8484 3612
rect 8428 3502 8430 3554
rect 8482 3502 8484 3554
rect 8428 3490 8484 3502
rect 7644 3390 7646 3442
rect 7698 3390 7700 3442
rect 7644 3378 7700 3390
rect 8764 3442 8820 5852
rect 8876 5796 8932 7308
rect 8988 7140 9044 7980
rect 9772 8036 9828 8046
rect 9772 7476 9828 7980
rect 9884 7476 9940 7486
rect 9772 7474 9940 7476
rect 9772 7422 9886 7474
rect 9938 7422 9940 7474
rect 9772 7420 9940 7422
rect 8988 7074 9044 7084
rect 9100 7362 9156 7374
rect 9100 7310 9102 7362
rect 9154 7310 9156 7362
rect 9100 7028 9156 7310
rect 9100 6962 9156 6972
rect 9772 6916 9828 6926
rect 9324 6804 9380 6814
rect 9772 6804 9828 6860
rect 9324 6802 9828 6804
rect 9324 6750 9326 6802
rect 9378 6750 9828 6802
rect 9324 6748 9828 6750
rect 9324 6738 9380 6748
rect 8876 5730 8932 5740
rect 8876 4900 8932 4910
rect 8876 4450 8932 4844
rect 8876 4398 8878 4450
rect 8930 4398 8932 4450
rect 8876 4386 8932 4398
rect 9660 4338 9716 6748
rect 9772 6690 9828 6748
rect 9884 6804 9940 7420
rect 9884 6738 9940 6748
rect 9772 6638 9774 6690
rect 9826 6638 9828 6690
rect 9772 6626 9828 6638
rect 10108 6692 10164 10444
rect 10332 10050 10388 10668
rect 10556 10836 10612 10846
rect 10556 10610 10612 10780
rect 10556 10558 10558 10610
rect 10610 10558 10612 10610
rect 10556 10546 10612 10558
rect 10668 10500 10724 11118
rect 10780 10724 10836 12236
rect 11228 12198 11284 12236
rect 11340 11788 11396 13692
rect 11452 13074 11508 13918
rect 11452 13022 11454 13074
rect 11506 13022 11508 13074
rect 11452 13010 11508 13022
rect 12012 13636 12068 13646
rect 12124 13636 12180 16604
rect 12236 16098 12292 16110
rect 12236 16046 12238 16098
rect 12290 16046 12292 16098
rect 12236 15538 12292 16046
rect 12236 15486 12238 15538
rect 12290 15486 12292 15538
rect 12236 15474 12292 15486
rect 12236 15316 12292 15326
rect 12348 15316 12404 19404
rect 12796 18676 12852 19966
rect 12908 19908 12964 21084
rect 12908 19236 12964 19852
rect 13020 20132 13076 22316
rect 13020 19346 13076 20076
rect 13020 19294 13022 19346
rect 13074 19294 13076 19346
rect 13020 19282 13076 19294
rect 13132 22260 13188 22270
rect 12908 19170 12964 19180
rect 12796 18610 12852 18620
rect 12908 18564 12964 18574
rect 13132 18564 13188 22204
rect 13244 21924 13300 22540
rect 13244 21858 13300 21868
rect 13356 21140 13412 24892
rect 13692 23938 13748 24892
rect 13692 23886 13694 23938
rect 13746 23886 13748 23938
rect 13692 23874 13748 23886
rect 13804 26292 13860 26302
rect 13916 26292 13972 26684
rect 13804 26290 13972 26292
rect 13804 26238 13806 26290
rect 13858 26238 13972 26290
rect 13804 26236 13972 26238
rect 14028 26516 14084 26526
rect 13580 23828 13636 23838
rect 13580 23734 13636 23772
rect 13804 23604 13860 26236
rect 13916 24722 13972 24734
rect 13916 24670 13918 24722
rect 13970 24670 13972 24722
rect 13916 24500 13972 24670
rect 13916 24434 13972 24444
rect 13580 23548 13860 23604
rect 13916 24276 13972 24286
rect 13468 22260 13524 22270
rect 13468 22166 13524 22204
rect 13580 21252 13636 23548
rect 13916 23378 13972 24220
rect 13916 23326 13918 23378
rect 13970 23326 13972 23378
rect 13916 23314 13972 23326
rect 14028 23044 14084 26460
rect 14140 25620 14196 26684
rect 14252 26178 14308 27692
rect 14252 26126 14254 26178
rect 14306 26126 14308 26178
rect 14252 26114 14308 26126
rect 14476 28308 14532 28318
rect 14252 25620 14308 25630
rect 14140 25618 14308 25620
rect 14140 25566 14254 25618
rect 14306 25566 14308 25618
rect 14140 25564 14308 25566
rect 14252 25554 14308 25564
rect 14476 25284 14532 28252
rect 15036 28084 15092 28094
rect 14812 27858 14868 27870
rect 14812 27806 14814 27858
rect 14866 27806 14868 27858
rect 14812 27524 14868 27806
rect 14812 27458 14868 27468
rect 14924 27746 14980 27758
rect 14924 27694 14926 27746
rect 14978 27694 14980 27746
rect 14924 27300 14980 27694
rect 15036 27412 15092 28028
rect 15036 27346 15092 27356
rect 15260 27860 15316 28476
rect 14924 27234 14980 27244
rect 15036 27188 15092 27198
rect 15260 27188 15316 27804
rect 15372 27858 15428 29484
rect 15484 28644 15540 30716
rect 15708 30660 15764 30670
rect 15708 30210 15764 30604
rect 16044 30548 16100 31052
rect 16156 30994 16212 31500
rect 16156 30942 16158 30994
rect 16210 30942 16212 30994
rect 16156 30930 16212 30942
rect 16492 30996 16548 35980
rect 16604 35812 16660 35822
rect 16604 34914 16660 35756
rect 16604 34862 16606 34914
rect 16658 34862 16660 34914
rect 16604 34850 16660 34862
rect 16716 35698 16772 35710
rect 16716 35646 16718 35698
rect 16770 35646 16772 35698
rect 16716 34580 16772 35646
rect 16828 35700 16884 36540
rect 16828 35634 16884 35644
rect 16716 32786 16772 34524
rect 16828 35474 16884 35486
rect 16828 35422 16830 35474
rect 16882 35422 16884 35474
rect 16828 33346 16884 35422
rect 16940 34356 16996 39116
rect 17164 38052 17220 39452
rect 17612 39284 17668 40238
rect 17724 39620 17780 40908
rect 17948 40898 18004 40908
rect 18060 40628 18116 41804
rect 18060 40562 18116 40572
rect 17948 40292 18004 40302
rect 17724 39554 17780 39564
rect 17836 40290 18004 40292
rect 17836 40238 17950 40290
rect 18002 40238 18004 40290
rect 17836 40236 18004 40238
rect 17612 39218 17668 39228
rect 17388 38724 17444 38734
rect 17836 38722 17892 40236
rect 17948 40226 18004 40236
rect 18172 40180 18228 43596
rect 18284 43586 18340 43596
rect 18284 42084 18340 42094
rect 18284 41990 18340 42028
rect 18396 41298 18452 44940
rect 18732 44548 18788 45614
rect 19292 45444 19348 45724
rect 19404 45714 19460 45724
rect 19292 45378 19348 45388
rect 18732 44482 18788 44492
rect 19292 44996 19348 45006
rect 18508 44212 18564 44222
rect 18508 44210 18900 44212
rect 18508 44158 18510 44210
rect 18562 44158 18900 44210
rect 18508 44156 18900 44158
rect 18508 44146 18564 44156
rect 18620 43764 18676 43774
rect 18620 43652 18676 43708
rect 18508 43650 18676 43652
rect 18508 43598 18622 43650
rect 18674 43598 18676 43650
rect 18508 43596 18676 43598
rect 18508 41972 18564 43596
rect 18620 43586 18676 43596
rect 18844 43316 18900 44156
rect 19068 43876 19124 43886
rect 19068 43650 19124 43820
rect 19292 43764 19348 44940
rect 19292 43698 19348 43708
rect 19068 43598 19070 43650
rect 19122 43598 19124 43650
rect 19068 43586 19124 43598
rect 18956 43540 19012 43550
rect 18956 43446 19012 43484
rect 19292 43540 19348 43550
rect 19292 43538 19460 43540
rect 19292 43486 19294 43538
rect 19346 43486 19460 43538
rect 19292 43484 19460 43486
rect 19292 43474 19348 43484
rect 18844 43260 19124 43316
rect 19068 42866 19124 43260
rect 19068 42814 19070 42866
rect 19122 42814 19124 42866
rect 19068 42802 19124 42814
rect 18620 42754 18676 42766
rect 18620 42702 18622 42754
rect 18674 42702 18676 42754
rect 18620 42644 18676 42702
rect 18620 42578 18676 42588
rect 19404 42642 19460 43484
rect 19404 42590 19406 42642
rect 19458 42590 19460 42642
rect 19404 42578 19460 42590
rect 19516 42644 19572 42654
rect 18956 42532 19012 42542
rect 18508 41878 18564 41916
rect 18844 42530 19012 42532
rect 18844 42478 18958 42530
rect 19010 42478 19012 42530
rect 18844 42476 19012 42478
rect 18844 41300 18900 42476
rect 18956 42466 19012 42476
rect 19068 42532 19124 42542
rect 19068 42308 19124 42476
rect 19180 42530 19236 42542
rect 19180 42478 19182 42530
rect 19234 42478 19236 42530
rect 19180 42420 19236 42478
rect 19180 42354 19236 42364
rect 18956 42252 19124 42308
rect 18956 42082 19012 42252
rect 18956 42030 18958 42082
rect 19010 42030 19012 42082
rect 18956 42018 19012 42030
rect 18396 41246 18398 41298
rect 18450 41246 18452 41298
rect 18396 41234 18452 41246
rect 18732 41244 18900 41300
rect 18508 41186 18564 41198
rect 18508 41134 18510 41186
rect 18562 41134 18564 41186
rect 18284 41076 18340 41086
rect 18284 40982 18340 41020
rect 18284 40628 18340 40638
rect 18284 40534 18340 40572
rect 18508 40404 18564 41134
rect 18508 40338 18564 40348
rect 18620 40516 18676 40526
rect 18060 39394 18116 39406
rect 18060 39342 18062 39394
rect 18114 39342 18116 39394
rect 18060 38836 18116 39342
rect 18060 38770 18116 38780
rect 18172 38946 18228 40124
rect 18172 38894 18174 38946
rect 18226 38894 18228 38946
rect 17836 38670 17838 38722
rect 17890 38670 17892 38722
rect 17836 38668 17892 38670
rect 18172 38668 18228 38894
rect 17388 38612 17892 38668
rect 17948 38612 18228 38668
rect 18396 39618 18452 39630
rect 18396 39566 18398 39618
rect 18450 39566 18452 39618
rect 18396 38668 18452 39566
rect 18620 39618 18676 40460
rect 18620 39566 18622 39618
rect 18674 39566 18676 39618
rect 18620 39060 18676 39566
rect 18620 38994 18676 39004
rect 18732 38668 18788 41244
rect 18844 41076 18900 41086
rect 18844 41074 19012 41076
rect 18844 41022 18846 41074
rect 18898 41022 19012 41074
rect 18844 41020 19012 41022
rect 18844 41010 18900 41020
rect 18844 40852 18900 40862
rect 18844 40402 18900 40796
rect 18844 40350 18846 40402
rect 18898 40350 18900 40402
rect 18844 40338 18900 40350
rect 18956 39730 19012 41020
rect 19404 40962 19460 40974
rect 19404 40910 19406 40962
rect 19458 40910 19460 40962
rect 19180 40404 19236 40414
rect 19180 40310 19236 40348
rect 19292 40290 19348 40302
rect 19292 40238 19294 40290
rect 19346 40238 19348 40290
rect 19292 40180 19348 40238
rect 19292 40114 19348 40124
rect 19404 39732 19460 40910
rect 19516 40404 19572 42588
rect 19628 40628 19684 45838
rect 20076 45892 20132 45902
rect 20188 45892 20244 49200
rect 20076 45890 20244 45892
rect 20076 45838 20078 45890
rect 20130 45838 20244 45890
rect 20076 45836 20244 45838
rect 20076 45668 20132 45836
rect 20076 45602 20132 45612
rect 20972 45666 21028 45678
rect 20972 45614 20974 45666
rect 21026 45614 21028 45666
rect 19836 45500 20100 45510
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 19836 45434 20100 45444
rect 20748 45108 20804 45118
rect 20972 45108 21028 45614
rect 20748 45106 21028 45108
rect 20748 45054 20750 45106
rect 20802 45054 21028 45106
rect 20748 45052 21028 45054
rect 22876 45108 22932 49200
rect 23548 46340 23604 49200
rect 23548 46284 23828 46340
rect 22988 45666 23044 45678
rect 22988 45614 22990 45666
rect 23042 45614 23044 45666
rect 22988 45332 23044 45614
rect 22988 45266 23044 45276
rect 20412 44996 20468 45006
rect 20412 44902 20468 44940
rect 20636 44436 20692 44446
rect 20188 44434 20692 44436
rect 20188 44382 20638 44434
rect 20690 44382 20692 44434
rect 20188 44380 20692 44382
rect 19836 43932 20100 43942
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 19836 43866 20100 43876
rect 19740 43426 19796 43438
rect 19740 43374 19742 43426
rect 19794 43374 19796 43426
rect 19740 42756 19796 43374
rect 20188 42868 20244 44380
rect 20636 44370 20692 44380
rect 19740 42690 19796 42700
rect 19964 42812 20244 42868
rect 19964 42754 20020 42812
rect 19964 42702 19966 42754
rect 20018 42702 20020 42754
rect 19964 42532 20020 42702
rect 19964 42466 20020 42476
rect 19836 42364 20100 42374
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 19836 42298 20100 42308
rect 19852 42084 19908 42094
rect 19852 41186 19908 42028
rect 19852 41134 19854 41186
rect 19906 41134 19908 41186
rect 19852 41122 19908 41134
rect 19964 41972 20020 41982
rect 19964 41074 20020 41916
rect 19964 41022 19966 41074
rect 20018 41022 20020 41074
rect 19964 41010 20020 41022
rect 20188 40852 20244 42812
rect 20412 43764 20468 43774
rect 20412 42754 20468 43708
rect 20412 42702 20414 42754
rect 20466 42702 20468 42754
rect 20412 42196 20468 42702
rect 20636 43428 20692 43438
rect 20748 43428 20804 45052
rect 22876 45042 22932 45052
rect 23100 45220 23156 45230
rect 21532 44996 21588 45006
rect 21420 44994 21588 44996
rect 21420 44942 21534 44994
rect 21586 44942 21588 44994
rect 21420 44940 21588 44942
rect 21420 43762 21476 44940
rect 21532 44930 21588 44940
rect 22652 44996 22708 45006
rect 21980 44436 22036 44446
rect 21868 44324 21924 44334
rect 21868 44230 21924 44268
rect 21532 44100 21588 44110
rect 21532 44098 21700 44100
rect 21532 44046 21534 44098
rect 21586 44046 21700 44098
rect 21532 44044 21700 44046
rect 21532 44034 21588 44044
rect 21420 43710 21422 43762
rect 21474 43710 21476 43762
rect 21420 43698 21476 43710
rect 21644 43538 21700 44044
rect 21644 43486 21646 43538
rect 21698 43486 21700 43538
rect 21644 43474 21700 43486
rect 20636 43426 20804 43428
rect 20636 43374 20638 43426
rect 20690 43374 20804 43426
rect 20636 43372 20804 43374
rect 21084 43428 21140 43438
rect 20636 42644 20692 43372
rect 21084 43334 21140 43372
rect 20636 42578 20692 42588
rect 20412 42130 20468 42140
rect 20636 41972 20692 41982
rect 21980 41972 22036 44380
rect 22092 44210 22148 44222
rect 22092 44158 22094 44210
rect 22146 44158 22148 44210
rect 22092 43428 22148 44158
rect 22652 44210 22708 44940
rect 23100 44434 23156 45164
rect 23660 44996 23716 45006
rect 23660 44902 23716 44940
rect 23100 44382 23102 44434
rect 23154 44382 23156 44434
rect 23100 44370 23156 44382
rect 22652 44158 22654 44210
rect 22706 44158 22708 44210
rect 22092 43362 22148 43372
rect 22428 43540 22484 43550
rect 20300 41970 21028 41972
rect 20300 41918 20638 41970
rect 20690 41918 21028 41970
rect 20300 41916 21028 41918
rect 20300 41074 20356 41916
rect 20636 41906 20692 41916
rect 20972 41860 21028 41916
rect 21980 41906 22036 41916
rect 21644 41860 21700 41870
rect 20972 41858 21364 41860
rect 20972 41806 20974 41858
rect 21026 41806 21364 41858
rect 20972 41804 21364 41806
rect 20972 41794 21028 41804
rect 20860 41748 20916 41758
rect 20300 41022 20302 41074
rect 20354 41022 20356 41074
rect 20300 41010 20356 41022
rect 20412 41186 20468 41198
rect 20412 41134 20414 41186
rect 20466 41134 20468 41186
rect 20412 40852 20468 41134
rect 20636 40964 20692 40974
rect 20692 40908 20804 40964
rect 20636 40898 20692 40908
rect 19836 40796 20100 40806
rect 20188 40796 20468 40852
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 19836 40730 20100 40740
rect 19740 40628 19796 40638
rect 19628 40626 19796 40628
rect 19628 40574 19742 40626
rect 19794 40574 19796 40626
rect 19628 40572 19796 40574
rect 19516 40348 19684 40404
rect 18956 39678 18958 39730
rect 19010 39678 19012 39730
rect 18956 39666 19012 39678
rect 19292 39676 19460 39732
rect 19516 40178 19572 40190
rect 19516 40126 19518 40178
rect 19570 40126 19572 40178
rect 18844 39508 18900 39518
rect 18844 39414 18900 39452
rect 19068 39508 19124 39518
rect 19068 39414 19124 39452
rect 18396 38612 18676 38668
rect 18732 38612 18900 38668
rect 17388 38162 17444 38612
rect 17388 38110 17390 38162
rect 17442 38110 17444 38162
rect 17388 38098 17444 38110
rect 17164 37986 17220 37996
rect 17500 37940 17556 37950
rect 17500 37846 17556 37884
rect 17948 37938 18004 38612
rect 18508 38276 18564 38286
rect 18396 38220 18508 38276
rect 17948 37886 17950 37938
rect 18002 37886 18004 37938
rect 17948 37874 18004 37886
rect 18060 37940 18116 37950
rect 18060 37846 18116 37884
rect 17724 37828 17780 37838
rect 17724 37734 17780 37772
rect 17276 37492 17332 37502
rect 17052 36372 17108 36382
rect 17052 36278 17108 36316
rect 17164 36260 17220 36270
rect 17164 36166 17220 36204
rect 17276 36036 17332 37436
rect 17612 37378 17668 37390
rect 17612 37326 17614 37378
rect 17666 37326 17668 37378
rect 17388 37268 17444 37278
rect 17388 37174 17444 37212
rect 16940 34290 16996 34300
rect 17052 35980 17332 36036
rect 17612 36036 17668 37326
rect 17724 37380 17780 37390
rect 17724 37286 17780 37324
rect 18284 37154 18340 37166
rect 18284 37102 18286 37154
rect 18338 37102 18340 37154
rect 18284 36596 18340 37102
rect 18284 36530 18340 36540
rect 18396 36484 18452 38220
rect 18508 38210 18564 38220
rect 18620 38162 18676 38612
rect 18620 38110 18622 38162
rect 18674 38110 18676 38162
rect 18620 38098 18676 38110
rect 18732 38500 18788 38510
rect 18508 37940 18564 37950
rect 18732 37940 18788 38444
rect 18508 37846 18564 37884
rect 18620 37938 18788 37940
rect 18620 37886 18734 37938
rect 18786 37886 18788 37938
rect 18620 37884 18788 37886
rect 18620 37380 18676 37884
rect 18732 37874 18788 37884
rect 18508 37324 18676 37380
rect 18732 37604 18788 37614
rect 18508 36708 18564 37324
rect 18620 37154 18676 37166
rect 18620 37102 18622 37154
rect 18674 37102 18676 37154
rect 18620 37042 18676 37102
rect 18620 36990 18622 37042
rect 18674 36990 18676 37042
rect 18620 36978 18676 36990
rect 18732 37156 18788 37548
rect 18508 36652 18676 36708
rect 18508 36484 18564 36494
rect 18396 36482 18564 36484
rect 18396 36430 18510 36482
rect 18562 36430 18564 36482
rect 18396 36428 18564 36430
rect 18508 36418 18564 36428
rect 16828 33294 16830 33346
rect 16882 33294 16884 33346
rect 16828 33236 16884 33294
rect 16828 33170 16884 33180
rect 16716 32734 16718 32786
rect 16770 32734 16772 32786
rect 16716 32722 16772 32734
rect 16828 32788 16884 32798
rect 16716 31778 16772 31790
rect 16716 31726 16718 31778
rect 16770 31726 16772 31778
rect 16716 31218 16772 31726
rect 16716 31166 16718 31218
rect 16770 31166 16772 31218
rect 16716 31154 16772 31166
rect 16604 30996 16660 31006
rect 16492 30994 16660 30996
rect 16492 30942 16606 30994
rect 16658 30942 16660 30994
rect 16492 30940 16660 30942
rect 16604 30930 16660 30940
rect 16044 30492 16436 30548
rect 16380 30322 16436 30492
rect 16380 30270 16382 30322
rect 16434 30270 16436 30322
rect 16380 30258 16436 30270
rect 15708 30158 15710 30210
rect 15762 30158 15764 30210
rect 15708 30146 15764 30158
rect 16268 30212 16324 30222
rect 16268 30118 16324 30156
rect 16604 30212 16660 30222
rect 16044 30098 16100 30110
rect 16492 30100 16548 30110
rect 16044 30046 16046 30098
rect 16098 30046 16100 30098
rect 15596 29988 15652 29998
rect 16044 29988 16100 30046
rect 15596 29986 16100 29988
rect 15596 29934 15598 29986
rect 15650 29934 16100 29986
rect 15596 29932 16100 29934
rect 16380 30098 16548 30100
rect 16380 30046 16494 30098
rect 16546 30046 16548 30098
rect 16380 30044 16548 30046
rect 15596 28868 15652 29932
rect 16380 29876 16436 30044
rect 16492 30034 16548 30044
rect 16604 29986 16660 30156
rect 16604 29934 16606 29986
rect 16658 29934 16660 29986
rect 16380 29820 16548 29876
rect 16492 29764 16548 29820
rect 16492 29698 16548 29708
rect 16380 29652 16436 29662
rect 16044 29540 16100 29550
rect 16044 29446 16100 29484
rect 16380 29538 16436 29596
rect 16380 29486 16382 29538
rect 16434 29486 16436 29538
rect 16380 29474 16436 29486
rect 15596 28802 15652 28812
rect 16268 29316 16324 29326
rect 15484 28588 15764 28644
rect 15708 27970 15764 28588
rect 16044 28642 16100 28654
rect 16044 28590 16046 28642
rect 16098 28590 16100 28642
rect 16044 28532 16100 28590
rect 16044 28466 16100 28476
rect 15708 27918 15710 27970
rect 15762 27918 15764 27970
rect 15708 27906 15764 27918
rect 15820 28084 15876 28094
rect 15372 27806 15374 27858
rect 15426 27806 15428 27858
rect 15372 27794 15428 27806
rect 15820 27636 15876 28028
rect 16044 27748 16100 27758
rect 16044 27654 16100 27692
rect 16156 27636 16212 27646
rect 15820 27634 15988 27636
rect 15820 27582 15822 27634
rect 15874 27582 15988 27634
rect 15820 27580 15988 27582
rect 15820 27570 15876 27580
rect 15036 27186 15316 27188
rect 15036 27134 15038 27186
rect 15090 27134 15316 27186
rect 15036 27132 15316 27134
rect 15708 27188 15764 27198
rect 15036 27122 15092 27132
rect 15372 27076 15428 27086
rect 15372 26982 15428 27020
rect 15708 26962 15764 27132
rect 15820 27076 15876 27086
rect 15820 26982 15876 27020
rect 15708 26910 15710 26962
rect 15762 26910 15764 26962
rect 15484 26852 15540 26862
rect 15148 26850 15540 26852
rect 15148 26798 15486 26850
rect 15538 26798 15540 26850
rect 15148 26796 15540 26798
rect 14476 25218 14532 25228
rect 14588 26740 14644 26750
rect 14476 23938 14532 23950
rect 14476 23886 14478 23938
rect 14530 23886 14532 23938
rect 14252 23826 14308 23838
rect 14252 23774 14254 23826
rect 14306 23774 14308 23826
rect 14252 23604 14308 23774
rect 14252 23538 14308 23548
rect 14364 23714 14420 23726
rect 14364 23662 14366 23714
rect 14418 23662 14420 23714
rect 14028 22978 14084 22988
rect 14140 23266 14196 23278
rect 14140 23214 14142 23266
rect 14194 23214 14196 23266
rect 14140 22708 14196 23214
rect 14140 22642 14196 22652
rect 14028 22372 14084 22382
rect 14028 22278 14084 22316
rect 13692 22258 13748 22270
rect 13692 22206 13694 22258
rect 13746 22206 13748 22258
rect 13692 22148 13748 22206
rect 13692 22082 13748 22092
rect 13804 22146 13860 22158
rect 13804 22094 13806 22146
rect 13858 22094 13860 22146
rect 13804 21700 13860 22094
rect 13804 21634 13860 21644
rect 13580 21186 13636 21196
rect 13244 21084 13412 21140
rect 13244 20804 13300 21084
rect 13580 21026 13636 21038
rect 13580 20974 13582 21026
rect 13634 20974 13636 21026
rect 13468 20804 13524 20814
rect 13244 20802 13524 20804
rect 13244 20750 13470 20802
rect 13522 20750 13524 20802
rect 13244 20748 13524 20750
rect 13468 20738 13524 20748
rect 13580 20132 13636 20974
rect 13916 20804 13972 20814
rect 13916 20710 13972 20748
rect 14140 20690 14196 20702
rect 14140 20638 14142 20690
rect 14194 20638 14196 20690
rect 13580 20066 13636 20076
rect 13692 20578 13748 20590
rect 13692 20526 13694 20578
rect 13746 20526 13748 20578
rect 13692 20018 13748 20526
rect 14140 20580 14196 20638
rect 14140 20514 14196 20524
rect 14364 20356 14420 23662
rect 14476 23716 14532 23886
rect 14476 23650 14532 23660
rect 14476 23154 14532 23166
rect 14476 23102 14478 23154
rect 14530 23102 14532 23154
rect 14476 22820 14532 23102
rect 14476 22754 14532 22764
rect 14476 22484 14532 22494
rect 14588 22484 14644 26684
rect 14812 26740 14868 26750
rect 14812 24836 14868 26684
rect 15148 26628 15204 26796
rect 15484 26786 15540 26796
rect 15708 26740 15764 26910
rect 15708 26674 15764 26684
rect 15372 26628 15428 26638
rect 14924 26572 15204 26628
rect 15260 26572 15372 26628
rect 14924 26290 14980 26572
rect 15260 26404 15316 26572
rect 14924 26238 14926 26290
rect 14978 26238 14980 26290
rect 14924 26226 14980 26238
rect 15148 26348 15316 26404
rect 15148 26290 15204 26348
rect 15148 26238 15150 26290
rect 15202 26238 15204 26290
rect 15148 26226 15204 26238
rect 15260 26178 15316 26190
rect 15260 26126 15262 26178
rect 15314 26126 15316 26178
rect 15260 25620 15316 26126
rect 15260 25554 15316 25564
rect 15036 24836 15092 24846
rect 14812 24834 15092 24836
rect 14812 24782 15038 24834
rect 15090 24782 15092 24834
rect 14812 24780 15092 24782
rect 15036 24770 15092 24780
rect 14924 24276 14980 24286
rect 15372 24276 15428 26572
rect 15820 26516 15876 26526
rect 15484 26514 15876 26516
rect 15484 26462 15822 26514
rect 15874 26462 15876 26514
rect 15484 26460 15876 26462
rect 15484 26290 15540 26460
rect 15820 26450 15876 26460
rect 15484 26238 15486 26290
rect 15538 26238 15540 26290
rect 15484 26226 15540 26238
rect 15596 26290 15652 26302
rect 15596 26238 15598 26290
rect 15650 26238 15652 26290
rect 15596 26180 15652 26238
rect 15596 26114 15652 26124
rect 15932 25956 15988 27580
rect 16156 27542 16212 27580
rect 16268 27412 16324 29260
rect 16604 29316 16660 29934
rect 16828 29538 16884 32732
rect 16828 29486 16830 29538
rect 16882 29486 16884 29538
rect 16828 29474 16884 29486
rect 16940 32676 16996 32686
rect 16604 28980 16660 29260
rect 16716 29204 16772 29214
rect 16716 29110 16772 29148
rect 16940 28980 16996 32620
rect 17052 30772 17108 35980
rect 17612 35970 17668 35980
rect 18284 36036 18340 36046
rect 17612 35810 17668 35822
rect 17612 35758 17614 35810
rect 17666 35758 17668 35810
rect 17612 35308 17668 35758
rect 17724 35812 17780 35822
rect 17724 35718 17780 35756
rect 18060 35812 18116 35822
rect 17276 35252 17668 35308
rect 17836 35700 17892 35710
rect 17276 35026 17332 35252
rect 17276 34974 17278 35026
rect 17330 34974 17332 35026
rect 17276 34962 17332 34974
rect 17724 35028 17780 35038
rect 17724 34934 17780 34972
rect 17612 34916 17668 34926
rect 17388 34020 17444 34030
rect 17388 33684 17444 33964
rect 17388 33618 17444 33628
rect 17500 33796 17556 33806
rect 17500 32674 17556 33740
rect 17500 32622 17502 32674
rect 17554 32622 17556 32674
rect 17500 32610 17556 32622
rect 17164 32452 17220 32462
rect 17164 31778 17220 32396
rect 17388 32340 17444 32350
rect 17388 32246 17444 32284
rect 17164 31726 17166 31778
rect 17218 31726 17220 31778
rect 17164 31714 17220 31726
rect 17500 32116 17556 32126
rect 17052 30716 17444 30772
rect 17164 30212 17220 30222
rect 17164 30118 17220 30156
rect 16044 27356 16324 27412
rect 16492 28924 16660 28980
rect 16716 28924 16996 28980
rect 16492 28196 16548 28924
rect 16716 28530 16772 28924
rect 16940 28868 16996 28924
rect 16940 28802 16996 28812
rect 17052 29652 17108 29662
rect 17052 28644 17108 29596
rect 16716 28478 16718 28530
rect 16770 28478 16772 28530
rect 16716 28466 16772 28478
rect 16828 28642 17108 28644
rect 16828 28590 17054 28642
rect 17106 28590 17108 28642
rect 16828 28588 17108 28590
rect 17276 29540 17332 29550
rect 17276 28644 17332 29484
rect 17388 29426 17444 30716
rect 17500 30322 17556 32060
rect 17500 30270 17502 30322
rect 17554 30270 17556 30322
rect 17500 30258 17556 30270
rect 17388 29374 17390 29426
rect 17442 29374 17444 29426
rect 17388 29362 17444 29374
rect 17388 28644 17444 28654
rect 17276 28642 17444 28644
rect 17276 28590 17390 28642
rect 17442 28590 17444 28642
rect 17276 28588 17444 28590
rect 16044 26964 16100 27356
rect 16492 27300 16548 28140
rect 16828 28084 16884 28588
rect 17052 28308 17108 28588
rect 17388 28578 17444 28588
rect 17052 28252 17556 28308
rect 16604 28028 16884 28084
rect 17276 28084 17332 28094
rect 16604 27970 16660 28028
rect 16604 27918 16606 27970
rect 16658 27918 16660 27970
rect 16604 27906 16660 27918
rect 16828 27860 16884 27870
rect 16044 26402 16100 26908
rect 16044 26350 16046 26402
rect 16098 26350 16100 26402
rect 16044 26338 16100 26350
rect 16268 27244 16548 27300
rect 16716 27634 16772 27646
rect 16716 27582 16718 27634
rect 16770 27582 16772 27634
rect 16716 27524 16772 27582
rect 16156 26292 16212 26302
rect 16156 26198 16212 26236
rect 15596 25900 15988 25956
rect 15484 24948 15540 24958
rect 15596 24948 15652 25900
rect 16268 25620 16324 27244
rect 16492 26962 16548 26974
rect 16492 26910 16494 26962
rect 16546 26910 16548 26962
rect 16492 26740 16548 26910
rect 16716 26740 16772 27468
rect 16828 26962 16884 27804
rect 16828 26910 16830 26962
rect 16882 26910 16884 26962
rect 16828 26898 16884 26910
rect 17164 26962 17220 26974
rect 17164 26910 17166 26962
rect 17218 26910 17220 26962
rect 17164 26740 17220 26910
rect 16716 26684 16884 26740
rect 16492 26516 16548 26684
rect 16492 26450 16548 26460
rect 16828 26514 16884 26684
rect 17164 26674 17220 26684
rect 16828 26462 16830 26514
rect 16882 26462 16884 26514
rect 16828 26450 16884 26462
rect 16716 26292 16772 26302
rect 15932 25564 16324 25620
rect 16380 25620 16436 25630
rect 15484 24946 15652 24948
rect 15484 24894 15486 24946
rect 15538 24894 15652 24946
rect 15484 24892 15652 24894
rect 15708 25508 15764 25518
rect 15484 24882 15540 24892
rect 15708 24836 15764 25452
rect 15708 24388 15764 24780
rect 14980 24220 15316 24276
rect 14924 24210 14980 24220
rect 15260 23938 15316 24220
rect 15260 23886 15262 23938
rect 15314 23886 15316 23938
rect 15260 23874 15316 23886
rect 15372 23828 15428 24220
rect 15372 23762 15428 23772
rect 15596 24332 15764 24388
rect 15820 25396 15876 25406
rect 15036 23268 15092 23278
rect 14924 23156 14980 23166
rect 14924 23062 14980 23100
rect 15036 22820 15092 23212
rect 15596 22930 15652 24332
rect 15708 23828 15764 23838
rect 15708 23378 15764 23772
rect 15708 23326 15710 23378
rect 15762 23326 15764 23378
rect 15708 23314 15764 23326
rect 15596 22878 15598 22930
rect 15650 22878 15652 22930
rect 15596 22866 15652 22878
rect 14924 22764 15092 22820
rect 15148 22820 15204 22830
rect 14476 22482 14868 22484
rect 14476 22430 14478 22482
rect 14530 22430 14868 22482
rect 14476 22428 14868 22430
rect 14476 22418 14532 22428
rect 14812 22370 14868 22428
rect 14812 22318 14814 22370
rect 14866 22318 14868 22370
rect 14476 21924 14532 21934
rect 14476 20802 14532 21868
rect 14812 21588 14868 22318
rect 14812 21522 14868 21532
rect 14476 20750 14478 20802
rect 14530 20750 14532 20802
rect 14476 20738 14532 20750
rect 14700 21476 14756 21486
rect 14700 20802 14756 21420
rect 14924 21028 14980 22764
rect 15148 22036 15204 22764
rect 15036 21980 15204 22036
rect 15372 22596 15428 22606
rect 15036 21474 15092 21980
rect 15036 21422 15038 21474
rect 15090 21422 15092 21474
rect 15036 21410 15092 21422
rect 15036 21028 15092 21038
rect 14924 21026 15092 21028
rect 14924 20974 15038 21026
rect 15090 20974 15092 21026
rect 14924 20972 15092 20974
rect 15036 20962 15092 20972
rect 15372 20916 15428 22540
rect 15596 22258 15652 22270
rect 15596 22206 15598 22258
rect 15650 22206 15652 22258
rect 15596 22148 15652 22206
rect 15596 22082 15652 22092
rect 15484 21588 15540 21598
rect 15484 21494 15540 21532
rect 15372 20860 15652 20916
rect 14700 20750 14702 20802
rect 14754 20750 14756 20802
rect 14700 20692 14756 20750
rect 14700 20626 14756 20636
rect 15372 20692 15428 20702
rect 15484 20692 15540 20702
rect 15372 20690 15540 20692
rect 15372 20638 15374 20690
rect 15426 20638 15486 20690
rect 15538 20638 15540 20690
rect 15372 20636 15540 20638
rect 14140 20300 14420 20356
rect 14588 20580 14644 20590
rect 13692 19966 13694 20018
rect 13746 19966 13748 20018
rect 13356 19796 13412 19806
rect 13356 19702 13412 19740
rect 13692 19236 13748 19966
rect 13916 20020 13972 20030
rect 13916 19926 13972 19964
rect 14028 20018 14084 20030
rect 14028 19966 14030 20018
rect 14082 19966 14084 20018
rect 14028 19908 14084 19966
rect 13916 19236 13972 19246
rect 14028 19236 14084 19852
rect 13692 19122 13748 19180
rect 13692 19070 13694 19122
rect 13746 19070 13748 19122
rect 13468 19012 13524 19022
rect 13692 19012 13748 19070
rect 13524 18956 13748 19012
rect 13804 19234 14084 19236
rect 13804 19182 13918 19234
rect 13970 19182 14084 19234
rect 13804 19180 14084 19182
rect 14140 19234 14196 20300
rect 14476 19794 14532 19806
rect 14476 19742 14478 19794
rect 14530 19742 14532 19794
rect 14252 19684 14308 19694
rect 14252 19458 14308 19628
rect 14252 19406 14254 19458
rect 14306 19406 14308 19458
rect 14252 19394 14308 19406
rect 14476 19460 14532 19742
rect 14476 19394 14532 19404
rect 14140 19182 14142 19234
rect 14194 19182 14196 19234
rect 13468 18946 13524 18956
rect 13804 18900 13860 19180
rect 13916 19170 13972 19180
rect 14140 19170 14196 19182
rect 14364 19236 14420 19246
rect 14588 19236 14644 20524
rect 14924 20578 14980 20590
rect 15260 20580 15316 20590
rect 14924 20526 14926 20578
rect 14978 20526 14980 20578
rect 14924 19460 14980 20526
rect 15148 20578 15316 20580
rect 15148 20526 15262 20578
rect 15314 20526 15316 20578
rect 15148 20524 15316 20526
rect 15148 20018 15204 20524
rect 15260 20514 15316 20524
rect 15372 20132 15428 20636
rect 15484 20626 15540 20636
rect 15148 19966 15150 20018
rect 15202 19966 15204 20018
rect 15148 19954 15204 19966
rect 15260 20076 15428 20132
rect 15484 20468 15540 20478
rect 15260 19796 15316 20076
rect 15372 19908 15428 19918
rect 15372 19814 15428 19852
rect 15148 19740 15316 19796
rect 14924 19404 15092 19460
rect 14364 19234 14644 19236
rect 14364 19182 14366 19234
rect 14418 19182 14644 19234
rect 14364 19180 14644 19182
rect 14700 19234 14756 19246
rect 14700 19182 14702 19234
rect 14754 19182 14756 19234
rect 14364 19170 14420 19180
rect 13580 18844 13860 18900
rect 12908 18562 13188 18564
rect 12908 18510 12910 18562
rect 12962 18510 13188 18562
rect 12908 18508 13188 18510
rect 13244 18564 13300 18574
rect 12572 18452 12628 18462
rect 12572 17892 12628 18396
rect 12572 17826 12628 17836
rect 12684 18004 12740 18014
rect 12684 17666 12740 17948
rect 12684 17614 12686 17666
rect 12738 17614 12740 17666
rect 12684 17602 12740 17614
rect 12908 17554 12964 18508
rect 13244 18470 13300 18508
rect 13468 18562 13524 18574
rect 13468 18510 13470 18562
rect 13522 18510 13524 18562
rect 12908 17502 12910 17554
rect 12962 17502 12964 17554
rect 12572 17442 12628 17454
rect 12572 17390 12574 17442
rect 12626 17390 12628 17442
rect 12572 16324 12628 17390
rect 12572 16258 12628 16268
rect 12684 17332 12740 17342
rect 12684 16098 12740 17276
rect 12684 16046 12686 16098
rect 12738 16046 12740 16098
rect 12684 16034 12740 16046
rect 12796 16436 12852 16446
rect 12572 15876 12628 15886
rect 12572 15782 12628 15820
rect 12796 15652 12852 16380
rect 12908 15988 12964 17502
rect 13468 16884 13524 18510
rect 13580 18338 13636 18844
rect 14700 18788 14756 19182
rect 14924 19236 14980 19246
rect 14924 19142 14980 19180
rect 14476 18732 14756 18788
rect 13580 18286 13582 18338
rect 13634 18286 13636 18338
rect 13580 18274 13636 18286
rect 13692 18450 13748 18462
rect 13692 18398 13694 18450
rect 13746 18398 13748 18450
rect 13580 18004 13636 18014
rect 13580 17778 13636 17948
rect 13580 17726 13582 17778
rect 13634 17726 13636 17778
rect 13580 17714 13636 17726
rect 13468 16818 13524 16828
rect 13692 15988 13748 18398
rect 13804 18228 13860 18238
rect 13804 16994 13860 18172
rect 14028 17668 14084 17678
rect 14028 17574 14084 17612
rect 14476 17332 14532 18732
rect 14588 18562 14644 18574
rect 14588 18510 14590 18562
rect 14642 18510 14644 18562
rect 14588 18452 14644 18510
rect 14588 18386 14644 18396
rect 14700 18338 14756 18350
rect 14700 18286 14702 18338
rect 14754 18286 14756 18338
rect 14700 17778 14756 18286
rect 14812 18228 14868 18238
rect 14812 18134 14868 18172
rect 14700 17726 14702 17778
rect 14754 17726 14756 17778
rect 14700 17714 14756 17726
rect 14476 17266 14532 17276
rect 14588 17668 14644 17678
rect 14476 17108 14532 17118
rect 14476 17014 14532 17052
rect 13804 16942 13806 16994
rect 13858 16942 13860 16994
rect 13804 16884 13860 16942
rect 13804 16818 13860 16828
rect 14140 16882 14196 16894
rect 14140 16830 14142 16882
rect 14194 16830 14196 16882
rect 14140 16660 14196 16830
rect 14140 16594 14196 16604
rect 14476 16324 14532 16334
rect 12908 15986 13188 15988
rect 12908 15934 12910 15986
rect 12962 15934 13188 15986
rect 12908 15932 13188 15934
rect 12908 15922 12964 15932
rect 12796 15596 13076 15652
rect 12348 15260 12516 15316
rect 12236 15148 12292 15260
rect 12236 15092 12404 15148
rect 12236 14530 12292 14542
rect 12236 14478 12238 14530
rect 12290 14478 12292 14530
rect 12236 13860 12292 14478
rect 12236 13746 12292 13804
rect 12236 13694 12238 13746
rect 12290 13694 12292 13746
rect 12236 13682 12292 13694
rect 12012 13634 12180 13636
rect 12012 13582 12014 13634
rect 12066 13582 12180 13634
rect 12012 13580 12180 13582
rect 12012 13076 12068 13580
rect 12012 13010 12068 13020
rect 11116 11732 11396 11788
rect 12124 12066 12180 12078
rect 12124 12014 12126 12066
rect 12178 12014 12180 12066
rect 11004 11620 11060 11630
rect 11004 11526 11060 11564
rect 10780 10658 10836 10668
rect 10892 10612 10948 10622
rect 10892 10518 10948 10556
rect 10780 10500 10836 10510
rect 10668 10444 10780 10500
rect 10780 10406 10836 10444
rect 10332 9998 10334 10050
rect 10386 9998 10388 10050
rect 10332 9986 10388 9998
rect 10444 10386 10500 10398
rect 10444 10334 10446 10386
rect 10498 10334 10500 10386
rect 10444 10050 10500 10334
rect 10444 9998 10446 10050
rect 10498 9998 10500 10050
rect 10444 9986 10500 9998
rect 10556 10388 10612 10398
rect 10444 9042 10500 9054
rect 10444 8990 10446 9042
rect 10498 8990 10500 9042
rect 10444 8932 10500 8990
rect 10444 8866 10500 8876
rect 10332 8258 10388 8270
rect 10332 8206 10334 8258
rect 10386 8206 10388 8258
rect 10332 6916 10388 8206
rect 10332 6850 10388 6860
rect 10220 6692 10276 6702
rect 10108 6690 10276 6692
rect 10108 6638 10222 6690
rect 10274 6638 10276 6690
rect 10108 6636 10276 6638
rect 9772 6356 9828 6366
rect 9772 6130 9828 6300
rect 9772 6078 9774 6130
rect 9826 6078 9828 6130
rect 9772 4564 9828 6078
rect 10108 6132 10164 6142
rect 10220 6132 10276 6636
rect 10164 6076 10276 6132
rect 10108 6066 10164 6076
rect 9996 5908 10052 5918
rect 9996 5814 10052 5852
rect 10444 5908 10500 5918
rect 10444 5814 10500 5852
rect 10332 5236 10388 5246
rect 10556 5236 10612 10332
rect 11116 10388 11172 11732
rect 11676 11620 11732 11630
rect 11228 11396 11284 11406
rect 11284 11340 11620 11396
rect 11228 11302 11284 11340
rect 11564 10500 11620 11340
rect 11676 11394 11732 11564
rect 12124 11396 12180 12014
rect 11676 11342 11678 11394
rect 11730 11342 11732 11394
rect 11676 11330 11732 11342
rect 11900 11340 12180 11396
rect 12236 11396 12292 11406
rect 11788 11172 11844 11182
rect 11900 11172 11956 11340
rect 12236 11302 12292 11340
rect 11788 11170 11956 11172
rect 11788 11118 11790 11170
rect 11842 11118 11956 11170
rect 11788 11116 11956 11118
rect 12012 11172 12068 11182
rect 11676 10500 11732 10510
rect 11564 10498 11732 10500
rect 11564 10446 11678 10498
rect 11730 10446 11732 10498
rect 11564 10444 11732 10446
rect 11676 10434 11732 10444
rect 11116 10322 11172 10332
rect 11788 10276 11844 11116
rect 12012 11078 12068 11116
rect 11788 10220 12180 10276
rect 11900 9940 11956 9950
rect 11788 9884 11900 9940
rect 10668 9828 10724 9838
rect 10668 9734 10724 9772
rect 10892 9826 10948 9838
rect 10892 9774 10894 9826
rect 10946 9774 10948 9826
rect 10668 9154 10724 9166
rect 10668 9102 10670 9154
rect 10722 9102 10724 9154
rect 10668 9044 10724 9102
rect 10668 8978 10724 8988
rect 10892 9044 10948 9774
rect 11452 9828 11508 9838
rect 11004 9716 11060 9726
rect 11340 9716 11396 9726
rect 11004 9714 11396 9716
rect 11004 9662 11006 9714
rect 11058 9662 11342 9714
rect 11394 9662 11396 9714
rect 11004 9660 11396 9662
rect 11004 9650 11060 9660
rect 11340 9650 11396 9660
rect 11452 9156 11508 9772
rect 11676 9716 11732 9726
rect 11676 9622 11732 9660
rect 10892 8978 10948 8988
rect 11340 9100 11508 9156
rect 10780 8484 10836 8494
rect 10780 8390 10836 8428
rect 11340 8372 11396 9100
rect 11452 8932 11508 8942
rect 11676 8932 11732 8942
rect 11788 8932 11844 9884
rect 11900 9874 11956 9884
rect 12124 9604 12180 10220
rect 12236 9604 12292 9614
rect 12124 9602 12292 9604
rect 12124 9550 12238 9602
rect 12290 9550 12292 9602
rect 12124 9548 12292 9550
rect 12236 9492 12292 9548
rect 12236 9426 12292 9436
rect 11452 8930 11620 8932
rect 11452 8878 11454 8930
rect 11506 8878 11620 8930
rect 11452 8876 11620 8878
rect 11452 8866 11508 8876
rect 11452 8372 11508 8382
rect 11340 8370 11508 8372
rect 11340 8318 11454 8370
rect 11506 8318 11508 8370
rect 11340 8316 11508 8318
rect 10780 8260 10836 8270
rect 10780 8166 10836 8204
rect 11452 7700 11508 8316
rect 11452 7634 11508 7644
rect 11564 7588 11620 8876
rect 11676 8930 11844 8932
rect 11676 8878 11678 8930
rect 11730 8878 11844 8930
rect 11676 8876 11844 8878
rect 11900 8932 11956 8942
rect 12348 8932 12404 15092
rect 12460 11508 12516 15260
rect 12572 15302 12740 15316
rect 12572 15250 12574 15302
rect 12626 15260 12740 15302
rect 12626 15250 12628 15260
rect 12572 15238 12628 15250
rect 12684 15204 12740 15260
rect 12684 15138 12740 15148
rect 12908 14644 12964 14654
rect 12908 14530 12964 14588
rect 12908 14478 12910 14530
rect 12962 14478 12964 14530
rect 12908 14466 12964 14478
rect 12684 14308 12740 14318
rect 12460 11442 12516 11452
rect 12572 14306 12740 14308
rect 12572 14254 12686 14306
rect 12738 14254 12740 14306
rect 12572 14252 12740 14254
rect 12460 11172 12516 11182
rect 12460 11078 12516 11116
rect 12572 9940 12628 14252
rect 12684 14242 12740 14252
rect 12796 14308 12852 14318
rect 12796 14214 12852 14252
rect 12796 13972 12852 13982
rect 12796 13878 12852 13916
rect 12908 13972 12964 13982
rect 13020 13972 13076 15596
rect 13132 15304 13188 15932
rect 13692 15922 13748 15932
rect 14028 16098 14084 16110
rect 14028 16046 14030 16098
rect 14082 16046 14084 16098
rect 13244 15876 13300 15886
rect 13244 15426 13300 15820
rect 14028 15876 14084 16046
rect 14028 15810 14084 15820
rect 13244 15374 13246 15426
rect 13298 15374 13300 15426
rect 13244 15362 13300 15374
rect 13132 15248 13300 15304
rect 12908 13970 13076 13972
rect 12908 13918 12910 13970
rect 12962 13918 13076 13970
rect 12908 13916 13076 13918
rect 12908 13906 12964 13916
rect 12684 13748 12740 13758
rect 12684 13654 12740 13692
rect 13020 13074 13076 13916
rect 13020 13022 13022 13074
rect 13074 13022 13076 13074
rect 13020 13010 13076 13022
rect 13132 13300 13188 13310
rect 13132 12404 13188 13244
rect 12908 12402 13188 12404
rect 12908 12350 13134 12402
rect 13186 12350 13188 12402
rect 12908 12348 13188 12350
rect 12796 11506 12852 11518
rect 12796 11454 12798 11506
rect 12850 11454 12852 11506
rect 12796 11396 12852 11454
rect 12796 11330 12852 11340
rect 12908 11394 12964 12348
rect 13132 12338 13188 12348
rect 13244 11788 13300 15248
rect 13468 14644 13524 14654
rect 13468 13970 13524 14588
rect 13468 13918 13470 13970
rect 13522 13918 13524 13970
rect 13468 13906 13524 13918
rect 13916 14642 13972 14654
rect 13916 14590 13918 14642
rect 13970 14590 13972 14642
rect 13804 13748 13860 13758
rect 13916 13748 13972 14590
rect 14476 13858 14532 16268
rect 14588 16210 14644 17612
rect 14924 16996 14980 17006
rect 14924 16902 14980 16940
rect 14588 16158 14590 16210
rect 14642 16158 14644 16210
rect 14588 15204 14644 16158
rect 14588 15138 14644 15148
rect 14476 13806 14478 13858
rect 14530 13806 14532 13858
rect 14476 13794 14532 13806
rect 13804 13746 14420 13748
rect 13804 13694 13806 13746
rect 13858 13694 14420 13746
rect 13804 13692 14420 13694
rect 13804 13682 13860 13692
rect 13692 13186 13748 13198
rect 13692 13134 13694 13186
rect 13746 13134 13748 13186
rect 13468 13076 13524 13086
rect 13468 12982 13524 13020
rect 13244 11732 13636 11788
rect 12908 11342 12910 11394
rect 12962 11342 12964 11394
rect 12908 11330 12964 11342
rect 13020 11508 13076 11518
rect 12684 11284 12740 11294
rect 12684 11190 12740 11228
rect 12908 9940 12964 9950
rect 12572 9884 12852 9940
rect 11956 8876 12404 8932
rect 12572 9714 12628 9726
rect 12572 9662 12574 9714
rect 12626 9662 12628 9714
rect 12572 9492 12628 9662
rect 12684 9604 12740 9614
rect 12684 9510 12740 9548
rect 11676 8866 11732 8876
rect 11900 8036 11956 8876
rect 12572 8820 12628 9436
rect 12572 8754 12628 8764
rect 12236 8146 12292 8158
rect 12236 8094 12238 8146
rect 12290 8094 12292 8146
rect 11900 7970 11956 7980
rect 12012 8034 12068 8046
rect 12012 7982 12014 8034
rect 12066 7982 12068 8034
rect 11564 7522 11620 7532
rect 10668 7364 10724 7374
rect 10668 7362 11620 7364
rect 10668 7310 10670 7362
rect 10722 7310 11620 7362
rect 10668 7308 11620 7310
rect 10668 7298 10724 7308
rect 11564 6914 11620 7308
rect 11564 6862 11566 6914
rect 11618 6862 11620 6914
rect 11564 6850 11620 6862
rect 11676 6916 11732 6926
rect 10668 6804 10724 6814
rect 10668 6690 10724 6748
rect 10668 6638 10670 6690
rect 10722 6638 10724 6690
rect 10668 6626 10724 6638
rect 11452 6804 11508 6814
rect 11004 6580 11060 6590
rect 11004 6486 11060 6524
rect 11116 6468 11172 6478
rect 11116 6466 11284 6468
rect 11116 6414 11118 6466
rect 11170 6414 11284 6466
rect 11116 6412 11284 6414
rect 11116 6402 11172 6412
rect 10780 6020 10836 6030
rect 10780 5926 10836 5964
rect 11228 6020 11284 6412
rect 11228 5954 11284 5964
rect 11340 6466 11396 6478
rect 11340 6414 11342 6466
rect 11394 6414 11396 6466
rect 11116 5908 11172 5918
rect 11116 5814 11172 5852
rect 11004 5348 11060 5358
rect 11060 5292 11172 5348
rect 11004 5282 11060 5292
rect 10332 5234 10612 5236
rect 10332 5182 10334 5234
rect 10386 5182 10612 5234
rect 10332 5180 10612 5182
rect 10332 5170 10388 5180
rect 9772 4498 9828 4508
rect 9660 4286 9662 4338
rect 9714 4286 9716 4338
rect 9660 4274 9716 4286
rect 8988 4228 9044 4238
rect 8988 4134 9044 4172
rect 9436 4116 9492 4126
rect 8764 3390 8766 3442
rect 8818 3390 8820 3442
rect 8764 3378 8820 3390
rect 9324 3780 9380 3790
rect 9324 3442 9380 3724
rect 9324 3390 9326 3442
rect 9378 3390 9380 3442
rect 9324 3378 9380 3390
rect 9436 800 9492 4060
rect 9548 3892 9604 3902
rect 9548 3554 9604 3836
rect 9548 3502 9550 3554
rect 9602 3502 9604 3554
rect 9548 3490 9604 3502
rect 10108 3668 10164 3678
rect 10108 800 10164 3612
rect 10444 3554 10500 5180
rect 10556 5124 10612 5180
rect 10668 5124 10724 5134
rect 10556 5122 10724 5124
rect 10556 5070 10670 5122
rect 10722 5070 10724 5122
rect 10556 5068 10724 5070
rect 10668 5058 10724 5068
rect 11116 5122 11172 5292
rect 11116 5070 11118 5122
rect 11170 5070 11172 5122
rect 11116 5058 11172 5070
rect 11340 5122 11396 6414
rect 11452 6468 11508 6748
rect 11676 6802 11732 6860
rect 11676 6750 11678 6802
rect 11730 6750 11732 6802
rect 11676 6738 11732 6750
rect 11452 6412 11620 6468
rect 11452 6244 11508 6254
rect 11452 6130 11508 6188
rect 11452 6078 11454 6130
rect 11506 6078 11508 6130
rect 11452 6066 11508 6078
rect 11340 5070 11342 5122
rect 11394 5070 11396 5122
rect 11340 5058 11396 5070
rect 10892 5012 10948 5022
rect 10892 4918 10948 4956
rect 10780 4898 10836 4910
rect 10780 4846 10782 4898
rect 10834 4846 10836 4898
rect 10780 4452 10836 4846
rect 11564 4788 11620 6412
rect 12012 6132 12068 7982
rect 12124 6916 12180 6926
rect 12124 6802 12180 6860
rect 12124 6750 12126 6802
rect 12178 6750 12180 6802
rect 12124 6738 12180 6750
rect 12236 6132 12292 8094
rect 12348 8034 12404 8046
rect 12348 7982 12350 8034
rect 12402 7982 12404 8034
rect 12348 6916 12404 7982
rect 12796 7924 12852 9884
rect 12908 9826 12964 9884
rect 12908 9774 12910 9826
rect 12962 9774 12964 9826
rect 12908 9762 12964 9774
rect 13020 8596 13076 11452
rect 13468 11396 13524 11406
rect 13468 11302 13524 11340
rect 13580 11284 13636 11732
rect 13692 11732 13748 13134
rect 14364 13076 14420 13692
rect 14364 13020 14868 13076
rect 14364 12850 14420 12862
rect 14364 12798 14366 12850
rect 14418 12798 14420 12850
rect 14028 12740 14084 12750
rect 14028 12646 14084 12684
rect 14028 12068 14084 12078
rect 14364 12068 14420 12798
rect 14476 12852 14532 12862
rect 14476 12758 14532 12796
rect 14476 12404 14532 12414
rect 14588 12404 14644 13020
rect 14812 12962 14868 13020
rect 14812 12910 14814 12962
rect 14866 12910 14868 12962
rect 14812 12898 14868 12910
rect 15036 12852 15092 19404
rect 15148 16884 15204 19740
rect 15260 19460 15316 19470
rect 15484 19460 15540 20412
rect 15260 19458 15540 19460
rect 15260 19406 15262 19458
rect 15314 19406 15540 19458
rect 15260 19404 15540 19406
rect 15260 19394 15316 19404
rect 15596 19012 15652 20860
rect 15820 20692 15876 25340
rect 15932 21812 15988 25564
rect 16380 25526 16436 25564
rect 16716 25508 16772 26236
rect 17276 26068 17332 28028
rect 17500 28082 17556 28252
rect 17500 28030 17502 28082
rect 17554 28030 17556 28082
rect 17276 26002 17332 26012
rect 17388 26964 17444 26974
rect 16716 25442 16772 25452
rect 17052 25506 17108 25518
rect 17052 25454 17054 25506
rect 17106 25454 17108 25506
rect 16940 25396 16996 25406
rect 16828 25340 16940 25396
rect 16716 25284 16772 25294
rect 16716 24946 16772 25228
rect 16716 24894 16718 24946
rect 16770 24894 16772 24946
rect 16716 24882 16772 24894
rect 16156 24836 16212 24846
rect 16156 24742 16212 24780
rect 16044 24722 16100 24734
rect 16044 24670 16046 24722
rect 16098 24670 16100 24722
rect 16044 24164 16100 24670
rect 16380 24722 16436 24734
rect 16380 24670 16382 24722
rect 16434 24670 16436 24722
rect 16044 24108 16324 24164
rect 16044 23938 16100 23950
rect 16044 23886 16046 23938
rect 16098 23886 16100 23938
rect 16044 23828 16100 23886
rect 16044 22932 16100 23772
rect 16156 23826 16212 23838
rect 16156 23774 16158 23826
rect 16210 23774 16212 23826
rect 16156 23268 16212 23774
rect 16268 23548 16324 24108
rect 16380 23940 16436 24670
rect 16604 24724 16660 24734
rect 16828 24724 16884 25340
rect 16940 25330 16996 25340
rect 17052 25284 17108 25454
rect 17052 25218 17108 25228
rect 17276 25508 17332 25518
rect 17276 25060 17332 25452
rect 17276 24994 17332 25004
rect 16604 24722 16884 24724
rect 16604 24670 16606 24722
rect 16658 24670 16884 24722
rect 16604 24668 16884 24670
rect 16940 24724 16996 24734
rect 17388 24724 17444 26908
rect 17500 26962 17556 28030
rect 17500 26910 17502 26962
rect 17554 26910 17556 26962
rect 17500 26898 17556 26910
rect 17612 26404 17668 34860
rect 17724 33458 17780 33470
rect 17724 33406 17726 33458
rect 17778 33406 17780 33458
rect 17724 31666 17780 33406
rect 17724 31614 17726 31666
rect 17778 31614 17780 31666
rect 17724 31602 17780 31614
rect 17724 31220 17780 31230
rect 17836 31220 17892 35644
rect 17948 35698 18004 35710
rect 17948 35646 17950 35698
rect 18002 35646 18004 35698
rect 17948 35140 18004 35646
rect 18060 35252 18116 35756
rect 18284 35698 18340 35980
rect 18284 35646 18286 35698
rect 18338 35646 18340 35698
rect 18284 35588 18340 35646
rect 18284 35522 18340 35532
rect 18060 35196 18228 35252
rect 17948 35074 18004 35084
rect 17948 34914 18004 34926
rect 17948 34862 17950 34914
rect 18002 34862 18004 34914
rect 17948 34804 18004 34862
rect 17948 34738 18004 34748
rect 17948 34132 18004 34142
rect 17948 34038 18004 34076
rect 17724 31218 17892 31220
rect 17724 31166 17726 31218
rect 17778 31166 17892 31218
rect 17724 31164 17892 31166
rect 17724 31154 17780 31164
rect 17836 30996 17892 31164
rect 18060 32450 18116 32462
rect 18060 32398 18062 32450
rect 18114 32398 18116 32450
rect 17836 30930 17892 30940
rect 17948 30994 18004 31006
rect 17948 30942 17950 30994
rect 18002 30942 18004 30994
rect 17836 29876 17892 29886
rect 17724 28756 17780 28766
rect 17724 27972 17780 28700
rect 17836 28754 17892 29820
rect 17948 29428 18004 30942
rect 18060 30212 18116 32398
rect 18060 30146 18116 30156
rect 18172 32340 18228 35196
rect 18508 35140 18564 35150
rect 18508 34914 18564 35084
rect 18508 34862 18510 34914
rect 18562 34862 18564 34914
rect 18508 34850 18564 34862
rect 18508 34692 18564 34702
rect 18508 33572 18564 34636
rect 18396 33516 18564 33572
rect 18396 33124 18452 33516
rect 18508 33348 18564 33358
rect 18508 33254 18564 33292
rect 18396 33068 18564 33124
rect 18396 32450 18452 32462
rect 18396 32398 18398 32450
rect 18450 32398 18452 32450
rect 18396 32340 18452 32398
rect 18172 32284 18452 32340
rect 18060 29986 18116 29998
rect 18060 29934 18062 29986
rect 18114 29934 18116 29986
rect 18060 29652 18116 29934
rect 18060 29586 18116 29596
rect 17948 29426 18116 29428
rect 17948 29374 17950 29426
rect 18002 29374 18116 29426
rect 17948 29372 18116 29374
rect 17948 29362 18004 29372
rect 17836 28702 17838 28754
rect 17890 28702 17892 28754
rect 17836 28690 17892 28702
rect 17948 28644 18004 28654
rect 17948 28420 18004 28588
rect 18060 28420 18116 29372
rect 18172 28644 18228 32284
rect 18508 30324 18564 33068
rect 18620 32788 18676 36652
rect 18732 35698 18788 37100
rect 18732 35646 18734 35698
rect 18786 35646 18788 35698
rect 18732 35028 18788 35646
rect 18844 35364 18900 38612
rect 18956 38164 19012 38174
rect 18956 36036 19012 38108
rect 19292 37492 19348 39676
rect 19404 39508 19460 39518
rect 19404 39414 19460 39452
rect 19516 39172 19572 40126
rect 19404 39116 19572 39172
rect 19404 38388 19460 39116
rect 19516 38948 19572 38958
rect 19516 38854 19572 38892
rect 19404 38332 19572 38388
rect 19404 38164 19460 38174
rect 19404 38070 19460 38108
rect 19516 37940 19572 38332
rect 19292 37426 19348 37436
rect 19404 37884 19572 37940
rect 19404 37378 19460 37884
rect 19516 37492 19572 37502
rect 19516 37398 19572 37436
rect 19404 37326 19406 37378
rect 19458 37326 19460 37378
rect 19068 37268 19124 37278
rect 19404 37268 19460 37326
rect 19068 37266 19460 37268
rect 19068 37214 19070 37266
rect 19122 37214 19460 37266
rect 19068 37212 19460 37214
rect 19068 37042 19124 37212
rect 19068 36990 19070 37042
rect 19122 36990 19124 37042
rect 19068 36978 19124 36990
rect 18956 35970 19012 35980
rect 19180 36820 19236 36830
rect 18844 35308 19124 35364
rect 18732 34356 18788 34972
rect 18956 35028 19012 35038
rect 18956 34916 19012 34972
rect 18732 34290 18788 34300
rect 18844 34860 19012 34916
rect 19068 34914 19124 35308
rect 19180 35140 19236 36764
rect 19404 36148 19460 37212
rect 19516 36820 19572 36830
rect 19516 36370 19572 36764
rect 19516 36318 19518 36370
rect 19570 36318 19572 36370
rect 19516 36306 19572 36318
rect 19404 36092 19572 36148
rect 19180 35074 19236 35084
rect 19292 35922 19348 35934
rect 19292 35870 19294 35922
rect 19346 35870 19348 35922
rect 19292 35028 19348 35870
rect 19404 35812 19460 35822
rect 19404 35718 19460 35756
rect 19516 35028 19572 36092
rect 19628 35308 19684 40348
rect 19740 40178 19796 40572
rect 20412 40514 20468 40526
rect 20412 40462 20414 40514
rect 20466 40462 20468 40514
rect 20188 40402 20244 40414
rect 20188 40350 20190 40402
rect 20242 40350 20244 40402
rect 19740 40126 19742 40178
rect 19794 40126 19796 40178
rect 19740 40114 19796 40126
rect 19852 40180 19908 40190
rect 19852 39618 19908 40124
rect 19852 39566 19854 39618
rect 19906 39566 19908 39618
rect 19852 39554 19908 39566
rect 19836 39228 20100 39238
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 19836 39162 20100 39172
rect 20188 38948 20244 40350
rect 20300 39620 20356 39630
rect 20412 39620 20468 40462
rect 20636 40402 20692 40414
rect 20636 40350 20638 40402
rect 20690 40350 20692 40402
rect 20636 40292 20692 40350
rect 20300 39618 20468 39620
rect 20300 39566 20302 39618
rect 20354 39566 20468 39618
rect 20300 39564 20468 39566
rect 20300 39554 20356 39564
rect 19852 38722 19908 38734
rect 19852 38670 19854 38722
rect 19906 38670 19908 38722
rect 19852 38276 19908 38670
rect 20188 38722 20244 38892
rect 20300 39396 20356 39406
rect 20300 39058 20356 39340
rect 20300 39006 20302 39058
rect 20354 39006 20356 39058
rect 20300 38836 20356 39006
rect 20300 38770 20356 38780
rect 20188 38670 20190 38722
rect 20242 38670 20244 38722
rect 20188 38658 20244 38670
rect 20412 38668 20468 39564
rect 20524 40236 20636 40292
rect 20524 38946 20580 40236
rect 20636 40226 20692 40236
rect 20524 38894 20526 38946
rect 20578 38894 20580 38946
rect 20524 38882 20580 38894
rect 20748 38668 20804 40908
rect 20300 38612 20468 38668
rect 20300 38388 20356 38612
rect 19852 38210 19908 38220
rect 20076 38332 20356 38388
rect 20076 38274 20132 38332
rect 20076 38222 20078 38274
rect 20130 38222 20132 38274
rect 20076 38210 20132 38222
rect 19852 38052 19908 38062
rect 19852 38050 20244 38052
rect 19852 37998 19854 38050
rect 19906 37998 20244 38050
rect 19852 37996 20244 37998
rect 19852 37986 19908 37996
rect 19836 37660 20100 37670
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 19836 37594 20100 37604
rect 20188 37492 20244 37996
rect 20188 37266 20244 37436
rect 20188 37214 20190 37266
rect 20242 37214 20244 37266
rect 20188 37202 20244 37214
rect 20300 38050 20356 38062
rect 20300 37998 20302 38050
rect 20354 37998 20356 38050
rect 20300 37268 20356 37998
rect 20412 37940 20468 38612
rect 20412 37268 20468 37884
rect 20636 38612 20804 38668
rect 20860 40514 20916 41692
rect 21308 41186 21364 41804
rect 21308 41134 21310 41186
rect 21362 41134 21364 41186
rect 21308 41122 21364 41134
rect 20860 40462 20862 40514
rect 20914 40462 20916 40514
rect 20524 37268 20580 37278
rect 20412 37266 20580 37268
rect 20412 37214 20526 37266
rect 20578 37214 20580 37266
rect 20412 37212 20580 37214
rect 20300 37202 20356 37212
rect 20524 37202 20580 37212
rect 20636 36820 20692 38612
rect 20300 36764 20692 36820
rect 20748 37826 20804 37838
rect 20748 37774 20750 37826
rect 20802 37774 20804 37826
rect 20748 36820 20804 37774
rect 20860 37380 20916 40462
rect 20972 40402 21028 40414
rect 20972 40350 20974 40402
rect 21026 40350 21028 40402
rect 20972 40292 21028 40350
rect 20972 40226 21028 40236
rect 21644 39508 21700 41804
rect 21756 41298 21812 41310
rect 21756 41246 21758 41298
rect 21810 41246 21812 41298
rect 21756 40292 21812 41246
rect 22316 41076 22372 41086
rect 22428 41076 22484 43484
rect 22540 43540 22596 43550
rect 22652 43540 22708 44158
rect 23660 43652 23716 43662
rect 23772 43652 23828 46284
rect 23884 45890 23940 45902
rect 23884 45838 23886 45890
rect 23938 45838 23940 45890
rect 23884 45220 23940 45838
rect 25452 45890 25508 45902
rect 25452 45838 25454 45890
rect 25506 45838 25508 45890
rect 24556 45780 24612 45790
rect 24556 45686 24612 45724
rect 25340 45780 25396 45790
rect 24892 45668 24948 45678
rect 24892 45666 25284 45668
rect 24892 45614 24894 45666
rect 24946 45614 25284 45666
rect 24892 45612 25284 45614
rect 24892 45602 24948 45612
rect 23884 45154 23940 45164
rect 24444 45108 24500 45118
rect 24444 45014 24500 45052
rect 24108 44996 24164 45006
rect 24108 44994 24388 44996
rect 24108 44942 24110 44994
rect 24162 44942 24388 44994
rect 24108 44940 24388 44942
rect 24108 44930 24164 44940
rect 23660 43650 23828 43652
rect 23660 43598 23662 43650
rect 23714 43598 23828 43650
rect 23660 43596 23828 43598
rect 23660 43586 23716 43596
rect 22540 43538 22708 43540
rect 22540 43486 22542 43538
rect 22594 43486 22708 43538
rect 22540 43484 22708 43486
rect 22540 43474 22596 43484
rect 23212 42756 23268 42766
rect 23100 41860 23156 41870
rect 23100 41766 23156 41804
rect 23212 41748 23268 42700
rect 23324 42756 23380 42766
rect 23324 42754 23492 42756
rect 23324 42702 23326 42754
rect 23378 42702 23492 42754
rect 23324 42700 23492 42702
rect 23324 42690 23380 42700
rect 23436 41972 23492 42700
rect 23996 42644 24052 42654
rect 23996 42642 24276 42644
rect 23996 42590 23998 42642
rect 24050 42590 24276 42642
rect 23996 42588 24276 42590
rect 23996 42578 24052 42588
rect 24220 42194 24276 42588
rect 24220 42142 24222 42194
rect 24274 42142 24276 42194
rect 24220 42130 24276 42142
rect 23436 41916 23716 41972
rect 23660 41860 23716 41916
rect 23772 41970 23828 41982
rect 23772 41918 23774 41970
rect 23826 41918 23828 41970
rect 23772 41860 23828 41918
rect 23660 41804 24164 41860
rect 23548 41748 23604 41758
rect 23212 41692 23548 41748
rect 23548 41682 23604 41692
rect 24108 41298 24164 41804
rect 24108 41246 24110 41298
rect 24162 41246 24164 41298
rect 22652 41076 22708 41086
rect 22428 41074 22708 41076
rect 22428 41022 22654 41074
rect 22706 41022 22708 41074
rect 22428 41020 22708 41022
rect 22316 40514 22372 41020
rect 22652 41010 22708 41020
rect 22988 40962 23044 40974
rect 22988 40910 22990 40962
rect 23042 40910 23044 40962
rect 22316 40462 22318 40514
rect 22370 40462 22372 40514
rect 22316 40450 22372 40462
rect 22876 40628 22932 40638
rect 22764 40402 22820 40414
rect 22764 40350 22766 40402
rect 22818 40350 22820 40402
rect 21812 40236 21924 40292
rect 21756 40226 21812 40236
rect 21644 39452 21812 39508
rect 21420 39396 21476 39406
rect 21084 39394 21476 39396
rect 21084 39342 21422 39394
rect 21474 39342 21476 39394
rect 21084 39340 21476 39342
rect 21084 38668 21140 39340
rect 21420 39330 21476 39340
rect 21196 39116 21476 39172
rect 21196 38946 21252 39116
rect 21420 39060 21476 39116
rect 21644 39060 21700 39070
rect 21420 39058 21700 39060
rect 21420 39006 21646 39058
rect 21698 39006 21700 39058
rect 21420 39004 21700 39006
rect 21644 38994 21700 39004
rect 21196 38894 21198 38946
rect 21250 38894 21252 38946
rect 21196 38882 21252 38894
rect 21308 38946 21364 38958
rect 21308 38894 21310 38946
rect 21362 38894 21364 38946
rect 21084 38612 21252 38668
rect 20860 37314 20916 37324
rect 21196 38050 21252 38612
rect 21196 37998 21198 38050
rect 21250 37998 21252 38050
rect 21084 37268 21140 37278
rect 21084 37174 21140 37212
rect 19836 36092 20100 36102
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 19836 36026 20100 36036
rect 19964 35924 20020 35934
rect 19964 35830 20020 35868
rect 19628 35252 19908 35308
rect 19740 35140 19796 35150
rect 19516 34972 19684 35028
rect 19292 34962 19348 34972
rect 19068 34862 19070 34914
rect 19122 34862 19124 34914
rect 18844 34804 18900 34860
rect 19068 34850 19124 34862
rect 19628 34916 19684 34972
rect 19628 34822 19684 34860
rect 18844 34244 18900 34748
rect 19516 34802 19572 34814
rect 19516 34750 19518 34802
rect 19570 34750 19572 34802
rect 18956 34692 19012 34702
rect 19180 34692 19236 34702
rect 18956 34598 19012 34636
rect 19068 34690 19236 34692
rect 19068 34638 19182 34690
rect 19234 34638 19236 34690
rect 19068 34636 19236 34638
rect 18956 34244 19012 34254
rect 18844 34188 18956 34244
rect 18956 34150 19012 34188
rect 19068 33684 19124 34636
rect 19180 34626 19236 34636
rect 19292 34692 19348 34702
rect 19180 34132 19236 34142
rect 19292 34132 19348 34636
rect 19236 34076 19348 34132
rect 19180 34038 19236 34076
rect 19516 33796 19572 34750
rect 19740 34692 19796 35084
rect 19852 34804 19908 35252
rect 20076 34916 20132 34926
rect 20076 34822 20132 34860
rect 19852 34738 19908 34748
rect 20188 34804 20244 34814
rect 19740 34626 19796 34636
rect 19836 34524 20100 34534
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 19836 34458 20100 34468
rect 19852 34356 19908 34366
rect 19516 33730 19572 33740
rect 19628 34244 19684 34254
rect 19292 33684 19348 33694
rect 19068 33628 19292 33684
rect 19292 33346 19348 33628
rect 19292 33294 19294 33346
rect 19346 33294 19348 33346
rect 18956 32788 19012 32798
rect 18620 32732 18956 32788
rect 18956 32694 19012 32732
rect 18844 32228 18900 32238
rect 18508 30258 18564 30268
rect 18620 31668 18676 31678
rect 18284 30100 18340 30110
rect 18284 29650 18340 30044
rect 18284 29598 18286 29650
rect 18338 29598 18340 29650
rect 18284 29586 18340 29598
rect 18396 29986 18452 29998
rect 18396 29934 18398 29986
rect 18450 29934 18452 29986
rect 18396 29652 18452 29934
rect 18396 29586 18452 29596
rect 18508 29988 18564 29998
rect 18508 29426 18564 29932
rect 18508 29374 18510 29426
rect 18562 29374 18564 29426
rect 18508 29362 18564 29374
rect 18172 28578 18228 28588
rect 18396 28420 18452 28430
rect 18060 28418 18452 28420
rect 18060 28366 18398 28418
rect 18450 28366 18452 28418
rect 18060 28364 18452 28366
rect 17948 28354 18004 28364
rect 17836 28084 17892 28094
rect 17836 27990 17892 28028
rect 17724 27906 17780 27916
rect 18396 27860 18452 28364
rect 18396 27766 18452 27804
rect 18060 27524 18116 27534
rect 18060 27074 18116 27468
rect 18060 27022 18062 27074
rect 18114 27022 18116 27074
rect 18060 27010 18116 27022
rect 17836 26964 17892 27002
rect 17836 26898 17892 26908
rect 18396 26852 18452 26862
rect 18396 26850 18564 26852
rect 18396 26798 18398 26850
rect 18450 26798 18564 26850
rect 18396 26796 18564 26798
rect 18396 26786 18452 26796
rect 17612 26402 17780 26404
rect 17612 26350 17614 26402
rect 17666 26350 17780 26402
rect 17612 26348 17780 26350
rect 17612 26338 17668 26348
rect 17500 26290 17556 26302
rect 17500 26238 17502 26290
rect 17554 26238 17556 26290
rect 17500 25396 17556 26238
rect 17500 25330 17556 25340
rect 17612 25282 17668 25294
rect 17612 25230 17614 25282
rect 17666 25230 17668 25282
rect 17612 25172 17668 25230
rect 17500 25116 17612 25172
rect 17500 24948 17556 25116
rect 17612 25106 17668 25116
rect 17500 24882 17556 24892
rect 17612 24948 17668 24958
rect 17724 24948 17780 26348
rect 18060 26402 18116 26414
rect 18060 26350 18062 26402
rect 18114 26350 18116 26402
rect 17836 26292 17892 26302
rect 17836 26290 18004 26292
rect 17836 26238 17838 26290
rect 17890 26238 18004 26290
rect 17836 26236 18004 26238
rect 17836 26226 17892 26236
rect 17836 25508 17892 25546
rect 17836 25442 17892 25452
rect 17948 25396 18004 26236
rect 18060 25620 18116 26350
rect 18284 26404 18340 26414
rect 18284 26310 18340 26348
rect 18508 26402 18564 26796
rect 18508 26350 18510 26402
rect 18562 26350 18564 26402
rect 18508 26338 18564 26350
rect 18620 26850 18676 31612
rect 18844 27746 18900 32172
rect 19292 32004 19348 33294
rect 19628 33460 19684 34188
rect 19852 34130 19908 34300
rect 19852 34078 19854 34130
rect 19906 34078 19908 34130
rect 19852 34066 19908 34078
rect 19740 33460 19796 33470
rect 19628 33458 19796 33460
rect 19628 33406 19742 33458
rect 19794 33406 19796 33458
rect 19628 33404 19796 33406
rect 19628 32788 19684 33404
rect 19740 33394 19796 33404
rect 20188 33460 20244 34748
rect 20188 33394 20244 33404
rect 19836 32956 20100 32966
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 19836 32890 20100 32900
rect 19628 32732 19796 32788
rect 19516 32676 19572 32686
rect 19516 32564 19572 32620
rect 19628 32564 19684 32574
rect 19516 32562 19684 32564
rect 19516 32510 19630 32562
rect 19682 32510 19684 32562
rect 19516 32508 19684 32510
rect 19628 32498 19684 32508
rect 19292 31938 19348 31948
rect 19628 31780 19684 31790
rect 19740 31780 19796 32732
rect 20188 32452 20244 32462
rect 20076 32396 20188 32452
rect 19628 31778 19796 31780
rect 19628 31726 19630 31778
rect 19682 31726 19796 31778
rect 19628 31724 19796 31726
rect 19852 32004 19908 32014
rect 19852 31778 19908 31948
rect 19852 31726 19854 31778
rect 19906 31726 19908 31778
rect 19628 31714 19684 31724
rect 19852 31714 19908 31726
rect 19292 31554 19348 31566
rect 19292 31502 19294 31554
rect 19346 31502 19348 31554
rect 19292 31220 19348 31502
rect 19404 31554 19460 31566
rect 19404 31502 19406 31554
rect 19458 31502 19460 31554
rect 19404 31332 19460 31502
rect 19516 31556 19572 31566
rect 20076 31556 20132 32396
rect 20188 32358 20244 32396
rect 20300 32228 20356 36764
rect 20748 36754 20804 36764
rect 20860 37042 20916 37054
rect 20860 36990 20862 37042
rect 20914 36990 20916 37042
rect 20412 36596 20468 36606
rect 20468 36540 20580 36596
rect 20412 36530 20468 36540
rect 20524 35810 20580 36540
rect 20524 35758 20526 35810
rect 20578 35758 20580 35810
rect 20524 35746 20580 35758
rect 20748 36482 20804 36494
rect 20748 36430 20750 36482
rect 20802 36430 20804 36482
rect 20188 32172 20356 32228
rect 20412 35698 20468 35710
rect 20412 35646 20414 35698
rect 20466 35646 20468 35698
rect 20188 31778 20244 32172
rect 20412 32004 20468 35646
rect 20748 34130 20804 36430
rect 20860 35700 20916 36990
rect 20860 35634 20916 35644
rect 20748 34078 20750 34130
rect 20802 34078 20804 34130
rect 20748 34066 20804 34078
rect 21084 34242 21140 34254
rect 21084 34190 21086 34242
rect 21138 34190 21140 34242
rect 20524 34018 20580 34030
rect 20524 33966 20526 34018
rect 20578 33966 20580 34018
rect 20524 33908 20580 33966
rect 21084 33908 21140 34190
rect 20524 33852 21140 33908
rect 20972 32452 21028 32462
rect 20972 32358 21028 32396
rect 21196 32228 21252 37998
rect 21308 36260 21364 38894
rect 21532 38836 21588 38846
rect 21756 38836 21812 39452
rect 21532 38834 21812 38836
rect 21532 38782 21534 38834
rect 21586 38782 21812 38834
rect 21532 38780 21812 38782
rect 21868 39058 21924 40236
rect 21868 39006 21870 39058
rect 21922 39006 21924 39058
rect 21532 38770 21588 38780
rect 21532 38612 21588 38622
rect 21532 37492 21588 38556
rect 21868 38052 21924 39006
rect 22092 39618 22148 39630
rect 22092 39566 22094 39618
rect 22146 39566 22148 39618
rect 21980 38834 22036 38846
rect 21980 38782 21982 38834
rect 22034 38782 22036 38834
rect 21980 38612 22036 38782
rect 22092 38836 22148 39566
rect 22652 39620 22708 39630
rect 22764 39620 22820 40350
rect 22876 39732 22932 40572
rect 22988 40516 23044 40910
rect 23212 40516 23268 40526
rect 22988 40514 23268 40516
rect 22988 40462 23214 40514
rect 23266 40462 23268 40514
rect 22988 40460 23268 40462
rect 23212 40068 23268 40460
rect 23212 40002 23268 40012
rect 23436 40402 23492 40414
rect 23436 40350 23438 40402
rect 23490 40350 23492 40402
rect 22988 39732 23044 39742
rect 22876 39730 23044 39732
rect 22876 39678 22990 39730
rect 23042 39678 23044 39730
rect 22876 39676 23044 39678
rect 22988 39666 23044 39676
rect 23436 39620 23492 40350
rect 22652 39618 22820 39620
rect 22652 39566 22654 39618
rect 22706 39566 22820 39618
rect 22652 39564 22820 39566
rect 22652 39554 22708 39564
rect 22652 39060 22708 39070
rect 22652 38966 22708 39004
rect 22092 38770 22148 38780
rect 21980 38546 22036 38556
rect 22764 38052 22820 39564
rect 23100 39618 23492 39620
rect 23100 39566 23438 39618
rect 23490 39566 23492 39618
rect 23100 39564 23492 39566
rect 22988 39060 23044 39070
rect 23100 39060 23156 39564
rect 23436 39554 23492 39564
rect 23660 40068 23716 40078
rect 22988 39058 23156 39060
rect 22988 39006 22990 39058
rect 23042 39006 23156 39058
rect 22988 39004 23156 39006
rect 23660 39058 23716 40012
rect 23996 39620 24052 39630
rect 24108 39620 24164 41246
rect 23996 39618 24108 39620
rect 23996 39566 23998 39618
rect 24050 39566 24108 39618
rect 23996 39564 24108 39566
rect 23996 39554 24052 39564
rect 24108 39526 24164 39564
rect 23660 39006 23662 39058
rect 23714 39006 23716 39058
rect 22988 38668 23044 39004
rect 23660 38994 23716 39006
rect 23324 38946 23380 38958
rect 23324 38894 23326 38946
rect 23378 38894 23380 38946
rect 22988 38612 23156 38668
rect 21868 37996 22036 38052
rect 21644 37940 21700 37950
rect 21644 37846 21700 37884
rect 21420 37436 21588 37492
rect 21756 37826 21812 37838
rect 21756 37774 21758 37826
rect 21810 37774 21812 37826
rect 21420 36482 21476 37436
rect 21644 37380 21700 37390
rect 21532 37266 21588 37278
rect 21532 37214 21534 37266
rect 21586 37214 21588 37266
rect 21532 37156 21588 37214
rect 21532 37090 21588 37100
rect 21420 36430 21422 36482
rect 21474 36430 21476 36482
rect 21420 36418 21476 36430
rect 21308 36204 21476 36260
rect 21308 35028 21364 35038
rect 21308 34914 21364 34972
rect 21420 35026 21476 36204
rect 21532 35812 21588 35822
rect 21644 35812 21700 37324
rect 21756 36484 21812 37774
rect 21868 37826 21924 37838
rect 21868 37774 21870 37826
rect 21922 37774 21924 37826
rect 21868 37268 21924 37774
rect 21980 37268 22036 37996
rect 22764 37986 22820 37996
rect 22876 38388 22932 38398
rect 22652 37938 22708 37950
rect 22652 37886 22654 37938
rect 22706 37886 22708 37938
rect 22316 37828 22372 37838
rect 22316 37826 22596 37828
rect 22316 37774 22318 37826
rect 22370 37774 22596 37826
rect 22316 37772 22596 37774
rect 22316 37762 22372 37772
rect 22540 37380 22596 37772
rect 22428 37268 22484 37278
rect 21980 37266 22484 37268
rect 21980 37214 22430 37266
rect 22482 37214 22484 37266
rect 21980 37212 22484 37214
rect 21868 37154 21924 37212
rect 21868 37102 21870 37154
rect 21922 37102 21924 37154
rect 21868 37090 21924 37102
rect 21756 36428 22148 36484
rect 21588 35756 21700 35812
rect 21756 36258 21812 36270
rect 21756 36206 21758 36258
rect 21810 36206 21812 36258
rect 21532 35746 21588 35756
rect 21420 34974 21422 35026
rect 21474 34974 21476 35026
rect 21420 34962 21476 34974
rect 21532 35252 21588 35262
rect 21308 34862 21310 34914
rect 21362 34862 21364 34914
rect 21308 34850 21364 34862
rect 21532 34802 21588 35196
rect 21756 35252 21812 36206
rect 21868 36260 21924 36270
rect 21868 36166 21924 36204
rect 21980 36258 22036 36270
rect 21980 36206 21982 36258
rect 22034 36206 22036 36258
rect 21756 35186 21812 35196
rect 21756 34916 21812 34926
rect 21756 34914 21924 34916
rect 21756 34862 21758 34914
rect 21810 34862 21924 34914
rect 21756 34860 21924 34862
rect 21756 34850 21812 34860
rect 21532 34750 21534 34802
rect 21586 34750 21588 34802
rect 21532 34468 21588 34750
rect 21532 34412 21812 34468
rect 21644 34244 21700 34254
rect 21308 34242 21700 34244
rect 21308 34190 21646 34242
rect 21698 34190 21700 34242
rect 21308 34188 21700 34190
rect 21308 33458 21364 34188
rect 21644 34178 21700 34188
rect 21756 33796 21812 34412
rect 21868 34356 21924 34860
rect 21980 34356 22036 36206
rect 22092 34914 22148 36428
rect 22316 36372 22372 36382
rect 22204 36370 22372 36372
rect 22204 36318 22318 36370
rect 22370 36318 22372 36370
rect 22204 36316 22372 36318
rect 22204 35698 22260 36316
rect 22316 36306 22372 36316
rect 22204 35646 22206 35698
rect 22258 35646 22260 35698
rect 22204 35634 22260 35646
rect 22092 34862 22094 34914
rect 22146 34862 22148 34914
rect 22092 34850 22148 34862
rect 22428 34916 22484 37212
rect 22540 35140 22596 37324
rect 22652 36594 22708 37886
rect 22764 37828 22820 37838
rect 22876 37828 22932 38332
rect 22764 37826 22876 37828
rect 22764 37774 22766 37826
rect 22818 37774 22876 37826
rect 22764 37772 22876 37774
rect 22764 37762 22820 37772
rect 22876 37734 22932 37772
rect 22988 37826 23044 37838
rect 22988 37774 22990 37826
rect 23042 37774 23044 37826
rect 22652 36542 22654 36594
rect 22706 36542 22708 36594
rect 22652 36260 22708 36542
rect 22652 36194 22708 36204
rect 22764 37492 22820 37502
rect 22540 35074 22596 35084
rect 22428 34850 22484 34860
rect 22540 34804 22596 34814
rect 22540 34710 22596 34748
rect 22764 34580 22820 37436
rect 22988 37266 23044 37774
rect 22988 37214 22990 37266
rect 23042 37214 23044 37266
rect 22988 37202 23044 37214
rect 22988 36820 23044 36830
rect 22988 35810 23044 36764
rect 22988 35758 22990 35810
rect 23042 35758 23044 35810
rect 22988 35746 23044 35758
rect 22988 35252 23044 35262
rect 22876 35026 22932 35038
rect 22876 34974 22878 35026
rect 22930 34974 22932 35026
rect 22876 34916 22932 34974
rect 22876 34850 22932 34860
rect 22988 34914 23044 35196
rect 22988 34862 22990 34914
rect 23042 34862 23044 34914
rect 22988 34850 23044 34862
rect 22764 34514 22820 34524
rect 23100 34468 23156 38612
rect 23324 38612 23380 38894
rect 24108 38722 24164 38734
rect 24108 38670 24110 38722
rect 24162 38670 24164 38722
rect 24108 38668 24164 38670
rect 24108 38612 24276 38668
rect 23324 37268 23380 38556
rect 23660 38274 23716 38286
rect 23660 38222 23662 38274
rect 23714 38222 23716 38274
rect 23660 38164 23716 38222
rect 24108 38274 24164 38286
rect 24108 38222 24110 38274
rect 24162 38222 24164 38274
rect 23660 38162 23828 38164
rect 23660 38110 23662 38162
rect 23714 38110 23828 38162
rect 23660 38108 23828 38110
rect 23660 38098 23716 38108
rect 23772 37604 23828 38108
rect 24108 38162 24164 38222
rect 24108 38110 24110 38162
rect 24162 38110 24164 38162
rect 24108 38098 24164 38110
rect 24220 37828 24276 38612
rect 24332 38274 24388 44940
rect 25228 44434 25284 45612
rect 25340 45330 25396 45724
rect 25340 45278 25342 45330
rect 25394 45278 25396 45330
rect 25340 45266 25396 45278
rect 25228 44382 25230 44434
rect 25282 44382 25284 44434
rect 25228 44370 25284 44382
rect 25340 45108 25396 45118
rect 25340 43650 25396 45052
rect 25340 43598 25342 43650
rect 25394 43598 25396 43650
rect 25340 43586 25396 43598
rect 24892 43428 24948 43438
rect 24556 41970 24612 41982
rect 24556 41918 24558 41970
rect 24610 41918 24612 41970
rect 24556 41860 24612 41918
rect 24556 41794 24612 41804
rect 24892 41748 24948 43372
rect 24892 41298 24948 41692
rect 24892 41246 24894 41298
rect 24946 41246 24948 41298
rect 24892 41234 24948 41246
rect 25116 41972 25172 41982
rect 25452 41972 25508 45838
rect 25564 45332 25620 49200
rect 26236 46116 26292 49200
rect 26236 46050 26292 46060
rect 26908 46002 26964 49200
rect 29372 46116 29428 46126
rect 29372 46022 29428 46060
rect 30268 46116 30324 49200
rect 30268 46050 30324 46060
rect 26908 45950 26910 46002
rect 26962 45950 26964 46002
rect 26908 45938 26964 45950
rect 25564 45266 25620 45276
rect 28588 45890 28644 45902
rect 28588 45838 28590 45890
rect 28642 45838 28644 45890
rect 25676 45220 25732 45230
rect 25676 45106 25732 45164
rect 26460 45218 26516 45230
rect 26460 45166 26462 45218
rect 26514 45166 26516 45218
rect 25676 45054 25678 45106
rect 25730 45054 25732 45106
rect 25676 45042 25732 45054
rect 26348 45106 26404 45118
rect 26348 45054 26350 45106
rect 26402 45054 26404 45106
rect 25900 44322 25956 44334
rect 25900 44270 25902 44322
rect 25954 44270 25956 44322
rect 25900 43538 25956 44270
rect 25900 43486 25902 43538
rect 25954 43486 25956 43538
rect 25900 42532 25956 43486
rect 25900 42466 25956 42476
rect 26124 43764 26180 43774
rect 26124 42866 26180 43708
rect 26124 42814 26126 42866
rect 26178 42814 26180 42866
rect 26124 42084 26180 42814
rect 26348 42196 26404 45054
rect 26460 44996 26516 45166
rect 27356 45108 27412 45118
rect 26908 44996 26964 45006
rect 26460 44994 26964 44996
rect 26460 44942 26910 44994
rect 26962 44942 26964 44994
rect 26460 44940 26964 44942
rect 26572 44772 26628 44782
rect 26460 44098 26516 44110
rect 26460 44046 26462 44098
rect 26514 44046 26516 44098
rect 26460 42532 26516 44046
rect 26572 43764 26628 44716
rect 26908 44548 26964 44940
rect 26908 44482 26964 44492
rect 27356 44546 27412 45052
rect 28588 44772 28644 45838
rect 30156 45332 30212 45342
rect 29036 45330 30212 45332
rect 29036 45278 30158 45330
rect 30210 45278 30212 45330
rect 29036 45276 30212 45278
rect 29036 45218 29092 45276
rect 30156 45266 30212 45276
rect 29036 45166 29038 45218
rect 29090 45166 29092 45218
rect 29036 45154 29092 45166
rect 28588 44706 28644 44716
rect 29820 45106 29876 45118
rect 29820 45054 29822 45106
rect 29874 45054 29876 45106
rect 27356 44494 27358 44546
rect 27410 44494 27412 44546
rect 27356 44482 27412 44494
rect 27692 44548 27748 44558
rect 27692 44454 27748 44492
rect 28364 44322 28420 44334
rect 28364 44270 28366 44322
rect 28418 44270 28420 44322
rect 28364 44100 28420 44270
rect 28700 44324 28756 44334
rect 29820 44324 29876 45054
rect 30380 45108 30436 45118
rect 30380 45014 30436 45052
rect 29932 44324 29988 44334
rect 29820 44268 29932 44324
rect 28364 44034 28420 44044
rect 28476 44210 28532 44222
rect 28476 44158 28478 44210
rect 28530 44158 28532 44210
rect 26572 43698 26628 43708
rect 26572 43428 26628 43438
rect 26572 43426 27076 43428
rect 26572 43374 26574 43426
rect 26626 43374 27076 43426
rect 26572 43372 27076 43374
rect 26572 43362 26628 43372
rect 27020 42642 27076 43372
rect 28476 42756 28532 44158
rect 28700 43426 28756 44268
rect 29372 44100 29428 44110
rect 29372 44006 29428 44044
rect 29148 43764 29204 43802
rect 29820 43764 29876 43774
rect 29932 43708 29988 44268
rect 30380 44324 30436 44334
rect 30380 44230 30436 44268
rect 29148 43698 29204 43708
rect 28700 43374 28702 43426
rect 28754 43374 28756 43426
rect 28700 42980 28756 43374
rect 29708 43652 29988 43708
rect 30268 44100 30324 44110
rect 29708 43538 29764 43652
rect 29708 43486 29710 43538
rect 29762 43486 29764 43538
rect 29596 42980 29652 42990
rect 28700 42978 29652 42980
rect 28700 42926 29598 42978
rect 29650 42926 29652 42978
rect 28700 42924 29652 42926
rect 29596 42914 29652 42924
rect 28476 42690 28532 42700
rect 27020 42590 27022 42642
rect 27074 42590 27076 42642
rect 27020 42578 27076 42590
rect 27356 42644 27412 42654
rect 27356 42550 27412 42588
rect 29260 42644 29316 42654
rect 29260 42550 29316 42588
rect 26572 42532 26628 42542
rect 26460 42476 26572 42532
rect 26628 42476 26740 42532
rect 26572 42438 26628 42476
rect 26348 42140 26516 42196
rect 26236 42084 26292 42094
rect 26124 42082 26292 42084
rect 26124 42030 26238 42082
rect 26290 42030 26292 42082
rect 26124 42028 26292 42030
rect 26236 42018 26292 42028
rect 25452 41916 26068 41972
rect 24668 39508 24724 39518
rect 24668 39414 24724 39452
rect 24332 38222 24334 38274
rect 24386 38222 24388 38274
rect 24332 38210 24388 38222
rect 24220 37762 24276 37772
rect 24668 37826 24724 37838
rect 24668 37774 24670 37826
rect 24722 37774 24724 37826
rect 23436 37492 23492 37502
rect 23436 37378 23492 37436
rect 23436 37326 23438 37378
rect 23490 37326 23492 37378
rect 23436 37314 23492 37326
rect 23548 37380 23604 37390
rect 23548 37286 23604 37324
rect 23772 37378 23828 37548
rect 24668 37492 24724 37774
rect 24668 37426 24724 37436
rect 24220 37380 24276 37390
rect 23772 37326 23774 37378
rect 23826 37326 23828 37378
rect 23772 37314 23828 37326
rect 23996 37378 24276 37380
rect 23996 37326 24222 37378
rect 24274 37326 24276 37378
rect 23996 37324 24276 37326
rect 23324 37202 23380 37212
rect 23436 37154 23492 37166
rect 23436 37102 23438 37154
rect 23490 37102 23492 37154
rect 23212 36482 23268 36494
rect 23212 36430 23214 36482
rect 23266 36430 23268 36482
rect 23212 35028 23268 36430
rect 23436 35924 23492 37102
rect 23436 35858 23492 35868
rect 23884 37156 23940 37166
rect 23324 35700 23380 35710
rect 23548 35700 23604 35710
rect 23380 35698 23604 35700
rect 23380 35646 23550 35698
rect 23602 35646 23604 35698
rect 23380 35644 23604 35646
rect 23324 35634 23380 35644
rect 23548 35634 23604 35644
rect 23772 35364 23828 35374
rect 23772 35028 23828 35308
rect 23212 34972 23828 35028
rect 23212 34916 23268 34972
rect 23212 34850 23268 34860
rect 23100 34412 23380 34468
rect 21980 34300 23268 34356
rect 21868 34290 21924 34300
rect 21308 33406 21310 33458
rect 21362 33406 21364 33458
rect 21308 33394 21364 33406
rect 21420 33740 21812 33796
rect 21868 34130 21924 34142
rect 21868 34078 21870 34130
rect 21922 34078 21924 34130
rect 21196 32162 21252 32172
rect 21308 32450 21364 32462
rect 21308 32398 21310 32450
rect 21362 32398 21364 32450
rect 20412 31948 20580 32004
rect 20188 31726 20190 31778
rect 20242 31726 20244 31778
rect 20188 31714 20244 31726
rect 20300 31780 20356 31790
rect 20300 31686 20356 31724
rect 20412 31778 20468 31790
rect 20412 31726 20414 31778
rect 20466 31726 20468 31778
rect 20076 31500 20244 31556
rect 19516 31462 19572 31500
rect 19836 31388 20100 31398
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 19404 31276 19572 31332
rect 19836 31322 20100 31332
rect 19516 31220 19572 31276
rect 19292 31164 19460 31220
rect 19516 31164 19796 31220
rect 18956 31108 19012 31118
rect 19404 31108 19460 31164
rect 19404 31052 19684 31108
rect 18956 30994 19012 31052
rect 18956 30942 18958 30994
rect 19010 30942 19012 30994
rect 18956 30930 19012 30942
rect 19516 30884 19572 30894
rect 19292 30828 19516 30884
rect 18956 30324 19012 30334
rect 19180 30324 19236 30334
rect 18956 30210 19012 30268
rect 18956 30158 18958 30210
rect 19010 30158 19012 30210
rect 18956 30146 19012 30158
rect 19068 30268 19180 30324
rect 19068 29650 19124 30268
rect 19180 30258 19236 30268
rect 19068 29598 19070 29650
rect 19122 29598 19124 29650
rect 19068 29586 19124 29598
rect 19180 29988 19236 29998
rect 18956 29316 19012 29326
rect 18956 29222 19012 29260
rect 18956 28644 19012 28654
rect 18956 28550 19012 28588
rect 19180 28084 19236 29932
rect 19180 28018 19236 28028
rect 18844 27694 18846 27746
rect 18898 27694 18900 27746
rect 18620 26798 18622 26850
rect 18674 26798 18676 26850
rect 18508 26180 18564 26190
rect 18396 26068 18452 26078
rect 18396 25974 18452 26012
rect 18060 25554 18116 25564
rect 18172 25732 18228 25742
rect 18172 25618 18228 25676
rect 18172 25566 18174 25618
rect 18226 25566 18228 25618
rect 18172 25554 18228 25566
rect 18396 25508 18452 25518
rect 17948 25340 18228 25396
rect 17836 25284 17892 25294
rect 17836 25172 17892 25228
rect 18172 25282 18228 25340
rect 18172 25230 18174 25282
rect 18226 25230 18228 25282
rect 18172 25218 18228 25230
rect 18396 25282 18452 25452
rect 18396 25230 18398 25282
rect 18450 25230 18452 25282
rect 17836 25116 18004 25172
rect 17612 24946 17780 24948
rect 17612 24894 17614 24946
rect 17666 24894 17780 24946
rect 17612 24892 17780 24894
rect 17612 24882 17668 24892
rect 17388 24668 17668 24724
rect 16604 24658 16660 24668
rect 16940 24630 16996 24668
rect 16940 24052 16996 24062
rect 16828 23940 16884 23950
rect 16380 23938 16884 23940
rect 16380 23886 16830 23938
rect 16882 23886 16884 23938
rect 16380 23884 16884 23886
rect 16828 23874 16884 23884
rect 16268 23492 16884 23548
rect 16156 23202 16212 23212
rect 16044 22866 16100 22876
rect 16156 23042 16212 23054
rect 16156 22990 16158 23042
rect 16210 22990 16212 23042
rect 16156 22930 16212 22990
rect 16156 22878 16158 22930
rect 16210 22878 16212 22930
rect 16156 22866 16212 22878
rect 15932 21810 16324 21812
rect 15932 21758 15934 21810
rect 15986 21758 16324 21810
rect 15932 21756 16324 21758
rect 15932 21746 15988 21756
rect 16156 21362 16212 21374
rect 16156 21310 16158 21362
rect 16210 21310 16212 21362
rect 16156 20802 16212 21310
rect 16156 20750 16158 20802
rect 16210 20750 16212 20802
rect 16156 20738 16212 20750
rect 16268 20802 16324 21756
rect 16380 21362 16436 23492
rect 16828 23378 16884 23492
rect 16828 23326 16830 23378
rect 16882 23326 16884 23378
rect 16828 23314 16884 23326
rect 16604 23156 16660 23166
rect 16940 23156 16996 23996
rect 17276 23940 17332 23950
rect 17276 23846 17332 23884
rect 17388 23716 17444 23726
rect 17388 23622 17444 23660
rect 17612 23378 17668 24668
rect 17836 24722 17892 24734
rect 17836 24670 17838 24722
rect 17890 24670 17892 24722
rect 17836 24052 17892 24670
rect 17836 23986 17892 23996
rect 17612 23326 17614 23378
rect 17666 23326 17668 23378
rect 17612 23314 17668 23326
rect 17836 23826 17892 23838
rect 17836 23774 17838 23826
rect 17890 23774 17892 23826
rect 17836 23380 17892 23774
rect 17836 23314 17892 23324
rect 16604 23154 16996 23156
rect 16604 23102 16606 23154
rect 16658 23102 16996 23154
rect 16604 23100 16996 23102
rect 17948 23156 18004 25116
rect 18284 25060 18340 25070
rect 18172 25004 18284 25060
rect 18172 24946 18228 25004
rect 18284 24994 18340 25004
rect 18172 24894 18174 24946
rect 18226 24894 18228 24946
rect 18172 24882 18228 24894
rect 18060 24724 18116 24734
rect 18396 24724 18452 25230
rect 18060 23938 18116 24668
rect 18060 23886 18062 23938
rect 18114 23886 18116 23938
rect 18060 23874 18116 23886
rect 18172 24668 18452 24724
rect 18172 23492 18228 24668
rect 18284 23828 18340 23838
rect 18284 23734 18340 23772
rect 18396 23714 18452 23726
rect 18396 23662 18398 23714
rect 18450 23662 18452 23714
rect 18172 23436 18340 23492
rect 18060 23156 18116 23166
rect 17948 23154 18116 23156
rect 17948 23102 18062 23154
rect 18114 23102 18116 23154
rect 17948 23100 18116 23102
rect 16604 23090 16660 23100
rect 16492 21476 16548 21486
rect 16492 21382 16548 21420
rect 16380 21310 16382 21362
rect 16434 21310 16436 21362
rect 16380 21252 16436 21310
rect 16716 21364 16772 23100
rect 17836 22708 17892 22718
rect 17836 22482 17892 22652
rect 17836 22430 17838 22482
rect 17890 22430 17892 22482
rect 17836 22418 17892 22430
rect 17500 21588 17556 21598
rect 18060 21588 18116 23100
rect 17500 21586 18116 21588
rect 17500 21534 17502 21586
rect 17554 21534 18116 21586
rect 17500 21532 18116 21534
rect 16716 21308 16996 21364
rect 16380 21196 16884 21252
rect 16268 20750 16270 20802
rect 16322 20750 16324 20802
rect 16268 20738 16324 20750
rect 15708 20244 15764 20254
rect 15708 20150 15764 20188
rect 15820 19346 15876 20636
rect 15932 20692 15988 20702
rect 16604 20692 16660 20702
rect 15932 20690 16100 20692
rect 15932 20638 15934 20690
rect 15986 20638 16100 20690
rect 15932 20636 16100 20638
rect 15932 20626 15988 20636
rect 16044 20468 16100 20636
rect 16380 20580 16436 20590
rect 16380 20486 16436 20524
rect 16492 20578 16548 20590
rect 16492 20526 16494 20578
rect 16546 20526 16548 20578
rect 16044 20412 16324 20468
rect 16044 20244 16100 20254
rect 16044 20242 16212 20244
rect 16044 20190 16046 20242
rect 16098 20190 16212 20242
rect 16044 20188 16212 20190
rect 16044 20178 16100 20188
rect 16044 20020 16100 20030
rect 16044 19926 16100 19964
rect 15820 19294 15822 19346
rect 15874 19294 15876 19346
rect 15820 19282 15876 19294
rect 16044 19012 16100 19022
rect 15596 18956 16044 19012
rect 15932 18676 15988 18686
rect 15820 17444 15876 17454
rect 15820 17106 15876 17388
rect 15820 17054 15822 17106
rect 15874 17054 15876 17106
rect 15820 17042 15876 17054
rect 15148 16818 15204 16828
rect 15372 16772 15428 16782
rect 15372 15202 15428 16716
rect 15372 15150 15374 15202
rect 15426 15150 15428 15202
rect 15372 15138 15428 15150
rect 15820 15204 15876 15242
rect 15820 15138 15876 15148
rect 15932 15148 15988 18620
rect 16044 18674 16100 18956
rect 16044 18622 16046 18674
rect 16098 18622 16100 18674
rect 16044 18610 16100 18622
rect 16044 16772 16100 16782
rect 16044 16678 16100 16716
rect 15932 15092 16100 15148
rect 15036 12786 15092 12796
rect 15372 12852 15428 12862
rect 14476 12402 14644 12404
rect 14476 12350 14478 12402
rect 14530 12350 14644 12402
rect 14476 12348 14644 12350
rect 14476 12338 14532 12348
rect 14084 12012 14420 12068
rect 14028 11974 14084 12012
rect 13692 11666 13748 11676
rect 13804 11506 13860 11518
rect 13804 11454 13806 11506
rect 13858 11454 13860 11506
rect 13692 11284 13748 11294
rect 13580 11282 13748 11284
rect 13580 11230 13694 11282
rect 13746 11230 13748 11282
rect 13580 11228 13748 11230
rect 13692 11218 13748 11228
rect 13804 10722 13860 11454
rect 14364 11172 14420 11182
rect 14364 11170 14532 11172
rect 14364 11118 14366 11170
rect 14418 11118 14532 11170
rect 14364 11116 14532 11118
rect 14364 11106 14420 11116
rect 13804 10670 13806 10722
rect 13858 10670 13860 10722
rect 13804 10658 13860 10670
rect 13580 9826 13636 9838
rect 13580 9774 13582 9826
rect 13634 9774 13636 9826
rect 12908 8540 13188 8596
rect 12908 8260 12964 8540
rect 13020 8372 13076 8382
rect 13020 8278 13076 8316
rect 12908 8194 12964 8204
rect 12796 7868 12964 7924
rect 12572 7588 12628 7598
rect 12628 7532 12740 7588
rect 12572 7522 12628 7532
rect 12348 6850 12404 6860
rect 12572 7028 12628 7038
rect 12460 6578 12516 6590
rect 12460 6526 12462 6578
rect 12514 6526 12516 6578
rect 12348 6132 12404 6142
rect 12012 6076 12180 6132
rect 12236 6130 12404 6132
rect 12236 6078 12350 6130
rect 12402 6078 12404 6130
rect 12236 6076 12404 6078
rect 11900 6020 11956 6030
rect 11956 5964 12068 6020
rect 11900 5926 11956 5964
rect 11788 5906 11844 5918
rect 11788 5854 11790 5906
rect 11842 5854 11844 5906
rect 11788 5236 11844 5854
rect 11900 5684 11956 5694
rect 11900 5590 11956 5628
rect 11788 5170 11844 5180
rect 12012 5122 12068 5964
rect 12012 5070 12014 5122
rect 12066 5070 12068 5122
rect 12012 5058 12068 5070
rect 11788 5012 11844 5022
rect 11788 4918 11844 4956
rect 11564 4722 11620 4732
rect 10780 4386 10836 4396
rect 10668 4116 10724 4126
rect 10668 4022 10724 4060
rect 10444 3502 10446 3554
rect 10498 3502 10500 3554
rect 10444 3490 10500 3502
rect 10780 3892 10836 3902
rect 10780 800 10836 3836
rect 12124 3556 12180 6076
rect 12348 6066 12404 6076
rect 12460 6132 12516 6526
rect 12572 6580 12628 6972
rect 12684 6692 12740 7532
rect 12796 7364 12852 7374
rect 12908 7364 12964 7868
rect 13132 7812 13188 8540
rect 13468 8372 13524 8382
rect 13468 8258 13524 8316
rect 13468 8206 13470 8258
rect 13522 8206 13524 8258
rect 13468 8194 13524 8206
rect 13580 8260 13636 9774
rect 14364 9714 14420 9726
rect 14364 9662 14366 9714
rect 14418 9662 14420 9714
rect 13692 9604 13748 9614
rect 13692 8482 13748 9548
rect 14364 9268 14420 9662
rect 14364 9202 14420 9212
rect 14476 9156 14532 11116
rect 14476 9090 14532 9100
rect 14588 10836 14644 12348
rect 15148 12740 15204 12750
rect 15148 12290 15204 12684
rect 15148 12238 15150 12290
rect 15202 12238 15204 12290
rect 15148 11956 15204 12238
rect 15372 12290 15428 12796
rect 15596 12850 15652 12862
rect 15596 12798 15598 12850
rect 15650 12798 15652 12850
rect 15596 12402 15652 12798
rect 15596 12350 15598 12402
rect 15650 12350 15652 12402
rect 15596 12338 15652 12350
rect 15372 12238 15374 12290
rect 15426 12238 15428 12290
rect 15372 12226 15428 12238
rect 15932 12180 15988 12190
rect 15932 12086 15988 12124
rect 15148 11890 15204 11900
rect 15708 12068 15764 12078
rect 15708 11954 15764 12012
rect 15708 11902 15710 11954
rect 15762 11902 15764 11954
rect 15708 11890 15764 11902
rect 15036 10836 15092 10846
rect 14588 10834 15204 10836
rect 14588 10782 15038 10834
rect 15090 10782 15204 10834
rect 14588 10780 15204 10782
rect 14588 10610 14644 10780
rect 15036 10742 15092 10780
rect 14588 10558 14590 10610
rect 14642 10558 14644 10610
rect 14588 9042 14644 10558
rect 15148 10500 15204 10780
rect 15484 10500 15540 10510
rect 15148 10498 15540 10500
rect 15148 10446 15486 10498
rect 15538 10446 15540 10498
rect 15148 10444 15540 10446
rect 15484 10164 15540 10444
rect 15484 10098 15540 10108
rect 15932 10498 15988 10510
rect 15932 10446 15934 10498
rect 15986 10446 15988 10498
rect 14924 9380 14980 9390
rect 14588 8990 14590 9042
rect 14642 8990 14644 9042
rect 14588 8978 14644 8990
rect 14812 9156 14868 9166
rect 13804 8932 13860 8942
rect 13804 8930 13972 8932
rect 13804 8878 13806 8930
rect 13858 8878 13972 8930
rect 13804 8876 13972 8878
rect 13804 8866 13860 8876
rect 13692 8430 13694 8482
rect 13746 8430 13748 8482
rect 13692 8418 13748 8430
rect 13132 7746 13188 7756
rect 13244 7588 13300 7598
rect 13244 7586 13412 7588
rect 13244 7534 13246 7586
rect 13298 7534 13412 7586
rect 13244 7532 13412 7534
rect 13244 7522 13300 7532
rect 12796 7362 12964 7364
rect 12796 7310 12798 7362
rect 12850 7310 12964 7362
rect 12796 7308 12964 7310
rect 12796 7298 12852 7308
rect 12908 6692 12964 7308
rect 13132 7474 13188 7486
rect 13132 7422 13134 7474
rect 13186 7422 13188 7474
rect 12684 6636 12852 6692
rect 12572 6486 12628 6524
rect 12684 6468 12740 6478
rect 12684 6356 12740 6412
rect 12460 6066 12516 6076
rect 12572 6300 12740 6356
rect 12124 3490 12180 3500
rect 12236 5796 12292 5806
rect 11564 3442 11620 3454
rect 11564 3390 11566 3442
rect 11618 3390 11620 3442
rect 11564 3388 11620 3390
rect 12236 3388 12292 5740
rect 12572 5348 12628 6300
rect 12684 5906 12740 5918
rect 12684 5854 12686 5906
rect 12738 5854 12740 5906
rect 12684 5796 12740 5854
rect 12684 5730 12740 5740
rect 12572 5292 12740 5348
rect 12572 5124 12628 5134
rect 12572 5010 12628 5068
rect 12572 4958 12574 5010
rect 12626 4958 12628 5010
rect 12572 4946 12628 4958
rect 12684 5012 12740 5292
rect 12684 4946 12740 4956
rect 12796 5122 12852 6636
rect 12908 6598 12964 6636
rect 13020 6916 13076 6926
rect 12908 6132 12964 6142
rect 12908 6038 12964 6076
rect 13020 5796 13076 6860
rect 13132 6468 13188 7422
rect 13132 6402 13188 6412
rect 13244 7250 13300 7262
rect 13244 7198 13246 7250
rect 13298 7198 13300 7250
rect 13244 6132 13300 7198
rect 13244 6066 13300 6076
rect 13132 6020 13188 6030
rect 13132 5926 13188 5964
rect 13244 5906 13300 5918
rect 13244 5854 13246 5906
rect 13298 5854 13300 5906
rect 13244 5796 13300 5854
rect 13020 5740 13300 5796
rect 12796 5070 12798 5122
rect 12850 5070 12852 5122
rect 11452 3332 11620 3388
rect 12124 3332 12292 3388
rect 11452 800 11508 3332
rect 12124 800 12180 3332
rect 12796 800 12852 5070
rect 12908 4788 12964 4798
rect 12908 4338 12964 4732
rect 12908 4286 12910 4338
rect 12962 4286 12964 4338
rect 12908 4274 12964 4286
rect 13132 3444 13188 3454
rect 13356 3444 13412 7532
rect 13580 7476 13636 8204
rect 13916 8034 13972 8876
rect 14028 8148 14084 8158
rect 14028 8054 14084 8092
rect 14252 8146 14308 8158
rect 14252 8094 14254 8146
rect 14306 8094 14308 8146
rect 13916 7982 13918 8034
rect 13970 7982 13972 8034
rect 13916 7970 13972 7982
rect 14252 7700 14308 8094
rect 14700 8036 14756 8046
rect 14252 7634 14308 7644
rect 14588 8034 14756 8036
rect 14588 7982 14702 8034
rect 14754 7982 14756 8034
rect 14588 7980 14756 7982
rect 14588 7924 14644 7980
rect 14700 7970 14756 7980
rect 13692 7476 13748 7486
rect 13580 7474 13748 7476
rect 13580 7422 13694 7474
rect 13746 7422 13748 7474
rect 13580 7420 13748 7422
rect 13580 6804 13636 7420
rect 13692 7410 13748 7420
rect 13580 6738 13636 6748
rect 14476 7362 14532 7374
rect 14476 7310 14478 7362
rect 14530 7310 14532 7362
rect 13692 6692 13748 6702
rect 13692 6598 13748 6636
rect 13692 6468 13748 6478
rect 13580 6018 13636 6030
rect 13580 5966 13582 6018
rect 13634 5966 13636 6018
rect 13468 5684 13524 5694
rect 13468 5122 13524 5628
rect 13580 5348 13636 5966
rect 13580 5282 13636 5292
rect 13468 5070 13470 5122
rect 13522 5070 13524 5122
rect 13468 5058 13524 5070
rect 13692 4900 13748 6412
rect 13916 5906 13972 5918
rect 13916 5854 13918 5906
rect 13970 5854 13972 5906
rect 13916 5796 13972 5854
rect 13916 5730 13972 5740
rect 13804 5348 13860 5358
rect 13804 5122 13860 5292
rect 14476 5236 14532 7310
rect 14476 5170 14532 5180
rect 13804 5070 13806 5122
rect 13858 5070 13860 5122
rect 13804 5058 13860 5070
rect 13580 4844 13748 4900
rect 13916 5012 13972 5022
rect 13916 4900 13972 4956
rect 14028 4900 14084 4910
rect 13916 4898 14084 4900
rect 13916 4846 14030 4898
rect 14082 4846 14084 4898
rect 13916 4844 14084 4846
rect 13468 3556 13524 3566
rect 13468 3462 13524 3500
rect 13132 3442 13412 3444
rect 13132 3390 13134 3442
rect 13186 3390 13412 3442
rect 13132 3388 13412 3390
rect 13132 3378 13188 3388
rect 13580 3220 13636 4844
rect 14028 4834 14084 4844
rect 14140 4900 14196 4910
rect 14140 4806 14196 4844
rect 14252 4898 14308 4910
rect 14252 4846 14254 4898
rect 14306 4846 14308 4898
rect 13692 4228 13748 4238
rect 13692 4134 13748 4172
rect 14252 4228 14308 4846
rect 14252 4162 14308 4172
rect 13468 3164 13636 3220
rect 14140 3556 14196 3566
rect 13468 800 13524 3164
rect 14140 800 14196 3500
rect 14252 3556 14308 3566
rect 14588 3556 14644 7868
rect 14700 6468 14756 6478
rect 14700 6374 14756 6412
rect 14812 6244 14868 9100
rect 14924 9042 14980 9324
rect 15932 9380 15988 10446
rect 15932 9314 15988 9324
rect 15036 9268 15092 9278
rect 15036 9174 15092 9212
rect 16044 9268 16100 15092
rect 16156 14308 16212 20188
rect 16268 19794 16324 20412
rect 16268 19742 16270 19794
rect 16322 19742 16324 19794
rect 16268 19730 16324 19742
rect 16380 20356 16436 20366
rect 16268 19122 16324 19134
rect 16268 19070 16270 19122
rect 16322 19070 16324 19122
rect 16268 18676 16324 19070
rect 16380 19012 16436 20300
rect 16492 19234 16548 20526
rect 16604 20130 16660 20636
rect 16716 20690 16772 20702
rect 16716 20638 16718 20690
rect 16770 20638 16772 20690
rect 16716 20580 16772 20638
rect 16716 20514 16772 20524
rect 16604 20078 16606 20130
rect 16658 20078 16660 20130
rect 16604 20066 16660 20078
rect 16828 20130 16884 21196
rect 16940 20356 16996 21308
rect 17276 20580 17332 20590
rect 17276 20486 17332 20524
rect 16940 20290 16996 20300
rect 16828 20078 16830 20130
rect 16882 20078 16884 20130
rect 16828 19572 16884 20078
rect 16828 19506 16884 19516
rect 17388 19460 17444 19470
rect 16716 19348 16772 19358
rect 16716 19346 17332 19348
rect 16716 19294 16718 19346
rect 16770 19294 17332 19346
rect 16716 19292 17332 19294
rect 16716 19282 16772 19292
rect 16492 19182 16494 19234
rect 16546 19182 16548 19234
rect 16492 19124 16548 19182
rect 17276 19234 17332 19292
rect 17276 19182 17278 19234
rect 17330 19182 17332 19234
rect 17276 19170 17332 19182
rect 16492 19068 16660 19124
rect 16380 18956 16548 19012
rect 16268 18610 16324 18620
rect 16268 18452 16324 18462
rect 16268 18450 16436 18452
rect 16268 18398 16270 18450
rect 16322 18398 16436 18450
rect 16268 18396 16436 18398
rect 16268 18386 16324 18396
rect 16268 18228 16324 18238
rect 16268 18134 16324 18172
rect 16380 17780 16436 18396
rect 16380 17714 16436 17724
rect 16268 17444 16324 17454
rect 16268 16882 16324 17388
rect 16268 16830 16270 16882
rect 16322 16830 16324 16882
rect 16268 16818 16324 16830
rect 16492 16660 16548 18956
rect 16604 18562 16660 19068
rect 16828 19122 16884 19134
rect 16828 19070 16830 19122
rect 16882 19070 16884 19122
rect 16716 19012 16772 19022
rect 16828 19012 16884 19070
rect 17388 19122 17444 19404
rect 17500 19236 17556 21532
rect 18172 21474 18228 21486
rect 18172 21422 18174 21474
rect 18226 21422 18228 21474
rect 18060 20580 18116 20590
rect 17836 19236 17892 19246
rect 17500 19234 17892 19236
rect 17500 19182 17838 19234
rect 17890 19182 17892 19234
rect 17500 19180 17892 19182
rect 17836 19170 17892 19180
rect 17388 19070 17390 19122
rect 17442 19070 17444 19122
rect 17388 19058 17444 19070
rect 16940 19012 16996 19022
rect 16828 18956 16940 19012
rect 16716 18918 16772 18956
rect 16940 18946 16996 18956
rect 17612 19010 17668 19022
rect 17612 18958 17614 19010
rect 17666 18958 17668 19010
rect 16604 18510 16606 18562
rect 16658 18510 16660 18562
rect 16604 17106 16660 18510
rect 17276 18788 17332 18798
rect 16604 17054 16606 17106
rect 16658 17054 16660 17106
rect 16604 17042 16660 17054
rect 16828 17780 16884 17790
rect 16828 16884 16884 17724
rect 16940 17556 16996 17566
rect 16996 17500 17108 17556
rect 16940 17490 16996 17500
rect 16828 16818 16884 16828
rect 16268 16604 16548 16660
rect 16940 16772 16996 16782
rect 16268 15202 16324 16604
rect 16940 16100 16996 16716
rect 16604 16098 16996 16100
rect 16604 16046 16942 16098
rect 16994 16046 16996 16098
rect 16604 16044 16996 16046
rect 16492 15876 16548 15886
rect 16380 15428 16436 15438
rect 16380 15334 16436 15372
rect 16268 15150 16270 15202
rect 16322 15150 16324 15202
rect 16268 15138 16324 15150
rect 16268 14532 16324 14542
rect 16492 14532 16548 15820
rect 16604 15426 16660 16044
rect 16940 16034 16996 16044
rect 17052 15876 17108 17500
rect 17276 16212 17332 18732
rect 17500 18338 17556 18350
rect 17500 18286 17502 18338
rect 17554 18286 17556 18338
rect 17500 17668 17556 18286
rect 17500 17602 17556 17612
rect 17500 17444 17556 17454
rect 17500 17350 17556 17388
rect 17612 17220 17668 18958
rect 17836 17556 17892 17566
rect 17836 17462 17892 17500
rect 17612 17154 17668 17164
rect 17948 17444 18004 17454
rect 17500 16882 17556 16894
rect 17500 16830 17502 16882
rect 17554 16830 17556 16882
rect 17500 16772 17556 16830
rect 17948 16882 18004 17388
rect 17948 16830 17950 16882
rect 18002 16830 18004 16882
rect 17948 16818 18004 16830
rect 17500 16706 17556 16716
rect 17276 15986 17332 16156
rect 17276 15934 17278 15986
rect 17330 15934 17332 15986
rect 17276 15922 17332 15934
rect 17388 15988 17444 15998
rect 16604 15374 16606 15426
rect 16658 15374 16660 15426
rect 16604 15362 16660 15374
rect 16828 15820 17108 15876
rect 16268 14530 16492 14532
rect 16268 14478 16270 14530
rect 16322 14478 16492 14530
rect 16268 14476 16492 14478
rect 16268 14466 16324 14476
rect 16492 14466 16548 14476
rect 16604 14530 16660 14542
rect 16604 14478 16606 14530
rect 16658 14478 16660 14530
rect 16604 14308 16660 14478
rect 16156 14252 16660 14308
rect 16716 14308 16772 14318
rect 16716 14214 16772 14252
rect 16604 13634 16660 13646
rect 16604 13582 16606 13634
rect 16658 13582 16660 13634
rect 16604 13524 16660 13582
rect 16604 13458 16660 13468
rect 16268 13076 16324 13086
rect 16268 10612 16324 13020
rect 16716 12852 16772 12862
rect 16716 12402 16772 12796
rect 16716 12350 16718 12402
rect 16770 12350 16772 12402
rect 16716 12338 16772 12350
rect 16604 12068 16660 12078
rect 16604 11974 16660 12012
rect 16492 11956 16548 11966
rect 16492 11862 16548 11900
rect 16380 10836 16436 10846
rect 16828 10836 16884 15820
rect 17276 15652 17332 15662
rect 16940 15204 16996 15214
rect 16940 14530 16996 15148
rect 16940 14478 16942 14530
rect 16994 14478 16996 14530
rect 16940 14466 16996 14478
rect 17276 14530 17332 15596
rect 17388 15316 17444 15932
rect 17388 15222 17444 15260
rect 17724 15428 17780 15438
rect 17724 14644 17780 15372
rect 18060 15148 18116 20524
rect 17724 14578 17780 14588
rect 17836 15092 18116 15148
rect 17276 14478 17278 14530
rect 17330 14478 17332 14530
rect 17276 14466 17332 14478
rect 17500 14532 17556 14542
rect 17500 13970 17556 14476
rect 17500 13918 17502 13970
rect 17554 13918 17556 13970
rect 17500 13906 17556 13918
rect 17836 13300 17892 15092
rect 17948 14418 18004 14430
rect 17948 14366 17950 14418
rect 18002 14366 18004 14418
rect 17948 13970 18004 14366
rect 17948 13918 17950 13970
rect 18002 13918 18004 13970
rect 17948 13906 18004 13918
rect 17500 13244 17892 13300
rect 16940 10836 16996 10846
rect 17500 10836 17556 13244
rect 17724 13074 17780 13086
rect 17724 13022 17726 13074
rect 17778 13022 17780 13074
rect 17724 12964 17780 13022
rect 18172 13076 18228 21422
rect 18284 20468 18340 23436
rect 18396 22932 18452 23662
rect 18396 22866 18452 22876
rect 18284 20402 18340 20412
rect 18508 20244 18564 26124
rect 18620 24948 18676 26798
rect 18732 26962 18788 26974
rect 18732 26910 18734 26962
rect 18786 26910 18788 26962
rect 18732 25506 18788 26910
rect 18844 26180 18900 27694
rect 18844 26114 18900 26124
rect 19180 27074 19236 27086
rect 19180 27022 19182 27074
rect 19234 27022 19236 27074
rect 18732 25454 18734 25506
rect 18786 25454 18788 25506
rect 18732 25396 18788 25454
rect 19180 25396 19236 27022
rect 19292 26290 19348 30828
rect 19516 30790 19572 30828
rect 19628 30434 19684 31052
rect 19628 30382 19630 30434
rect 19682 30382 19684 30434
rect 19404 30322 19460 30334
rect 19404 30270 19406 30322
rect 19458 30270 19460 30322
rect 19404 30212 19460 30270
rect 19628 30324 19684 30382
rect 19628 30258 19684 30268
rect 19740 30884 19796 31164
rect 19404 30146 19460 30156
rect 19740 30100 19796 30828
rect 19964 30212 20020 30222
rect 19964 30118 20020 30156
rect 19516 30044 19796 30100
rect 19404 29988 19460 29998
rect 19404 29894 19460 29932
rect 19404 29652 19460 29662
rect 19404 29558 19460 29596
rect 19516 29538 19572 30044
rect 19836 29820 20100 29830
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 19836 29754 20100 29764
rect 19516 29486 19518 29538
rect 19570 29486 19572 29538
rect 19516 29474 19572 29486
rect 20188 29428 20244 31500
rect 20300 30436 20356 30446
rect 20300 30342 20356 30380
rect 20412 29652 20468 31726
rect 20524 31220 20580 31948
rect 20524 31154 20580 31164
rect 20636 31778 20692 31790
rect 20636 31726 20638 31778
rect 20690 31726 20692 31778
rect 20524 30996 20580 31006
rect 20524 30210 20580 30940
rect 20636 30322 20692 31726
rect 21308 31108 21364 32398
rect 21420 31892 21476 33740
rect 21756 33572 21812 33582
rect 21756 33346 21812 33516
rect 21756 33294 21758 33346
rect 21810 33294 21812 33346
rect 21756 33282 21812 33294
rect 21420 31798 21476 31836
rect 21756 31892 21812 31902
rect 21364 31052 21476 31108
rect 21308 31042 21364 31052
rect 21308 30882 21364 30894
rect 21308 30830 21310 30882
rect 21362 30830 21364 30882
rect 20636 30270 20638 30322
rect 20690 30270 20692 30322
rect 20636 30258 20692 30270
rect 20748 30548 20804 30558
rect 20524 30158 20526 30210
rect 20578 30158 20580 30210
rect 20524 29988 20580 30158
rect 20748 30210 20804 30492
rect 21308 30548 21364 30830
rect 21308 30482 21364 30492
rect 21420 30212 21476 31052
rect 21532 30994 21588 31006
rect 21532 30942 21534 30994
rect 21586 30942 21588 30994
rect 21532 30884 21588 30942
rect 21756 30994 21812 31836
rect 21756 30942 21758 30994
rect 21810 30942 21812 30994
rect 21756 30930 21812 30942
rect 21532 30818 21588 30828
rect 21868 30660 21924 34078
rect 22540 34132 22596 34142
rect 22316 34018 22372 34030
rect 22316 33966 22318 34018
rect 22370 33966 22372 34018
rect 22316 33572 22372 33966
rect 22316 33506 22372 33516
rect 22204 33346 22260 33358
rect 22204 33294 22206 33346
rect 22258 33294 22260 33346
rect 21980 32676 22036 32686
rect 21980 32582 22036 32620
rect 22092 32564 22148 32574
rect 22092 32470 22148 32508
rect 21980 32340 22036 32350
rect 22204 32340 22260 33294
rect 21980 32338 22260 32340
rect 21980 32286 21982 32338
rect 22034 32286 22260 32338
rect 21980 32284 22260 32286
rect 22316 32676 22372 32686
rect 21980 32274 22036 32284
rect 22204 31780 22260 31790
rect 22316 31780 22372 32620
rect 22204 31778 22372 31780
rect 22204 31726 22206 31778
rect 22258 31726 22372 31778
rect 22204 31724 22372 31726
rect 22428 31892 22484 31902
rect 22204 30660 22260 31724
rect 22428 31666 22484 31836
rect 22428 31614 22430 31666
rect 22482 31614 22484 31666
rect 22428 31602 22484 31614
rect 20748 30158 20750 30210
rect 20802 30158 20804 30210
rect 20748 30146 20804 30158
rect 21196 30156 21476 30212
rect 21532 30604 21924 30660
rect 22092 30604 22204 30660
rect 20524 29922 20580 29932
rect 20636 30100 20692 30110
rect 20412 29586 20468 29596
rect 20524 29652 20580 29662
rect 20636 29652 20692 30044
rect 20524 29650 20692 29652
rect 20524 29598 20526 29650
rect 20578 29598 20692 29650
rect 20524 29596 20692 29598
rect 20524 29586 20580 29596
rect 20188 29362 20244 29372
rect 20076 29316 20132 29326
rect 20076 29222 20132 29260
rect 20636 29092 20692 29596
rect 20636 29026 20692 29036
rect 21084 29316 21140 29326
rect 19740 28980 19796 28990
rect 19740 28754 19796 28924
rect 20412 28980 20468 28990
rect 19740 28702 19742 28754
rect 19794 28702 19796 28754
rect 19740 28690 19796 28702
rect 20188 28868 20244 28878
rect 20188 28642 20244 28812
rect 20412 28754 20468 28924
rect 20412 28702 20414 28754
rect 20466 28702 20468 28754
rect 20412 28690 20468 28702
rect 20188 28590 20190 28642
rect 20242 28590 20244 28642
rect 20188 28578 20244 28590
rect 20748 28532 20804 28542
rect 20636 28530 20804 28532
rect 20636 28478 20750 28530
rect 20802 28478 20804 28530
rect 20636 28476 20804 28478
rect 19836 28252 20100 28262
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 19836 28186 20100 28196
rect 20300 27746 20356 27758
rect 20300 27694 20302 27746
rect 20354 27694 20356 27746
rect 20188 27074 20244 27086
rect 20188 27022 20190 27074
rect 20242 27022 20244 27074
rect 19404 26852 19460 26862
rect 19404 26850 19684 26852
rect 19404 26798 19406 26850
rect 19458 26798 19684 26850
rect 19404 26796 19684 26798
rect 19404 26786 19460 26796
rect 19628 26516 19684 26796
rect 19836 26684 20100 26694
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 19836 26618 20100 26628
rect 19628 26460 20020 26516
rect 19964 26402 20020 26460
rect 19964 26350 19966 26402
rect 20018 26350 20020 26402
rect 19964 26338 20020 26350
rect 19292 26238 19294 26290
rect 19346 26238 19348 26290
rect 19292 25620 19348 26238
rect 20188 26180 20244 27022
rect 19292 25554 19348 25564
rect 19852 25844 19908 25854
rect 19852 25508 19908 25788
rect 19516 25396 19572 25406
rect 19180 25394 19572 25396
rect 19180 25342 19518 25394
rect 19570 25342 19572 25394
rect 19180 25340 19572 25342
rect 18732 25330 18788 25340
rect 19516 25330 19572 25340
rect 18844 25282 18900 25294
rect 18844 25230 18846 25282
rect 18898 25230 18900 25282
rect 18844 25172 18900 25230
rect 19068 25284 19124 25294
rect 19852 25284 19908 25452
rect 20188 25396 20244 26124
rect 20188 25330 20244 25340
rect 19068 25282 19236 25284
rect 19068 25230 19070 25282
rect 19122 25230 19236 25282
rect 19068 25228 19236 25230
rect 19068 25218 19124 25228
rect 18844 25106 18900 25116
rect 19068 24948 19124 24958
rect 18620 24946 19124 24948
rect 18620 24894 19070 24946
rect 19122 24894 19124 24946
rect 18620 24892 19124 24894
rect 19068 24882 19124 24892
rect 19180 24724 19236 25228
rect 19628 25228 19908 25284
rect 20300 25284 20356 27694
rect 20524 27074 20580 27086
rect 20524 27022 20526 27074
rect 20578 27022 20580 27074
rect 20524 26852 20580 27022
rect 20412 26796 20580 26852
rect 20412 25844 20468 26796
rect 20412 25778 20468 25788
rect 20636 25508 20692 28476
rect 20748 28466 20804 28476
rect 20748 27188 20804 27198
rect 20748 27094 20804 27132
rect 20524 25506 20692 25508
rect 20524 25454 20638 25506
rect 20690 25454 20692 25506
rect 20524 25452 20692 25454
rect 20412 25396 20468 25406
rect 20412 25302 20468 25340
rect 19404 25172 19460 25182
rect 19628 25172 19684 25228
rect 20300 25218 20356 25228
rect 20524 25172 20580 25452
rect 20636 25442 20692 25452
rect 19460 25116 19684 25172
rect 19836 25116 20100 25126
rect 19404 24946 19460 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20412 25116 20580 25172
rect 20412 25060 20468 25116
rect 19836 25050 20100 25060
rect 19404 24894 19406 24946
rect 19458 24894 19460 24946
rect 19404 24882 19460 24894
rect 20300 25004 20468 25060
rect 18956 24668 19236 24724
rect 18732 23716 18788 23726
rect 18732 23714 18900 23716
rect 18732 23662 18734 23714
rect 18786 23662 18900 23714
rect 18732 23660 18900 23662
rect 18732 23650 18788 23660
rect 18844 23266 18900 23660
rect 18844 23214 18846 23266
rect 18898 23214 18900 23266
rect 18844 23202 18900 23214
rect 18956 20804 19012 24668
rect 19852 24612 19908 24622
rect 19852 24164 19908 24556
rect 19628 24162 19908 24164
rect 19628 24110 19854 24162
rect 19906 24110 19908 24162
rect 19628 24108 19908 24110
rect 19068 23828 19124 23838
rect 19516 23828 19572 23838
rect 19068 23826 19572 23828
rect 19068 23774 19070 23826
rect 19122 23774 19518 23826
rect 19570 23774 19572 23826
rect 19068 23772 19572 23774
rect 19068 23762 19124 23772
rect 19516 23762 19572 23772
rect 19068 22596 19124 22606
rect 19628 22596 19684 24108
rect 19852 24098 19908 24108
rect 20300 23938 20356 25004
rect 20300 23886 20302 23938
rect 20354 23886 20356 23938
rect 20300 23874 20356 23886
rect 20412 24722 20468 24734
rect 20412 24670 20414 24722
rect 20466 24670 20468 24722
rect 20412 23828 20468 24670
rect 20748 24722 20804 24734
rect 20748 24670 20750 24722
rect 20802 24670 20804 24722
rect 20748 24612 20804 24670
rect 20748 24546 20804 24556
rect 20636 23828 20692 23838
rect 20412 23826 20692 23828
rect 20412 23774 20638 23826
rect 20690 23774 20692 23826
rect 20412 23772 20692 23774
rect 19836 23548 20100 23558
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 19836 23482 20100 23492
rect 20636 23044 20692 23772
rect 20972 23044 21028 23054
rect 20636 23042 21028 23044
rect 20636 22990 20974 23042
rect 21026 22990 21028 23042
rect 20636 22988 21028 22990
rect 20972 22978 21028 22988
rect 19124 22540 19684 22596
rect 19068 22482 19124 22540
rect 19068 22430 19070 22482
rect 19122 22430 19124 22482
rect 19068 22418 19124 22430
rect 21084 22372 21140 29260
rect 21196 28532 21252 30156
rect 21420 29986 21476 29998
rect 21420 29934 21422 29986
rect 21474 29934 21476 29986
rect 21308 29428 21364 29438
rect 21420 29428 21476 29934
rect 21364 29372 21476 29428
rect 21308 29314 21364 29372
rect 21308 29262 21310 29314
rect 21362 29262 21364 29314
rect 21308 29250 21364 29262
rect 21196 27860 21252 28476
rect 21308 29092 21364 29102
rect 21308 28530 21364 29036
rect 21308 28478 21310 28530
rect 21362 28478 21364 28530
rect 21308 28466 21364 28478
rect 21532 28418 21588 30604
rect 21756 30324 21812 30362
rect 21756 30258 21812 30268
rect 21868 30212 21924 30222
rect 21980 30212 22036 30222
rect 21868 30210 21980 30212
rect 21868 30158 21870 30210
rect 21922 30158 21980 30210
rect 21868 30156 21980 30158
rect 21868 30146 21924 30156
rect 21644 30100 21700 30110
rect 21644 30006 21700 30044
rect 21756 29428 21812 29438
rect 21756 29334 21812 29372
rect 21532 28366 21534 28418
rect 21586 28366 21588 28418
rect 21532 28354 21588 28366
rect 21308 27860 21364 27870
rect 21196 27804 21308 27860
rect 21308 27766 21364 27804
rect 21196 27300 21252 27310
rect 21196 26516 21252 27244
rect 21980 27076 22036 30156
rect 22092 29428 22148 30604
rect 22204 30566 22260 30604
rect 22204 30212 22260 30222
rect 22428 30212 22484 30222
rect 22204 30210 22484 30212
rect 22204 30158 22206 30210
rect 22258 30158 22430 30210
rect 22482 30158 22484 30210
rect 22204 30156 22484 30158
rect 22204 30146 22260 30156
rect 22428 30146 22484 30156
rect 22540 30212 22596 34076
rect 22652 32788 22708 34300
rect 22988 34132 23044 34142
rect 22876 34076 22988 34132
rect 22876 32900 22932 34076
rect 22988 34038 23044 34076
rect 23100 34018 23156 34030
rect 23100 33966 23102 34018
rect 23154 33966 23156 34018
rect 23100 33684 23156 33966
rect 23100 33618 23156 33628
rect 23100 33348 23156 33358
rect 23100 33254 23156 33292
rect 23212 33346 23268 34300
rect 23212 33294 23214 33346
rect 23266 33294 23268 33346
rect 23212 33282 23268 33294
rect 22988 33124 23044 33134
rect 22988 33030 23044 33068
rect 22876 32844 23268 32900
rect 22764 32788 22820 32798
rect 22652 32786 22820 32788
rect 22652 32734 22766 32786
rect 22818 32734 22820 32786
rect 22652 32732 22820 32734
rect 22764 32722 22820 32732
rect 23212 32674 23268 32844
rect 23324 32788 23380 34412
rect 23884 34356 23940 37100
rect 23996 35364 24052 37324
rect 24220 37314 24276 37324
rect 24332 37268 24388 37278
rect 24388 37212 24500 37268
rect 24332 37174 24388 37212
rect 24220 37042 24276 37054
rect 24220 36990 24222 37042
rect 24274 36990 24276 37042
rect 24108 36484 24164 36494
rect 24108 36390 24164 36428
rect 24220 35810 24276 36990
rect 24332 35924 24388 35934
rect 24332 35830 24388 35868
rect 24220 35758 24222 35810
rect 24274 35758 24276 35810
rect 24220 35746 24276 35758
rect 23996 35298 24052 35308
rect 24444 35308 24500 37212
rect 24780 36372 24836 36382
rect 24556 36370 24836 36372
rect 24556 36318 24782 36370
rect 24834 36318 24836 36370
rect 24556 36316 24836 36318
rect 24556 35922 24612 36316
rect 24780 36306 24836 36316
rect 24556 35870 24558 35922
rect 24610 35870 24612 35922
rect 24556 35858 24612 35870
rect 24444 35252 24724 35308
rect 24668 34802 24724 35252
rect 24668 34750 24670 34802
rect 24722 34750 24724 34802
rect 24108 34692 24164 34702
rect 24108 34598 24164 34636
rect 24668 34692 24724 34750
rect 24668 34626 24724 34636
rect 24780 34690 24836 34702
rect 25004 34692 25060 34702
rect 24780 34638 24782 34690
rect 24834 34638 24836 34690
rect 24780 34356 24836 34638
rect 23884 34300 24276 34356
rect 24220 34244 24276 34300
rect 24668 34300 24836 34356
rect 24892 34690 25060 34692
rect 24892 34638 25006 34690
rect 25058 34638 25060 34690
rect 24892 34636 25060 34638
rect 24220 34188 24388 34244
rect 24108 34130 24164 34142
rect 24108 34078 24110 34130
rect 24162 34078 24164 34130
rect 23772 34018 23828 34030
rect 23772 33966 23774 34018
rect 23826 33966 23828 34018
rect 23772 33908 23828 33966
rect 23772 33852 24052 33908
rect 23772 33684 23828 33694
rect 23660 33346 23716 33358
rect 23660 33294 23662 33346
rect 23714 33294 23716 33346
rect 23324 32732 23604 32788
rect 23212 32622 23214 32674
rect 23266 32622 23268 32674
rect 22988 32340 23044 32350
rect 22764 31892 22820 31902
rect 22652 31836 22764 31892
rect 22652 31444 22708 31836
rect 22764 31826 22820 31836
rect 22764 31668 22820 31678
rect 22764 31666 22932 31668
rect 22764 31614 22766 31666
rect 22818 31614 22932 31666
rect 22764 31612 22932 31614
rect 22764 31602 22820 31612
rect 22652 31388 22820 31444
rect 22652 31106 22708 31118
rect 22652 31054 22654 31106
rect 22706 31054 22708 31106
rect 22652 30884 22708 31054
rect 22652 30818 22708 30828
rect 22540 30146 22596 30156
rect 22764 30210 22820 31388
rect 22876 30884 22932 31612
rect 22988 31554 23044 32284
rect 23100 31892 23156 31902
rect 23100 31778 23156 31836
rect 23100 31726 23102 31778
rect 23154 31726 23156 31778
rect 23100 31714 23156 31726
rect 23212 31778 23268 32622
rect 23212 31726 23214 31778
rect 23266 31726 23268 31778
rect 23212 31714 23268 31726
rect 23324 32562 23380 32574
rect 23324 32510 23326 32562
rect 23378 32510 23380 32562
rect 23324 32452 23380 32510
rect 23436 32564 23492 32574
rect 23436 32470 23492 32508
rect 22988 31502 22990 31554
rect 23042 31502 23044 31554
rect 22988 31490 23044 31502
rect 22988 31220 23044 31230
rect 23324 31220 23380 32396
rect 23548 31220 23604 32732
rect 23660 32228 23716 33294
rect 23660 32162 23716 32172
rect 23772 33124 23828 33628
rect 23884 33348 23940 33358
rect 23884 33254 23940 33292
rect 23996 33236 24052 33852
rect 24108 33460 24164 34078
rect 24332 34130 24388 34188
rect 24332 34078 24334 34130
rect 24386 34078 24388 34130
rect 24220 34020 24276 34030
rect 24220 33926 24276 33964
rect 24332 33684 24388 34078
rect 24668 34132 24724 34300
rect 24668 34066 24724 34076
rect 24780 34132 24836 34142
rect 24892 34132 24948 34636
rect 25004 34626 25060 34636
rect 24780 34130 24948 34132
rect 24780 34078 24782 34130
rect 24834 34078 24948 34130
rect 24780 34076 24948 34078
rect 24780 34066 24836 34076
rect 24332 33618 24388 33628
rect 24892 33684 24948 33694
rect 24332 33460 24388 33470
rect 24108 33458 24388 33460
rect 24108 33406 24334 33458
rect 24386 33406 24388 33458
rect 24108 33404 24388 33406
rect 24332 33394 24388 33404
rect 24220 33236 24276 33246
rect 23996 33180 24220 33236
rect 24220 33142 24276 33180
rect 23772 31556 23828 33068
rect 24444 33124 24500 33134
rect 24444 33030 24500 33068
rect 24892 33122 24948 33628
rect 24892 33070 24894 33122
rect 24946 33070 24948 33122
rect 23884 32676 23940 32686
rect 23884 32582 23940 32620
rect 23996 32674 24052 32686
rect 23996 32622 23998 32674
rect 24050 32622 24052 32674
rect 23996 31892 24052 32622
rect 24220 32564 24276 32574
rect 24220 32562 24500 32564
rect 24220 32510 24222 32562
rect 24274 32510 24500 32562
rect 24220 32508 24500 32510
rect 24220 32498 24276 32508
rect 23996 31826 24052 31836
rect 24220 31892 24276 31902
rect 23996 31556 24052 31566
rect 23772 31554 23940 31556
rect 23772 31502 23774 31554
rect 23826 31502 23940 31554
rect 23772 31500 23940 31502
rect 23772 31490 23828 31500
rect 22988 31218 23380 31220
rect 22988 31166 22990 31218
rect 23042 31166 23380 31218
rect 22988 31164 23380 31166
rect 22988 31154 23044 31164
rect 22876 30818 22932 30828
rect 22764 30158 22766 30210
rect 22818 30158 22820 30210
rect 22764 30146 22820 30158
rect 23212 30210 23268 30222
rect 23212 30158 23214 30210
rect 23266 30158 23268 30210
rect 22652 29988 22708 29998
rect 22652 29894 22708 29932
rect 22764 29650 22820 29662
rect 22764 29598 22766 29650
rect 22818 29598 22820 29650
rect 22092 29362 22148 29372
rect 22652 29538 22708 29550
rect 22652 29486 22654 29538
rect 22706 29486 22708 29538
rect 22652 29204 22708 29486
rect 22652 29138 22708 29148
rect 22764 28532 22820 29598
rect 22764 28466 22820 28476
rect 22876 28812 23156 28868
rect 22204 27972 22260 27982
rect 22876 27972 22932 28812
rect 22204 27878 22260 27916
rect 22764 27916 22932 27972
rect 22988 28644 23044 28654
rect 22764 27858 22820 27916
rect 22988 27860 23044 28588
rect 23100 28642 23156 28812
rect 23100 28590 23102 28642
rect 23154 28590 23156 28642
rect 23100 28578 23156 28590
rect 22764 27806 22766 27858
rect 22818 27806 22820 27858
rect 22764 27188 22820 27806
rect 22764 27122 22820 27132
rect 22876 27858 23044 27860
rect 22876 27806 22990 27858
rect 23042 27806 23044 27858
rect 22876 27804 23044 27806
rect 22092 27076 22148 27086
rect 21980 27020 22092 27076
rect 21420 26964 21476 26974
rect 21756 26964 21812 26974
rect 21308 26962 21812 26964
rect 21308 26910 21422 26962
rect 21474 26910 21758 26962
rect 21810 26910 21812 26962
rect 21308 26908 21812 26910
rect 22092 26962 22148 27020
rect 22092 26910 22094 26962
rect 22146 26910 22148 26962
rect 21308 26852 21364 26908
rect 21420 26898 21476 26908
rect 21756 26852 22036 26908
rect 22092 26898 22148 26910
rect 22428 26962 22484 26974
rect 22428 26910 22430 26962
rect 22482 26910 22484 26962
rect 22428 26908 22484 26910
rect 22428 26852 22708 26908
rect 21308 26786 21364 26796
rect 21980 26628 22036 26852
rect 21980 26572 22484 26628
rect 21196 26450 21252 26460
rect 22428 26514 22484 26572
rect 22428 26462 22430 26514
rect 22482 26462 22484 26514
rect 22428 26450 22484 26462
rect 22652 26290 22708 26852
rect 22652 26238 22654 26290
rect 22706 26238 22708 26290
rect 22092 26180 22148 26190
rect 22092 26086 22148 26124
rect 21420 25844 21476 25854
rect 21308 25788 21420 25844
rect 21308 24834 21364 25788
rect 21420 25778 21476 25788
rect 22316 25620 22372 25630
rect 22316 25526 22372 25564
rect 21420 25508 21476 25518
rect 21420 25414 21476 25452
rect 21308 24782 21310 24834
rect 21362 24782 21364 24834
rect 21308 24770 21364 24782
rect 22428 25284 22484 25294
rect 21868 24612 21924 24622
rect 21868 24518 21924 24556
rect 22428 23938 22484 25228
rect 22428 23886 22430 23938
rect 22482 23886 22484 23938
rect 22428 23492 22484 23886
rect 22428 23426 22484 23436
rect 22316 23154 22372 23166
rect 22316 23102 22318 23154
rect 22370 23102 22372 23154
rect 22316 22594 22372 23102
rect 22316 22542 22318 22594
rect 22370 22542 22372 22594
rect 22316 22530 22372 22542
rect 22092 22372 22148 22382
rect 21084 22306 21140 22316
rect 21868 22370 22484 22372
rect 21868 22318 22094 22370
rect 22146 22318 22484 22370
rect 21868 22316 22484 22318
rect 21756 22260 21812 22270
rect 21756 22166 21812 22204
rect 20188 22148 20244 22158
rect 19836 21980 20100 21990
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 19836 21914 20100 21924
rect 18956 20738 19012 20748
rect 19836 20412 20100 20422
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 19836 20346 20100 20356
rect 18508 20188 18900 20244
rect 18396 20132 18452 20142
rect 18396 20130 18676 20132
rect 18396 20078 18398 20130
rect 18450 20078 18676 20130
rect 18396 20076 18676 20078
rect 18396 20066 18452 20076
rect 18620 19346 18676 20076
rect 18620 19294 18622 19346
rect 18674 19294 18676 19346
rect 18620 19282 18676 19294
rect 18732 20018 18788 20030
rect 18732 19966 18734 20018
rect 18786 19966 18788 20018
rect 18620 18676 18676 18686
rect 18732 18676 18788 19966
rect 18844 19348 18900 20188
rect 18844 19282 18900 19292
rect 18956 20132 19012 20142
rect 19740 20132 19796 20142
rect 18620 18674 18788 18676
rect 18620 18622 18622 18674
rect 18674 18622 18788 18674
rect 18620 18620 18788 18622
rect 18620 18610 18676 18620
rect 18956 18450 19012 20076
rect 19628 20076 19740 20132
rect 19516 18676 19572 18686
rect 19516 18562 19572 18620
rect 19516 18510 19518 18562
rect 19570 18510 19572 18562
rect 19516 18498 19572 18510
rect 18956 18398 18958 18450
rect 19010 18398 19012 18450
rect 18956 18386 19012 18398
rect 19628 18452 19684 20076
rect 19740 20066 19796 20076
rect 19836 18844 20100 18854
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 19836 18778 20100 18788
rect 20188 18676 20244 22092
rect 20636 21812 20692 21822
rect 20636 21718 20692 21756
rect 21756 21700 21812 21710
rect 21868 21700 21924 22316
rect 22092 22306 22148 22316
rect 22428 22260 22484 22316
rect 22540 22260 22596 22270
rect 22428 22204 22540 22260
rect 22540 22166 22596 22204
rect 21756 21698 21924 21700
rect 21756 21646 21758 21698
rect 21810 21646 21924 21698
rect 21756 21644 21924 21646
rect 21980 22146 22036 22158
rect 22316 22148 22372 22158
rect 21980 22094 21982 22146
rect 22034 22094 22036 22146
rect 21756 21634 21812 21644
rect 20300 21588 20356 21598
rect 20300 21474 20356 21532
rect 20300 21422 20302 21474
rect 20354 21422 20356 21474
rect 20300 21410 20356 21422
rect 20860 21588 20916 21598
rect 21420 21588 21476 21598
rect 20860 21586 21476 21588
rect 20860 21534 20862 21586
rect 20914 21534 21422 21586
rect 21474 21534 21476 21586
rect 20860 21532 21476 21534
rect 20412 19794 20468 19806
rect 20412 19742 20414 19794
rect 20466 19742 20468 19794
rect 20412 19236 20468 19742
rect 20748 19796 20804 19806
rect 20748 19702 20804 19740
rect 20412 19170 20468 19180
rect 20748 19346 20804 19358
rect 20748 19294 20750 19346
rect 20802 19294 20804 19346
rect 20748 18676 20804 19294
rect 20188 18620 20356 18676
rect 19628 18450 20132 18452
rect 19628 18398 19630 18450
rect 19682 18398 20132 18450
rect 19628 18396 20132 18398
rect 19628 18386 19684 18396
rect 20076 17778 20132 18396
rect 20076 17726 20078 17778
rect 20130 17726 20132 17778
rect 19740 17668 19796 17678
rect 19628 17612 19740 17668
rect 18956 17554 19012 17566
rect 18956 17502 18958 17554
rect 19010 17502 19012 17554
rect 18284 17444 18340 17454
rect 18284 17350 18340 17388
rect 18732 16884 18788 16894
rect 18396 16882 18788 16884
rect 18396 16830 18734 16882
rect 18786 16830 18788 16882
rect 18396 16828 18788 16830
rect 18284 16100 18340 16110
rect 18284 15428 18340 16044
rect 18396 15652 18452 16828
rect 18732 16818 18788 16828
rect 18956 16322 19012 17502
rect 19292 17444 19348 17454
rect 19292 17442 19572 17444
rect 19292 17390 19294 17442
rect 19346 17390 19572 17442
rect 19292 17388 19572 17390
rect 19292 17378 19348 17388
rect 18956 16270 18958 16322
rect 19010 16270 19012 16322
rect 18956 16258 19012 16270
rect 19292 17220 19348 17230
rect 19292 16322 19348 17164
rect 19516 16994 19572 17388
rect 19628 17108 19684 17612
rect 19740 17574 19796 17612
rect 20076 17444 20132 17726
rect 20076 17388 20244 17444
rect 19836 17276 20100 17286
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 19836 17210 20100 17220
rect 20188 17108 20244 17388
rect 19628 17042 19684 17052
rect 20076 17052 20244 17108
rect 19516 16942 19518 16994
rect 19570 16942 19572 16994
rect 19516 16930 19572 16942
rect 19292 16270 19294 16322
rect 19346 16270 19348 16322
rect 19292 16258 19348 16270
rect 20076 16212 20132 17052
rect 19404 16156 20132 16212
rect 19404 16100 19460 16156
rect 18396 15586 18452 15596
rect 19292 16044 19460 16100
rect 20076 16098 20132 16156
rect 20076 16046 20078 16098
rect 20130 16046 20132 16098
rect 18284 15372 18452 15428
rect 18284 15090 18340 15102
rect 18284 15038 18286 15090
rect 18338 15038 18340 15090
rect 18284 13858 18340 15038
rect 18284 13806 18286 13858
rect 18338 13806 18340 13858
rect 18284 13794 18340 13806
rect 18172 13010 18228 13020
rect 17724 12898 17780 12908
rect 18172 12740 18228 12750
rect 16380 10834 16996 10836
rect 16380 10782 16382 10834
rect 16434 10782 16942 10834
rect 16994 10782 16996 10834
rect 16380 10780 16996 10782
rect 16380 10770 16436 10780
rect 16940 10770 16996 10780
rect 17388 10834 17556 10836
rect 17388 10782 17502 10834
rect 17554 10782 17556 10834
rect 17388 10780 17556 10782
rect 16268 10556 16548 10612
rect 16492 9940 16548 10556
rect 16492 9938 16660 9940
rect 16492 9886 16494 9938
rect 16546 9886 16660 9938
rect 16492 9884 16660 9886
rect 16492 9874 16548 9884
rect 16044 9202 16100 9212
rect 14924 8990 14926 9042
rect 14978 8990 14980 9042
rect 14924 8428 14980 8990
rect 15148 9042 15204 9054
rect 15148 8990 15150 9042
rect 15202 8990 15204 9042
rect 15148 8596 15204 8990
rect 15708 9044 15764 9054
rect 16380 9044 16436 9054
rect 15708 8950 15764 8988
rect 16156 9042 16436 9044
rect 16156 8990 16382 9042
rect 16434 8990 16436 9042
rect 16156 8988 16436 8990
rect 15484 8820 15540 8830
rect 16156 8820 16212 8988
rect 16380 8978 16436 8988
rect 16492 9044 16548 9054
rect 15484 8818 16212 8820
rect 15484 8766 15486 8818
rect 15538 8766 16212 8818
rect 15484 8764 16212 8766
rect 16268 8820 16324 8830
rect 15484 8754 15540 8764
rect 16268 8726 16324 8764
rect 15148 8530 15204 8540
rect 16492 8596 16548 8988
rect 16604 9042 16660 9884
rect 16940 9826 16996 9838
rect 16940 9774 16942 9826
rect 16994 9774 16996 9826
rect 16940 9604 16996 9774
rect 16940 9538 16996 9548
rect 16604 8990 16606 9042
rect 16658 8990 16660 9042
rect 16604 8978 16660 8990
rect 16716 9268 16772 9278
rect 14924 8372 15204 8428
rect 14924 7700 14980 8372
rect 15148 8370 15204 8372
rect 15148 8318 15150 8370
rect 15202 8318 15204 8370
rect 15148 8306 15204 8318
rect 16268 8260 16324 8270
rect 16156 8204 16268 8260
rect 15596 8148 15652 8158
rect 15484 8036 15540 8046
rect 14924 7634 14980 7644
rect 15260 8034 15540 8036
rect 15260 7982 15486 8034
rect 15538 7982 15540 8034
rect 15260 7980 15540 7982
rect 14812 6188 14980 6244
rect 14700 6132 14756 6142
rect 14756 6076 14868 6132
rect 14700 6066 14756 6076
rect 14252 3554 14644 3556
rect 14252 3502 14254 3554
rect 14306 3502 14644 3554
rect 14252 3500 14644 3502
rect 14700 5794 14756 5806
rect 14700 5742 14702 5794
rect 14754 5742 14756 5794
rect 14252 3490 14308 3500
rect 14700 2884 14756 5742
rect 14812 5122 14868 6076
rect 14924 5796 14980 6188
rect 14924 5730 14980 5740
rect 14812 5070 14814 5122
rect 14866 5070 14868 5122
rect 14812 5058 14868 5070
rect 15036 5348 15092 5358
rect 15036 5122 15092 5292
rect 15148 5236 15204 5246
rect 15148 5142 15204 5180
rect 15036 5070 15038 5122
rect 15090 5070 15092 5122
rect 15036 5058 15092 5070
rect 15260 5010 15316 7980
rect 15484 7970 15540 7980
rect 15596 7924 15652 8092
rect 15596 7858 15652 7868
rect 15260 4958 15262 5010
rect 15314 4958 15316 5010
rect 15260 4946 15316 4958
rect 15484 6132 15540 6142
rect 15484 4898 15540 6076
rect 16156 5122 16212 8204
rect 16268 8194 16324 8204
rect 16268 8036 16324 8046
rect 16492 8036 16548 8540
rect 16268 8034 16548 8036
rect 16268 7982 16270 8034
rect 16322 7982 16548 8034
rect 16268 7980 16548 7982
rect 16604 8148 16660 8158
rect 16268 7970 16324 7980
rect 16604 7362 16660 8092
rect 16604 7310 16606 7362
rect 16658 7310 16660 7362
rect 16604 7298 16660 7310
rect 16156 5070 16158 5122
rect 16210 5070 16212 5122
rect 16156 5058 16212 5070
rect 16268 6580 16324 6590
rect 15484 4846 15486 4898
rect 15538 4846 15540 4898
rect 15484 4564 15540 4846
rect 15484 4498 15540 4508
rect 15820 4228 15876 4238
rect 15820 4134 15876 4172
rect 16268 4226 16324 6524
rect 16716 5906 16772 9212
rect 16828 8258 16884 8270
rect 16828 8206 16830 8258
rect 16882 8206 16884 8258
rect 16828 7812 16884 8206
rect 17388 8148 17444 10780
rect 17500 10770 17556 10780
rect 17724 12738 18228 12740
rect 17724 12686 18174 12738
rect 18226 12686 18228 12738
rect 17724 12684 18228 12686
rect 17724 10052 17780 12684
rect 18172 12674 18228 12684
rect 18172 12180 18228 12190
rect 18172 12086 18228 12124
rect 17612 9716 17668 9726
rect 17612 9622 17668 9660
rect 17724 9380 17780 9996
rect 17948 11394 18004 11406
rect 17948 11342 17950 11394
rect 18002 11342 18004 11394
rect 17948 9604 18004 11342
rect 17948 9538 18004 9548
rect 18396 9380 18452 15372
rect 19292 15314 19348 16044
rect 20076 16034 20132 16046
rect 19964 15988 20020 15998
rect 19964 15894 20020 15932
rect 19836 15708 20100 15718
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 19836 15642 20100 15652
rect 19292 15262 19294 15314
rect 19346 15262 19348 15314
rect 19292 15250 19348 15262
rect 19404 15426 19460 15438
rect 19404 15374 19406 15426
rect 19458 15374 19460 15426
rect 18620 15204 18676 15242
rect 18620 15138 18676 15148
rect 19404 15148 19460 15374
rect 19404 15092 20132 15148
rect 20076 14642 20132 15092
rect 20076 14590 20078 14642
rect 20130 14590 20132 14642
rect 20076 14308 20132 14590
rect 20076 14252 20244 14308
rect 19836 14140 20100 14150
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 19836 14074 20100 14084
rect 18732 13972 18788 13982
rect 20188 13972 20244 14252
rect 18732 13878 18788 13916
rect 20076 13916 20244 13972
rect 20076 13860 20132 13916
rect 20076 13794 20132 13804
rect 19180 13636 19236 13646
rect 19180 13542 19236 13580
rect 19628 13634 19684 13646
rect 19628 13582 19630 13634
rect 19682 13582 19684 13634
rect 19068 13524 19124 13534
rect 19068 12740 19124 13468
rect 19404 13524 19460 13534
rect 19404 13430 19460 13468
rect 19628 13076 19684 13582
rect 20076 13636 20132 13646
rect 20076 13186 20132 13580
rect 20076 13134 20078 13186
rect 20130 13134 20132 13186
rect 20076 13122 20132 13134
rect 19628 12982 19684 13020
rect 20076 12852 20132 12862
rect 19628 12850 20132 12852
rect 19628 12798 20078 12850
rect 20130 12798 20132 12850
rect 19628 12796 20132 12798
rect 19180 12740 19236 12750
rect 19068 12684 19180 12740
rect 19180 12646 19236 12684
rect 18620 12402 18676 12414
rect 18620 12350 18622 12402
rect 18674 12350 18676 12402
rect 18508 12068 18564 12078
rect 18508 11974 18564 12012
rect 18620 11506 18676 12350
rect 18620 11454 18622 11506
rect 18674 11454 18676 11506
rect 18620 11442 18676 11454
rect 18732 12404 18788 12414
rect 18732 12178 18788 12348
rect 19516 12292 19572 12302
rect 19404 12290 19572 12292
rect 19404 12238 19518 12290
rect 19570 12238 19572 12290
rect 19404 12236 19572 12238
rect 18732 12126 18734 12178
rect 18786 12126 18788 12178
rect 17500 9324 17780 9380
rect 17500 9266 17556 9324
rect 17500 9214 17502 9266
rect 17554 9214 17556 9266
rect 17500 9202 17556 9214
rect 17724 9268 17780 9324
rect 17948 9324 18452 9380
rect 17780 9212 17892 9268
rect 17724 9202 17780 9212
rect 17836 8372 17892 9212
rect 17948 9266 18004 9324
rect 17948 9214 17950 9266
rect 18002 9214 18004 9266
rect 17948 8820 18004 9214
rect 18396 9156 18452 9166
rect 18396 9062 18452 9100
rect 17948 8754 18004 8764
rect 17948 8372 18004 8382
rect 17892 8370 18004 8372
rect 17892 8318 17950 8370
rect 18002 8318 18004 8370
rect 17892 8316 18004 8318
rect 17836 8278 17892 8316
rect 17948 8306 18004 8316
rect 17388 8082 17444 8092
rect 18732 8148 18788 12126
rect 18956 12180 19012 12190
rect 19292 12180 19348 12190
rect 18956 12178 19348 12180
rect 18956 12126 18958 12178
rect 19010 12126 19294 12178
rect 19346 12126 19348 12178
rect 18956 12124 19348 12126
rect 18956 11956 19012 12124
rect 19292 12114 19348 12124
rect 18956 11890 19012 11900
rect 19404 11396 19460 12236
rect 19516 12226 19572 12236
rect 19516 12068 19572 12078
rect 19516 11974 19572 12012
rect 19516 11396 19572 11406
rect 19404 11340 19516 11396
rect 19516 11330 19572 11340
rect 19628 9940 19684 12796
rect 20076 12786 20132 12796
rect 20188 12850 20244 12862
rect 20188 12798 20190 12850
rect 20242 12798 20244 12850
rect 20188 12740 20244 12798
rect 19836 12572 20100 12582
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 19836 12506 20100 12516
rect 20076 12404 20132 12414
rect 20076 12310 20132 12348
rect 20188 11844 20244 12684
rect 20188 11778 20244 11788
rect 20300 11620 20356 18620
rect 20748 18610 20804 18620
rect 20748 16436 20804 16446
rect 20748 16212 20804 16380
rect 20748 16118 20804 16156
rect 20412 15652 20468 15662
rect 20412 15316 20468 15596
rect 20412 14418 20468 15260
rect 20860 15148 20916 21532
rect 21420 21522 21476 21532
rect 21644 21586 21700 21598
rect 21644 21534 21646 21586
rect 21698 21534 21700 21586
rect 21644 21364 21700 21534
rect 21644 21298 21700 21308
rect 21420 20802 21476 20814
rect 21420 20750 21422 20802
rect 21474 20750 21476 20802
rect 20972 20132 21028 20142
rect 20972 20038 21028 20076
rect 21308 19236 21364 19246
rect 21308 19142 21364 19180
rect 20412 14366 20414 14418
rect 20466 14366 20468 14418
rect 20412 14354 20468 14366
rect 20524 15092 20916 15148
rect 21084 18452 21140 18462
rect 21084 15540 21140 18396
rect 21420 18004 21476 20750
rect 21980 20804 22036 22094
rect 21980 20710 22036 20748
rect 22092 22146 22372 22148
rect 22092 22094 22318 22146
rect 22370 22094 22372 22146
rect 22092 22092 22372 22094
rect 21532 20130 21588 20142
rect 21532 20078 21534 20130
rect 21586 20078 21588 20130
rect 21532 18340 21588 20078
rect 21644 19012 21700 19022
rect 21980 19012 22036 19022
rect 21644 19010 21812 19012
rect 21644 18958 21646 19010
rect 21698 18958 21812 19010
rect 21644 18956 21812 18958
rect 21644 18946 21700 18956
rect 21756 18562 21812 18956
rect 21756 18510 21758 18562
rect 21810 18510 21812 18562
rect 21756 18498 21812 18510
rect 21532 18274 21588 18284
rect 21420 17938 21476 17948
rect 21868 17666 21924 17678
rect 21868 17614 21870 17666
rect 21922 17614 21924 17666
rect 21644 16770 21700 16782
rect 21644 16718 21646 16770
rect 21698 16718 21700 16770
rect 21644 15988 21700 16718
rect 21868 16772 21924 17614
rect 21980 17556 22036 18956
rect 22092 17668 22148 22092
rect 22316 22082 22372 22092
rect 22652 21924 22708 26238
rect 22764 25956 22820 25966
rect 22764 22482 22820 25900
rect 22876 25844 22932 27804
rect 22988 27794 23044 27804
rect 23100 27972 23156 27982
rect 22988 27076 23044 27114
rect 22988 27010 23044 27020
rect 23100 26908 23156 27916
rect 22876 25778 22932 25788
rect 22988 26852 23156 26908
rect 23212 27076 23268 30158
rect 23324 29428 23380 31164
rect 23436 31218 23604 31220
rect 23436 31166 23550 31218
rect 23602 31166 23604 31218
rect 23436 31164 23604 31166
rect 23436 30098 23492 31164
rect 23548 31154 23604 31164
rect 23436 30046 23438 30098
rect 23490 30046 23492 30098
rect 23436 30034 23492 30046
rect 23772 30660 23828 30670
rect 23772 30098 23828 30604
rect 23772 30046 23774 30098
rect 23826 30046 23828 30098
rect 23772 30034 23828 30046
rect 23772 29428 23828 29438
rect 23324 29426 23828 29428
rect 23324 29374 23774 29426
rect 23826 29374 23828 29426
rect 23324 29372 23828 29374
rect 23772 29362 23828 29372
rect 23884 29204 23940 31500
rect 23996 30882 24052 31500
rect 23996 30830 23998 30882
rect 24050 30830 24052 30882
rect 23996 30436 24052 30830
rect 23996 30370 24052 30380
rect 24108 30548 24164 30558
rect 24108 30210 24164 30492
rect 24108 30158 24110 30210
rect 24162 30158 24164 30210
rect 24108 29538 24164 30158
rect 24108 29486 24110 29538
rect 24162 29486 24164 29538
rect 24108 29474 24164 29486
rect 24108 29316 24164 29326
rect 24220 29316 24276 31836
rect 24444 31220 24500 32508
rect 24556 32450 24612 32462
rect 24556 32398 24558 32450
rect 24610 32398 24612 32450
rect 24556 32228 24612 32398
rect 24556 32162 24612 32172
rect 24892 31892 24948 33070
rect 24892 31826 24948 31836
rect 24556 31778 24612 31790
rect 24556 31726 24558 31778
rect 24610 31726 24612 31778
rect 24556 31556 24612 31726
rect 24556 31490 24612 31500
rect 25004 31778 25060 31790
rect 25004 31726 25006 31778
rect 25058 31726 25060 31778
rect 24556 31220 24612 31230
rect 24444 31218 24612 31220
rect 24444 31166 24558 31218
rect 24610 31166 24612 31218
rect 24444 31164 24612 31166
rect 24556 31154 24612 31164
rect 24444 30994 24500 31006
rect 24444 30942 24446 30994
rect 24498 30942 24500 30994
rect 24444 30324 24500 30942
rect 24780 30994 24836 31006
rect 24780 30942 24782 30994
rect 24834 30942 24836 30994
rect 24780 30884 24836 30942
rect 25004 30996 25060 31726
rect 25004 30930 25060 30940
rect 24780 30818 24836 30828
rect 24444 30258 24500 30268
rect 24556 30212 24612 30222
rect 24556 30118 24612 30156
rect 24164 29260 24276 29316
rect 24108 29250 24164 29260
rect 23772 29148 23940 29204
rect 23436 28644 23492 28654
rect 23436 28550 23492 28588
rect 23660 28644 23716 28654
rect 23436 27860 23492 27870
rect 23324 27076 23380 27086
rect 23212 27074 23380 27076
rect 23212 27022 23326 27074
rect 23378 27022 23380 27074
rect 23212 27020 23380 27022
rect 22988 25060 23044 26852
rect 23212 25956 23268 27020
rect 23324 27010 23380 27020
rect 23436 26292 23492 27804
rect 23212 25890 23268 25900
rect 23324 26236 23492 26292
rect 23548 26964 23604 26974
rect 23212 25506 23268 25518
rect 23212 25454 23214 25506
rect 23266 25454 23268 25506
rect 23212 25284 23268 25454
rect 23212 25218 23268 25228
rect 22876 25004 23044 25060
rect 22876 23492 22932 25004
rect 23324 24948 23380 26236
rect 23548 26180 23604 26908
rect 23436 26124 23604 26180
rect 23436 26066 23492 26124
rect 23436 26014 23438 26066
rect 23490 26014 23492 26066
rect 23436 26002 23492 26014
rect 23324 24892 23492 24948
rect 22988 24836 23044 24846
rect 22988 24834 23268 24836
rect 22988 24782 22990 24834
rect 23042 24782 23268 24834
rect 22988 24780 23268 24782
rect 22988 24770 23044 24780
rect 23212 24050 23268 24780
rect 23212 23998 23214 24050
rect 23266 23998 23268 24050
rect 23212 23986 23268 23998
rect 23324 24722 23380 24734
rect 23324 24670 23326 24722
rect 23378 24670 23380 24722
rect 22876 23436 23156 23492
rect 22876 23268 22932 23278
rect 22876 23174 22932 23212
rect 22764 22430 22766 22482
rect 22818 22430 22820 22482
rect 22764 22418 22820 22430
rect 22876 22260 22932 22270
rect 22204 21868 22708 21924
rect 22764 22146 22820 22158
rect 22764 22094 22766 22146
rect 22818 22094 22820 22146
rect 22204 21810 22260 21868
rect 22204 21758 22206 21810
rect 22258 21758 22260 21810
rect 22204 21746 22260 21758
rect 22428 21364 22484 21374
rect 22428 20914 22484 21308
rect 22428 20862 22430 20914
rect 22482 20862 22484 20914
rect 22428 20850 22484 20862
rect 22764 20804 22820 22094
rect 22876 21810 22932 22204
rect 22876 21758 22878 21810
rect 22930 21758 22932 21810
rect 22876 21746 22932 21758
rect 22988 22146 23044 22158
rect 22988 22094 22990 22146
rect 23042 22094 23044 22146
rect 22988 21812 23044 22094
rect 22988 21746 23044 21756
rect 23100 21588 23156 23436
rect 23324 23378 23380 24670
rect 23436 23604 23492 24892
rect 23436 23538 23492 23548
rect 23324 23326 23326 23378
rect 23378 23326 23380 23378
rect 23324 23314 23380 23326
rect 23660 23156 23716 28588
rect 23772 26292 23828 29148
rect 23884 28980 23940 28990
rect 23884 27186 23940 28924
rect 23996 28532 24052 28542
rect 23996 28438 24052 28476
rect 24444 27858 24500 27870
rect 24444 27806 24446 27858
rect 24498 27806 24500 27858
rect 23996 27746 24052 27758
rect 23996 27694 23998 27746
rect 24050 27694 24052 27746
rect 23996 27300 24052 27694
rect 23996 27234 24052 27244
rect 23884 27134 23886 27186
rect 23938 27134 23940 27186
rect 23884 27122 23940 27134
rect 24444 27076 24500 27806
rect 24444 27010 24500 27020
rect 24556 26964 24612 27002
rect 24556 26898 24612 26908
rect 24220 26852 24276 26862
rect 23772 26226 23828 26236
rect 23996 26850 24276 26852
rect 23996 26798 24222 26850
rect 24274 26798 24276 26850
rect 23996 26796 24276 26798
rect 23772 26066 23828 26078
rect 23772 26014 23774 26066
rect 23826 26014 23828 26066
rect 23772 25732 23828 26014
rect 23772 25666 23828 25676
rect 23996 25618 24052 26796
rect 24220 26786 24276 26796
rect 24444 26404 24500 26414
rect 24444 26292 24500 26348
rect 23996 25566 23998 25618
rect 24050 25566 24052 25618
rect 23996 25554 24052 25566
rect 24220 26290 24500 26292
rect 24220 26238 24446 26290
rect 24498 26238 24500 26290
rect 24220 26236 24500 26238
rect 24220 23268 24276 26236
rect 24444 26226 24500 26236
rect 24556 26402 24612 26414
rect 24556 26350 24558 26402
rect 24610 26350 24612 26402
rect 24556 25620 24612 26350
rect 24556 25554 24612 25564
rect 24668 24724 24724 24734
rect 25116 24724 25172 41916
rect 25340 41860 25396 41870
rect 25340 41766 25396 41804
rect 25676 41746 25732 41758
rect 25676 41694 25678 41746
rect 25730 41694 25732 41746
rect 25676 41298 25732 41694
rect 26012 41748 26068 41916
rect 26348 41970 26404 41982
rect 26348 41918 26350 41970
rect 26402 41918 26404 41970
rect 26348 41748 26404 41918
rect 26012 41692 26292 41748
rect 25676 41246 25678 41298
rect 25730 41246 25732 41298
rect 25676 41076 25732 41246
rect 25676 41020 26068 41076
rect 25900 40180 25956 40190
rect 25564 40178 25956 40180
rect 25564 40126 25902 40178
rect 25954 40126 25956 40178
rect 25564 40124 25956 40126
rect 25228 39508 25284 39518
rect 25228 39058 25284 39452
rect 25228 39006 25230 39058
rect 25282 39006 25284 39058
rect 25228 38994 25284 39006
rect 25564 38946 25620 40124
rect 25900 40114 25956 40124
rect 26012 40180 26068 41020
rect 26236 40292 26292 41692
rect 26348 41682 26404 41692
rect 26460 40628 26516 42140
rect 26460 40514 26516 40572
rect 26460 40462 26462 40514
rect 26514 40462 26516 40514
rect 26460 40450 26516 40462
rect 26684 40292 26740 42476
rect 27692 42082 27748 42094
rect 27692 42030 27694 42082
rect 27746 42030 27748 42082
rect 27468 41972 27524 41982
rect 27468 41970 27636 41972
rect 27468 41918 27470 41970
rect 27522 41918 27636 41970
rect 27468 41916 27636 41918
rect 27468 41906 27524 41916
rect 27580 41076 27636 41916
rect 27692 41300 27748 42030
rect 28812 41858 28868 41870
rect 28812 41806 28814 41858
rect 28866 41806 28868 41858
rect 27804 41300 27860 41310
rect 27692 41298 27860 41300
rect 27692 41246 27806 41298
rect 27858 41246 27860 41298
rect 27692 41244 27860 41246
rect 27804 41234 27860 41244
rect 28588 41188 28644 41198
rect 28812 41188 28868 41806
rect 28588 41186 28868 41188
rect 28588 41134 28590 41186
rect 28642 41134 28868 41186
rect 28588 41132 28868 41134
rect 29372 41188 29428 41198
rect 29708 41188 29764 43486
rect 30268 42980 30324 44044
rect 30940 43652 30996 49200
rect 31500 45892 31556 45902
rect 31388 45890 31556 45892
rect 31388 45838 31502 45890
rect 31554 45838 31556 45890
rect 31388 45836 31556 45838
rect 31276 45668 31332 45678
rect 31052 45666 31332 45668
rect 31052 45614 31278 45666
rect 31330 45614 31332 45666
rect 31052 45612 31332 45614
rect 31052 44434 31108 45612
rect 31276 45602 31332 45612
rect 31276 45332 31332 45342
rect 31388 45332 31444 45836
rect 31500 45826 31556 45836
rect 31276 45330 31444 45332
rect 31276 45278 31278 45330
rect 31330 45278 31444 45330
rect 31276 45276 31444 45278
rect 31276 45266 31332 45276
rect 31612 45108 31668 49200
rect 32172 45890 32228 45902
rect 32172 45838 32174 45890
rect 32226 45838 32228 45890
rect 31948 45218 32004 45230
rect 31948 45166 31950 45218
rect 32002 45166 32004 45218
rect 31612 45052 31780 45108
rect 31052 44382 31054 44434
rect 31106 44382 31108 44434
rect 31052 44370 31108 44382
rect 31612 44882 31668 44894
rect 31612 44830 31614 44882
rect 31666 44830 31668 44882
rect 31612 44436 31668 44830
rect 31724 44548 31780 45052
rect 31724 44482 31780 44492
rect 31612 44370 31668 44380
rect 31948 43764 32004 45166
rect 32172 44772 32228 45838
rect 31948 43698 32004 43708
rect 32060 44716 32228 44772
rect 30940 43586 30996 43596
rect 30380 43428 30436 43438
rect 30380 43426 31332 43428
rect 30380 43374 30382 43426
rect 30434 43374 31332 43426
rect 30380 43372 31332 43374
rect 30380 43362 30436 43372
rect 30268 42924 30548 42980
rect 30268 42756 30324 42766
rect 29372 41186 29764 41188
rect 29372 41134 29374 41186
rect 29426 41134 29764 41186
rect 29372 41132 29764 41134
rect 29932 42642 29988 42654
rect 29932 42590 29934 42642
rect 29986 42590 29988 42642
rect 29932 41860 29988 42590
rect 30268 42642 30324 42700
rect 30268 42590 30270 42642
rect 30322 42590 30324 42642
rect 30268 42578 30324 42590
rect 30380 42082 30436 42094
rect 30380 42030 30382 42082
rect 30434 42030 30436 42082
rect 30044 41860 30100 41870
rect 29932 41858 30100 41860
rect 29932 41806 30046 41858
rect 30098 41806 30100 41858
rect 29932 41804 30100 41806
rect 27580 41020 28308 41076
rect 28252 40626 28308 41020
rect 28252 40574 28254 40626
rect 28306 40574 28308 40626
rect 28252 40562 28308 40574
rect 27020 40514 27076 40526
rect 27020 40462 27022 40514
rect 27074 40462 27076 40514
rect 26236 40290 26628 40292
rect 26236 40238 26238 40290
rect 26290 40238 26628 40290
rect 26236 40236 26628 40238
rect 26684 40236 26964 40292
rect 26236 40226 26292 40236
rect 26572 40180 26628 40236
rect 26572 40124 26852 40180
rect 26012 40114 26068 40124
rect 26796 39730 26852 40124
rect 26796 39678 26798 39730
rect 26850 39678 26852 39730
rect 26796 39666 26852 39678
rect 25564 38894 25566 38946
rect 25618 38894 25620 38946
rect 25564 38882 25620 38894
rect 26124 39620 26180 39630
rect 26124 39396 26180 39564
rect 26124 38834 26180 39340
rect 26796 39396 26852 39406
rect 26908 39396 26964 40236
rect 26852 39340 26964 39396
rect 26796 39330 26852 39340
rect 27020 39284 27076 40462
rect 28588 40404 28644 41132
rect 29260 40514 29316 40526
rect 29260 40462 29262 40514
rect 29314 40462 29316 40514
rect 28476 40348 28644 40404
rect 29148 40404 29204 40414
rect 27244 39396 27300 39406
rect 27244 39302 27300 39340
rect 28476 39396 28532 40348
rect 29148 40310 29204 40348
rect 28588 40180 28644 40190
rect 28588 40086 28644 40124
rect 29260 39620 29316 40462
rect 29260 39554 29316 39564
rect 28476 39330 28532 39340
rect 29260 39396 29316 39406
rect 29372 39396 29428 41132
rect 29316 39340 29428 39396
rect 29932 40404 29988 41804
rect 30044 41794 30100 41804
rect 30156 41300 30212 41310
rect 30380 41300 30436 42030
rect 30156 41298 30436 41300
rect 30156 41246 30158 41298
rect 30210 41246 30436 41298
rect 30156 41244 30436 41246
rect 30156 41234 30212 41244
rect 27020 39218 27076 39228
rect 29036 39284 29092 39294
rect 26124 38782 26126 38834
rect 26178 38782 26180 38834
rect 26124 38770 26180 38782
rect 26908 38724 26964 38734
rect 27692 38724 27748 38734
rect 26908 38722 27412 38724
rect 26908 38670 26910 38722
rect 26962 38670 27412 38722
rect 26908 38668 27412 38670
rect 26908 38658 26964 38668
rect 26012 38052 26068 38062
rect 25340 37380 25396 37390
rect 25340 35922 25396 37324
rect 25340 35870 25342 35922
rect 25394 35870 25396 35922
rect 25340 35858 25396 35870
rect 26012 35810 26068 37996
rect 27356 37938 27412 38668
rect 27692 38050 27748 38668
rect 29036 38722 29092 39228
rect 29036 38670 29038 38722
rect 29090 38670 29092 38722
rect 29036 38658 29092 38670
rect 27692 37998 27694 38050
rect 27746 37998 27748 38050
rect 27692 37986 27748 37998
rect 29260 38052 29316 39340
rect 29820 39284 29876 39294
rect 29820 38834 29876 39228
rect 29820 38782 29822 38834
rect 29874 38782 29876 38834
rect 29820 38770 29876 38782
rect 29484 38724 29540 38734
rect 29484 38630 29540 38668
rect 29372 38052 29428 38062
rect 29260 38050 29428 38052
rect 29260 37998 29374 38050
rect 29426 37998 29428 38050
rect 29260 37996 29428 37998
rect 27356 37886 27358 37938
rect 27410 37886 27412 37938
rect 27356 37874 27412 37886
rect 29148 37380 29204 37390
rect 28700 37378 29204 37380
rect 28700 37326 29150 37378
rect 29202 37326 29204 37378
rect 28700 37324 29204 37326
rect 26908 36594 26964 36606
rect 26908 36542 26910 36594
rect 26962 36542 26964 36594
rect 26908 36484 26964 36542
rect 28028 36596 28084 36606
rect 28028 36502 28084 36540
rect 27468 36484 27524 36494
rect 26908 36482 27524 36484
rect 26908 36430 27470 36482
rect 27522 36430 27524 36482
rect 26908 36428 27524 36430
rect 26012 35758 26014 35810
rect 26066 35758 26068 35810
rect 26012 35746 26068 35758
rect 26124 36260 26180 36270
rect 25900 35588 25956 35598
rect 25900 35138 25956 35532
rect 25900 35086 25902 35138
rect 25954 35086 25956 35138
rect 25900 35074 25956 35086
rect 26124 35252 26180 36204
rect 26908 36036 26964 36428
rect 27468 36418 27524 36428
rect 27244 36260 27300 36270
rect 27244 36166 27300 36204
rect 26236 35980 26964 36036
rect 26236 35698 26292 35980
rect 26348 35812 26404 35822
rect 26348 35810 26516 35812
rect 26348 35758 26350 35810
rect 26402 35758 26516 35810
rect 26348 35756 26516 35758
rect 26348 35746 26404 35756
rect 26236 35646 26238 35698
rect 26290 35646 26292 35698
rect 26236 35634 26292 35646
rect 26124 34914 26180 35196
rect 26124 34862 26126 34914
rect 26178 34862 26180 34914
rect 26124 34850 26180 34862
rect 26460 34804 26516 35756
rect 28700 35810 28756 37324
rect 29148 37314 29204 37324
rect 29372 36596 29428 37996
rect 29932 37940 29988 40348
rect 30380 39620 30436 39630
rect 30044 38948 30100 38958
rect 30044 38162 30100 38892
rect 30380 38946 30436 39564
rect 30380 38894 30382 38946
rect 30434 38894 30436 38946
rect 30380 38724 30436 38894
rect 30492 39060 30548 42924
rect 31164 42754 31220 42766
rect 31164 42702 31166 42754
rect 31218 42702 31220 42754
rect 30716 41972 30772 41982
rect 30716 41970 30996 41972
rect 30716 41918 30718 41970
rect 30770 41918 30996 41970
rect 30716 41916 30996 41918
rect 30716 41906 30772 41916
rect 30940 40626 30996 41916
rect 30940 40574 30942 40626
rect 30994 40574 30996 40626
rect 30940 40562 30996 40574
rect 31164 39172 31220 42702
rect 31276 42194 31332 43372
rect 31836 42756 31892 42766
rect 31276 42142 31278 42194
rect 31330 42142 31332 42194
rect 31276 42130 31332 42142
rect 31612 42532 31668 42542
rect 31612 42082 31668 42476
rect 31612 42030 31614 42082
rect 31666 42030 31668 42082
rect 31612 42018 31668 42030
rect 31836 41972 31892 42700
rect 31836 41916 32004 41972
rect 31276 41300 31332 41310
rect 31276 40290 31332 41244
rect 31276 40238 31278 40290
rect 31330 40238 31332 40290
rect 31276 40226 31332 40238
rect 31500 40514 31556 40526
rect 31500 40462 31502 40514
rect 31554 40462 31556 40514
rect 30492 38834 30548 39004
rect 30492 38782 30494 38834
rect 30546 38782 30548 38834
rect 30492 38770 30548 38782
rect 30940 39116 31220 39172
rect 30380 38658 30436 38668
rect 30044 38110 30046 38162
rect 30098 38110 30100 38162
rect 30044 38098 30100 38110
rect 29932 37884 30100 37940
rect 29484 37266 29540 37278
rect 29484 37214 29486 37266
rect 29538 37214 29540 37266
rect 29484 36820 29540 37214
rect 29484 36754 29540 36764
rect 29484 36596 29540 36606
rect 29372 36540 29484 36596
rect 29484 36530 29540 36540
rect 29820 36596 29876 36606
rect 29820 36502 29876 36540
rect 29260 36484 29316 36494
rect 29316 36428 29428 36484
rect 29260 36390 29316 36428
rect 28700 35758 28702 35810
rect 28754 35758 28756 35810
rect 28700 35746 28756 35758
rect 25340 34690 25396 34702
rect 25340 34638 25342 34690
rect 25394 34638 25396 34690
rect 25340 34356 25396 34638
rect 25340 34290 25396 34300
rect 25228 34130 25284 34142
rect 25228 34078 25230 34130
rect 25282 34078 25284 34130
rect 25228 30996 25284 34078
rect 25788 34132 25844 34142
rect 25844 34076 25956 34132
rect 25788 34066 25844 34076
rect 25452 33236 25508 33246
rect 25900 33236 25956 34076
rect 26012 34020 26068 34030
rect 26012 33926 26068 33964
rect 26348 33348 26404 33358
rect 26460 33348 26516 34748
rect 26348 33346 26516 33348
rect 26348 33294 26350 33346
rect 26402 33294 26516 33346
rect 26348 33292 26516 33294
rect 26684 35698 26740 35710
rect 26684 35646 26686 35698
rect 26738 35646 26740 35698
rect 26684 34802 26740 35646
rect 27356 35698 27412 35710
rect 27356 35646 27358 35698
rect 27410 35646 27412 35698
rect 26684 34750 26686 34802
rect 26738 34750 26740 34802
rect 26348 33282 26404 33292
rect 26012 33236 26068 33246
rect 25900 33234 26068 33236
rect 25900 33182 26014 33234
rect 26066 33182 26068 33234
rect 25900 33180 26068 33182
rect 25340 33124 25396 33134
rect 25340 33030 25396 33068
rect 25340 30996 25396 31006
rect 25228 30940 25340 30996
rect 25340 30324 25396 30940
rect 25340 27076 25396 30268
rect 25452 29876 25508 33180
rect 26012 33170 26068 33180
rect 26236 32674 26292 32686
rect 26236 32622 26238 32674
rect 26290 32622 26292 32674
rect 26236 32452 26292 32622
rect 26236 32386 26292 32396
rect 26572 32564 26628 32574
rect 26684 32564 26740 34750
rect 26572 32562 26740 32564
rect 26572 32510 26574 32562
rect 26626 32510 26740 32562
rect 26572 32508 26740 32510
rect 26908 34916 26964 34926
rect 27356 34916 27412 35646
rect 28028 35698 28084 35710
rect 28028 35646 28030 35698
rect 28082 35646 28084 35698
rect 28028 35028 28084 35646
rect 28028 34962 28084 34972
rect 29148 35028 29204 35038
rect 26908 34914 27412 34916
rect 26908 34862 26910 34914
rect 26962 34862 27412 34914
rect 26908 34860 27412 34862
rect 29148 34916 29204 34972
rect 29148 34914 29316 34916
rect 29148 34862 29150 34914
rect 29202 34862 29316 34914
rect 29148 34860 29316 34862
rect 26572 31892 26628 32508
rect 26572 31826 26628 31836
rect 25788 31780 25844 31790
rect 25788 31686 25844 31724
rect 26012 30884 26068 30894
rect 26012 30790 26068 30828
rect 26908 30548 26964 34860
rect 29148 34850 29204 34860
rect 28140 34804 28196 34814
rect 28140 34018 28196 34748
rect 28812 34244 28868 34254
rect 28812 34150 28868 34188
rect 28140 33966 28142 34018
rect 28194 33966 28196 34018
rect 28140 33954 28196 33966
rect 28588 34130 28644 34142
rect 28588 34078 28590 34130
rect 28642 34078 28644 34130
rect 28364 33908 28420 33918
rect 27916 31892 27972 31902
rect 27916 31798 27972 31836
rect 26908 30482 26964 30492
rect 28140 30882 28196 30894
rect 28140 30830 28142 30882
rect 28194 30830 28196 30882
rect 28140 30548 28196 30830
rect 28140 30482 28196 30492
rect 26796 30100 26852 30110
rect 26684 30098 26852 30100
rect 26684 30046 26798 30098
rect 26850 30046 26852 30098
rect 26684 30044 26852 30046
rect 25452 29810 25508 29820
rect 26236 29988 26292 29998
rect 25900 29540 25956 29550
rect 25900 28866 25956 29484
rect 25900 28814 25902 28866
rect 25954 28814 25956 28866
rect 25900 28802 25956 28814
rect 25788 28642 25844 28654
rect 25788 28590 25790 28642
rect 25842 28590 25844 28642
rect 25788 28532 25844 28590
rect 26236 28644 26292 29932
rect 26572 29652 26628 29662
rect 26236 28550 26292 28588
rect 26460 29650 26628 29652
rect 26460 29598 26574 29650
rect 26626 29598 26628 29650
rect 26460 29596 26628 29598
rect 25788 27972 25844 28476
rect 25788 27906 25844 27916
rect 26460 28530 26516 29596
rect 26572 29586 26628 29596
rect 26572 29426 26628 29438
rect 26572 29374 26574 29426
rect 26626 29374 26628 29426
rect 26572 28644 26628 29374
rect 26572 28578 26628 28588
rect 26460 28478 26462 28530
rect 26514 28478 26516 28530
rect 26460 27636 26516 28478
rect 26684 28308 26740 30044
rect 26796 30034 26852 30044
rect 26908 29988 26964 29998
rect 26908 29894 26964 29932
rect 27132 29988 27188 29998
rect 27132 29894 27188 29932
rect 26796 29650 26852 29662
rect 26796 29598 26798 29650
rect 26850 29598 26852 29650
rect 26796 29538 26852 29598
rect 27020 29540 27076 29550
rect 26796 29486 26798 29538
rect 26850 29486 26852 29538
rect 26796 29474 26852 29486
rect 26908 29484 27020 29540
rect 26908 28756 26964 29484
rect 27020 29446 27076 29484
rect 27692 29540 27748 29550
rect 27692 29446 27748 29484
rect 26572 28252 26740 28308
rect 26796 28700 26964 28756
rect 26572 28082 26628 28252
rect 26572 28030 26574 28082
rect 26626 28030 26628 28082
rect 26572 28018 26628 28030
rect 26684 28084 26740 28094
rect 26796 28084 26852 28700
rect 26908 28532 26964 28542
rect 26908 28438 26964 28476
rect 27468 28532 27524 28542
rect 27468 28438 27524 28476
rect 26684 28082 26852 28084
rect 26684 28030 26686 28082
rect 26738 28030 26852 28082
rect 26684 28028 26852 28030
rect 26684 28018 26740 28028
rect 27132 27970 27188 27982
rect 27132 27918 27134 27970
rect 27186 27918 27188 27970
rect 26348 27634 26516 27636
rect 26348 27582 26462 27634
rect 26514 27582 26516 27634
rect 26348 27580 26516 27582
rect 25676 27076 25732 27086
rect 25340 27074 25732 27076
rect 25340 27022 25678 27074
rect 25730 27022 25732 27074
rect 25340 27020 25732 27022
rect 25676 27010 25732 27020
rect 26124 25620 26180 25630
rect 25228 24724 25284 24734
rect 24668 24722 25284 24724
rect 24668 24670 24670 24722
rect 24722 24670 25230 24722
rect 25282 24670 25284 24722
rect 24668 24668 25284 24670
rect 24668 24658 24724 24668
rect 25228 24658 25284 24668
rect 25340 24050 25396 24062
rect 25676 24052 25732 24062
rect 25340 23998 25342 24050
rect 25394 23998 25396 24050
rect 24332 23604 24388 23614
rect 24388 23548 24500 23604
rect 24332 23538 24388 23548
rect 23660 23100 23828 23156
rect 23660 22932 23716 22942
rect 23660 22838 23716 22876
rect 23436 22708 23492 22718
rect 23324 22146 23380 22158
rect 23324 22094 23326 22146
rect 23378 22094 23380 22146
rect 23100 21494 23156 21532
rect 23212 21812 23268 21822
rect 22764 20738 22820 20748
rect 22988 21474 23044 21486
rect 22988 21422 22990 21474
rect 23042 21422 23044 21474
rect 22988 20916 23044 21422
rect 23212 21364 23268 21756
rect 22988 20802 23044 20860
rect 22988 20750 22990 20802
rect 23042 20750 23044 20802
rect 22988 20738 23044 20750
rect 23100 21308 23268 21364
rect 23100 20802 23156 21308
rect 23100 20750 23102 20802
rect 23154 20750 23156 20802
rect 23100 20738 23156 20750
rect 23212 20804 23268 20814
rect 23324 20804 23380 22094
rect 23436 21586 23492 22652
rect 23436 21534 23438 21586
rect 23490 21534 23492 21586
rect 23436 21522 23492 21534
rect 23660 22258 23716 22270
rect 23660 22206 23662 22258
rect 23714 22206 23716 22258
rect 23660 21364 23716 22206
rect 23660 21298 23716 21308
rect 23660 21028 23716 21038
rect 23772 21028 23828 23100
rect 24220 23154 24276 23212
rect 24220 23102 24222 23154
rect 24274 23102 24276 23154
rect 24220 23090 24276 23102
rect 24332 23266 24388 23278
rect 24332 23214 24334 23266
rect 24386 23214 24388 23266
rect 24332 23156 24388 23214
rect 24332 23090 24388 23100
rect 24220 22146 24276 22158
rect 24220 22094 24222 22146
rect 24274 22094 24276 22146
rect 24220 21364 24276 22094
rect 24220 21298 24276 21308
rect 23660 21026 23828 21028
rect 23660 20974 23662 21026
rect 23714 20974 23828 21026
rect 23660 20972 23828 20974
rect 23660 20962 23716 20972
rect 23996 20916 24052 20926
rect 23996 20822 24052 20860
rect 23268 20748 23380 20804
rect 23212 20710 23268 20748
rect 24108 20690 24164 20702
rect 24108 20638 24110 20690
rect 24162 20638 24164 20690
rect 23100 20244 23156 20254
rect 22652 19234 22708 19246
rect 22652 19182 22654 19234
rect 22706 19182 22708 19234
rect 22652 18564 22708 19182
rect 22652 18498 22708 18508
rect 22092 17602 22148 17612
rect 21980 17490 22036 17500
rect 22092 17442 22148 17454
rect 22092 17390 22094 17442
rect 22146 17390 22148 17442
rect 22092 17108 22148 17390
rect 22092 17042 22148 17052
rect 22540 17442 22596 17454
rect 22540 17390 22542 17442
rect 22594 17390 22596 17442
rect 22540 17332 22596 17390
rect 22316 16884 22372 16894
rect 22316 16790 22372 16828
rect 22540 16882 22596 17276
rect 22540 16830 22542 16882
rect 22594 16830 22596 16882
rect 22540 16818 22596 16830
rect 21756 16212 21812 16222
rect 21756 16118 21812 16156
rect 21868 15988 21924 16716
rect 21644 15922 21700 15932
rect 21756 15932 21924 15988
rect 22204 16772 22260 16782
rect 22204 16100 22260 16716
rect 22876 16660 22932 16670
rect 22876 16566 22932 16604
rect 22204 15986 22260 16044
rect 22428 16436 22484 16446
rect 22428 16098 22484 16380
rect 22428 16046 22430 16098
rect 22482 16046 22484 16098
rect 22428 16034 22484 16046
rect 22204 15934 22206 15986
rect 22258 15934 22260 15986
rect 21308 15876 21364 15886
rect 20188 11564 20356 11620
rect 19836 11004 20100 11014
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 19836 10938 20100 10948
rect 19740 9940 19796 9950
rect 19628 9938 19796 9940
rect 19628 9886 19742 9938
rect 19794 9886 19796 9938
rect 19628 9884 19796 9886
rect 19740 9874 19796 9884
rect 20188 9940 20244 11564
rect 20524 11508 20580 15092
rect 20636 14644 20692 14654
rect 20636 14530 20692 14588
rect 20636 14478 20638 14530
rect 20690 14478 20692 14530
rect 20636 13972 20692 14478
rect 20636 13906 20692 13916
rect 20636 13524 20692 13534
rect 20636 12738 20692 13468
rect 20636 12686 20638 12738
rect 20690 12686 20692 12738
rect 20636 12628 20692 12686
rect 20636 12562 20692 12572
rect 21084 12964 21140 15484
rect 21196 15874 21364 15876
rect 21196 15822 21310 15874
rect 21362 15822 21364 15874
rect 21196 15820 21364 15822
rect 21196 14644 21252 15820
rect 21308 15810 21364 15820
rect 21196 14578 21252 14588
rect 21308 15314 21364 15326
rect 21308 15262 21310 15314
rect 21362 15262 21364 15314
rect 21308 14532 21364 15262
rect 21756 14754 21812 15932
rect 22204 15922 22260 15934
rect 22876 15876 22932 15886
rect 22764 15874 22932 15876
rect 22764 15822 22878 15874
rect 22930 15822 22932 15874
rect 22764 15820 22932 15822
rect 22764 15652 22820 15820
rect 22876 15810 22932 15820
rect 23100 15652 23156 20188
rect 24108 20244 24164 20638
rect 24108 20178 24164 20188
rect 23436 19122 23492 19134
rect 23436 19070 23438 19122
rect 23490 19070 23492 19122
rect 23436 18452 23492 19070
rect 23436 18386 23492 18396
rect 23996 18676 24052 18686
rect 23884 18340 23940 18350
rect 23772 17108 23828 17118
rect 23772 17014 23828 17052
rect 23324 16996 23380 17006
rect 23212 16940 23324 16996
rect 23212 16882 23268 16940
rect 23212 16830 23214 16882
rect 23266 16830 23268 16882
rect 23212 16818 23268 16830
rect 23212 15988 23268 15998
rect 23212 15894 23268 15932
rect 22764 15586 22820 15596
rect 22876 15596 23156 15652
rect 21868 15540 21924 15550
rect 21868 15202 21924 15484
rect 21868 15150 21870 15202
rect 21922 15150 21924 15202
rect 21868 15138 21924 15150
rect 21756 14702 21758 14754
rect 21810 14702 21812 14754
rect 21756 14690 21812 14702
rect 21980 14642 22036 14654
rect 21980 14590 21982 14642
rect 22034 14590 22036 14642
rect 21308 14466 21364 14476
rect 21868 14530 21924 14542
rect 21868 14478 21870 14530
rect 21922 14478 21924 14530
rect 21420 13634 21476 13646
rect 21420 13582 21422 13634
rect 21474 13582 21476 13634
rect 21308 12964 21364 12974
rect 21084 12962 21364 12964
rect 21084 12910 21310 12962
rect 21362 12910 21364 12962
rect 21084 12908 21364 12910
rect 20188 9874 20244 9884
rect 20300 11452 20580 11508
rect 20748 11506 20804 11518
rect 20748 11454 20750 11506
rect 20802 11454 20804 11506
rect 19628 9604 19684 9614
rect 18844 9268 18900 9278
rect 18844 9174 18900 9212
rect 19628 9042 19684 9548
rect 20188 9604 20244 9614
rect 20188 9510 20244 9548
rect 19836 9436 20100 9446
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 19836 9370 20100 9380
rect 19628 8990 19630 9042
rect 19682 8990 19684 9042
rect 19628 8978 19684 8990
rect 20188 9044 20244 9054
rect 20188 8950 20244 8988
rect 19628 8372 20020 8428
rect 19404 8260 19460 8270
rect 19628 8260 19684 8372
rect 19964 8370 20020 8372
rect 19964 8318 19966 8370
rect 20018 8318 20020 8370
rect 19404 8258 19684 8260
rect 19404 8206 19406 8258
rect 19458 8206 19684 8258
rect 19404 8204 19684 8206
rect 19740 8258 19796 8270
rect 19740 8206 19742 8258
rect 19794 8206 19796 8258
rect 19404 8194 19460 8204
rect 18732 8082 18788 8092
rect 19292 8146 19348 8158
rect 19292 8094 19294 8146
rect 19346 8094 19348 8146
rect 16828 7746 16884 7756
rect 17052 8034 17108 8046
rect 17052 7982 17054 8034
rect 17106 7982 17108 8034
rect 17052 7700 17108 7982
rect 17052 7634 17108 7644
rect 17500 8034 17556 8046
rect 17500 7982 17502 8034
rect 17554 7982 17556 8034
rect 17500 7812 17556 7982
rect 17500 7362 17556 7756
rect 18396 8034 18452 8046
rect 18396 7982 18398 8034
rect 18450 7982 18452 8034
rect 18396 7700 18452 7982
rect 18844 8036 18900 8046
rect 19292 8036 19348 8094
rect 19740 8036 19796 8206
rect 18844 7942 18900 7980
rect 19180 7980 19796 8036
rect 19964 8036 20020 8318
rect 20300 8370 20356 11452
rect 20748 11396 20804 11454
rect 20748 11330 20804 11340
rect 20524 10612 20580 10622
rect 21084 10612 21140 12908
rect 21308 12898 21364 12908
rect 20524 10610 21140 10612
rect 20524 10558 20526 10610
rect 20578 10558 21140 10610
rect 20524 10556 21140 10558
rect 21420 11170 21476 13582
rect 21868 13076 21924 14478
rect 21980 13636 22036 14590
rect 21980 13570 22036 13580
rect 22204 14530 22260 14542
rect 22204 14478 22206 14530
rect 22258 14478 22260 14530
rect 22204 13524 22260 14478
rect 22540 14532 22596 14542
rect 22540 13746 22596 14476
rect 22540 13694 22542 13746
rect 22594 13694 22596 13746
rect 22540 13682 22596 13694
rect 22764 13524 22820 13534
rect 22204 13522 22820 13524
rect 22204 13470 22766 13522
rect 22818 13470 22820 13522
rect 22204 13468 22820 13470
rect 21868 12292 21924 13020
rect 22092 12852 22148 12862
rect 22092 12850 22708 12852
rect 22092 12798 22094 12850
rect 22146 12798 22708 12850
rect 22092 12796 22708 12798
rect 22092 12786 22148 12796
rect 21980 12292 22036 12302
rect 21868 12236 21980 12292
rect 21980 12226 22036 12236
rect 22652 12066 22708 12796
rect 22764 12628 22820 13468
rect 22764 12562 22820 12572
rect 22764 12404 22820 12414
rect 22764 12310 22820 12348
rect 22652 12014 22654 12066
rect 22706 12014 22708 12066
rect 22652 12002 22708 12014
rect 21420 11118 21422 11170
rect 21474 11118 21476 11170
rect 20524 10546 20580 10556
rect 21196 10498 21252 10510
rect 21196 10446 21198 10498
rect 21250 10446 21252 10498
rect 21196 9716 21252 10446
rect 21196 9650 21252 9660
rect 21420 9604 21476 11118
rect 22428 10500 22484 10510
rect 22428 9826 22484 10444
rect 22876 10276 22932 15596
rect 23324 15540 23380 16940
rect 23884 16884 23940 18284
rect 23884 16818 23940 16828
rect 23660 16660 23716 16670
rect 23660 16100 23716 16604
rect 23660 16006 23716 16044
rect 23884 16100 23940 16110
rect 23996 16100 24052 18620
rect 24220 18452 24276 18462
rect 24220 18358 24276 18396
rect 24332 18340 24388 18350
rect 24332 18246 24388 18284
rect 24444 18116 24500 23548
rect 25228 23492 25284 23502
rect 25228 22370 25284 23436
rect 25340 23156 25396 23998
rect 25564 24050 25732 24052
rect 25564 23998 25678 24050
rect 25730 23998 25732 24050
rect 25564 23996 25732 23998
rect 25340 23090 25396 23100
rect 25452 23492 25508 23502
rect 25452 23266 25508 23436
rect 25452 23214 25454 23266
rect 25506 23214 25508 23266
rect 25228 22318 25230 22370
rect 25282 22318 25284 22370
rect 25228 22306 25284 22318
rect 25452 20804 25508 23214
rect 25564 23268 25620 23996
rect 25676 23986 25732 23996
rect 25676 23380 25732 23390
rect 25676 23378 25956 23380
rect 25676 23326 25678 23378
rect 25730 23326 25956 23378
rect 25676 23324 25956 23326
rect 25676 23314 25732 23324
rect 25564 23202 25620 23212
rect 25676 23156 25732 23166
rect 25676 23062 25732 23100
rect 25900 21812 25956 23324
rect 26012 23154 26068 23166
rect 26012 23102 26014 23154
rect 26066 23102 26068 23154
rect 26012 22596 26068 23102
rect 26012 22530 26068 22540
rect 26124 22484 26180 25564
rect 26348 22708 26404 27580
rect 26460 27570 26516 27580
rect 26684 27860 26740 27870
rect 26460 27188 26516 27198
rect 26460 27094 26516 27132
rect 26684 26514 26740 27804
rect 27132 27188 27188 27918
rect 27356 27860 27412 27870
rect 27356 27766 27412 27804
rect 27132 27122 27188 27132
rect 26684 26462 26686 26514
rect 26738 26462 26740 26514
rect 26684 26450 26740 26462
rect 27804 26404 27860 26414
rect 27804 26310 27860 26348
rect 27468 26292 27524 26302
rect 27020 26068 27076 26078
rect 27020 25974 27076 26012
rect 26460 25394 26516 25406
rect 26460 25342 26462 25394
rect 26514 25342 26516 25394
rect 26460 23378 26516 25342
rect 26796 25282 26852 25294
rect 26796 25230 26798 25282
rect 26850 25230 26852 25282
rect 26796 24052 26852 25230
rect 26796 23986 26852 23996
rect 26460 23326 26462 23378
rect 26514 23326 26516 23378
rect 26460 23314 26516 23326
rect 26572 23380 26628 23390
rect 26628 23324 26852 23380
rect 26572 23314 26628 23324
rect 26796 23154 26852 23324
rect 26796 23102 26798 23154
rect 26850 23102 26852 23154
rect 26796 23090 26852 23102
rect 27468 23154 27524 26236
rect 27804 24052 27860 24062
rect 27804 23958 27860 23996
rect 27580 23268 27636 23278
rect 27580 23174 27636 23212
rect 27468 23102 27470 23154
rect 27522 23102 27524 23154
rect 27468 23090 27524 23102
rect 28364 22820 28420 33852
rect 28588 33348 28644 34078
rect 28588 33282 28644 33292
rect 29260 34020 29316 34860
rect 29260 33346 29316 33964
rect 29260 33294 29262 33346
rect 29314 33294 29316 33346
rect 28588 33124 28644 33134
rect 28644 33068 28756 33124
rect 28588 33030 28644 33068
rect 28588 31780 28644 31790
rect 28588 30212 28644 31724
rect 28476 29428 28532 29438
rect 28588 29428 28644 30156
rect 28476 29426 28588 29428
rect 28476 29374 28478 29426
rect 28530 29374 28588 29426
rect 28476 29372 28588 29374
rect 28476 29362 28532 29372
rect 28588 29334 28644 29372
rect 28588 27186 28644 27198
rect 28588 27134 28590 27186
rect 28642 27134 28644 27186
rect 28588 26404 28644 27134
rect 28588 26338 28644 26348
rect 28700 24834 28756 33068
rect 29260 31948 29316 33294
rect 29372 34130 29428 36428
rect 29932 34804 29988 34814
rect 29932 34710 29988 34748
rect 29372 34078 29374 34130
rect 29426 34078 29428 34130
rect 29372 33124 29428 34078
rect 29932 34244 29988 34254
rect 29932 33458 29988 34188
rect 29932 33406 29934 33458
rect 29986 33406 29988 33458
rect 29932 33394 29988 33406
rect 29372 33058 29428 33068
rect 29820 32674 29876 32686
rect 29820 32622 29822 32674
rect 29874 32622 29876 32674
rect 29148 31892 29316 31948
rect 29596 32562 29652 32574
rect 29596 32510 29598 32562
rect 29650 32510 29652 32562
rect 29148 31780 29204 31892
rect 29148 31686 29204 31724
rect 29596 31220 29652 32510
rect 29820 31948 29876 32622
rect 29820 31892 29988 31948
rect 29932 31890 29988 31892
rect 29932 31838 29934 31890
rect 29986 31838 29988 31890
rect 29932 31826 29988 31838
rect 29596 31154 29652 31164
rect 29372 31108 29428 31118
rect 29148 31106 29428 31108
rect 29148 31054 29374 31106
rect 29426 31054 29428 31106
rect 29148 31052 29428 31054
rect 29148 29538 29204 31052
rect 29372 31042 29428 31052
rect 29708 30994 29764 31006
rect 29708 30942 29710 30994
rect 29762 30942 29764 30994
rect 29148 29486 29150 29538
rect 29202 29486 29204 29538
rect 29148 29474 29204 29486
rect 29260 29988 29316 29998
rect 29260 28642 29316 29932
rect 29596 29988 29652 29998
rect 29596 29894 29652 29932
rect 29260 28590 29262 28642
rect 29314 28590 29316 28642
rect 29260 28578 29316 28590
rect 29484 29428 29540 29438
rect 29484 27858 29540 29372
rect 29596 29092 29652 29102
rect 29596 28754 29652 29036
rect 29708 28868 29764 30942
rect 30044 29092 30100 37884
rect 30828 35700 30884 35710
rect 30828 35586 30884 35644
rect 30828 35534 30830 35586
rect 30882 35534 30884 35586
rect 30828 35522 30884 35534
rect 30268 34020 30324 34030
rect 30268 33926 30324 33964
rect 30940 31948 30996 39116
rect 31052 38948 31108 38958
rect 31052 38854 31108 38892
rect 31276 38836 31332 38846
rect 31164 38834 31332 38836
rect 31164 38782 31278 38834
rect 31330 38782 31332 38834
rect 31164 38780 31332 38782
rect 31052 37492 31108 37502
rect 31164 37492 31220 38780
rect 31276 38770 31332 38780
rect 31052 37490 31220 37492
rect 31052 37438 31054 37490
rect 31106 37438 31220 37490
rect 31052 37436 31220 37438
rect 31388 38612 31444 38622
rect 31052 37426 31108 37436
rect 31388 37266 31444 38556
rect 31500 37380 31556 40462
rect 31948 40514 32004 41916
rect 31948 40462 31950 40514
rect 32002 40462 32004 40514
rect 31948 40450 32004 40462
rect 31612 39732 31668 39742
rect 31948 39732 32004 39742
rect 31612 39730 31948 39732
rect 31612 39678 31614 39730
rect 31666 39678 31948 39730
rect 31612 39676 31948 39678
rect 31612 39666 31668 39676
rect 31948 39618 32004 39676
rect 31948 39566 31950 39618
rect 32002 39566 32004 39618
rect 31948 39554 32004 39566
rect 31836 39060 31892 39070
rect 31836 38966 31892 39004
rect 31612 37380 31668 37390
rect 31500 37378 31780 37380
rect 31500 37326 31614 37378
rect 31666 37326 31780 37378
rect 31500 37324 31780 37326
rect 31612 37314 31668 37324
rect 31388 37214 31390 37266
rect 31442 37214 31444 37266
rect 31388 37202 31444 37214
rect 31276 36820 31332 36830
rect 31276 35922 31332 36764
rect 31612 36484 31668 36494
rect 31612 36390 31668 36428
rect 31276 35870 31278 35922
rect 31330 35870 31332 35922
rect 31276 35858 31332 35870
rect 31388 36260 31444 36270
rect 31388 35140 31444 36204
rect 31724 35812 31780 37324
rect 31948 35812 32004 35822
rect 31724 35810 32004 35812
rect 31724 35758 31950 35810
rect 32002 35758 32004 35810
rect 31724 35756 32004 35758
rect 31612 35700 31668 35710
rect 31612 35606 31668 35644
rect 31276 35084 31444 35140
rect 31164 33348 31220 33358
rect 31164 32786 31220 33292
rect 31164 32734 31166 32786
rect 31218 32734 31220 32786
rect 31164 32722 31220 32734
rect 30940 31892 31108 31948
rect 30716 31220 30772 31230
rect 30716 31126 30772 31164
rect 31052 30994 31108 31836
rect 31052 30942 31054 30994
rect 31106 30942 31108 30994
rect 31052 30930 31108 30942
rect 30044 29026 30100 29036
rect 30156 30098 30212 30110
rect 30156 30046 30158 30098
rect 30210 30046 30212 30098
rect 29708 28802 29764 28812
rect 29596 28702 29598 28754
rect 29650 28702 29652 28754
rect 29596 28690 29652 28702
rect 30156 28756 30212 30046
rect 31276 29540 31332 35084
rect 31388 34916 31444 34926
rect 31388 31948 31444 34860
rect 31948 34132 32004 35756
rect 32060 35700 32116 44716
rect 32172 43652 32228 43662
rect 32172 42978 32228 43596
rect 32284 43428 32340 49200
rect 32956 47012 33012 49200
rect 32956 46946 33012 46956
rect 33180 46116 33236 46126
rect 33180 46022 33236 46060
rect 32396 45218 32452 45230
rect 32396 45166 32398 45218
rect 32450 45166 32452 45218
rect 32396 43708 32452 45166
rect 33292 44994 33348 45006
rect 33292 44942 33294 44994
rect 33346 44942 33348 44994
rect 33068 44436 33124 44446
rect 33180 44436 33236 44446
rect 33124 44434 33236 44436
rect 33124 44382 33182 44434
rect 33234 44382 33236 44434
rect 33124 44380 33236 44382
rect 33068 44370 33124 44380
rect 33180 44212 33236 44380
rect 33180 44146 33236 44156
rect 33292 44436 33348 44942
rect 33628 44660 33684 49200
rect 34972 46116 35028 49200
rect 36316 46564 36372 49200
rect 36988 47012 37044 47022
rect 36316 46508 36484 46564
rect 35196 46284 35460 46294
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35196 46218 35460 46228
rect 34972 46060 35252 46116
rect 35084 45668 35140 45678
rect 34636 45666 35140 45668
rect 34636 45614 35086 45666
rect 35138 45614 35140 45666
rect 34636 45612 35140 45614
rect 34636 45218 34692 45612
rect 35084 45602 35140 45612
rect 35196 45332 35252 46060
rect 35980 45892 36036 45902
rect 35868 45890 36036 45892
rect 35868 45838 35982 45890
rect 36034 45838 36036 45890
rect 35868 45836 36036 45838
rect 35196 45266 35252 45276
rect 35420 45778 35476 45790
rect 35420 45726 35422 45778
rect 35474 45726 35476 45778
rect 34636 45166 34638 45218
rect 34690 45166 34692 45218
rect 34636 45154 34692 45166
rect 33964 45108 34020 45118
rect 33964 45014 34020 45052
rect 35420 44884 35476 45726
rect 35420 44818 35476 44828
rect 35196 44716 35460 44726
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 33628 44604 34020 44660
rect 35196 44650 35460 44660
rect 33292 43708 33348 44380
rect 32396 43652 32564 43708
rect 32284 43362 32340 43372
rect 32508 43426 32564 43652
rect 32508 43374 32510 43426
rect 32562 43374 32564 43426
rect 32172 42926 32174 42978
rect 32226 42926 32228 42978
rect 32172 42914 32228 42926
rect 32508 42980 32564 43374
rect 32508 42914 32564 42924
rect 33180 43652 33348 43708
rect 33740 44322 33796 44334
rect 33740 44270 33742 44322
rect 33794 44270 33796 44322
rect 32284 41972 32340 41982
rect 32284 41300 32340 41916
rect 32508 41972 32564 41982
rect 33180 41972 33236 43652
rect 32508 41970 33236 41972
rect 32508 41918 32510 41970
rect 32562 41918 33182 41970
rect 33234 41918 33236 41970
rect 32508 41916 33236 41918
rect 32508 41906 32564 41916
rect 32284 41206 32340 41244
rect 32732 41298 32788 41916
rect 33180 41906 33236 41916
rect 33292 43538 33348 43550
rect 33292 43486 33294 43538
rect 33346 43486 33348 43538
rect 32732 41246 32734 41298
rect 32786 41246 32788 41298
rect 32732 39732 32788 41246
rect 32620 39676 32732 39732
rect 32284 38724 32340 38734
rect 32172 38612 32228 38622
rect 32172 38162 32228 38556
rect 32172 38110 32174 38162
rect 32226 38110 32228 38162
rect 32172 38098 32228 38110
rect 32172 37492 32228 37502
rect 32284 37492 32340 38668
rect 32228 37436 32340 37492
rect 32620 38162 32676 39676
rect 32732 39666 32788 39676
rect 33180 40402 33236 40414
rect 33180 40350 33182 40402
rect 33234 40350 33236 40402
rect 32732 39508 32788 39518
rect 32732 39506 33124 39508
rect 32732 39454 32734 39506
rect 32786 39454 33124 39506
rect 32732 39452 33124 39454
rect 32732 39442 32788 39452
rect 33068 39058 33124 39452
rect 33068 39006 33070 39058
rect 33122 39006 33124 39058
rect 33068 38994 33124 39006
rect 32620 38110 32622 38162
rect 32674 38110 32676 38162
rect 32172 37378 32228 37436
rect 32172 37326 32174 37378
rect 32226 37326 32228 37378
rect 32172 37314 32228 37326
rect 32620 36482 32676 38110
rect 32620 36430 32622 36482
rect 32674 36430 32676 36482
rect 32620 35924 32676 36430
rect 32620 35858 32676 35868
rect 32060 35634 32116 35644
rect 32396 35810 32452 35822
rect 32396 35758 32398 35810
rect 32450 35758 32452 35810
rect 32060 35028 32116 35038
rect 32396 35028 32452 35758
rect 32844 35028 32900 35038
rect 32060 35026 32900 35028
rect 32060 34974 32062 35026
rect 32114 34974 32846 35026
rect 32898 34974 32900 35026
rect 32060 34972 32900 34974
rect 32060 34962 32116 34972
rect 32844 34962 32900 34972
rect 32060 34804 32116 34814
rect 32060 34354 32116 34748
rect 32508 34692 32564 34702
rect 32060 34302 32062 34354
rect 32114 34302 32116 34354
rect 32060 34290 32116 34302
rect 32396 34690 32564 34692
rect 32396 34638 32510 34690
rect 32562 34638 32564 34690
rect 32396 34636 32564 34638
rect 32396 34242 32452 34636
rect 32508 34626 32564 34636
rect 32396 34190 32398 34242
rect 32450 34190 32452 34242
rect 32396 34178 32452 34190
rect 31948 34076 32228 34132
rect 32060 33908 32116 33918
rect 32060 33460 32116 33852
rect 31500 33458 32116 33460
rect 31500 33406 32062 33458
rect 32114 33406 32116 33458
rect 31500 33404 32116 33406
rect 31500 32562 31556 33404
rect 32060 33366 32116 33404
rect 31500 32510 31502 32562
rect 31554 32510 31556 32562
rect 31500 32498 31556 32510
rect 32172 33124 32228 34076
rect 33180 34130 33236 40350
rect 33292 38612 33348 43486
rect 33628 41186 33684 41198
rect 33628 41134 33630 41186
rect 33682 41134 33684 41186
rect 33628 41076 33684 41134
rect 33628 41010 33684 41020
rect 33516 40852 33572 40862
rect 33516 40290 33572 40796
rect 33516 40238 33518 40290
rect 33570 40238 33572 40290
rect 33516 40226 33572 40238
rect 33404 38836 33460 38846
rect 33404 38742 33460 38780
rect 33292 38546 33348 38556
rect 33740 36484 33796 44270
rect 33964 43652 34020 44604
rect 34524 44548 34580 44558
rect 34524 44454 34580 44492
rect 33964 43586 34020 43596
rect 34412 43764 34468 43774
rect 34076 43428 34132 43438
rect 34076 43334 34132 43372
rect 34188 42532 34244 42542
rect 34188 42438 34244 42476
rect 33852 41858 33908 41870
rect 33852 41806 33854 41858
rect 33906 41806 33908 41858
rect 33852 41074 33908 41806
rect 33852 41022 33854 41074
rect 33906 41022 33908 41074
rect 33852 41010 33908 41022
rect 34300 41076 34356 41086
rect 34300 40982 34356 41020
rect 33964 40402 34020 40414
rect 33964 40350 33966 40402
rect 34018 40350 34020 40402
rect 33964 40292 34020 40350
rect 34412 40292 34468 43708
rect 35196 43148 35460 43158
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35196 43082 35460 43092
rect 34524 42980 34580 42990
rect 34524 42886 34580 42924
rect 35084 42756 35140 42766
rect 34748 42642 34804 42654
rect 34748 42590 34750 42642
rect 34802 42590 34804 42642
rect 34636 41860 34692 41870
rect 34636 41410 34692 41804
rect 34636 41358 34638 41410
rect 34690 41358 34692 41410
rect 34636 41346 34692 41358
rect 34748 40852 34804 42590
rect 34748 40786 34804 40796
rect 35084 42642 35140 42700
rect 35084 42590 35086 42642
rect 35138 42590 35140 42642
rect 33964 40068 34020 40236
rect 33964 40002 34020 40012
rect 34300 40290 34468 40292
rect 34300 40238 34414 40290
rect 34466 40238 34468 40290
rect 34300 40236 34468 40238
rect 34076 38836 34132 38846
rect 34076 38742 34132 38780
rect 34300 38612 34356 40236
rect 34412 40226 34468 40236
rect 34972 40628 35028 40638
rect 34860 40180 34916 40190
rect 34860 39732 34916 40124
rect 34412 39730 34916 39732
rect 34412 39678 34862 39730
rect 34914 39678 34916 39730
rect 34412 39676 34916 39678
rect 34412 38834 34468 39676
rect 34860 39666 34916 39676
rect 34972 39508 35028 40572
rect 34412 38782 34414 38834
rect 34466 38782 34468 38834
rect 34412 38770 34468 38782
rect 34524 39452 35028 39508
rect 35084 39508 35140 42590
rect 35868 41972 35924 45836
rect 35980 45826 36036 45836
rect 36316 45108 36372 45118
rect 35980 44212 36036 44222
rect 35980 43538 36036 44156
rect 35980 43486 35982 43538
rect 36034 43486 36036 43538
rect 35980 43474 36036 43486
rect 35868 41906 35924 41916
rect 36204 42754 36260 42766
rect 36204 42702 36206 42754
rect 36258 42702 36260 42754
rect 35980 41860 36036 41870
rect 35980 41766 36036 41804
rect 35196 41580 35460 41590
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35196 41514 35460 41524
rect 36204 41412 36260 42702
rect 36316 41972 36372 45052
rect 36428 42980 36484 46508
rect 36988 46114 37044 46956
rect 36988 46062 36990 46114
rect 37042 46062 37044 46114
rect 36988 46050 37044 46062
rect 37324 45892 37380 45902
rect 37100 45108 37156 45118
rect 37100 45014 37156 45052
rect 36764 44994 36820 45006
rect 36764 44942 36766 44994
rect 36818 44942 36820 44994
rect 36764 43540 36820 44942
rect 37100 44436 37156 44446
rect 37100 44342 37156 44380
rect 36764 43474 36820 43484
rect 36988 43652 37044 43662
rect 36988 43426 37044 43596
rect 36988 43374 36990 43426
rect 37042 43374 37044 43426
rect 36988 43362 37044 43374
rect 36428 42914 36484 42924
rect 37212 42980 37268 42990
rect 37212 42886 37268 42924
rect 36428 42532 36484 42542
rect 36428 42530 36932 42532
rect 36428 42478 36430 42530
rect 36482 42478 36932 42530
rect 36428 42476 36932 42478
rect 36428 42466 36484 42476
rect 36876 41972 36932 42476
rect 37100 41972 37156 41982
rect 36316 41970 36708 41972
rect 36316 41918 36318 41970
rect 36370 41918 36708 41970
rect 36316 41916 36708 41918
rect 36876 41970 37156 41972
rect 36876 41918 37102 41970
rect 37154 41918 37156 41970
rect 36876 41916 37156 41918
rect 36316 41906 36372 41916
rect 36204 41346 36260 41356
rect 35196 41186 35252 41198
rect 35196 41134 35198 41186
rect 35250 41134 35252 41186
rect 35196 40852 35252 41134
rect 36204 41188 36260 41198
rect 36204 41094 36260 41132
rect 35420 41076 35476 41086
rect 35420 41074 35588 41076
rect 35420 41022 35422 41074
rect 35474 41022 35588 41074
rect 35420 41020 35588 41022
rect 35420 41010 35476 41020
rect 35196 40786 35252 40796
rect 35196 40402 35252 40414
rect 35196 40350 35198 40402
rect 35250 40350 35252 40402
rect 35196 40292 35252 40350
rect 35196 40226 35252 40236
rect 35196 40012 35460 40022
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35196 39946 35460 39956
rect 35532 39620 35588 41020
rect 36428 40964 36484 40974
rect 36428 40870 36484 40908
rect 36316 40628 36372 40638
rect 36316 40534 36372 40572
rect 35644 40516 35700 40526
rect 35644 40422 35700 40460
rect 36652 40404 36708 41916
rect 37100 41906 37156 41916
rect 37212 41412 37268 41422
rect 37212 41318 37268 41356
rect 36428 40402 36708 40404
rect 36428 40350 36654 40402
rect 36706 40350 36708 40402
rect 36428 40348 36708 40350
rect 35420 39564 35588 39620
rect 35868 39732 35924 39742
rect 35196 39508 35252 39518
rect 35084 39506 35252 39508
rect 35084 39454 35198 39506
rect 35250 39454 35252 39506
rect 35084 39452 35252 39454
rect 34524 39060 34580 39452
rect 35196 39442 35252 39452
rect 34412 38612 34468 38622
rect 34300 38556 34412 38612
rect 34412 38546 34468 38556
rect 34524 38162 34580 39004
rect 34524 38110 34526 38162
rect 34578 38110 34580 38162
rect 34524 38098 34580 38110
rect 35084 38946 35140 38958
rect 35084 38894 35086 38946
rect 35138 38894 35140 38946
rect 34860 38050 34916 38062
rect 34860 37998 34862 38050
rect 34914 37998 34916 38050
rect 33740 36428 33908 36484
rect 33292 36372 33348 36382
rect 33292 36370 33796 36372
rect 33292 36318 33294 36370
rect 33346 36318 33796 36370
rect 33292 36316 33796 36318
rect 33292 36306 33348 36316
rect 33292 35924 33348 35934
rect 33292 35830 33348 35868
rect 33740 35922 33796 36316
rect 33740 35870 33742 35922
rect 33794 35870 33796 35922
rect 33740 35858 33796 35870
rect 33516 34914 33572 34926
rect 33516 34862 33518 34914
rect 33570 34862 33572 34914
rect 33404 34804 33460 34814
rect 33404 34710 33460 34748
rect 33180 34078 33182 34130
rect 33234 34078 33236 34130
rect 32956 33460 33012 33470
rect 32956 33348 33012 33404
rect 32732 33346 33012 33348
rect 32732 33294 32958 33346
rect 33010 33294 33012 33346
rect 32732 33292 33012 33294
rect 32396 33234 32452 33246
rect 32396 33182 32398 33234
rect 32450 33182 32452 33234
rect 32396 33124 32452 33182
rect 32172 33068 32452 33124
rect 32172 32562 32228 33068
rect 32284 32676 32340 32686
rect 32284 32582 32340 32620
rect 32172 32510 32174 32562
rect 32226 32510 32228 32562
rect 32172 32498 32228 32510
rect 31388 31892 31668 31948
rect 31388 31108 31444 31118
rect 31388 31014 31444 31052
rect 31612 31106 31668 31892
rect 32060 31892 32116 31902
rect 32060 31798 32116 31836
rect 32396 31780 32452 31790
rect 32396 31686 32452 31724
rect 31612 31054 31614 31106
rect 31666 31054 31668 31106
rect 31276 29474 31332 29484
rect 31276 29316 31332 29326
rect 31164 29314 31332 29316
rect 31164 29262 31278 29314
rect 31330 29262 31332 29314
rect 31164 29260 31332 29262
rect 30716 28868 30772 28878
rect 30716 28774 30772 28812
rect 30268 28756 30324 28766
rect 30156 28700 30268 28756
rect 30268 28662 30324 28700
rect 29484 27806 29486 27858
rect 29538 27806 29540 27858
rect 29484 27794 29540 27806
rect 31052 28644 31108 28654
rect 31164 28644 31220 29260
rect 31276 29250 31332 29260
rect 31052 28642 31220 28644
rect 31052 28590 31054 28642
rect 31106 28590 31220 28642
rect 31052 28588 31220 28590
rect 30268 27746 30324 27758
rect 30268 27694 30270 27746
rect 30322 27694 30324 27746
rect 30268 26962 30324 27694
rect 31052 27300 31108 28588
rect 31612 28530 31668 31054
rect 31836 30100 31892 30110
rect 31836 28756 31892 30044
rect 32732 28980 32788 33292
rect 32956 33282 33012 33292
rect 33180 31948 33236 34078
rect 33516 34020 33572 34862
rect 33516 33926 33572 33964
rect 33852 33908 33908 36428
rect 34860 36260 34916 37998
rect 34860 36194 34916 36204
rect 35084 36708 35140 38894
rect 35196 38834 35252 38846
rect 35196 38782 35198 38834
rect 35250 38782 35252 38834
rect 35196 38612 35252 38782
rect 35420 38612 35476 39564
rect 35532 39396 35588 39406
rect 35532 39394 35700 39396
rect 35532 39342 35534 39394
rect 35586 39342 35700 39394
rect 35532 39340 35700 39342
rect 35532 39330 35588 39340
rect 35420 38556 35588 38612
rect 35196 38546 35252 38556
rect 35196 38444 35460 38454
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35196 38378 35460 38388
rect 35420 37492 35476 37502
rect 35532 37492 35588 38556
rect 35476 37436 35588 37492
rect 35420 37398 35476 37436
rect 35196 36876 35460 36886
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35196 36810 35460 36820
rect 35084 36652 35476 36708
rect 34076 35700 34132 35710
rect 34636 35700 34692 35710
rect 34076 35698 34692 35700
rect 34076 35646 34078 35698
rect 34130 35646 34638 35698
rect 34690 35646 34692 35698
rect 34076 35644 34692 35646
rect 34076 35634 34132 35644
rect 34636 35634 34692 35644
rect 34972 35700 35028 35710
rect 35084 35700 35140 36652
rect 35420 36594 35476 36652
rect 35420 36542 35422 36594
rect 35474 36542 35476 36594
rect 35420 36530 35476 36542
rect 35308 36484 35364 36494
rect 35308 35810 35364 36428
rect 35308 35758 35310 35810
rect 35362 35758 35364 35810
rect 35308 35746 35364 35758
rect 35532 35810 35588 35822
rect 35532 35758 35534 35810
rect 35586 35758 35588 35810
rect 34972 35698 35140 35700
rect 34972 35646 34974 35698
rect 35026 35646 35140 35698
rect 34972 35644 35140 35646
rect 34972 35634 35028 35644
rect 35196 35308 35460 35318
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35196 35242 35460 35252
rect 34636 34916 34692 34926
rect 34636 34914 34804 34916
rect 34636 34862 34638 34914
rect 34690 34862 34804 34914
rect 34636 34860 34804 34862
rect 34636 34850 34692 34860
rect 33852 33842 33908 33852
rect 33964 34018 34020 34030
rect 33964 33966 33966 34018
rect 34018 33966 34020 34018
rect 33404 33460 33460 33470
rect 33404 33366 33460 33404
rect 33964 33348 34020 33966
rect 34748 33572 34804 34860
rect 35532 34804 35588 35758
rect 34860 34692 34916 34702
rect 34860 34598 34916 34636
rect 35532 33908 35588 34748
rect 35532 33842 35588 33852
rect 35196 33740 35460 33750
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35196 33674 35460 33684
rect 34860 33572 34916 33582
rect 34748 33570 34916 33572
rect 34748 33518 34862 33570
rect 34914 33518 34916 33570
rect 34748 33516 34916 33518
rect 34860 33506 34916 33516
rect 33964 32676 34020 33292
rect 35196 33348 35252 33358
rect 35196 33254 35252 33292
rect 33964 32610 34020 32620
rect 35532 33236 35588 33246
rect 35196 32172 35460 32182
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35196 32106 35460 32116
rect 32732 28914 32788 28924
rect 32844 31892 33236 31948
rect 31836 28642 31892 28700
rect 31836 28590 31838 28642
rect 31890 28590 31892 28642
rect 31836 28578 31892 28590
rect 31612 28478 31614 28530
rect 31666 28478 31668 28530
rect 31612 28466 31668 28478
rect 32844 28532 32900 31892
rect 35308 31890 35364 31902
rect 35308 31838 35310 31890
rect 35362 31838 35364 31890
rect 33180 31668 33236 31678
rect 34636 31668 34692 31678
rect 33180 31666 33460 31668
rect 33180 31614 33182 31666
rect 33234 31614 33460 31666
rect 33180 31612 33460 31614
rect 33180 31602 33236 31612
rect 33404 31218 33460 31612
rect 33404 31166 33406 31218
rect 33458 31166 33460 31218
rect 33404 31154 33460 31166
rect 33740 30996 33796 31006
rect 34300 30996 34356 31006
rect 33740 30994 34356 30996
rect 33740 30942 33742 30994
rect 33794 30942 34302 30994
rect 34354 30942 34356 30994
rect 33740 30940 34356 30942
rect 33740 30930 33796 30940
rect 34300 30930 34356 30940
rect 34636 30994 34692 31612
rect 35308 31668 35364 31838
rect 35308 31602 35364 31612
rect 34860 31108 34916 31118
rect 34860 31014 34916 31052
rect 35420 31108 35476 31118
rect 35532 31108 35588 33180
rect 35644 31948 35700 39340
rect 35868 38834 35924 39676
rect 36428 39732 36484 40348
rect 36652 40338 36708 40348
rect 37324 40180 37380 45836
rect 37660 45220 37716 49200
rect 37660 45154 37716 45164
rect 37884 45668 37940 45678
rect 37884 45218 37940 45612
rect 37884 45166 37886 45218
rect 37938 45166 37940 45218
rect 37884 45154 37940 45166
rect 37772 45108 37828 45118
rect 37772 44322 37828 45052
rect 38332 45108 38388 49200
rect 39676 46116 39732 49200
rect 39676 46060 40180 46116
rect 39788 45892 39844 45902
rect 39788 45798 39844 45836
rect 39228 45778 39284 45790
rect 39228 45726 39230 45778
rect 39282 45726 39284 45778
rect 38892 45668 38948 45678
rect 38892 45574 38948 45612
rect 38332 45042 38388 45052
rect 37772 44270 37774 44322
rect 37826 44270 37828 44322
rect 37772 44258 37828 44270
rect 39004 44884 39060 44894
rect 38556 44210 38612 44222
rect 38556 44158 38558 44210
rect 38610 44158 38612 44210
rect 38556 43652 38612 44158
rect 38556 43586 38612 43596
rect 38668 43876 38724 43886
rect 37548 41972 37604 41982
rect 37548 41410 37604 41916
rect 38668 41636 38724 43820
rect 39004 43650 39060 44828
rect 39228 44548 39284 45726
rect 39228 44482 39284 44492
rect 40012 44994 40068 45006
rect 40012 44942 40014 44994
rect 40066 44942 40068 44994
rect 40012 43988 40068 44942
rect 40012 43922 40068 43932
rect 39004 43598 39006 43650
rect 39058 43598 39060 43650
rect 39004 43586 39060 43598
rect 39564 43764 39620 43774
rect 39564 43650 39620 43708
rect 39564 43598 39566 43650
rect 39618 43598 39620 43650
rect 39564 43586 39620 43598
rect 39900 43650 39956 43662
rect 39900 43598 39902 43650
rect 39954 43598 39956 43650
rect 39340 43540 39396 43550
rect 39340 42754 39396 43484
rect 39340 42702 39342 42754
rect 39394 42702 39396 42754
rect 39340 42690 39396 42702
rect 39228 41972 39284 41982
rect 39228 41858 39284 41916
rect 39228 41806 39230 41858
rect 39282 41806 39284 41858
rect 39228 41748 39284 41806
rect 39228 41682 39284 41692
rect 39676 41972 39732 41982
rect 37548 41358 37550 41410
rect 37602 41358 37604 41410
rect 37548 41346 37604 41358
rect 38332 41580 38724 41636
rect 37772 41074 37828 41086
rect 37772 41022 37774 41074
rect 37826 41022 37828 41074
rect 37436 40964 37492 40974
rect 37436 40514 37492 40908
rect 37436 40462 37438 40514
rect 37490 40462 37492 40514
rect 37436 40450 37492 40462
rect 37772 40516 37828 41022
rect 38220 41076 38276 41086
rect 38220 40982 38276 41020
rect 37772 40450 37828 40460
rect 37324 40114 37380 40124
rect 37772 40180 37828 40190
rect 36428 39638 36484 39676
rect 37100 39732 37156 39742
rect 37100 39638 37156 39676
rect 37772 39506 37828 40124
rect 38332 39842 38388 41580
rect 38892 41188 38948 41198
rect 38892 41094 38948 41132
rect 39228 41186 39284 41198
rect 39228 41134 39230 41186
rect 39282 41134 39284 41186
rect 39228 41076 39284 41134
rect 39676 41186 39732 41916
rect 39900 41860 39956 43598
rect 40124 42978 40180 46060
rect 42924 45892 42980 45902
rect 42812 45890 42980 45892
rect 42812 45838 42926 45890
rect 42978 45838 42980 45890
rect 42812 45836 42980 45838
rect 40796 45666 40852 45678
rect 42700 45668 42756 45678
rect 40796 45614 40798 45666
rect 40850 45614 40852 45666
rect 40796 45332 40852 45614
rect 40796 45266 40852 45276
rect 42588 45666 42756 45668
rect 42588 45614 42702 45666
rect 42754 45614 42756 45666
rect 42588 45612 42756 45614
rect 42028 45220 42084 45230
rect 41804 45106 41860 45118
rect 41804 45054 41806 45106
rect 41858 45054 41860 45106
rect 41132 44996 41188 45006
rect 41580 44996 41636 45006
rect 41804 44996 41860 45054
rect 41132 44994 41860 44996
rect 41132 44942 41134 44994
rect 41186 44942 41582 44994
rect 41634 44942 41860 44994
rect 41132 44940 41860 44942
rect 40684 44436 40740 44446
rect 40684 44342 40740 44380
rect 41020 44324 41076 44334
rect 40124 42926 40126 42978
rect 40178 42926 40180 42978
rect 40124 42914 40180 42926
rect 40796 44322 41076 44324
rect 40796 44270 41022 44322
rect 41074 44270 41076 44322
rect 40796 44268 41076 44270
rect 39900 41794 39956 41804
rect 40124 41860 40180 41870
rect 39676 41134 39678 41186
rect 39730 41134 39732 41186
rect 39284 41020 39396 41076
rect 39228 41010 39284 41020
rect 39340 40852 39396 41020
rect 39340 40796 39620 40852
rect 39340 40628 39396 40638
rect 38780 40404 38836 40414
rect 38332 39790 38334 39842
rect 38386 39790 38388 39842
rect 38332 39778 38388 39790
rect 38668 39844 38724 39854
rect 38668 39750 38724 39788
rect 37772 39454 37774 39506
rect 37826 39454 37828 39506
rect 37772 39442 37828 39454
rect 38108 39506 38164 39518
rect 38108 39454 38110 39506
rect 38162 39454 38164 39506
rect 38108 38948 38164 39454
rect 38108 38882 38164 38892
rect 35868 38782 35870 38834
rect 35922 38782 35924 38834
rect 35868 38770 35924 38782
rect 36540 38724 36596 38734
rect 36428 38722 36596 38724
rect 36428 38670 36542 38722
rect 36594 38670 36596 38722
rect 36428 38668 36596 38670
rect 36204 38050 36260 38062
rect 36204 37998 36206 38050
rect 36258 37998 36260 38050
rect 36204 37940 36260 37998
rect 36204 37874 36260 37884
rect 36428 37938 36484 38668
rect 36540 38658 36596 38668
rect 37548 38724 37604 38734
rect 37548 38274 37604 38668
rect 38668 38724 38724 38762
rect 38668 38658 38724 38668
rect 37548 38222 37550 38274
rect 37602 38222 37604 38274
rect 37548 38210 37604 38222
rect 37772 38612 37828 38622
rect 36428 37886 36430 37938
rect 36482 37886 36484 37938
rect 36428 37874 36484 37886
rect 37212 37940 37268 37950
rect 37212 37846 37268 37884
rect 37772 37938 37828 38556
rect 37772 37886 37774 37938
rect 37826 37886 37828 37938
rect 37772 37874 37828 37886
rect 38220 37938 38276 37950
rect 38220 37886 38222 37938
rect 38274 37886 38276 37938
rect 37772 37378 37828 37390
rect 37772 37326 37774 37378
rect 37826 37326 37828 37378
rect 35756 37266 35812 37278
rect 35756 37214 35758 37266
rect 35810 37214 35812 37266
rect 35756 37156 35812 37214
rect 37548 37268 37604 37278
rect 37548 37266 37716 37268
rect 37548 37214 37550 37266
rect 37602 37214 37716 37266
rect 37548 37212 37716 37214
rect 37548 37202 37604 37212
rect 36204 37156 36260 37166
rect 35756 37154 36484 37156
rect 35756 37102 36206 37154
rect 36258 37102 36484 37154
rect 35756 37100 36484 37102
rect 36204 37090 36260 37100
rect 36316 36484 36372 36494
rect 36316 36390 36372 36428
rect 35756 36260 35812 36270
rect 35756 36166 35812 36204
rect 36092 34692 36148 34702
rect 36092 34242 36148 34636
rect 36092 34190 36094 34242
rect 36146 34190 36148 34242
rect 36092 34178 36148 34190
rect 35756 34020 35812 34030
rect 35756 33346 35812 33964
rect 35756 33294 35758 33346
rect 35810 33294 35812 33346
rect 35756 32676 35812 33294
rect 35980 33236 36036 33246
rect 35980 33142 36036 33180
rect 35756 32610 35812 32620
rect 35644 31892 36148 31948
rect 35420 31106 35588 31108
rect 35420 31054 35422 31106
rect 35474 31054 35588 31106
rect 35420 31052 35588 31054
rect 35420 31042 35476 31052
rect 34636 30942 34638 30994
rect 34690 30942 34692 30994
rect 34636 30930 34692 30942
rect 35196 30604 35460 30614
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35196 30538 35460 30548
rect 34860 30322 34916 30334
rect 34860 30270 34862 30322
rect 34914 30270 34916 30322
rect 33180 29988 33236 29998
rect 33068 29314 33124 29326
rect 33068 29262 33070 29314
rect 33122 29262 33124 29314
rect 33068 29204 33124 29262
rect 33068 29138 33124 29148
rect 33180 28642 33236 29932
rect 34076 29986 34132 29998
rect 34076 29934 34078 29986
rect 34130 29934 34132 29986
rect 34076 29764 34132 29934
rect 34524 29988 34580 29998
rect 34524 29894 34580 29932
rect 34076 29698 34132 29708
rect 33180 28590 33182 28642
rect 33234 28590 33236 28642
rect 33180 28578 33236 28590
rect 33404 29316 33460 29326
rect 32844 28466 32900 28476
rect 33404 28530 33460 29260
rect 34860 29204 34916 30270
rect 35420 30100 35476 30110
rect 35532 30100 35588 31052
rect 35980 30994 36036 31006
rect 35980 30942 35982 30994
rect 36034 30942 36036 30994
rect 35420 30098 35588 30100
rect 35420 30046 35422 30098
rect 35474 30046 35588 30098
rect 35420 30044 35588 30046
rect 35644 30210 35700 30222
rect 35644 30158 35646 30210
rect 35698 30158 35700 30210
rect 35196 29316 35252 29326
rect 35196 29222 35252 29260
rect 35420 29316 35476 30044
rect 35644 29764 35700 30158
rect 35644 29698 35700 29708
rect 35980 29428 36036 30942
rect 35980 29334 36036 29372
rect 35420 29250 35476 29260
rect 34860 28868 34916 29148
rect 35196 29036 35460 29046
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35196 28970 35460 28980
rect 35420 28868 35476 28878
rect 34860 28866 35476 28868
rect 34860 28814 35422 28866
rect 35474 28814 35476 28866
rect 34860 28812 35476 28814
rect 35420 28802 35476 28812
rect 33404 28478 33406 28530
rect 33458 28478 33460 28530
rect 33404 28466 33460 28478
rect 35868 28642 35924 28654
rect 35868 28590 35870 28642
rect 35922 28590 35924 28642
rect 35084 28420 35140 28430
rect 34748 28418 35140 28420
rect 34748 28366 35086 28418
rect 35138 28366 35140 28418
rect 34748 28364 35140 28366
rect 33628 27858 33684 27870
rect 33628 27806 33630 27858
rect 33682 27806 33684 27858
rect 32396 27746 32452 27758
rect 32396 27694 32398 27746
rect 32450 27694 32452 27746
rect 31388 27300 31444 27310
rect 32396 27300 32452 27694
rect 31052 27298 31444 27300
rect 31052 27246 31390 27298
rect 31442 27246 31444 27298
rect 31052 27244 31444 27246
rect 31388 27234 31444 27244
rect 32172 27244 32396 27300
rect 31612 27076 31668 27086
rect 30268 26910 30270 26962
rect 30322 26910 30324 26962
rect 30268 26898 30324 26910
rect 30604 26964 30660 26974
rect 31052 26964 31108 26974
rect 30604 26962 31108 26964
rect 30604 26910 30606 26962
rect 30658 26910 31054 26962
rect 31106 26910 31108 26962
rect 30604 26908 31108 26910
rect 30604 26898 30660 26908
rect 31052 26898 31108 26908
rect 31612 26962 31668 27020
rect 31612 26910 31614 26962
rect 31666 26910 31668 26962
rect 31612 26898 31668 26910
rect 32172 26962 32228 27244
rect 32396 27234 32452 27244
rect 32172 26910 32174 26962
rect 32226 26910 32228 26962
rect 32172 26898 32228 26910
rect 29484 26404 29540 26414
rect 28700 24782 28702 24834
rect 28754 24782 28756 24834
rect 28588 23940 28644 23950
rect 28588 23846 28644 23884
rect 28700 23604 28756 24782
rect 29372 25508 29428 25518
rect 29260 24724 29316 24734
rect 29260 24050 29316 24668
rect 29260 23998 29262 24050
rect 29314 23998 29316 24050
rect 29260 23986 29316 23998
rect 28700 23538 28756 23548
rect 29036 23938 29092 23950
rect 29036 23886 29038 23938
rect 29090 23886 29092 23938
rect 29036 23492 29092 23886
rect 29372 23940 29428 25452
rect 29372 23874 29428 23884
rect 29484 23938 29540 26348
rect 33068 26292 33124 26302
rect 33628 26292 33684 27806
rect 34412 27746 34468 27758
rect 34412 27694 34414 27746
rect 34466 27694 34468 27746
rect 34412 26962 34468 27694
rect 34748 27074 34804 28364
rect 35084 28354 35140 28364
rect 35196 27468 35460 27478
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35196 27402 35460 27412
rect 34748 27022 34750 27074
rect 34802 27022 34804 27074
rect 34748 27010 34804 27022
rect 35868 27076 35924 28590
rect 35868 27010 35924 27020
rect 34412 26910 34414 26962
rect 34466 26910 34468 26962
rect 34412 26898 34468 26910
rect 33068 26290 33684 26292
rect 33068 26238 33070 26290
rect 33122 26238 33684 26290
rect 33068 26236 33684 26238
rect 30380 25620 30436 25630
rect 30044 25394 30100 25406
rect 30044 25342 30046 25394
rect 30098 25342 30100 25394
rect 30044 24948 30100 25342
rect 30044 24882 30100 24892
rect 29484 23886 29486 23938
rect 29538 23886 29540 23938
rect 29484 23874 29540 23886
rect 29596 23938 29652 23950
rect 29596 23886 29598 23938
rect 29650 23886 29652 23938
rect 29036 23154 29092 23436
rect 29372 23380 29428 23390
rect 29372 23286 29428 23324
rect 29484 23268 29540 23278
rect 29484 23174 29540 23212
rect 29036 23102 29038 23154
rect 29090 23102 29092 23154
rect 29036 23090 29092 23102
rect 28364 22754 28420 22764
rect 26348 22642 26404 22652
rect 28140 22484 28196 22494
rect 26124 22428 26516 22484
rect 26012 22260 26068 22270
rect 26012 22258 26292 22260
rect 26012 22206 26014 22258
rect 26066 22206 26292 22258
rect 26012 22204 26292 22206
rect 26012 22194 26068 22204
rect 26124 21812 26180 21822
rect 25900 21810 26180 21812
rect 25900 21758 26126 21810
rect 26178 21758 26180 21810
rect 25900 21756 26180 21758
rect 26124 21746 26180 21756
rect 26236 21810 26292 22204
rect 26236 21758 26238 21810
rect 26290 21758 26292 21810
rect 26236 21746 26292 21758
rect 26348 21588 26404 21598
rect 26236 21586 26404 21588
rect 26236 21534 26350 21586
rect 26402 21534 26404 21586
rect 26236 21532 26404 21534
rect 25900 20804 25956 20814
rect 25452 20802 25956 20804
rect 25452 20750 25902 20802
rect 25954 20750 25956 20802
rect 25452 20748 25956 20750
rect 25452 20690 25508 20748
rect 25900 20738 25956 20748
rect 25452 20638 25454 20690
rect 25506 20638 25508 20690
rect 25452 20626 25508 20638
rect 24220 18060 24500 18116
rect 24780 20580 24836 20590
rect 25116 20580 25172 20590
rect 24780 20578 25172 20580
rect 24780 20526 24782 20578
rect 24834 20526 25118 20578
rect 25170 20526 25172 20578
rect 24780 20524 25172 20526
rect 24220 17108 24276 18060
rect 24220 17106 24612 17108
rect 24220 17054 24222 17106
rect 24274 17054 24612 17106
rect 24220 17052 24612 17054
rect 24220 17042 24276 17052
rect 23884 16098 24052 16100
rect 23884 16046 23886 16098
rect 23938 16046 24052 16098
rect 23884 16044 24052 16046
rect 23884 16034 23940 16044
rect 23100 15484 23380 15540
rect 23436 15988 23492 15998
rect 22988 13634 23044 13646
rect 22988 13582 22990 13634
rect 23042 13582 23044 13634
rect 22988 13522 23044 13582
rect 22988 13470 22990 13522
rect 23042 13470 23044 13522
rect 22988 13458 23044 13470
rect 23100 13300 23156 15484
rect 23436 15148 23492 15932
rect 24332 15988 24388 15998
rect 24332 15894 24388 15932
rect 23996 15874 24052 15886
rect 23996 15822 23998 15874
rect 24050 15822 24052 15874
rect 23996 15316 24052 15822
rect 24108 15876 24164 15886
rect 24108 15782 24164 15820
rect 24444 15764 24500 15774
rect 24444 15538 24500 15708
rect 24444 15486 24446 15538
rect 24498 15486 24500 15538
rect 24444 15474 24500 15486
rect 23996 15250 24052 15260
rect 24108 15314 24164 15326
rect 24108 15262 24110 15314
rect 24162 15262 24164 15314
rect 23548 15204 23604 15214
rect 23324 15092 23604 15148
rect 24108 15204 24164 15262
rect 24220 15316 24276 15326
rect 24220 15222 24276 15260
rect 24444 15202 24500 15214
rect 24444 15150 24446 15202
rect 24498 15150 24500 15202
rect 24108 15092 24388 15148
rect 23324 13858 23380 15092
rect 23660 14644 23716 14654
rect 23660 14550 23716 14588
rect 23548 14530 23604 14542
rect 23548 14478 23550 14530
rect 23602 14478 23604 14530
rect 23548 14420 23604 14478
rect 24332 14530 24388 15092
rect 24332 14478 24334 14530
rect 24386 14478 24388 14530
rect 24332 14466 24388 14478
rect 23324 13806 23326 13858
rect 23378 13806 23380 13858
rect 23324 13794 23380 13806
rect 23436 14364 23604 14420
rect 23996 14418 24052 14430
rect 23996 14366 23998 14418
rect 24050 14366 24052 14418
rect 23436 13748 23492 14364
rect 23996 14084 24052 14366
rect 23548 14028 24052 14084
rect 24444 14084 24500 15150
rect 24556 14532 24612 17052
rect 24780 16436 24836 20524
rect 25116 20514 25172 20524
rect 26124 20578 26180 20590
rect 26124 20526 26126 20578
rect 26178 20526 26180 20578
rect 25564 20018 25620 20030
rect 25564 19966 25566 20018
rect 25618 19966 25620 20018
rect 25564 19572 25620 19966
rect 25564 19516 25844 19572
rect 25564 19348 25620 19358
rect 25564 19254 25620 19292
rect 25452 18676 25508 18686
rect 25452 18582 25508 18620
rect 25788 18564 25844 19516
rect 25340 18450 25396 18462
rect 25340 18398 25342 18450
rect 25394 18398 25396 18450
rect 25228 17668 25284 17678
rect 25228 17108 25284 17612
rect 25340 17220 25396 18398
rect 25676 18452 25732 18462
rect 25676 18358 25732 18396
rect 25564 18340 25620 18350
rect 25564 18246 25620 18284
rect 25788 17666 25844 18508
rect 25900 19348 25956 19358
rect 25900 18676 25956 19292
rect 26124 19236 26180 20526
rect 26236 20132 26292 21532
rect 26348 21522 26404 21532
rect 26348 20804 26404 20814
rect 26460 20804 26516 22428
rect 27916 22482 28196 22484
rect 27916 22430 28142 22482
rect 28194 22430 28196 22482
rect 27916 22428 28196 22430
rect 27916 21810 27972 22428
rect 28140 22418 28196 22428
rect 29596 22484 29652 23886
rect 30268 23826 30324 23838
rect 30268 23774 30270 23826
rect 30322 23774 30324 23826
rect 30268 23492 30324 23774
rect 30268 23426 30324 23436
rect 30380 23826 30436 25564
rect 32172 25620 32228 25630
rect 32172 25526 32228 25564
rect 33068 25508 33124 26236
rect 33852 26180 33908 26190
rect 35980 26180 36036 26190
rect 36092 26180 36148 31892
rect 36204 28532 36260 28542
rect 36204 28438 36260 28476
rect 33068 25442 33124 25452
rect 33740 26178 33908 26180
rect 33740 26126 33854 26178
rect 33906 26126 33908 26178
rect 33740 26124 33908 26126
rect 33740 25394 33796 26124
rect 33852 26114 33908 26124
rect 35644 26178 36148 26180
rect 35644 26126 35982 26178
rect 36034 26126 36148 26178
rect 35644 26124 36148 26126
rect 36316 26180 36372 26190
rect 35196 25900 35460 25910
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35196 25834 35460 25844
rect 35196 25618 35252 25630
rect 35196 25566 35198 25618
rect 35250 25566 35252 25618
rect 33740 25342 33742 25394
rect 33794 25342 33796 25394
rect 33740 25330 33796 25342
rect 34076 25396 34132 25406
rect 34076 25394 34580 25396
rect 34076 25342 34078 25394
rect 34130 25342 34580 25394
rect 34076 25340 34580 25342
rect 34076 25330 34132 25340
rect 30604 25116 31332 25172
rect 30604 23938 30660 25116
rect 30940 24948 30996 24958
rect 30940 24854 30996 24892
rect 31276 24946 31332 25116
rect 31276 24894 31278 24946
rect 31330 24894 31332 24946
rect 31276 24882 31332 24894
rect 34524 24946 34580 25340
rect 34524 24894 34526 24946
rect 34578 24894 34580 24946
rect 34524 24882 34580 24894
rect 35196 24948 35252 25566
rect 35644 25506 35700 26124
rect 35980 26114 36036 26124
rect 36316 26086 36372 26124
rect 35644 25454 35646 25506
rect 35698 25454 35700 25506
rect 35644 25442 35700 25454
rect 35196 24892 35476 24948
rect 35420 24836 35476 24892
rect 35420 24834 35588 24836
rect 35420 24782 35422 24834
rect 35474 24782 35588 24834
rect 35420 24780 35588 24782
rect 35420 24770 35476 24780
rect 30828 24724 30884 24734
rect 30828 24630 30884 24668
rect 31052 24724 31108 24734
rect 31052 24722 31332 24724
rect 31052 24670 31054 24722
rect 31106 24670 31332 24722
rect 31052 24668 31332 24670
rect 31052 24658 31108 24668
rect 30604 23886 30606 23938
rect 30658 23886 30660 23938
rect 30604 23874 30660 23886
rect 30828 23940 30884 23950
rect 30380 23774 30382 23826
rect 30434 23774 30436 23826
rect 29708 23156 29764 23166
rect 29708 23062 29764 23100
rect 29596 22418 29652 22428
rect 29260 22370 29316 22382
rect 29260 22318 29262 22370
rect 29314 22318 29316 22370
rect 27916 21758 27918 21810
rect 27970 21758 27972 21810
rect 26796 21588 26852 21598
rect 26796 21494 26852 21532
rect 27692 21588 27748 21598
rect 27692 21494 27748 21532
rect 26348 20802 26516 20804
rect 26348 20750 26350 20802
rect 26402 20750 26516 20802
rect 26348 20748 26516 20750
rect 26348 20738 26404 20748
rect 26572 20692 26628 20702
rect 26572 20598 26628 20636
rect 27580 20580 27636 20590
rect 26236 20076 26628 20132
rect 26236 19908 26292 19918
rect 26236 19906 26516 19908
rect 26236 19854 26238 19906
rect 26290 19854 26516 19906
rect 26236 19852 26516 19854
rect 26236 19842 26292 19852
rect 26460 19346 26516 19852
rect 26460 19294 26462 19346
rect 26514 19294 26516 19346
rect 26460 19282 26516 19294
rect 26348 19236 26404 19246
rect 26124 19234 26404 19236
rect 26124 19182 26350 19234
rect 26402 19182 26404 19234
rect 26124 19180 26404 19182
rect 26348 19170 26404 19180
rect 26572 19234 26628 20076
rect 26572 19182 26574 19234
rect 26626 19182 26628 19234
rect 25900 18562 25956 18620
rect 25900 18510 25902 18562
rect 25954 18510 25956 18562
rect 25900 18498 25956 18510
rect 26124 19010 26180 19022
rect 26572 19012 26628 19182
rect 27020 19796 27076 19806
rect 27020 19234 27076 19740
rect 27020 19182 27022 19234
rect 27074 19182 27076 19234
rect 27020 19170 27076 19182
rect 26124 18958 26126 19010
rect 26178 18958 26180 19010
rect 26124 18452 26180 18958
rect 26460 18956 26628 19012
rect 26348 18452 26404 18462
rect 26124 18450 26404 18452
rect 26124 18398 26350 18450
rect 26402 18398 26404 18450
rect 26124 18396 26404 18398
rect 25788 17614 25790 17666
rect 25842 17614 25844 17666
rect 25788 17602 25844 17614
rect 25340 17164 25620 17220
rect 25228 17014 25284 17052
rect 25564 17106 25620 17164
rect 25564 17054 25566 17106
rect 25618 17054 25620 17106
rect 24780 16370 24836 16380
rect 24668 16100 24724 16110
rect 24668 16006 24724 16044
rect 25004 15874 25060 15886
rect 25004 15822 25006 15874
rect 25058 15822 25060 15874
rect 24668 15316 24724 15326
rect 25004 15316 25060 15822
rect 25340 15428 25396 15438
rect 25340 15334 25396 15372
rect 24668 15314 25060 15316
rect 24668 15262 24670 15314
rect 24722 15262 25060 15314
rect 24668 15260 25060 15262
rect 24668 14532 24724 15260
rect 25564 14756 25620 17054
rect 26236 16772 26292 18396
rect 26348 18386 26404 18396
rect 26460 18452 26516 18956
rect 26572 18676 26628 18686
rect 26572 18562 26628 18620
rect 26572 18510 26574 18562
rect 26626 18510 26628 18562
rect 26572 18498 26628 18510
rect 27244 18562 27300 18574
rect 27244 18510 27246 18562
rect 27298 18510 27300 18562
rect 26460 18386 26516 18396
rect 27020 18450 27076 18462
rect 27020 18398 27022 18450
rect 27074 18398 27076 18450
rect 26796 18340 26852 18350
rect 26684 18338 26852 18340
rect 26684 18286 26798 18338
rect 26850 18286 26852 18338
rect 26684 18284 26852 18286
rect 26684 17780 26740 18284
rect 26796 18274 26852 18284
rect 27020 18340 27076 18398
rect 27020 18274 27076 18284
rect 27244 18452 27300 18510
rect 27244 18116 27300 18396
rect 27580 18450 27636 20524
rect 27916 19460 27972 21758
rect 29148 21924 29204 21934
rect 29148 21810 29204 21868
rect 29148 21758 29150 21810
rect 29202 21758 29204 21810
rect 29148 21746 29204 21758
rect 29260 21812 29316 22318
rect 29932 22260 29988 22270
rect 29260 21746 29316 21756
rect 29596 22258 29988 22260
rect 29596 22206 29934 22258
rect 29986 22206 29988 22258
rect 29596 22204 29988 22206
rect 29596 21810 29652 22204
rect 29932 22194 29988 22204
rect 29596 21758 29598 21810
rect 29650 21758 29652 21810
rect 29596 21746 29652 21758
rect 29708 21924 29764 21934
rect 29708 21810 29764 21868
rect 29708 21758 29710 21810
rect 29762 21758 29764 21810
rect 29708 21746 29764 21758
rect 28028 21586 28084 21598
rect 28028 21534 28030 21586
rect 28082 21534 28084 21586
rect 28028 20578 28084 21534
rect 28924 21586 28980 21598
rect 29484 21588 29540 21598
rect 28924 21534 28926 21586
rect 28978 21534 28980 21586
rect 28028 20526 28030 20578
rect 28082 20526 28084 20578
rect 28028 20020 28084 20526
rect 28028 19954 28084 19964
rect 28252 21364 28308 21374
rect 27916 19394 27972 19404
rect 28140 18452 28196 18462
rect 27580 18398 27582 18450
rect 27634 18398 27636 18450
rect 27580 18386 27636 18398
rect 27692 18450 28196 18452
rect 27692 18398 28142 18450
rect 28194 18398 28196 18450
rect 27692 18396 28196 18398
rect 26348 17724 26740 17780
rect 26796 18060 27300 18116
rect 26348 16882 26404 17724
rect 26460 17556 26516 17566
rect 26460 17554 26628 17556
rect 26460 17502 26462 17554
rect 26514 17502 26628 17554
rect 26460 17500 26628 17502
rect 26460 17490 26516 17500
rect 26572 16994 26628 17500
rect 26572 16942 26574 16994
rect 26626 16942 26628 16994
rect 26572 16930 26628 16942
rect 26348 16830 26350 16882
rect 26402 16830 26404 16882
rect 26348 16818 26404 16830
rect 26796 16882 26852 18060
rect 27692 17332 27748 18396
rect 28140 18386 28196 18396
rect 28252 18228 28308 21308
rect 28364 20690 28420 20702
rect 28364 20638 28366 20690
rect 28418 20638 28420 20690
rect 28364 20580 28420 20638
rect 28364 20514 28420 20524
rect 28812 20132 28868 20142
rect 28700 20130 28868 20132
rect 28700 20078 28814 20130
rect 28866 20078 28868 20130
rect 28700 20076 28868 20078
rect 28364 19908 28420 19918
rect 28700 19908 28756 20076
rect 28812 20066 28868 20076
rect 28364 19906 28756 19908
rect 28364 19854 28366 19906
rect 28418 19854 28756 19906
rect 28364 19852 28756 19854
rect 28364 19842 28420 19852
rect 28588 19012 28644 19022
rect 28588 18918 28644 18956
rect 28700 18788 28756 19852
rect 28924 20020 28980 21534
rect 28812 19796 28868 19806
rect 28812 19702 28868 19740
rect 28700 18722 28756 18732
rect 28364 18564 28420 18574
rect 28364 18340 28420 18508
rect 28476 18564 28532 18574
rect 28924 18564 28980 19964
rect 29372 21586 29540 21588
rect 29372 21534 29486 21586
rect 29538 21534 29540 21586
rect 29372 21532 29540 21534
rect 29260 19796 29316 19806
rect 29148 19124 29204 19134
rect 29036 19122 29204 19124
rect 29036 19070 29150 19122
rect 29202 19070 29204 19122
rect 29036 19068 29204 19070
rect 29036 18676 29092 19068
rect 29148 19058 29204 19068
rect 29260 19124 29316 19740
rect 29260 19030 29316 19068
rect 29372 18676 29428 21532
rect 29484 21522 29540 21532
rect 30156 21588 30212 21598
rect 30156 21494 30212 21532
rect 30380 20244 30436 23774
rect 30716 22372 30772 22382
rect 30716 21810 30772 22316
rect 30716 21758 30718 21810
rect 30770 21758 30772 21810
rect 30716 21746 30772 21758
rect 30828 21812 30884 23884
rect 31276 23548 31332 24668
rect 34860 24500 34916 24510
rect 34860 24498 35140 24500
rect 34860 24446 34862 24498
rect 34914 24446 35140 24498
rect 34860 24444 35140 24446
rect 34860 24434 34916 24444
rect 33740 24050 33796 24062
rect 33740 23998 33742 24050
rect 33794 23998 33796 24050
rect 31612 23828 31668 23838
rect 31500 23826 31668 23828
rect 31500 23774 31614 23826
rect 31666 23774 31668 23826
rect 31500 23772 31668 23774
rect 31164 23492 31444 23548
rect 30940 23380 30996 23390
rect 30940 23286 30996 23324
rect 31164 23378 31220 23492
rect 31164 23326 31166 23378
rect 31218 23326 31220 23378
rect 31164 23314 31220 23326
rect 31052 23268 31108 23278
rect 31052 23174 31108 23212
rect 31388 21924 31444 23492
rect 31500 23268 31556 23772
rect 31612 23762 31668 23772
rect 32732 23604 32788 23614
rect 32060 23492 32116 23502
rect 31724 23268 31780 23278
rect 31500 23202 31556 23212
rect 31612 23266 31780 23268
rect 31612 23214 31726 23266
rect 31778 23214 31780 23266
rect 31612 23212 31780 23214
rect 31612 23154 31668 23212
rect 31724 23202 31780 23212
rect 31948 23268 32004 23278
rect 31948 23174 32004 23212
rect 32060 23268 32116 23436
rect 32060 23266 32228 23268
rect 32060 23214 32062 23266
rect 32114 23214 32228 23266
rect 32060 23212 32228 23214
rect 32060 23202 32116 23212
rect 31612 23102 31614 23154
rect 31666 23102 31668 23154
rect 31612 23090 31668 23102
rect 32060 22482 32116 22494
rect 32060 22430 32062 22482
rect 32114 22430 32116 22482
rect 32060 22372 32116 22430
rect 32060 22306 32116 22316
rect 32172 22148 32228 23212
rect 32508 22596 32564 22606
rect 32564 22540 32676 22596
rect 32508 22530 32564 22540
rect 32284 22372 32340 22382
rect 32340 22316 32564 22372
rect 32284 22306 32340 22316
rect 30884 21756 30996 21812
rect 30828 21718 30884 21756
rect 30492 21588 30548 21598
rect 30492 21494 30548 21532
rect 30828 21588 30884 21598
rect 30716 20692 30772 20702
rect 30828 20692 30884 21532
rect 30940 20804 30996 21756
rect 31388 21810 31444 21868
rect 31388 21758 31390 21810
rect 31442 21758 31444 21810
rect 31388 21746 31444 21758
rect 32060 22092 32228 22148
rect 32060 21698 32116 22092
rect 32060 21646 32062 21698
rect 32114 21646 32116 21698
rect 30940 20738 30996 20748
rect 31164 21586 31220 21598
rect 31164 21534 31166 21586
rect 31218 21534 31220 21586
rect 30716 20690 30884 20692
rect 30716 20638 30718 20690
rect 30770 20638 30884 20690
rect 30716 20636 30884 20638
rect 30716 20626 30772 20636
rect 31052 20580 31108 20590
rect 31052 20486 31108 20524
rect 30380 20178 30436 20188
rect 30156 20132 30212 20142
rect 30156 20038 30212 20076
rect 30044 20018 30100 20030
rect 30044 19966 30046 20018
rect 30098 19966 30100 20018
rect 29596 19292 29988 19348
rect 29484 19236 29540 19246
rect 29596 19236 29652 19292
rect 29484 19234 29652 19236
rect 29484 19182 29486 19234
rect 29538 19182 29652 19234
rect 29484 19180 29652 19182
rect 29932 19234 29988 19292
rect 29932 19182 29934 19234
rect 29986 19182 29988 19234
rect 29484 19170 29540 19180
rect 29932 19170 29988 19182
rect 29708 19122 29764 19134
rect 29708 19070 29710 19122
rect 29762 19070 29764 19122
rect 29708 19012 29764 19070
rect 29708 18946 29764 18956
rect 29820 19124 29876 19134
rect 29036 18610 29092 18620
rect 29148 18620 29428 18676
rect 29484 18900 29540 18910
rect 28476 18562 28980 18564
rect 28476 18510 28478 18562
rect 28530 18510 28980 18562
rect 28476 18508 28980 18510
rect 28476 18498 28532 18508
rect 28364 18284 28644 18340
rect 28252 18172 28532 18228
rect 26908 17276 27748 17332
rect 26908 16994 26964 17276
rect 26908 16942 26910 16994
rect 26962 16942 26964 16994
rect 26908 16930 26964 16942
rect 26796 16830 26798 16882
rect 26850 16830 26852 16882
rect 26796 16818 26852 16830
rect 26236 16706 26292 16716
rect 26124 16660 26180 16670
rect 25900 16658 26180 16660
rect 25900 16606 26126 16658
rect 26178 16606 26180 16658
rect 25900 16604 26180 16606
rect 25900 16210 25956 16604
rect 26124 16594 26180 16604
rect 25900 16158 25902 16210
rect 25954 16158 25956 16210
rect 25900 16146 25956 16158
rect 27916 16436 27972 16446
rect 27916 16212 27972 16380
rect 27916 16210 28308 16212
rect 27916 16158 27918 16210
rect 27970 16158 28308 16210
rect 27916 16156 28308 16158
rect 27916 16146 27972 16156
rect 25676 16098 25732 16110
rect 25676 16046 25678 16098
rect 25730 16046 25732 16098
rect 25676 15764 25732 16046
rect 28252 16098 28308 16156
rect 28252 16046 28254 16098
rect 28306 16046 28308 16098
rect 28252 16034 28308 16046
rect 25676 15698 25732 15708
rect 26012 15986 26068 15998
rect 26012 15934 26014 15986
rect 26066 15934 26068 15986
rect 26012 15428 26068 15934
rect 27916 15876 27972 15886
rect 27916 15538 27972 15820
rect 27916 15486 27918 15538
rect 27970 15486 27972 15538
rect 27916 15474 27972 15486
rect 26012 15362 26068 15372
rect 26684 15428 26740 15438
rect 26124 15316 26180 15326
rect 26124 15222 26180 15260
rect 26572 15314 26628 15326
rect 26572 15262 26574 15314
rect 26626 15262 26628 15314
rect 25564 14690 25620 14700
rect 26012 15204 26068 15214
rect 26572 15148 26628 15262
rect 25004 14532 25060 14542
rect 25340 14532 25396 14542
rect 24668 14530 25172 14532
rect 24668 14478 25006 14530
rect 25058 14478 25172 14530
rect 24668 14476 25172 14478
rect 24556 14466 24612 14476
rect 25004 14466 25060 14476
rect 24556 14308 24612 14318
rect 24556 14214 24612 14252
rect 24668 14306 24724 14318
rect 24668 14254 24670 14306
rect 24722 14254 24724 14306
rect 24444 14028 24612 14084
rect 23548 13970 23604 14028
rect 23548 13918 23550 13970
rect 23602 13918 23604 13970
rect 23548 13906 23604 13918
rect 24444 13860 24500 13898
rect 24220 13804 24444 13860
rect 23772 13748 23828 13758
rect 23436 13692 23604 13748
rect 23324 13636 23380 13646
rect 23100 13234 23156 13244
rect 23212 13580 23324 13636
rect 23212 12740 23268 13580
rect 23324 13570 23380 13580
rect 23548 13076 23604 13692
rect 23772 13654 23828 13692
rect 23996 13746 24052 13758
rect 23996 13694 23998 13746
rect 24050 13694 24052 13746
rect 23660 13636 23716 13646
rect 23660 13542 23716 13580
rect 23996 13636 24052 13694
rect 23996 13570 24052 13580
rect 23548 13010 23604 13020
rect 23996 13300 24052 13310
rect 22988 12684 23268 12740
rect 22988 12290 23044 12684
rect 23996 12402 24052 13244
rect 23996 12350 23998 12402
rect 24050 12350 24052 12402
rect 23996 12338 24052 12350
rect 24220 12404 24276 13804
rect 24444 13794 24500 13804
rect 24444 13634 24500 13646
rect 24444 13582 24446 13634
rect 24498 13582 24500 13634
rect 24332 13076 24388 13086
rect 24332 12982 24388 13020
rect 22988 12238 22990 12290
rect 23042 12238 23044 12290
rect 22988 12226 23044 12238
rect 23436 12292 23492 12302
rect 23436 12198 23492 12236
rect 24220 12290 24276 12348
rect 24220 12238 24222 12290
rect 24274 12238 24276 12290
rect 24220 12226 24276 12238
rect 24108 12066 24164 12078
rect 24108 12014 24110 12066
rect 24162 12014 24164 12066
rect 24108 11506 24164 12014
rect 24108 11454 24110 11506
rect 24162 11454 24164 11506
rect 24108 11442 24164 11454
rect 23324 11394 23380 11406
rect 23324 11342 23326 11394
rect 23378 11342 23380 11394
rect 22988 11172 23044 11182
rect 23324 11172 23380 11342
rect 22988 11170 23380 11172
rect 22988 11118 22990 11170
rect 23042 11118 23380 11170
rect 22988 11116 23380 11118
rect 22988 10500 23044 11116
rect 23324 10500 23380 10510
rect 22988 10434 23044 10444
rect 23100 10498 23380 10500
rect 23100 10446 23326 10498
rect 23378 10446 23380 10498
rect 23100 10444 23380 10446
rect 23100 10276 23156 10444
rect 23324 10434 23380 10444
rect 22876 10220 23156 10276
rect 23212 10276 23268 10286
rect 23212 9938 23268 10220
rect 24444 10276 24500 13582
rect 24556 13188 24612 14028
rect 24668 13858 24724 14254
rect 24780 14306 24836 14318
rect 24780 14254 24782 14306
rect 24834 14254 24836 14306
rect 24780 14196 24836 14254
rect 24780 14130 24836 14140
rect 24668 13806 24670 13858
rect 24722 13806 24724 13858
rect 24668 13794 24724 13806
rect 25004 13860 25060 13870
rect 24780 13188 24836 13198
rect 24556 13186 24836 13188
rect 24556 13134 24782 13186
rect 24834 13134 24836 13186
rect 24556 13132 24836 13134
rect 24780 13122 24836 13132
rect 25004 12850 25060 13804
rect 25004 12798 25006 12850
rect 25058 12798 25060 12850
rect 25004 12786 25060 12798
rect 25116 13636 25172 14476
rect 25340 13970 25396 14476
rect 26012 14530 26068 15148
rect 26348 15092 26628 15148
rect 26684 15202 26740 15372
rect 27692 15428 27748 15438
rect 27580 15316 27636 15326
rect 27580 15222 27636 15260
rect 26684 15150 26686 15202
rect 26738 15150 26740 15202
rect 26236 14644 26292 14654
rect 26236 14550 26292 14588
rect 26012 14478 26014 14530
rect 26066 14478 26068 14530
rect 26012 14466 26068 14478
rect 25340 13918 25342 13970
rect 25394 13918 25396 13970
rect 25340 13906 25396 13918
rect 25676 14418 25732 14430
rect 25676 14366 25678 14418
rect 25730 14366 25732 14418
rect 24892 12738 24948 12750
rect 24892 12686 24894 12738
rect 24946 12686 24948 12738
rect 24892 10724 24948 12686
rect 25116 11060 25172 13580
rect 25676 12964 25732 14366
rect 25788 14306 25844 14318
rect 25788 14254 25790 14306
rect 25842 14254 25844 14306
rect 25788 14196 25844 14254
rect 26348 14306 26404 15092
rect 26572 14756 26628 14766
rect 26684 14756 26740 15150
rect 27692 15148 27748 15372
rect 27692 15092 27972 15148
rect 26572 14754 26740 14756
rect 26572 14702 26574 14754
rect 26626 14702 26740 14754
rect 26572 14700 26740 14702
rect 26572 14690 26628 14700
rect 27244 14420 27300 14430
rect 26348 14254 26350 14306
rect 26402 14254 26404 14306
rect 26124 14196 26180 14206
rect 25788 14140 26124 14196
rect 26124 13970 26180 14140
rect 26124 13918 26126 13970
rect 26178 13918 26180 13970
rect 26124 13906 26180 13918
rect 26348 13412 26404 14254
rect 27020 14306 27076 14318
rect 27020 14254 27022 14306
rect 27074 14254 27076 14306
rect 27020 13858 27076 14254
rect 27244 14196 27300 14364
rect 27356 14308 27412 14318
rect 27356 14214 27412 14252
rect 27468 14306 27524 14318
rect 27468 14254 27470 14306
rect 27522 14254 27524 14306
rect 27244 14130 27300 14140
rect 27468 14196 27524 14254
rect 27468 14130 27524 14140
rect 27916 13972 27972 15092
rect 28476 14644 28532 18172
rect 28588 17778 28644 18284
rect 28588 17726 28590 17778
rect 28642 17726 28644 17778
rect 28588 17714 28644 17726
rect 28924 16996 28980 17006
rect 28700 16212 28756 16222
rect 28588 15988 28644 15998
rect 28588 15894 28644 15932
rect 28476 14578 28532 14588
rect 28588 14644 28644 14654
rect 28700 14644 28756 16156
rect 28924 16100 28980 16940
rect 29148 16212 29204 18620
rect 29484 17106 29540 18844
rect 29596 18676 29652 18686
rect 29596 17666 29652 18620
rect 29708 18676 29764 18686
rect 29820 18676 29876 19068
rect 29708 18674 29876 18676
rect 29708 18622 29710 18674
rect 29762 18622 29876 18674
rect 29708 18620 29876 18622
rect 29708 18610 29764 18620
rect 29932 18564 29988 18602
rect 30044 18564 30100 19966
rect 30380 20020 30436 20030
rect 30380 20018 30772 20020
rect 30380 19966 30382 20018
rect 30434 19966 30772 20018
rect 30380 19964 30772 19966
rect 30380 19954 30436 19964
rect 30604 19794 30660 19806
rect 30604 19742 30606 19794
rect 30658 19742 30660 19794
rect 30156 19348 30212 19358
rect 30156 19254 30212 19292
rect 30268 19236 30324 19246
rect 30268 19142 30324 19180
rect 30604 19122 30660 19742
rect 30716 19236 30772 19964
rect 30828 19906 30884 19918
rect 30828 19854 30830 19906
rect 30882 19854 30884 19906
rect 30828 19794 30884 19854
rect 30828 19742 30830 19794
rect 30882 19742 30884 19794
rect 30828 19730 30884 19742
rect 30828 19236 30884 19246
rect 30716 19234 30884 19236
rect 30716 19182 30830 19234
rect 30882 19182 30884 19234
rect 30716 19180 30884 19182
rect 30828 19170 30884 19180
rect 30604 19070 30606 19122
rect 30658 19070 30660 19122
rect 30604 19012 30660 19070
rect 30604 18946 30660 18956
rect 30940 19012 30996 19050
rect 30940 18946 30996 18956
rect 31164 18900 31220 21534
rect 31836 21586 31892 21598
rect 31836 21534 31838 21586
rect 31890 21534 31892 21586
rect 31276 21474 31332 21486
rect 31276 21422 31278 21474
rect 31330 21422 31332 21474
rect 31276 20916 31332 21422
rect 31836 21364 31892 21534
rect 32060 21588 32116 21646
rect 32172 21700 32228 21710
rect 32172 21698 32452 21700
rect 32172 21646 32174 21698
rect 32226 21646 32452 21698
rect 32172 21644 32452 21646
rect 32172 21634 32228 21644
rect 32060 21522 32116 21532
rect 32172 21364 32228 21374
rect 31836 21362 32228 21364
rect 31836 21310 32174 21362
rect 32226 21310 32228 21362
rect 31836 21308 32228 21310
rect 32172 21298 32228 21308
rect 31276 20850 31332 20860
rect 32172 20916 32228 20926
rect 32172 20822 32228 20860
rect 31500 20804 31556 20814
rect 31500 20710 31556 20748
rect 31948 20692 32004 20702
rect 31948 20242 32004 20636
rect 31948 20190 31950 20242
rect 32002 20190 32004 20242
rect 31948 20178 32004 20190
rect 32396 20244 32452 21644
rect 32284 20132 32340 20142
rect 31612 20020 31668 20030
rect 31836 20020 31892 20030
rect 31388 20018 31668 20020
rect 31388 19966 31614 20018
rect 31666 19966 31668 20018
rect 31388 19964 31668 19966
rect 31276 19348 31332 19358
rect 31276 19234 31332 19292
rect 31276 19182 31278 19234
rect 31330 19182 31332 19234
rect 31276 19170 31332 19182
rect 31164 18834 31220 18844
rect 31276 19012 31332 19022
rect 30940 18788 30996 18798
rect 30380 18676 30436 18686
rect 30380 18582 30436 18620
rect 29988 18508 30100 18564
rect 29932 18498 29988 18508
rect 29820 18452 29876 18462
rect 29596 17614 29598 17666
rect 29650 17614 29652 17666
rect 29596 17602 29652 17614
rect 29708 18396 29820 18452
rect 29708 17668 29764 18396
rect 29820 18386 29876 18396
rect 29820 17668 29876 17678
rect 29708 17666 29876 17668
rect 29708 17614 29822 17666
rect 29874 17614 29876 17666
rect 29708 17612 29876 17614
rect 29820 17602 29876 17612
rect 30044 17666 30100 18508
rect 30156 18564 30212 18574
rect 30156 18470 30212 18508
rect 30604 18450 30660 18462
rect 30604 18398 30606 18450
rect 30658 18398 30660 18450
rect 30268 18338 30324 18350
rect 30268 18286 30270 18338
rect 30322 18286 30324 18338
rect 30044 17614 30046 17666
rect 30098 17614 30100 17666
rect 30044 17602 30100 17614
rect 30156 17780 30212 17790
rect 30156 17666 30212 17724
rect 30156 17614 30158 17666
rect 30210 17614 30212 17666
rect 30156 17602 30212 17614
rect 29932 17442 29988 17454
rect 29932 17390 29934 17442
rect 29986 17390 29988 17442
rect 29932 17108 29988 17390
rect 30268 17444 30324 18286
rect 30604 18340 30660 18398
rect 30604 18284 30884 18340
rect 30828 17780 30884 18284
rect 30940 18004 30996 18732
rect 31276 18788 31332 18956
rect 31276 18674 31332 18732
rect 31276 18622 31278 18674
rect 31330 18622 31332 18674
rect 31276 18610 31332 18622
rect 31164 18564 31220 18574
rect 31164 18470 31220 18508
rect 30940 17938 30996 17948
rect 31276 17892 31332 17902
rect 31276 17780 31332 17836
rect 30884 17778 31332 17780
rect 30884 17726 31278 17778
rect 31330 17726 31332 17778
rect 30884 17724 31332 17726
rect 30828 17686 30884 17724
rect 31276 17714 31332 17724
rect 31388 17668 31444 19964
rect 31612 19954 31668 19964
rect 31724 20018 31892 20020
rect 31724 19966 31838 20018
rect 31890 19966 31892 20018
rect 31724 19964 31892 19966
rect 31724 19124 31780 19964
rect 31836 19954 31892 19964
rect 32172 20018 32228 20030
rect 32172 19966 32174 20018
rect 32226 19966 32228 20018
rect 31500 19068 31780 19124
rect 31836 19460 31892 19470
rect 31836 19234 31892 19404
rect 32172 19346 32228 19966
rect 32172 19294 32174 19346
rect 32226 19294 32228 19346
rect 32172 19282 32228 19294
rect 31836 19182 31838 19234
rect 31890 19182 31892 19234
rect 31500 18450 31556 19068
rect 31836 19012 31892 19182
rect 32284 19234 32340 20076
rect 32284 19182 32286 19234
rect 32338 19182 32340 19234
rect 32284 19124 32340 19182
rect 32396 19234 32452 20188
rect 32396 19182 32398 19234
rect 32450 19182 32452 19234
rect 32396 19170 32452 19182
rect 32060 19012 32116 19022
rect 31724 18956 31892 19012
rect 31948 18956 32060 19012
rect 31500 18398 31502 18450
rect 31554 18398 31556 18450
rect 31500 18386 31556 18398
rect 31612 18788 31668 18798
rect 31500 17668 31556 17678
rect 31388 17612 31500 17668
rect 31500 17602 31556 17612
rect 31612 17444 31668 18732
rect 31724 18340 31780 18956
rect 31836 18788 31892 18798
rect 31836 18450 31892 18732
rect 31948 18674 32004 18956
rect 32060 18918 32116 18956
rect 31948 18622 31950 18674
rect 32002 18622 32004 18674
rect 31948 18610 32004 18622
rect 32172 18676 32228 18686
rect 32284 18676 32340 19068
rect 32172 18674 32340 18676
rect 32172 18622 32174 18674
rect 32226 18622 32340 18674
rect 32172 18620 32340 18622
rect 32508 18676 32564 22316
rect 32172 18610 32228 18620
rect 31836 18398 31838 18450
rect 31890 18398 31892 18450
rect 31836 18386 31892 18398
rect 32396 18452 32452 18462
rect 32508 18452 32564 18620
rect 32396 18450 32564 18452
rect 32396 18398 32398 18450
rect 32450 18398 32564 18450
rect 32396 18396 32564 18398
rect 32396 18386 32452 18396
rect 31724 18274 31780 18284
rect 32284 18338 32340 18350
rect 32284 18286 32286 18338
rect 32338 18286 32340 18338
rect 31836 18004 31892 18014
rect 31892 17948 32004 18004
rect 31836 17938 31892 17948
rect 31836 17668 31892 17678
rect 31836 17574 31892 17612
rect 30268 17388 30548 17444
rect 29484 17054 29486 17106
rect 29538 17054 29540 17106
rect 29484 17042 29540 17054
rect 29596 17052 29988 17108
rect 29260 16996 29316 17006
rect 29260 16902 29316 16940
rect 29484 16884 29540 16894
rect 29484 16790 29540 16828
rect 29260 16212 29316 16222
rect 29148 16210 29316 16212
rect 29148 16158 29262 16210
rect 29314 16158 29316 16210
rect 29148 16156 29316 16158
rect 29260 16146 29316 16156
rect 29036 16100 29092 16110
rect 28924 16098 29092 16100
rect 28924 16046 29038 16098
rect 29090 16046 29092 16098
rect 28924 16044 29092 16046
rect 28812 15540 28868 15550
rect 29036 15540 29092 16044
rect 28812 15538 29092 15540
rect 28812 15486 28814 15538
rect 28866 15486 29092 15538
rect 28812 15484 29092 15486
rect 28812 15474 28868 15484
rect 28588 14642 28756 14644
rect 28588 14590 28590 14642
rect 28642 14590 28756 14642
rect 28588 14588 28756 14590
rect 28588 14578 28644 14588
rect 28700 14532 28756 14588
rect 28700 14466 28756 14476
rect 27020 13806 27022 13858
rect 27074 13806 27076 13858
rect 27020 13794 27076 13806
rect 27468 13970 27972 13972
rect 27468 13918 27918 13970
rect 27970 13918 27972 13970
rect 27468 13916 27972 13918
rect 26908 13746 26964 13758
rect 26908 13694 26910 13746
rect 26962 13694 26964 13746
rect 26684 13524 26740 13534
rect 26684 13522 26852 13524
rect 26684 13470 26686 13522
rect 26738 13470 26852 13522
rect 26684 13468 26852 13470
rect 26684 13458 26740 13468
rect 26236 12964 26292 12974
rect 25676 12908 26236 12964
rect 26124 12738 26180 12750
rect 26124 12686 26126 12738
rect 26178 12686 26180 12738
rect 26124 12180 26180 12686
rect 26124 12114 26180 12124
rect 25116 10994 25172 11004
rect 25340 12068 25396 12078
rect 24892 10658 24948 10668
rect 25228 10610 25284 10622
rect 25228 10558 25230 10610
rect 25282 10558 25284 10610
rect 24668 10500 24724 10510
rect 24668 10406 24724 10444
rect 25228 10500 25284 10558
rect 25228 10434 25284 10444
rect 24444 10210 24500 10220
rect 23212 9886 23214 9938
rect 23266 9886 23268 9938
rect 23212 9874 23268 9886
rect 25340 9938 25396 12012
rect 26236 11506 26292 12908
rect 26348 12852 26404 13356
rect 26796 12962 26852 13468
rect 26796 12910 26798 12962
rect 26850 12910 26852 12962
rect 26460 12852 26516 12862
rect 26348 12850 26516 12852
rect 26348 12798 26462 12850
rect 26514 12798 26516 12850
rect 26348 12796 26516 12798
rect 26460 12786 26516 12796
rect 26796 12404 26852 12910
rect 26796 12338 26852 12348
rect 26908 13188 26964 13694
rect 27468 13746 27524 13916
rect 27916 13906 27972 13916
rect 28028 14420 28084 14430
rect 28028 14306 28084 14364
rect 28028 14254 28030 14306
rect 28082 14254 28084 14306
rect 27468 13694 27470 13746
rect 27522 13694 27524 13746
rect 27468 13682 27524 13694
rect 28028 13636 28084 14254
rect 28028 13570 28084 13580
rect 28476 13636 28532 13646
rect 28476 13542 28532 13580
rect 28924 13636 28980 13646
rect 28924 13542 28980 13580
rect 27244 13522 27300 13534
rect 27244 13470 27246 13522
rect 27298 13470 27300 13522
rect 27244 13412 27300 13470
rect 27020 13188 27076 13198
rect 26908 13186 27076 13188
rect 26908 13134 27022 13186
rect 27074 13134 27076 13186
rect 26908 13132 27076 13134
rect 26908 13076 26964 13132
rect 27020 13122 27076 13132
rect 27244 13186 27300 13356
rect 27244 13134 27246 13186
rect 27298 13134 27300 13186
rect 27244 13122 27300 13134
rect 28252 13522 28308 13534
rect 28252 13470 28254 13522
rect 28306 13470 28308 13522
rect 26684 12180 26740 12190
rect 26908 12180 26964 13020
rect 27468 12964 27524 12974
rect 27468 12870 27524 12908
rect 28252 12964 28308 13470
rect 28700 13076 28756 13086
rect 28700 12982 28756 13020
rect 27916 12740 27972 12750
rect 27692 12738 27972 12740
rect 27692 12686 27918 12738
rect 27970 12686 27972 12738
rect 27692 12684 27972 12686
rect 26684 12178 26964 12180
rect 26684 12126 26686 12178
rect 26738 12126 26964 12178
rect 26684 12124 26964 12126
rect 27244 12404 27300 12414
rect 27244 12290 27300 12348
rect 27244 12238 27246 12290
rect 27298 12238 27300 12290
rect 26684 12114 26740 12124
rect 27244 12068 27300 12238
rect 27244 12002 27300 12012
rect 26236 11454 26238 11506
rect 26290 11454 26292 11506
rect 26236 11442 26292 11454
rect 26012 10724 26068 10734
rect 26012 10630 26068 10668
rect 27468 10276 27524 10286
rect 25340 9886 25342 9938
rect 25394 9886 25396 9938
rect 25340 9874 25396 9886
rect 25676 9940 25732 9950
rect 25676 9846 25732 9884
rect 22428 9774 22430 9826
rect 22482 9774 22484 9826
rect 21420 9538 21476 9548
rect 22092 9604 22148 9614
rect 22428 9604 22484 9774
rect 22148 9548 22484 9604
rect 26236 9716 26292 9726
rect 20300 8318 20302 8370
rect 20354 8318 20356 8370
rect 20300 8306 20356 8318
rect 21196 9044 21252 9054
rect 20860 8036 20916 8046
rect 19964 7980 20244 8036
rect 18396 7588 18452 7644
rect 19068 7588 19124 7598
rect 18396 7532 18564 7588
rect 17500 7310 17502 7362
rect 17554 7310 17556 7362
rect 17500 7298 17556 7310
rect 17948 7474 18004 7486
rect 17948 7422 17950 7474
rect 18002 7422 18004 7474
rect 17948 7364 18004 7422
rect 18396 7364 18452 7374
rect 17948 7298 18004 7308
rect 18060 7362 18452 7364
rect 18060 7310 18398 7362
rect 18450 7310 18452 7362
rect 18060 7308 18452 7310
rect 16716 5854 16718 5906
rect 16770 5854 16772 5906
rect 16604 5796 16660 5806
rect 16604 4338 16660 5740
rect 16604 4286 16606 4338
rect 16658 4286 16660 4338
rect 16604 4274 16660 4286
rect 16268 4174 16270 4226
rect 16322 4174 16324 4226
rect 16268 4162 16324 4174
rect 16716 4228 16772 5854
rect 17052 6690 17108 6702
rect 17052 6638 17054 6690
rect 17106 6638 17108 6690
rect 16940 5684 16996 5694
rect 16940 5234 16996 5628
rect 16940 5182 16942 5234
rect 16994 5182 16996 5234
rect 16940 5170 16996 5182
rect 17052 5236 17108 6638
rect 17724 6578 17780 6590
rect 17724 6526 17726 6578
rect 17778 6526 17780 6578
rect 17724 6468 17780 6526
rect 17724 6402 17780 6412
rect 18060 6244 18116 7308
rect 18396 7298 18452 7308
rect 18508 7140 18564 7532
rect 19068 7494 19124 7532
rect 17052 5170 17108 5180
rect 17164 6188 18116 6244
rect 18172 7084 18564 7140
rect 18956 7364 19012 7374
rect 16716 4162 16772 4172
rect 16156 3666 16212 3678
rect 16156 3614 16158 3666
rect 16210 3614 16212 3666
rect 14700 2828 14868 2884
rect 14812 800 14868 2828
rect 16156 800 16212 3614
rect 17052 3556 17108 3566
rect 17164 3556 17220 6188
rect 17500 6020 17556 6030
rect 17500 5926 17556 5964
rect 17612 5908 17668 5918
rect 17948 5908 18004 5918
rect 17612 5906 18004 5908
rect 17612 5854 17614 5906
rect 17666 5854 17950 5906
rect 18002 5854 18004 5906
rect 17612 5852 18004 5854
rect 17612 5842 17668 5852
rect 17948 5842 18004 5852
rect 18060 5794 18116 5806
rect 18060 5742 18062 5794
rect 18114 5742 18116 5794
rect 17500 5682 17556 5694
rect 17500 5630 17502 5682
rect 17554 5630 17556 5682
rect 17500 4338 17556 5630
rect 18060 5572 18116 5742
rect 17500 4286 17502 4338
rect 17554 4286 17556 4338
rect 17500 4274 17556 4286
rect 17612 5516 18116 5572
rect 17612 4116 17668 5516
rect 17052 3554 17220 3556
rect 17052 3502 17054 3554
rect 17106 3502 17220 3554
rect 17052 3500 17220 3502
rect 17276 4060 17668 4116
rect 17724 5348 17780 5358
rect 17052 3388 17108 3500
rect 16828 3332 17108 3388
rect 17276 3442 17332 4060
rect 17276 3390 17278 3442
rect 17330 3390 17332 3442
rect 17276 3378 17332 3390
rect 17500 3668 17556 3678
rect 16828 800 16884 3332
rect 17500 800 17556 3612
rect 17724 3554 17780 5292
rect 17836 5124 17892 5134
rect 17836 4450 17892 5068
rect 18060 5124 18116 5134
rect 17948 4564 18004 4574
rect 17948 4470 18004 4508
rect 18060 4562 18116 5068
rect 18060 4510 18062 4562
rect 18114 4510 18116 4562
rect 18060 4498 18116 4510
rect 17836 4398 17838 4450
rect 17890 4398 17892 4450
rect 17836 4386 17892 4398
rect 18172 4338 18228 7084
rect 18508 5794 18564 5806
rect 18508 5742 18510 5794
rect 18562 5742 18564 5794
rect 18396 5684 18452 5694
rect 18396 5590 18452 5628
rect 18508 5124 18564 5742
rect 18956 5348 19012 7308
rect 19068 5908 19124 5918
rect 19180 5908 19236 7980
rect 19836 7868 20100 7878
rect 19404 7812 19460 7822
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 19836 7802 20100 7812
rect 19404 7698 19460 7756
rect 19404 7646 19406 7698
rect 19458 7646 19460 7698
rect 19404 7634 19460 7646
rect 20076 7700 20132 7710
rect 20188 7700 20244 7980
rect 20860 8034 21028 8036
rect 20860 7982 20862 8034
rect 20914 7982 21028 8034
rect 20860 7980 21028 7982
rect 20860 7970 20916 7980
rect 20076 7698 20244 7700
rect 20076 7646 20078 7698
rect 20130 7646 20244 7698
rect 20076 7644 20244 7646
rect 20076 7634 20132 7644
rect 19740 7588 19796 7598
rect 19740 7494 19796 7532
rect 20188 7362 20244 7374
rect 20188 7310 20190 7362
rect 20242 7310 20244 7362
rect 20188 7028 20244 7310
rect 19852 6972 20244 7028
rect 20860 7250 20916 7262
rect 20860 7198 20862 7250
rect 20914 7198 20916 7250
rect 19852 6802 19908 6972
rect 19852 6750 19854 6802
rect 19906 6750 19908 6802
rect 19852 6738 19908 6750
rect 20300 6468 20356 6478
rect 20300 6466 20468 6468
rect 20300 6414 20302 6466
rect 20354 6414 20468 6466
rect 20300 6412 20468 6414
rect 20300 6402 20356 6412
rect 19836 6300 20100 6310
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 19836 6234 20100 6244
rect 19292 6020 19348 6030
rect 19292 6018 19572 6020
rect 19292 5966 19294 6018
rect 19346 5966 19572 6018
rect 19292 5964 19572 5966
rect 19292 5954 19348 5964
rect 19068 5906 19236 5908
rect 19068 5854 19070 5906
rect 19122 5854 19236 5906
rect 19068 5852 19236 5854
rect 19068 5842 19124 5852
rect 19180 5796 19236 5852
rect 19180 5740 19460 5796
rect 19068 5348 19124 5358
rect 18956 5292 19068 5348
rect 18508 5058 18564 5068
rect 18732 5236 18788 5246
rect 18172 4286 18174 4338
rect 18226 4286 18228 4338
rect 18172 4274 18228 4286
rect 18732 4338 18788 5180
rect 19068 5234 19124 5292
rect 19068 5182 19070 5234
rect 19122 5182 19124 5234
rect 19068 5170 19124 5182
rect 18732 4286 18734 4338
rect 18786 4286 18788 4338
rect 18732 4274 18788 4286
rect 18844 5124 18900 5134
rect 18620 3668 18676 3678
rect 18620 3574 18676 3612
rect 17724 3502 17726 3554
rect 17778 3502 17780 3554
rect 17724 3490 17780 3502
rect 18844 800 18900 5068
rect 19404 5010 19460 5740
rect 19516 5684 19572 5964
rect 20076 6018 20132 6030
rect 20076 5966 20078 6018
rect 20130 5966 20132 6018
rect 19852 5908 19908 5918
rect 19852 5814 19908 5852
rect 19516 5618 19572 5628
rect 20076 5460 20132 5966
rect 20076 5404 20244 5460
rect 20188 5348 20244 5404
rect 20188 5292 20356 5348
rect 20076 5236 20132 5246
rect 19404 4958 19406 5010
rect 19458 4958 19460 5010
rect 19404 4946 19460 4958
rect 19516 5234 20132 5236
rect 19516 5182 20078 5234
rect 20130 5182 20132 5234
rect 19516 5180 20132 5182
rect 19404 4452 19460 4462
rect 19516 4452 19572 5180
rect 20076 5170 20132 5180
rect 20188 5122 20244 5134
rect 20188 5070 20190 5122
rect 20242 5070 20244 5122
rect 19740 5012 19796 5022
rect 19740 4918 19796 4956
rect 19836 4732 20100 4742
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 19836 4666 20100 4676
rect 20188 4564 20244 5070
rect 20188 4498 20244 4508
rect 19404 4450 19572 4452
rect 19404 4398 19406 4450
rect 19458 4398 19572 4450
rect 19404 4396 19572 4398
rect 19404 4386 19460 4396
rect 20300 3556 20356 5292
rect 20412 5124 20468 6412
rect 20748 6466 20804 6478
rect 20748 6414 20750 6466
rect 20802 6414 20804 6466
rect 20524 5908 20580 5918
rect 20524 5814 20580 5852
rect 20748 5796 20804 6414
rect 20860 5906 20916 7198
rect 20860 5854 20862 5906
rect 20914 5854 20916 5906
rect 20860 5842 20916 5854
rect 20748 5236 20804 5740
rect 20748 5142 20804 5180
rect 20972 5236 21028 7980
rect 21196 7474 21252 8988
rect 21644 9044 21700 9054
rect 21532 8484 21588 8494
rect 21420 7588 21476 7598
rect 21420 7494 21476 7532
rect 21196 7422 21198 7474
rect 21250 7422 21252 7474
rect 21196 7410 21252 7422
rect 21420 6468 21476 6478
rect 21532 6468 21588 8428
rect 21644 8146 21700 8988
rect 22092 8484 22148 9548
rect 22540 8932 22596 8942
rect 22092 8418 22148 8428
rect 22204 8930 22596 8932
rect 22204 8878 22542 8930
rect 22594 8878 22596 8930
rect 22204 8876 22596 8878
rect 21980 8260 22036 8270
rect 21980 8166 22036 8204
rect 21644 8094 21646 8146
rect 21698 8094 21700 8146
rect 21644 8082 21700 8094
rect 22204 7700 22260 8876
rect 22540 8866 22596 8876
rect 22988 8930 23044 8942
rect 22988 8878 22990 8930
rect 23042 8878 23044 8930
rect 22428 8484 22484 8494
rect 22428 8372 22484 8428
rect 22988 8372 23044 8878
rect 26236 8930 26292 9660
rect 26236 8878 26238 8930
rect 26290 8878 26292 8930
rect 26236 8866 26292 8878
rect 27468 8596 27524 10220
rect 27692 10052 27748 12684
rect 27916 12674 27972 12684
rect 28252 12516 28308 12908
rect 28252 12450 28308 12460
rect 28252 12180 28308 12190
rect 28700 12180 28756 12190
rect 28308 12178 28756 12180
rect 28308 12126 28702 12178
rect 28754 12126 28756 12178
rect 28308 12124 28756 12126
rect 28140 11508 28196 11518
rect 28140 11414 28196 11452
rect 28028 10612 28084 10622
rect 27916 10556 28028 10612
rect 27692 9986 27748 9996
rect 27804 10500 27860 10510
rect 27804 9938 27860 10444
rect 27804 9886 27806 9938
rect 27858 9886 27860 9938
rect 27804 9874 27860 9886
rect 27580 9604 27636 9614
rect 27580 9154 27636 9548
rect 27580 9102 27582 9154
rect 27634 9102 27636 9154
rect 27580 9090 27636 9102
rect 27916 8820 27972 10556
rect 28028 10546 28084 10556
rect 28140 10500 28196 10510
rect 28252 10500 28308 12124
rect 28700 12114 28756 12124
rect 29036 11508 29092 15484
rect 29484 15986 29540 15998
rect 29484 15934 29486 15986
rect 29538 15934 29540 15986
rect 29484 15148 29540 15934
rect 29596 15876 29652 17052
rect 30268 16994 30324 17006
rect 30268 16942 30270 16994
rect 30322 16942 30324 16994
rect 29820 16882 29876 16894
rect 29820 16830 29822 16882
rect 29874 16830 29876 16882
rect 29820 16772 29876 16830
rect 30156 16772 30212 16782
rect 29820 16770 30212 16772
rect 29820 16718 30158 16770
rect 30210 16718 30212 16770
rect 29820 16716 30212 16718
rect 30156 16706 30212 16716
rect 30156 16212 30212 16222
rect 29708 16210 30212 16212
rect 29708 16158 30158 16210
rect 30210 16158 30212 16210
rect 29708 16156 30212 16158
rect 29708 16098 29764 16156
rect 30156 16146 30212 16156
rect 29708 16046 29710 16098
rect 29762 16046 29764 16098
rect 29708 16034 29764 16046
rect 30044 15986 30100 15998
rect 30044 15934 30046 15986
rect 30098 15934 30100 15986
rect 30044 15876 30100 15934
rect 29596 15820 30100 15876
rect 30268 15988 30324 16942
rect 30492 16994 30548 17388
rect 31388 17388 31668 17444
rect 31388 17106 31444 17388
rect 31388 17054 31390 17106
rect 31442 17054 31444 17106
rect 31388 17042 31444 17054
rect 31500 17220 31556 17230
rect 30492 16942 30494 16994
rect 30546 16942 30548 16994
rect 30492 16930 30548 16942
rect 31500 16994 31556 17164
rect 31500 16942 31502 16994
rect 31554 16942 31556 16994
rect 31500 16930 31556 16942
rect 31724 17106 31780 17118
rect 31724 17054 31726 17106
rect 31778 17054 31780 17106
rect 31724 16996 31780 17054
rect 31724 16930 31780 16940
rect 31836 17108 31892 17118
rect 31612 16770 31668 16782
rect 31836 16772 31892 17052
rect 31612 16718 31614 16770
rect 31666 16718 31668 16770
rect 31612 16212 31668 16718
rect 29372 15092 29540 15148
rect 29820 15202 29876 15214
rect 29820 15150 29822 15202
rect 29874 15150 29876 15202
rect 29260 13860 29316 13870
rect 29260 13766 29316 13804
rect 29372 13748 29428 15092
rect 29484 14532 29540 14542
rect 29484 14438 29540 14476
rect 29820 14532 29876 15150
rect 30268 15148 30324 15932
rect 31500 16156 31668 16212
rect 31724 16716 31892 16772
rect 31948 16994 32004 17948
rect 32284 17892 32340 18286
rect 32284 17836 32564 17892
rect 32172 17666 32228 17678
rect 32172 17614 32174 17666
rect 32226 17614 32228 17666
rect 31948 16942 31950 16994
rect 32002 16942 32004 16994
rect 31164 15876 31220 15886
rect 31164 15782 31220 15820
rect 30044 15092 30324 15148
rect 31500 15148 31556 16156
rect 31724 16098 31780 16716
rect 31948 16548 32004 16942
rect 31724 16046 31726 16098
rect 31778 16046 31780 16098
rect 31724 16034 31780 16046
rect 31836 16492 32004 16548
rect 32060 17444 32116 17454
rect 32060 17220 32116 17388
rect 32172 17220 32228 17614
rect 32284 17668 32340 17678
rect 32284 17574 32340 17612
rect 32508 17666 32564 17836
rect 32508 17614 32510 17666
rect 32562 17614 32564 17666
rect 32508 17602 32564 17614
rect 32620 17668 32676 22540
rect 32732 22484 32788 23548
rect 33740 23268 33796 23998
rect 35084 23380 35140 24444
rect 35196 24332 35460 24342
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35196 24266 35460 24276
rect 35532 23716 35588 24780
rect 35644 24722 35700 24734
rect 35644 24670 35646 24722
rect 35698 24670 35700 24722
rect 35644 23940 35700 24670
rect 36316 24052 36372 24062
rect 35980 23940 36036 23950
rect 35644 23884 35924 23940
rect 35308 23660 35532 23716
rect 35196 23380 35252 23390
rect 35084 23378 35252 23380
rect 35084 23326 35198 23378
rect 35250 23326 35252 23378
rect 35084 23324 35252 23326
rect 35196 23314 35252 23324
rect 32732 22482 33124 22484
rect 32732 22430 32734 22482
rect 32786 22430 33124 22482
rect 32732 22428 33124 22430
rect 32732 22418 32788 22428
rect 33068 21586 33124 22428
rect 33068 21534 33070 21586
rect 33122 21534 33124 21586
rect 33068 20244 33124 21534
rect 33180 20244 33236 20254
rect 33068 20242 33236 20244
rect 33068 20190 33182 20242
rect 33234 20190 33236 20242
rect 33068 20188 33236 20190
rect 33180 19460 33236 20188
rect 33180 19394 33236 19404
rect 33292 20244 33348 20254
rect 33180 19236 33236 19246
rect 33180 19142 33236 19180
rect 33292 19234 33348 20188
rect 33740 20132 33796 23212
rect 35308 23156 35364 23660
rect 35532 23622 35588 23660
rect 35644 23714 35700 23726
rect 35644 23662 35646 23714
rect 35698 23662 35700 23714
rect 35084 23100 35364 23156
rect 35532 23156 35588 23166
rect 35644 23156 35700 23662
rect 35588 23100 35700 23156
rect 35084 22596 35140 23100
rect 35532 23062 35588 23100
rect 35196 22764 35460 22774
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35196 22698 35460 22708
rect 35196 22596 35252 22606
rect 35084 22594 35252 22596
rect 35084 22542 35198 22594
rect 35250 22542 35252 22594
rect 35084 22540 35252 22542
rect 35196 22530 35252 22540
rect 34076 22372 34132 22382
rect 34076 22370 34804 22372
rect 34076 22318 34078 22370
rect 34130 22318 34804 22370
rect 34076 22316 34804 22318
rect 34076 22306 34132 22316
rect 34300 22148 34356 22158
rect 34300 22146 34468 22148
rect 34300 22094 34302 22146
rect 34354 22094 34468 22146
rect 34300 22092 34468 22094
rect 34300 22082 34356 22092
rect 34300 20914 34356 20926
rect 34300 20862 34302 20914
rect 34354 20862 34356 20914
rect 34300 20244 34356 20862
rect 34412 20468 34468 22092
rect 34412 20402 34468 20412
rect 34636 21364 34692 21374
rect 34636 20804 34692 21308
rect 34748 21026 34804 22316
rect 35644 22260 35700 23100
rect 35868 23604 35924 23884
rect 35980 23826 36036 23884
rect 35980 23774 35982 23826
rect 36034 23774 36036 23826
rect 35980 23762 36036 23774
rect 35756 22260 35812 22270
rect 35644 22258 35812 22260
rect 35644 22206 35758 22258
rect 35810 22206 35812 22258
rect 35644 22204 35812 22206
rect 35756 22194 35812 22204
rect 34860 22148 34916 22158
rect 34860 22146 35140 22148
rect 34860 22094 34862 22146
rect 34914 22094 35140 22146
rect 34860 22092 35140 22094
rect 34860 22082 34916 22092
rect 34748 20974 34750 21026
rect 34802 20974 34804 21026
rect 34748 20962 34804 20974
rect 35084 21026 35140 22092
rect 35196 21474 35252 21486
rect 35196 21422 35198 21474
rect 35250 21422 35252 21474
rect 35196 21364 35252 21422
rect 35196 21298 35252 21308
rect 35196 21196 35460 21206
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35196 21130 35460 21140
rect 35084 20974 35086 21026
rect 35138 20974 35140 21026
rect 35084 20962 35140 20974
rect 34356 20188 34468 20244
rect 34300 20178 34356 20188
rect 33740 20076 34132 20132
rect 33964 19348 34020 19358
rect 33964 19254 34020 19292
rect 33292 19182 33294 19234
rect 33346 19182 33348 19234
rect 33292 19170 33348 19182
rect 33516 19236 33572 19246
rect 33852 19236 33908 19246
rect 33516 19234 33908 19236
rect 33516 19182 33518 19234
rect 33570 19182 33854 19234
rect 33906 19182 33908 19234
rect 33516 19180 33908 19182
rect 32844 19122 32900 19134
rect 32844 19070 32846 19122
rect 32898 19070 32900 19122
rect 32844 18676 32900 19070
rect 33068 19010 33124 19022
rect 33068 18958 33070 19010
rect 33122 18958 33124 19010
rect 33068 18788 33124 18958
rect 33068 18722 33124 18732
rect 33516 19012 33572 19180
rect 33852 19170 33908 19180
rect 34076 19012 34132 20076
rect 34412 19234 34468 20188
rect 34636 20018 34692 20748
rect 35756 20916 35812 20926
rect 35756 20690 35812 20860
rect 35868 20802 35924 23548
rect 36316 23266 36372 23996
rect 36316 23214 36318 23266
rect 36370 23214 36372 23266
rect 36316 23202 36372 23214
rect 36428 23828 36484 37100
rect 37100 36932 37156 36942
rect 37100 36482 37156 36876
rect 37100 36430 37102 36482
rect 37154 36430 37156 36482
rect 37100 36418 37156 36430
rect 37660 35924 37716 37212
rect 37772 36594 37828 37326
rect 37772 36542 37774 36594
rect 37826 36542 37828 36594
rect 37772 36530 37828 36542
rect 38220 36596 38276 37886
rect 38780 36708 38836 40348
rect 39004 39732 39060 39742
rect 39004 39620 39060 39676
rect 39116 39620 39172 39630
rect 39004 39618 39172 39620
rect 39004 39566 39118 39618
rect 39170 39566 39172 39618
rect 39004 39564 39172 39566
rect 39004 38668 39060 39564
rect 39116 39554 39172 39564
rect 39340 38946 39396 40572
rect 39564 40290 39620 40796
rect 39676 40740 39732 41134
rect 39676 40674 39732 40684
rect 39788 41076 39844 41086
rect 39788 40404 39844 41020
rect 39788 40338 39844 40348
rect 39564 40238 39566 40290
rect 39618 40238 39620 40290
rect 39564 40226 39620 40238
rect 40012 40290 40068 40302
rect 40012 40238 40014 40290
rect 40066 40238 40068 40290
rect 39900 39508 39956 39518
rect 39900 39414 39956 39452
rect 39340 38894 39342 38946
rect 39394 38894 39396 38946
rect 39340 38882 39396 38894
rect 39564 39060 39620 39070
rect 39564 38946 39620 39004
rect 40012 39060 40068 40238
rect 40124 39732 40180 41804
rect 40796 41412 40852 44268
rect 41020 44258 41076 44268
rect 40908 43652 40964 43662
rect 40908 43558 40964 43596
rect 41020 41860 41076 41870
rect 41132 41860 41188 44940
rect 41580 44930 41636 44940
rect 42028 44546 42084 45164
rect 42588 45218 42644 45612
rect 42700 45602 42756 45612
rect 42588 45166 42590 45218
rect 42642 45166 42644 45218
rect 42588 45154 42644 45166
rect 42028 44494 42030 44546
rect 42082 44494 42084 44546
rect 42028 44482 42084 44494
rect 42028 43988 42084 43998
rect 41244 43540 41300 43550
rect 41244 43446 41300 43484
rect 41804 43428 41860 43438
rect 41804 43426 41972 43428
rect 41804 43374 41806 43426
rect 41858 43374 41972 43426
rect 41804 43372 41972 43374
rect 41804 43362 41860 43372
rect 41076 41804 41188 41860
rect 41580 41858 41636 41870
rect 41580 41806 41582 41858
rect 41634 41806 41636 41858
rect 41020 41766 41076 41804
rect 40684 41356 40852 41412
rect 40124 39666 40180 39676
rect 40236 40404 40292 40414
rect 40012 38994 40068 39004
rect 40236 39058 40292 40348
rect 40236 39006 40238 39058
rect 40290 39006 40292 39058
rect 40236 38994 40292 39006
rect 40348 39060 40404 39070
rect 39564 38894 39566 38946
rect 39618 38894 39620 38946
rect 39564 38882 39620 38894
rect 39900 38836 39956 38846
rect 39900 38742 39956 38780
rect 38892 38612 39060 38668
rect 38892 38164 38948 38612
rect 38892 38162 39284 38164
rect 38892 38110 38894 38162
rect 38946 38110 39284 38162
rect 38892 38108 39284 38110
rect 38892 38098 38948 38108
rect 39228 38052 39284 38108
rect 39228 38050 39508 38052
rect 39228 37998 39230 38050
rect 39282 37998 39508 38050
rect 39228 37996 39508 37998
rect 39228 37986 39284 37996
rect 39452 37492 39508 37996
rect 40012 37940 40068 37950
rect 40012 37938 40292 37940
rect 40012 37886 40014 37938
rect 40066 37886 40292 37938
rect 40012 37884 40292 37886
rect 40012 37874 40068 37884
rect 39900 37492 39956 37502
rect 39452 37490 39900 37492
rect 39452 37438 39454 37490
rect 39506 37438 39900 37490
rect 39452 37436 39900 37438
rect 39956 37436 40180 37492
rect 39452 36932 39508 37436
rect 39900 37398 39956 37436
rect 39452 36866 39508 36876
rect 38780 36652 39172 36708
rect 37884 35924 37940 35934
rect 37660 35922 37940 35924
rect 37660 35870 37886 35922
rect 37938 35870 37940 35922
rect 37660 35868 37940 35870
rect 37884 35858 37940 35868
rect 38220 35698 38276 36540
rect 39004 36484 39060 36494
rect 38220 35646 38222 35698
rect 38274 35646 38276 35698
rect 38220 35634 38276 35646
rect 38780 35810 38836 35822
rect 38780 35758 38782 35810
rect 38834 35758 38836 35810
rect 37548 34914 37604 34926
rect 37548 34862 37550 34914
rect 37602 34862 37604 34914
rect 37100 34692 37156 34702
rect 37548 34692 37604 34862
rect 37100 34690 37604 34692
rect 37100 34638 37102 34690
rect 37154 34638 37604 34690
rect 37100 34636 37604 34638
rect 37100 34626 37156 34636
rect 36876 34132 36932 34142
rect 37436 34132 37492 34142
rect 36876 34130 37492 34132
rect 36876 34078 36878 34130
rect 36930 34078 37438 34130
rect 37490 34078 37492 34130
rect 36876 34076 37492 34078
rect 36876 34066 36932 34076
rect 37100 33908 37156 33918
rect 36988 32674 37044 32686
rect 36988 32622 36990 32674
rect 37042 32622 37044 32674
rect 36988 31948 37044 32622
rect 36652 31892 37044 31948
rect 37100 31948 37156 33852
rect 37436 33684 37492 34076
rect 37436 33618 37492 33628
rect 37548 33346 37604 34636
rect 37772 34692 37828 34702
rect 37772 33460 37828 34636
rect 37772 33394 37828 33404
rect 38108 34018 38164 34030
rect 38108 33966 38110 34018
rect 38162 33966 38164 34018
rect 37548 33294 37550 33346
rect 37602 33294 37604 33346
rect 37212 33124 37268 33134
rect 37548 33124 37604 33294
rect 37268 33068 37604 33124
rect 38108 33124 38164 33966
rect 38780 33236 38836 35758
rect 39004 35698 39060 36428
rect 39004 35646 39006 35698
rect 39058 35646 39060 35698
rect 39004 35634 39060 35646
rect 38780 33170 38836 33180
rect 37212 33030 37268 33068
rect 38108 33058 38164 33068
rect 38668 32674 38724 32686
rect 38668 32622 38670 32674
rect 38722 32622 38724 32674
rect 37324 32564 37380 32574
rect 37324 32562 37716 32564
rect 37324 32510 37326 32562
rect 37378 32510 37716 32562
rect 37324 32508 37716 32510
rect 37324 32498 37380 32508
rect 37660 32002 37716 32508
rect 37660 31950 37662 32002
rect 37714 31950 37716 32002
rect 37100 31892 37492 31948
rect 37660 31938 37716 31950
rect 38444 32562 38500 32574
rect 38444 32510 38446 32562
rect 38498 32510 38500 32562
rect 36652 31106 36708 31892
rect 36652 31054 36654 31106
rect 36706 31054 36708 31106
rect 36652 31042 36708 31054
rect 37212 31554 37268 31566
rect 37212 31502 37214 31554
rect 37266 31502 37268 31554
rect 37100 30210 37156 30222
rect 37100 30158 37102 30210
rect 37154 30158 37156 30210
rect 37100 29316 37156 30158
rect 37212 30212 37268 31502
rect 37212 29540 37268 30156
rect 37212 29474 37268 29484
rect 37324 29428 37380 29438
rect 37324 29316 37380 29372
rect 37100 29260 37380 29316
rect 36540 28532 36596 28542
rect 36540 27746 36596 28476
rect 37324 27860 37380 29260
rect 37436 29204 37492 31892
rect 37996 31778 38052 31790
rect 37996 31726 37998 31778
rect 38050 31726 38052 31778
rect 37996 30884 38052 31726
rect 37996 30818 38052 30828
rect 38220 31666 38276 31678
rect 38220 31614 38222 31666
rect 38274 31614 38276 31666
rect 38220 30212 38276 31614
rect 38444 31220 38500 32510
rect 38668 31892 38724 32622
rect 39116 32674 39172 36652
rect 39900 36596 39956 36606
rect 39900 36502 39956 36540
rect 40124 35924 40180 37436
rect 40236 36372 40292 37884
rect 40348 37492 40404 39004
rect 40684 38724 40740 41356
rect 40796 41188 40852 41198
rect 41468 41188 41524 41198
rect 40796 41186 41524 41188
rect 40796 41134 40798 41186
rect 40850 41134 41470 41186
rect 41522 41134 41524 41186
rect 40796 41132 41524 41134
rect 41580 41188 41636 41806
rect 41804 41188 41860 41198
rect 41580 41186 41860 41188
rect 41580 41134 41806 41186
rect 41858 41134 41860 41186
rect 41580 41132 41860 41134
rect 40796 41122 40852 41132
rect 41468 41122 41524 41132
rect 41020 40964 41076 40974
rect 41020 40870 41076 40908
rect 41804 40628 41860 41132
rect 41804 40562 41860 40572
rect 41692 40516 41748 40526
rect 41692 40422 41748 40460
rect 41020 40180 41076 40190
rect 41020 40178 41188 40180
rect 41020 40126 41022 40178
rect 41074 40126 41188 40178
rect 41020 40124 41188 40126
rect 41020 40114 41076 40124
rect 40908 39508 40964 39518
rect 40908 39058 40964 39452
rect 40908 39006 40910 39058
rect 40962 39006 40964 39058
rect 40908 38994 40964 39006
rect 41132 38834 41188 40124
rect 41356 40178 41412 40190
rect 41356 40126 41358 40178
rect 41410 40126 41412 40178
rect 41356 40068 41412 40126
rect 41804 40180 41860 40190
rect 41916 40180 41972 43372
rect 42028 42754 42084 43932
rect 42028 42702 42030 42754
rect 42082 42702 42084 42754
rect 42028 42690 42084 42702
rect 42028 41074 42084 41086
rect 42028 41022 42030 41074
rect 42082 41022 42084 41074
rect 42028 40852 42084 41022
rect 42364 41076 42420 41086
rect 42364 40982 42420 41020
rect 42028 40786 42084 40796
rect 42700 40852 42756 40862
rect 42028 40516 42084 40526
rect 42028 40514 42196 40516
rect 42028 40462 42030 40514
rect 42082 40462 42196 40514
rect 42028 40460 42196 40462
rect 42028 40450 42084 40460
rect 41860 40124 41972 40180
rect 41804 40114 41860 40124
rect 41356 40002 41412 40012
rect 42028 40068 42084 40078
rect 42028 39730 42084 40012
rect 42028 39678 42030 39730
rect 42082 39678 42084 39730
rect 42028 39666 42084 39678
rect 42140 39508 42196 40460
rect 42700 40402 42756 40796
rect 42700 40350 42702 40402
rect 42754 40350 42756 40402
rect 42700 40338 42756 40350
rect 42812 39844 42868 45836
rect 42924 45826 42980 45836
rect 44044 45892 44100 45902
rect 44044 45890 44324 45892
rect 44044 45838 44046 45890
rect 44098 45838 44324 45890
rect 44044 45836 44324 45838
rect 44044 45826 44100 45836
rect 43260 44436 43316 44446
rect 42924 43540 42980 43550
rect 42924 42978 42980 43484
rect 42924 42926 42926 42978
rect 42978 42926 42980 42978
rect 42924 42914 42980 42926
rect 43260 42978 43316 44380
rect 44156 44324 44212 44334
rect 44044 44322 44212 44324
rect 44044 44270 44158 44322
rect 44210 44270 44212 44322
rect 44044 44268 44212 44270
rect 43932 44098 43988 44110
rect 43932 44046 43934 44098
rect 43986 44046 43988 44098
rect 43932 43650 43988 44046
rect 43932 43598 43934 43650
rect 43986 43598 43988 43650
rect 43932 43586 43988 43598
rect 43260 42926 43262 42978
rect 43314 42926 43316 42978
rect 43260 42914 43316 42926
rect 43708 42754 43764 42766
rect 43708 42702 43710 42754
rect 43762 42702 43764 42754
rect 42812 39778 42868 39788
rect 42924 42644 42980 42654
rect 42924 40514 42980 42588
rect 43708 42084 43764 42702
rect 43820 42644 43876 42654
rect 43820 42550 43876 42588
rect 44044 42196 44100 44268
rect 44156 44258 44212 44268
rect 43596 42028 43764 42084
rect 43820 42140 44100 42196
rect 43596 41972 43652 42028
rect 43596 41906 43652 41916
rect 43708 41858 43764 41870
rect 43708 41806 43710 41858
rect 43762 41806 43764 41858
rect 43148 41076 43204 41086
rect 42924 40462 42926 40514
rect 42978 40462 42980 40514
rect 42028 39452 42196 39508
rect 41692 39060 41748 39070
rect 41692 38966 41748 39004
rect 41132 38782 41134 38834
rect 41186 38782 41188 38834
rect 41132 38770 41188 38782
rect 40684 38658 40740 38668
rect 42028 38164 42084 39452
rect 42476 39394 42532 39406
rect 42476 39342 42478 39394
rect 42530 39342 42532 39394
rect 42476 38834 42532 39342
rect 42476 38782 42478 38834
rect 42530 38782 42532 38834
rect 42140 38722 42196 38734
rect 42140 38670 42142 38722
rect 42194 38670 42196 38722
rect 42140 38668 42196 38670
rect 42476 38668 42532 38782
rect 42924 38668 42980 40462
rect 43036 41074 43204 41076
rect 43036 41022 43150 41074
rect 43202 41022 43204 41074
rect 43036 41020 43204 41022
rect 43036 39842 43092 41020
rect 43148 41010 43204 41020
rect 43484 40964 43540 40974
rect 43036 39790 43038 39842
rect 43090 39790 43092 39842
rect 43036 39778 43092 39790
rect 43260 40962 43540 40964
rect 43260 40910 43486 40962
rect 43538 40910 43540 40962
rect 43260 40908 43540 40910
rect 43260 38946 43316 40908
rect 43484 40898 43540 40908
rect 43708 40964 43764 41806
rect 43708 40898 43764 40908
rect 43820 40626 43876 42140
rect 43932 41860 43988 41870
rect 43932 41298 43988 41804
rect 44268 41748 44324 45836
rect 44380 45332 44436 49200
rect 45276 46452 45332 46462
rect 45164 46396 45276 46452
rect 45052 45780 45108 45790
rect 44940 45724 45052 45780
rect 44380 45266 44436 45276
rect 44604 45666 44660 45678
rect 44604 45614 44606 45666
rect 44658 45614 44660 45666
rect 44604 45108 44660 45614
rect 44604 45042 44660 45052
rect 44716 44996 44772 45006
rect 44716 43876 44772 44940
rect 44940 44772 44996 45724
rect 45052 45714 45108 45724
rect 45052 45106 45108 45118
rect 45052 45054 45054 45106
rect 45106 45054 45108 45106
rect 45052 44996 45108 45054
rect 45052 44930 45108 44940
rect 44940 44716 45108 44772
rect 44940 44548 44996 44558
rect 44940 44454 44996 44492
rect 44716 43810 44772 43820
rect 44604 43538 44660 43550
rect 44604 43486 44606 43538
rect 44658 43486 44660 43538
rect 44492 41970 44548 41982
rect 44492 41918 44494 41970
rect 44546 41918 44548 41970
rect 44492 41860 44548 41918
rect 44604 41860 44660 43486
rect 45052 43540 45108 44716
rect 45164 43764 45220 46396
rect 45276 46386 45332 46396
rect 46844 45666 46900 45678
rect 46844 45614 46846 45666
rect 46898 45614 46900 45666
rect 46060 45332 46116 45342
rect 46060 45238 46116 45276
rect 46844 45108 46900 45614
rect 46844 45042 46900 45052
rect 47740 45666 47796 45678
rect 47740 45614 47742 45666
rect 47794 45614 47796 45666
rect 45836 44436 45892 44446
rect 45276 44322 45332 44334
rect 45276 44270 45278 44322
rect 45330 44270 45332 44322
rect 45276 43988 45332 44270
rect 45276 43922 45332 43932
rect 45724 44322 45780 44334
rect 45724 44270 45726 44322
rect 45778 44270 45780 44322
rect 45276 43764 45332 43774
rect 45164 43762 45332 43764
rect 45164 43710 45278 43762
rect 45330 43710 45332 43762
rect 45164 43708 45332 43710
rect 45276 43698 45332 43708
rect 45052 43484 45332 43540
rect 45276 42642 45332 43484
rect 45276 42590 45278 42642
rect 45330 42590 45332 42642
rect 45276 42578 45332 42590
rect 45052 42196 45108 42206
rect 44828 41970 44884 41982
rect 44828 41918 44830 41970
rect 44882 41918 44884 41970
rect 44828 41860 44884 41918
rect 44548 41804 44884 41860
rect 44492 41794 44548 41804
rect 44268 41682 44324 41692
rect 43932 41246 43934 41298
rect 43986 41246 43988 41298
rect 43932 41234 43988 41246
rect 43820 40574 43822 40626
rect 43874 40574 43876 40626
rect 43820 40562 43876 40574
rect 44156 41188 44212 41198
rect 44156 40516 44212 41132
rect 44604 40626 44660 41804
rect 44604 40574 44606 40626
rect 44658 40574 44660 40626
rect 44604 40562 44660 40574
rect 44940 41074 44996 41086
rect 44940 41022 44942 41074
rect 44994 41022 44996 41074
rect 43484 40180 43540 40190
rect 43484 40086 43540 40124
rect 43372 39844 43428 39854
rect 43372 39750 43428 39788
rect 44156 39618 44212 40460
rect 44940 40404 44996 41022
rect 44940 40338 44996 40348
rect 45052 40402 45108 42140
rect 45612 41860 45668 41870
rect 45276 41858 45668 41860
rect 45276 41806 45614 41858
rect 45666 41806 45668 41858
rect 45276 41804 45668 41806
rect 45276 41074 45332 41804
rect 45612 41794 45668 41804
rect 45612 41188 45668 41198
rect 45276 41022 45278 41074
rect 45330 41022 45332 41074
rect 45276 41010 45332 41022
rect 45500 41186 45668 41188
rect 45500 41134 45614 41186
rect 45666 41134 45668 41186
rect 45500 41132 45668 41134
rect 45052 40350 45054 40402
rect 45106 40350 45108 40402
rect 45052 40338 45108 40350
rect 45276 40514 45332 40526
rect 45276 40462 45278 40514
rect 45330 40462 45332 40514
rect 45276 39732 45332 40462
rect 45276 39666 45332 39676
rect 45500 39844 45556 41132
rect 45612 41122 45668 41132
rect 45724 41188 45780 44270
rect 45836 44210 45892 44380
rect 47740 44436 47796 45614
rect 48188 45668 48244 45678
rect 48188 45666 48356 45668
rect 48188 45614 48190 45666
rect 48242 45614 48356 45666
rect 48188 45612 48356 45614
rect 48188 45602 48244 45612
rect 47740 44370 47796 44380
rect 48188 45218 48244 45230
rect 48188 45166 48190 45218
rect 48242 45166 48244 45218
rect 45836 44158 45838 44210
rect 45890 44158 45892 44210
rect 45836 44146 45892 44158
rect 47180 44322 47236 44334
rect 47180 44270 47182 44322
rect 47234 44270 47236 44322
rect 46844 44098 46900 44110
rect 46844 44046 46846 44098
rect 46898 44046 46900 44098
rect 45724 41122 45780 41132
rect 45836 43538 45892 43550
rect 45836 43486 45838 43538
rect 45890 43486 45892 43538
rect 45836 41860 45892 43486
rect 46844 42196 46900 44046
rect 46844 42130 46900 42140
rect 46956 42866 47012 42878
rect 46956 42814 46958 42866
rect 47010 42814 47012 42866
rect 45612 40402 45668 40414
rect 45612 40350 45614 40402
rect 45666 40350 45668 40402
rect 45612 40068 45668 40350
rect 45612 40002 45668 40012
rect 44156 39566 44158 39618
rect 44210 39566 44212 39618
rect 44156 39554 44212 39566
rect 45388 39618 45444 39630
rect 45388 39566 45390 39618
rect 45442 39566 45444 39618
rect 43260 38894 43262 38946
rect 43314 38894 43316 38946
rect 43260 38882 43316 38894
rect 43932 39506 43988 39518
rect 43932 39454 43934 39506
rect 43986 39454 43988 39506
rect 42140 38612 42644 38668
rect 42140 38164 42196 38174
rect 41804 38162 42196 38164
rect 41804 38110 42142 38162
rect 42194 38110 42196 38162
rect 41804 38108 42196 38110
rect 41692 37940 41748 37950
rect 41468 37828 41524 37838
rect 41020 37492 41076 37502
rect 40348 37490 40628 37492
rect 40348 37438 40350 37490
rect 40402 37438 40628 37490
rect 40348 37436 40628 37438
rect 40348 37426 40404 37436
rect 40348 36372 40404 36382
rect 40236 36370 40404 36372
rect 40236 36318 40350 36370
rect 40402 36318 40404 36370
rect 40236 36316 40404 36318
rect 40348 36306 40404 36316
rect 40572 36148 40628 37436
rect 41020 37398 41076 37436
rect 41468 37266 41524 37772
rect 41692 37490 41748 37884
rect 41692 37438 41694 37490
rect 41746 37438 41748 37490
rect 41692 37426 41748 37438
rect 41468 37214 41470 37266
rect 41522 37214 41524 37266
rect 41468 37202 41524 37214
rect 41692 36708 41748 36718
rect 41804 36708 41860 38108
rect 42140 38098 42196 38108
rect 42140 37492 42196 37502
rect 42252 37492 42308 38612
rect 42588 38162 42644 38612
rect 42588 38110 42590 38162
rect 42642 38110 42644 38162
rect 42588 38098 42644 38110
rect 42812 38612 42980 38668
rect 42196 37436 42308 37492
rect 42140 37426 42196 37436
rect 42028 37156 42084 37166
rect 42028 37062 42084 37100
rect 41692 36706 41860 36708
rect 41692 36654 41694 36706
rect 41746 36654 41860 36706
rect 41692 36652 41860 36654
rect 41692 36642 41748 36652
rect 42476 36484 42532 36494
rect 42476 36390 42532 36428
rect 40684 36372 40740 36382
rect 41356 36372 41412 36382
rect 40684 36370 41412 36372
rect 40684 36318 40686 36370
rect 40738 36318 41358 36370
rect 41410 36318 41412 36370
rect 40684 36316 41412 36318
rect 40684 36306 40740 36316
rect 41356 36306 41412 36316
rect 42252 36370 42308 36382
rect 42252 36318 42254 36370
rect 42306 36318 42308 36370
rect 40572 36092 41300 36148
rect 40124 35830 40180 35868
rect 41244 35922 41300 36092
rect 41244 35870 41246 35922
rect 41298 35870 41300 35922
rect 40236 35812 40292 35822
rect 39788 35364 39844 35374
rect 39788 35026 39844 35308
rect 39788 34974 39790 35026
rect 39842 34974 39844 35026
rect 39788 34962 39844 34974
rect 40236 34020 40292 35756
rect 41244 35474 41300 35870
rect 41692 35924 41748 35934
rect 41692 35830 41748 35868
rect 41244 35422 41246 35474
rect 41298 35422 41300 35474
rect 41244 35410 41300 35422
rect 41804 35474 41860 35486
rect 41804 35422 41806 35474
rect 41858 35422 41860 35474
rect 41356 35028 41412 35038
rect 41132 34916 41188 34926
rect 41132 34822 41188 34860
rect 40908 34692 40964 34702
rect 40908 34598 40964 34636
rect 41356 34580 41412 34972
rect 41804 35026 41860 35422
rect 41804 34974 41806 35026
rect 41858 34974 41860 35026
rect 41804 34962 41860 34974
rect 42252 35028 42308 36318
rect 42812 36260 42868 38612
rect 43148 38164 43204 38174
rect 43036 37828 43092 37838
rect 43036 37734 43092 37772
rect 43148 37604 43204 38108
rect 43372 38052 43428 38062
rect 43372 37958 43428 37996
rect 42252 34962 42308 34972
rect 42476 36204 42868 36260
rect 43036 37548 43204 37604
rect 43708 37938 43764 37950
rect 43708 37886 43710 37938
rect 43762 37886 43764 37938
rect 43036 36370 43092 37548
rect 43148 36484 43204 36494
rect 43148 36390 43204 36428
rect 43036 36318 43038 36370
rect 43090 36318 43092 36370
rect 42252 34804 42308 34814
rect 41468 34692 41524 34702
rect 41468 34690 41748 34692
rect 41468 34638 41470 34690
rect 41522 34638 41748 34690
rect 41468 34636 41748 34638
rect 41468 34626 41524 34636
rect 39900 34018 40292 34020
rect 39900 33966 40238 34018
rect 40290 33966 40292 34018
rect 39900 33964 40292 33966
rect 39116 32622 39118 32674
rect 39170 32622 39172 32674
rect 39116 31948 39172 32622
rect 39340 33684 39396 33694
rect 39340 33234 39396 33628
rect 39340 33182 39342 33234
rect 39394 33182 39396 33234
rect 39340 32116 39396 33182
rect 38668 31826 38724 31836
rect 38780 31892 39284 31948
rect 38780 31666 38836 31892
rect 38780 31614 38782 31666
rect 38834 31614 38836 31666
rect 38780 31602 38836 31614
rect 39228 31444 39284 31892
rect 39340 31778 39396 32060
rect 39676 32674 39732 32686
rect 39676 32622 39678 32674
rect 39730 32622 39732 32674
rect 39676 32004 39732 32622
rect 39900 32562 39956 33964
rect 40236 33954 40292 33964
rect 40908 34130 40964 34142
rect 40908 34078 40910 34130
rect 40962 34078 40964 34130
rect 40908 33684 40964 34078
rect 40908 33618 40964 33628
rect 40684 33348 40740 33358
rect 40236 33346 40740 33348
rect 40236 33294 40686 33346
rect 40738 33294 40740 33346
rect 40236 33292 40740 33294
rect 40236 32786 40292 33292
rect 40684 33282 40740 33292
rect 40460 33124 40516 33134
rect 40460 33030 40516 33068
rect 40236 32734 40238 32786
rect 40290 32734 40292 32786
rect 40236 32722 40292 32734
rect 41356 32674 41412 34524
rect 41692 34242 41748 34636
rect 41692 34190 41694 34242
rect 41746 34190 41748 34242
rect 41692 34178 41748 34190
rect 41692 33346 41748 33358
rect 41692 33294 41694 33346
rect 41746 33294 41748 33346
rect 41356 32622 41358 32674
rect 41410 32622 41412 32674
rect 41356 32610 41412 32622
rect 41580 32676 41636 32686
rect 41580 32582 41636 32620
rect 39900 32510 39902 32562
rect 39954 32510 39956 32562
rect 39900 32498 39956 32510
rect 40124 32564 40180 32574
rect 39676 31938 39732 31948
rect 39788 31892 39844 31902
rect 40012 31892 40068 31902
rect 39844 31890 40068 31892
rect 39844 31838 40014 31890
rect 40066 31838 40068 31890
rect 39844 31836 40068 31838
rect 39788 31826 39844 31836
rect 40012 31826 40068 31836
rect 39340 31726 39342 31778
rect 39394 31726 39396 31778
rect 39340 31714 39396 31726
rect 39228 31388 40068 31444
rect 38444 31154 38500 31164
rect 40012 31218 40068 31388
rect 40012 31166 40014 31218
rect 40066 31166 40068 31218
rect 40012 31154 40068 31166
rect 38780 30884 38836 30894
rect 38220 30146 38276 30156
rect 38556 30828 38780 30884
rect 37772 30098 37828 30110
rect 37772 30046 37774 30098
rect 37826 30046 37828 30098
rect 37772 29650 37828 30046
rect 37772 29598 37774 29650
rect 37826 29598 37828 29650
rect 37772 29586 37828 29598
rect 37548 29428 37604 29438
rect 38220 29428 38276 29438
rect 37548 29426 38276 29428
rect 37548 29374 37550 29426
rect 37602 29374 38222 29426
rect 38274 29374 38276 29426
rect 37548 29372 38276 29374
rect 37548 29362 37604 29372
rect 38220 29362 38276 29372
rect 38556 29426 38612 30828
rect 38780 30790 38836 30828
rect 39900 30324 39956 30334
rect 40124 30324 40180 32508
rect 41020 32116 41076 32126
rect 39340 30322 40180 30324
rect 39340 30270 39902 30322
rect 39954 30270 40180 30322
rect 39340 30268 40180 30270
rect 40236 30994 40292 31006
rect 40236 30942 40238 30994
rect 40290 30942 40292 30994
rect 39340 29538 39396 30268
rect 39900 30258 39956 30268
rect 39340 29486 39342 29538
rect 39394 29486 39396 29538
rect 39340 29474 39396 29486
rect 38556 29374 38558 29426
rect 38610 29374 38612 29426
rect 38556 29362 38612 29374
rect 39116 29426 39172 29438
rect 39116 29374 39118 29426
rect 39170 29374 39172 29426
rect 37436 29148 37604 29204
rect 37548 28530 37604 29148
rect 38332 28980 38388 28990
rect 37548 28478 37550 28530
rect 37602 28478 37604 28530
rect 37548 28466 37604 28478
rect 37772 28642 37828 28654
rect 37772 28590 37774 28642
rect 37826 28590 37828 28642
rect 37436 27860 37492 27870
rect 37324 27858 37492 27860
rect 37324 27806 37438 27858
rect 37490 27806 37492 27858
rect 37324 27804 37492 27806
rect 37436 27794 37492 27804
rect 36540 27694 36542 27746
rect 36594 27694 36596 27746
rect 36540 27682 36596 27694
rect 37772 27300 37828 28590
rect 37548 27244 37828 27300
rect 38220 27746 38276 27758
rect 38220 27694 38222 27746
rect 38274 27694 38276 27746
rect 37548 26180 37604 27244
rect 37772 27076 37828 27086
rect 37772 26982 37828 27020
rect 38220 26516 38276 27694
rect 38332 27186 38388 28924
rect 39116 28980 39172 29374
rect 39116 28914 39172 28924
rect 39340 29316 39396 29326
rect 39340 28530 39396 29260
rect 39900 29314 39956 29326
rect 39900 29262 39902 29314
rect 39954 29262 39956 29314
rect 39900 28980 39956 29262
rect 39900 28914 39956 28924
rect 40236 28644 40292 30942
rect 40684 30212 40740 30222
rect 40684 28754 40740 30156
rect 41020 29428 41076 32060
rect 41692 31948 41748 33294
rect 42252 32786 42308 34748
rect 42364 34692 42420 34702
rect 42364 34598 42420 34636
rect 42252 32734 42254 32786
rect 42306 32734 42308 32786
rect 42252 32722 42308 32734
rect 41916 32340 41972 32350
rect 41916 32246 41972 32284
rect 42476 31948 42532 36204
rect 42812 34916 42868 34926
rect 42812 34822 42868 34860
rect 42700 32562 42756 32574
rect 42700 32510 42702 32562
rect 42754 32510 42756 32562
rect 42700 31948 42756 32510
rect 41468 31892 42196 31948
rect 41132 31220 41188 31230
rect 41132 31126 41188 31164
rect 41468 30994 41524 31892
rect 42140 31890 42196 31892
rect 42140 31838 42142 31890
rect 42194 31838 42196 31890
rect 42140 31826 42196 31838
rect 42252 31892 42532 31948
rect 42588 31892 42756 31948
rect 41692 31780 41748 31790
rect 41692 31106 41748 31724
rect 41692 31054 41694 31106
rect 41746 31054 41748 31106
rect 41692 31042 41748 31054
rect 42252 31106 42308 31892
rect 42588 31668 42644 31892
rect 42588 31602 42644 31612
rect 42700 31556 42756 31566
rect 43036 31556 43092 36318
rect 43596 35476 43652 35486
rect 43484 35474 43652 35476
rect 43484 35422 43598 35474
rect 43650 35422 43652 35474
rect 43484 35420 43652 35422
rect 43260 35252 43316 35262
rect 43148 34916 43204 34926
rect 43260 34916 43316 35196
rect 43484 35140 43540 35420
rect 43596 35410 43652 35420
rect 43708 35140 43764 37886
rect 43932 37156 43988 39454
rect 45052 39394 45108 39406
rect 45052 39342 45054 39394
rect 45106 39342 45108 39394
rect 44156 38164 44212 38174
rect 44156 37938 44212 38108
rect 44940 38164 44996 38174
rect 45052 38164 45108 39342
rect 45388 38836 45444 39566
rect 44996 38108 45108 38164
rect 45276 38780 45444 38836
rect 44940 38070 44996 38108
rect 44156 37886 44158 37938
rect 44210 37886 44212 37938
rect 44156 37874 44212 37886
rect 45276 38050 45332 38780
rect 45500 38724 45556 39788
rect 45836 38836 45892 41804
rect 46956 40404 47012 42814
rect 47180 42756 47236 44270
rect 47516 44210 47572 44222
rect 47516 44158 47518 44210
rect 47570 44158 47572 44210
rect 47404 42756 47460 42766
rect 47180 42700 47404 42756
rect 47404 42690 47460 42700
rect 46956 40338 47012 40348
rect 46060 39732 46116 39742
rect 46060 39638 46116 39676
rect 47516 39060 47572 44158
rect 47964 44212 48020 44222
rect 47964 44210 48132 44212
rect 47964 44158 47966 44210
rect 48018 44158 48132 44210
rect 47964 44156 48132 44158
rect 47964 44146 48020 44156
rect 47964 43314 48020 43326
rect 47964 43262 47966 43314
rect 48018 43262 48020 43314
rect 47740 41860 47796 41870
rect 47740 41766 47796 41804
rect 47964 41748 48020 43262
rect 47964 41682 48020 41692
rect 47852 41298 47908 41310
rect 47852 41246 47854 41298
rect 47906 41246 47908 41298
rect 47852 39732 47908 41246
rect 47852 39666 47908 39676
rect 47964 40178 48020 40190
rect 47964 40126 47966 40178
rect 48018 40126 48020 40178
rect 45836 38770 45892 38780
rect 45948 38946 46004 38958
rect 45948 38894 45950 38946
rect 46002 38894 46004 38946
rect 45388 38695 45556 38724
rect 45388 38643 45390 38695
rect 45442 38668 45556 38695
rect 45948 38668 46004 38894
rect 46284 38836 46340 38846
rect 46732 38836 46788 38846
rect 46284 38834 46788 38836
rect 46284 38782 46286 38834
rect 46338 38782 46734 38834
rect 46786 38782 46788 38834
rect 46284 38780 46788 38782
rect 46284 38770 46340 38780
rect 46732 38770 46788 38780
rect 47516 38834 47572 39004
rect 47964 39060 48020 40126
rect 47964 38994 48020 39004
rect 47516 38782 47518 38834
rect 47570 38782 47572 38834
rect 47516 38770 47572 38782
rect 47852 38946 47908 38958
rect 47852 38894 47854 38946
rect 47906 38894 47908 38946
rect 45442 38643 45444 38668
rect 45388 38631 45444 38643
rect 45276 37998 45278 38050
rect 45330 37998 45332 38050
rect 44940 37268 44996 37278
rect 45276 37268 45332 37998
rect 44996 37212 45332 37268
rect 45724 38612 46004 38668
rect 47068 38722 47124 38734
rect 47068 38670 47070 38722
rect 47122 38670 47124 38722
rect 43820 36708 43876 36718
rect 43932 36708 43988 37100
rect 44156 37156 44212 37166
rect 44156 37154 44884 37156
rect 44156 37102 44158 37154
rect 44210 37102 44884 37154
rect 44156 37100 44884 37102
rect 44156 37090 44212 37100
rect 43820 36706 43988 36708
rect 43820 36654 43822 36706
rect 43874 36654 43988 36706
rect 43820 36652 43988 36654
rect 43820 36642 43876 36652
rect 44156 36372 44212 36382
rect 44156 36278 44212 36316
rect 44828 36370 44884 37100
rect 44828 36318 44830 36370
rect 44882 36318 44884 36370
rect 44828 36306 44884 36318
rect 44604 35700 44660 35710
rect 44940 35700 44996 37212
rect 45052 36482 45108 36494
rect 45052 36430 45054 36482
rect 45106 36430 45108 36482
rect 45052 36372 45108 36430
rect 45052 36306 45108 36316
rect 45612 36482 45668 36494
rect 45612 36430 45614 36482
rect 45666 36430 45668 36482
rect 45612 35924 45668 36430
rect 45612 35858 45668 35868
rect 45724 35810 45780 38612
rect 46060 37940 46116 37950
rect 46060 37846 46116 37884
rect 45724 35758 45726 35810
rect 45778 35758 45780 35810
rect 45724 35746 45780 35758
rect 45836 37266 45892 37278
rect 45836 37214 45838 37266
rect 45890 37214 45892 37266
rect 45052 35700 45108 35710
rect 44940 35698 45108 35700
rect 44940 35646 45054 35698
rect 45106 35646 45108 35698
rect 44940 35644 45108 35646
rect 44604 35606 44660 35644
rect 43484 35074 43540 35084
rect 43596 35084 43764 35140
rect 44268 35252 44324 35262
rect 43148 34914 43316 34916
rect 43148 34862 43150 34914
rect 43202 34862 43316 34914
rect 43148 34860 43316 34862
rect 43148 34850 43204 34860
rect 43596 34580 43652 35084
rect 43932 34916 43988 34926
rect 43932 34914 44212 34916
rect 43932 34862 43934 34914
rect 43986 34862 44212 34914
rect 43932 34860 44212 34862
rect 43932 34850 43988 34860
rect 43820 34802 43876 34814
rect 43820 34750 43822 34802
rect 43874 34750 43876 34802
rect 43820 34580 43876 34750
rect 43596 34524 43764 34580
rect 43148 34244 43204 34254
rect 43148 31780 43204 34188
rect 43484 33236 43540 33246
rect 43484 33142 43540 33180
rect 43708 32676 43764 34524
rect 43820 34244 43876 34524
rect 44156 34244 44212 34860
rect 43820 34188 43988 34244
rect 43820 34020 43876 34030
rect 43820 33926 43876 33964
rect 43708 32610 43764 32620
rect 43148 31686 43204 31724
rect 43820 31780 43876 31790
rect 43260 31666 43316 31678
rect 43260 31614 43262 31666
rect 43314 31614 43316 31666
rect 43260 31556 43316 31614
rect 42700 31554 43316 31556
rect 42700 31502 42702 31554
rect 42754 31502 43316 31554
rect 42700 31500 43316 31502
rect 42700 31490 42756 31500
rect 42252 31054 42254 31106
rect 42306 31054 42308 31106
rect 41468 30942 41470 30994
rect 41522 30942 41524 30994
rect 41468 30930 41524 30942
rect 41020 29334 41076 29372
rect 41244 30098 41300 30110
rect 41244 30046 41246 30098
rect 41298 30046 41300 30098
rect 41132 28868 41188 28878
rect 41244 28868 41300 30046
rect 41580 29988 41636 29998
rect 41580 29986 41748 29988
rect 41580 29934 41582 29986
rect 41634 29934 41748 29986
rect 41580 29932 41748 29934
rect 41580 29922 41636 29932
rect 41692 29538 41748 29932
rect 41692 29486 41694 29538
rect 41746 29486 41748 29538
rect 41692 29474 41748 29486
rect 41132 28866 41300 28868
rect 41132 28814 41134 28866
rect 41186 28814 41300 28866
rect 41132 28812 41300 28814
rect 41468 28868 41524 28878
rect 41132 28802 41188 28812
rect 41468 28774 41524 28812
rect 40684 28702 40686 28754
rect 40738 28702 40740 28754
rect 40684 28644 40740 28702
rect 40236 28588 40516 28644
rect 39340 28478 39342 28530
rect 39394 28478 39396 28530
rect 39340 28466 39396 28478
rect 39676 28418 39732 28430
rect 39676 28366 39678 28418
rect 39730 28366 39732 28418
rect 39676 27748 39732 28366
rect 40348 27748 40404 27758
rect 39732 27692 39956 27748
rect 39676 27682 39732 27692
rect 38332 27134 38334 27186
rect 38386 27134 38388 27186
rect 38332 27122 38388 27134
rect 38220 26450 38276 26460
rect 38332 26964 38388 26974
rect 37324 25956 37380 25966
rect 37100 24052 37156 24062
rect 37100 23938 37156 23996
rect 37100 23886 37102 23938
rect 37154 23886 37156 23938
rect 37100 23874 37156 23886
rect 35980 23154 36036 23166
rect 35980 23102 35982 23154
rect 36034 23102 36036 23154
rect 35980 22370 36036 23102
rect 35980 22318 35982 22370
rect 36034 22318 36036 22370
rect 35980 21028 36036 22318
rect 35980 20962 36036 20972
rect 36092 23044 36148 23054
rect 35868 20750 35870 20802
rect 35922 20750 35924 20802
rect 35868 20738 35924 20750
rect 35756 20638 35758 20690
rect 35810 20638 35812 20690
rect 35756 20626 35812 20638
rect 35308 20468 35364 20478
rect 35308 20130 35364 20412
rect 35308 20078 35310 20130
rect 35362 20078 35364 20130
rect 35308 20066 35364 20078
rect 34636 19966 34638 20018
rect 34690 19966 34692 20018
rect 34636 19954 34692 19966
rect 36092 19796 36148 22988
rect 36428 20916 36484 23772
rect 37324 23826 37380 25900
rect 37548 25396 37604 26124
rect 38332 25956 38388 26908
rect 39676 26964 39732 26974
rect 39676 26870 39732 26908
rect 39900 26962 39956 27692
rect 40348 27654 40404 27692
rect 39900 26910 39902 26962
rect 39954 26910 39956 26962
rect 39900 26898 39956 26910
rect 40012 27186 40068 27198
rect 40012 27134 40014 27186
rect 40066 27134 40068 27186
rect 39676 26516 39732 26526
rect 39676 26422 39732 26460
rect 39228 26292 39284 26302
rect 39228 26198 39284 26236
rect 39452 26290 39508 26302
rect 39452 26238 39454 26290
rect 39506 26238 39508 26290
rect 38220 25900 38388 25956
rect 38444 26178 38500 26190
rect 38444 26126 38446 26178
rect 38498 26126 38500 26178
rect 37660 25620 37716 25630
rect 37660 25618 38164 25620
rect 37660 25566 37662 25618
rect 37714 25566 38164 25618
rect 37660 25564 38164 25566
rect 37660 25554 37716 25564
rect 38108 25506 38164 25564
rect 38108 25454 38110 25506
rect 38162 25454 38164 25506
rect 38108 25442 38164 25454
rect 37548 25302 37604 25340
rect 37772 25394 37828 25406
rect 37772 25342 37774 25394
rect 37826 25342 37828 25394
rect 37772 25284 37828 25342
rect 38220 25284 38276 25900
rect 38332 25732 38388 25742
rect 38332 25506 38388 25676
rect 38332 25454 38334 25506
rect 38386 25454 38388 25506
rect 38332 25442 38388 25454
rect 37772 25228 38276 25284
rect 38444 25282 38500 26126
rect 39116 25732 39172 25742
rect 38780 25620 38836 25630
rect 38668 25564 38780 25620
rect 38668 25506 38724 25564
rect 38780 25554 38836 25564
rect 38668 25454 38670 25506
rect 38722 25454 38724 25506
rect 38668 25442 38724 25454
rect 38444 25230 38446 25282
rect 38498 25230 38500 25282
rect 37324 23774 37326 23826
rect 37378 23774 37380 23826
rect 37324 23762 37380 23774
rect 37996 24388 38052 25228
rect 38444 25218 38500 25230
rect 38780 25396 38836 25406
rect 38668 24724 38724 24734
rect 38780 24724 38836 25340
rect 38668 24722 38836 24724
rect 38668 24670 38670 24722
rect 38722 24670 38836 24722
rect 38668 24668 38836 24670
rect 38668 24658 38724 24668
rect 38444 24610 38500 24622
rect 38444 24558 38446 24610
rect 38498 24558 38500 24610
rect 38444 24500 38500 24558
rect 38668 24500 38724 24510
rect 38892 24500 38948 24510
rect 38444 24444 38668 24500
rect 38724 24498 38948 24500
rect 38724 24446 38894 24498
rect 38946 24446 38948 24498
rect 38724 24444 38948 24446
rect 38668 24406 38724 24444
rect 38892 24434 38948 24444
rect 37996 23826 38052 24332
rect 39116 24276 39172 25676
rect 39452 25618 39508 26238
rect 39788 26290 39844 26302
rect 39788 26238 39790 26290
rect 39842 26238 39844 26290
rect 39788 25732 39844 26238
rect 40012 26290 40068 27134
rect 40460 26908 40516 28588
rect 40684 28578 40740 28588
rect 41916 28644 41972 28654
rect 41916 28550 41972 28588
rect 41580 28532 41636 28542
rect 41580 28082 41636 28476
rect 42252 28532 42308 31054
rect 42812 30884 42868 30894
rect 42812 30790 42868 30828
rect 42700 30212 42756 30222
rect 43260 30212 43316 31500
rect 43820 30884 43876 31724
rect 43820 30818 43876 30828
rect 43260 30156 43652 30212
rect 42700 29428 42756 30156
rect 42252 28438 42308 28476
rect 42364 28980 42420 28990
rect 41580 28030 41582 28082
rect 41634 28030 41636 28082
rect 41580 28018 41636 28030
rect 42252 28084 42308 28094
rect 42364 28084 42420 28924
rect 42252 28082 42420 28084
rect 42252 28030 42254 28082
rect 42306 28030 42420 28082
rect 42252 28028 42420 28030
rect 42252 28018 42308 28028
rect 41244 27858 41300 27870
rect 41244 27806 41246 27858
rect 41298 27806 41300 27858
rect 40460 26852 40740 26908
rect 40012 26238 40014 26290
rect 40066 26238 40068 26290
rect 40012 26226 40068 26238
rect 39788 25666 39844 25676
rect 40124 26180 40180 26190
rect 39452 25566 39454 25618
rect 39506 25566 39508 25618
rect 39452 25554 39508 25566
rect 39564 25508 39620 25518
rect 39788 25508 39844 25518
rect 39564 25414 39620 25452
rect 39676 25506 39844 25508
rect 39676 25454 39790 25506
rect 39842 25454 39844 25506
rect 39676 25452 39844 25454
rect 39340 25394 39396 25406
rect 39340 25342 39342 25394
rect 39394 25342 39396 25394
rect 39340 25284 39396 25342
rect 39340 25218 39396 25228
rect 39676 25060 39732 25452
rect 39788 25442 39844 25452
rect 40012 25508 40068 25518
rect 40124 25508 40180 26124
rect 40348 25732 40404 25742
rect 40012 25506 40180 25508
rect 40012 25454 40014 25506
rect 40066 25454 40180 25506
rect 40012 25452 40180 25454
rect 40236 25676 40348 25732
rect 40236 25506 40292 25676
rect 40348 25666 40404 25676
rect 40572 25620 40628 25630
rect 40572 25526 40628 25564
rect 40236 25454 40238 25506
rect 40290 25454 40292 25506
rect 40012 25442 40068 25452
rect 40236 25442 40292 25454
rect 40460 25508 40516 25518
rect 39228 25004 39732 25060
rect 39788 25284 39844 25294
rect 39228 24946 39284 25004
rect 39228 24894 39230 24946
rect 39282 24894 39284 24946
rect 39228 24882 39284 24894
rect 39676 24612 39732 24622
rect 39788 24612 39844 25228
rect 39676 24610 39844 24612
rect 39676 24558 39678 24610
rect 39730 24558 39844 24610
rect 39676 24556 39844 24558
rect 40012 24612 40068 24622
rect 39676 24498 39732 24556
rect 39676 24446 39678 24498
rect 39730 24446 39732 24498
rect 39116 24220 39396 24276
rect 37996 23774 37998 23826
rect 38050 23774 38052 23826
rect 37996 23762 38052 23774
rect 38892 23938 38948 23950
rect 38892 23886 38894 23938
rect 38946 23886 38948 23938
rect 37436 23716 37492 23726
rect 37436 23380 37492 23660
rect 37436 23314 37492 23324
rect 37660 23714 37716 23726
rect 37660 23662 37662 23714
rect 37714 23662 37716 23714
rect 37660 23604 37716 23662
rect 38332 23714 38388 23726
rect 38332 23662 38334 23714
rect 38386 23662 38388 23714
rect 38332 23604 38388 23662
rect 37660 23548 38388 23604
rect 38892 23604 38948 23886
rect 37100 22148 37156 22158
rect 37548 22148 37604 22158
rect 37100 22146 37548 22148
rect 37100 22094 37102 22146
rect 37154 22094 37548 22146
rect 37100 22092 37548 22094
rect 37100 21700 37156 22092
rect 37548 22054 37604 22092
rect 36428 20822 36484 20860
rect 36764 21644 37156 21700
rect 37548 21700 37604 21710
rect 35196 19628 35460 19638
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35196 19562 35460 19572
rect 34412 19182 34414 19234
rect 34466 19182 34468 19234
rect 34412 19170 34468 19182
rect 35308 19460 35364 19470
rect 32844 18610 32900 18620
rect 32620 17602 32676 17612
rect 32956 18564 33012 18574
rect 32956 17556 33012 18508
rect 32956 17462 33012 17500
rect 33068 18340 33124 18350
rect 32620 17444 32676 17454
rect 32396 17442 32676 17444
rect 32396 17390 32622 17442
rect 32674 17390 32676 17442
rect 32396 17388 32676 17390
rect 32396 17220 32452 17388
rect 32620 17378 32676 17388
rect 32844 17442 32900 17454
rect 32844 17390 32846 17442
rect 32898 17390 32900 17442
rect 32172 17164 32452 17220
rect 31612 15988 31668 15998
rect 31612 15426 31668 15932
rect 31612 15374 31614 15426
rect 31666 15374 31668 15426
rect 31612 15362 31668 15374
rect 31724 15428 31780 15438
rect 31836 15428 31892 16492
rect 31724 15426 31892 15428
rect 31724 15374 31726 15426
rect 31778 15374 31892 15426
rect 31724 15372 31892 15374
rect 31948 16100 32004 16110
rect 32060 16100 32116 17164
rect 32844 16996 32900 17390
rect 32844 16930 32900 16940
rect 33068 17108 33124 18284
rect 33516 17554 33572 18956
rect 33516 17502 33518 17554
rect 33570 17502 33572 17554
rect 33516 17490 33572 17502
rect 33964 19010 34132 19012
rect 33964 18958 34078 19010
rect 34130 18958 34132 19010
rect 33964 18956 34132 18958
rect 33852 17442 33908 17454
rect 33852 17390 33854 17442
rect 33906 17390 33908 17442
rect 33068 16994 33124 17052
rect 33292 17108 33348 17118
rect 33292 17106 33684 17108
rect 33292 17054 33294 17106
rect 33346 17054 33684 17106
rect 33292 17052 33684 17054
rect 33292 17042 33348 17052
rect 33068 16942 33070 16994
rect 33122 16942 33124 16994
rect 33068 16930 33124 16942
rect 33516 16884 33572 16894
rect 33516 16790 33572 16828
rect 31948 16098 32116 16100
rect 31948 16046 31950 16098
rect 32002 16046 32116 16098
rect 31948 16044 32116 16046
rect 33068 16660 33124 16670
rect 31724 15362 31780 15372
rect 31948 15314 32004 16044
rect 33068 15988 33124 16604
rect 33068 15538 33124 15932
rect 33068 15486 33070 15538
rect 33122 15486 33124 15538
rect 33068 15474 33124 15486
rect 31948 15262 31950 15314
rect 32002 15262 32004 15314
rect 31948 15250 32004 15262
rect 33292 15314 33348 15326
rect 33292 15262 33294 15314
rect 33346 15262 33348 15314
rect 31164 15092 31220 15102
rect 31500 15092 31668 15148
rect 29820 14466 29876 14476
rect 29932 14756 29988 14766
rect 29708 14306 29764 14318
rect 29708 14254 29710 14306
rect 29762 14254 29764 14306
rect 29596 14196 29652 14206
rect 29372 13682 29428 13692
rect 29484 13860 29540 13870
rect 29484 13074 29540 13804
rect 29596 13746 29652 14140
rect 29596 13694 29598 13746
rect 29650 13694 29652 13746
rect 29596 13682 29652 13694
rect 29484 13022 29486 13074
rect 29538 13022 29540 13074
rect 29484 13010 29540 13022
rect 29596 12852 29652 12862
rect 29708 12852 29764 14254
rect 29820 12852 29876 12862
rect 29708 12796 29820 12852
rect 29372 12740 29428 12750
rect 28476 11396 28532 11406
rect 28476 11302 28532 11340
rect 29036 11394 29092 11452
rect 29036 11342 29038 11394
rect 29090 11342 29092 11394
rect 29036 11330 29092 11342
rect 29148 12738 29428 12740
rect 29148 12686 29374 12738
rect 29426 12686 29428 12738
rect 29148 12684 29428 12686
rect 28588 11172 28644 11182
rect 29148 11172 29204 12684
rect 29372 12674 29428 12684
rect 29260 12516 29316 12526
rect 29260 12290 29316 12460
rect 29372 12404 29428 12414
rect 29372 12310 29428 12348
rect 29260 12238 29262 12290
rect 29314 12238 29316 12290
rect 29260 12226 29316 12238
rect 29596 11508 29652 12796
rect 29820 12786 29876 12796
rect 29932 12404 29988 14700
rect 30044 13634 30100 15092
rect 30492 15090 31220 15092
rect 30492 15038 31166 15090
rect 31218 15038 31220 15090
rect 30492 15036 31220 15038
rect 30156 14532 30212 14542
rect 30156 14438 30212 14476
rect 30380 14418 30436 14430
rect 30380 14366 30382 14418
rect 30434 14366 30436 14418
rect 30380 14084 30436 14366
rect 30380 14018 30436 14028
rect 30044 13582 30046 13634
rect 30098 13582 30100 13634
rect 30044 12962 30100 13582
rect 30044 12910 30046 12962
rect 30098 12910 30100 12962
rect 30044 12898 30100 12910
rect 30380 13076 30436 13086
rect 30268 12852 30324 12862
rect 29932 12348 30212 12404
rect 30044 12180 30100 12190
rect 30044 11618 30100 12124
rect 30044 11566 30046 11618
rect 30098 11566 30100 11618
rect 30044 11554 30100 11566
rect 29596 11452 29988 11508
rect 29372 11396 29428 11406
rect 29372 11302 29428 11340
rect 29596 11282 29652 11452
rect 29932 11396 29988 11452
rect 29932 11340 30100 11396
rect 29596 11230 29598 11282
rect 29650 11230 29652 11282
rect 29596 11218 29652 11230
rect 29708 11284 29764 11294
rect 30044 11282 30100 11340
rect 29708 11190 29764 11228
rect 29932 11226 29988 11238
rect 28588 11170 29204 11172
rect 28588 11118 28590 11170
rect 28642 11118 29204 11170
rect 28588 11116 29204 11118
rect 29932 11174 29934 11226
rect 29986 11174 29988 11226
rect 30044 11230 30046 11282
rect 30098 11230 30100 11282
rect 30044 11218 30100 11230
rect 28588 11106 28644 11116
rect 29932 11060 29988 11174
rect 30156 11060 30212 12348
rect 29932 11004 30212 11060
rect 30268 12292 30324 12796
rect 30380 12850 30436 13020
rect 30380 12798 30382 12850
rect 30434 12798 30436 12850
rect 30380 12786 30436 12798
rect 29372 10836 29428 10846
rect 29036 10724 29092 10734
rect 29372 10724 29428 10780
rect 29036 10722 29428 10724
rect 29036 10670 29038 10722
rect 29090 10670 29374 10722
rect 29426 10670 29428 10722
rect 29036 10668 29428 10670
rect 29036 10658 29092 10668
rect 29372 10658 29428 10668
rect 28140 10498 28308 10500
rect 28140 10446 28142 10498
rect 28194 10446 28308 10498
rect 28140 10444 28308 10446
rect 28476 10610 28532 10622
rect 28476 10558 28478 10610
rect 28530 10558 28532 10610
rect 28140 10434 28196 10444
rect 28028 10388 28084 10398
rect 28028 9154 28084 10332
rect 28476 10052 28532 10558
rect 28700 10612 28756 10622
rect 28700 10518 28756 10556
rect 29484 10612 29540 10622
rect 28588 10500 28644 10510
rect 28588 10406 28644 10444
rect 28476 9996 29092 10052
rect 28588 9828 28644 9838
rect 28364 9772 28588 9828
rect 28028 9102 28030 9154
rect 28082 9102 28084 9154
rect 28028 9090 28084 9102
rect 28140 9156 28196 9166
rect 28140 9154 28308 9156
rect 28140 9102 28142 9154
rect 28194 9102 28308 9154
rect 28140 9100 28308 9102
rect 28140 9090 28196 9100
rect 28140 8820 28196 8830
rect 27916 8818 28196 8820
rect 27916 8766 28142 8818
rect 28194 8766 28196 8818
rect 27916 8764 28196 8766
rect 28140 8754 28196 8764
rect 28252 8708 28308 9100
rect 28252 8642 28308 8652
rect 27468 8530 27524 8540
rect 22428 8370 23044 8372
rect 22428 8318 22430 8370
rect 22482 8318 23044 8370
rect 22428 8316 23044 8318
rect 25676 8370 25732 8382
rect 25676 8318 25678 8370
rect 25730 8318 25732 8370
rect 22428 8306 22484 8316
rect 22764 8258 22820 8316
rect 22764 8206 22766 8258
rect 22818 8206 22820 8258
rect 22764 8194 22820 8206
rect 23548 8148 23604 8158
rect 21980 7644 22260 7700
rect 23212 8146 23604 8148
rect 23212 8094 23550 8146
rect 23602 8094 23604 8146
rect 23212 8092 23604 8094
rect 21980 7586 22036 7644
rect 21980 7534 21982 7586
rect 22034 7534 22036 7586
rect 21980 7522 22036 7534
rect 22764 7362 22820 7374
rect 22764 7310 22766 7362
rect 22818 7310 22820 7362
rect 22652 7250 22708 7262
rect 22652 7198 22654 7250
rect 22706 7198 22708 7250
rect 21980 6692 22036 6702
rect 22036 6636 22148 6692
rect 21980 6598 22036 6636
rect 21420 6466 21588 6468
rect 21420 6414 21422 6466
rect 21474 6414 21588 6466
rect 21420 6412 21588 6414
rect 21420 6402 21476 6412
rect 21308 6356 21364 6366
rect 21308 5906 21364 6300
rect 21308 5854 21310 5906
rect 21362 5854 21364 5906
rect 21308 5842 21364 5854
rect 21420 6020 21476 6030
rect 20972 5170 21028 5180
rect 21420 5234 21476 5964
rect 21532 5796 21588 6412
rect 21532 5730 21588 5740
rect 21644 6018 21700 6030
rect 21644 5966 21646 6018
rect 21698 5966 21700 6018
rect 21532 5348 21588 5358
rect 21532 5254 21588 5292
rect 21420 5182 21422 5234
rect 21474 5182 21476 5234
rect 21420 5170 21476 5182
rect 20412 5058 20468 5068
rect 21644 4564 21700 5966
rect 21980 5908 22036 5918
rect 21980 5346 22036 5852
rect 21980 5294 21982 5346
rect 22034 5294 22036 5346
rect 21980 5282 22036 5294
rect 22092 5346 22148 6636
rect 22204 6466 22260 6478
rect 22540 6468 22596 6478
rect 22204 6414 22206 6466
rect 22258 6414 22260 6466
rect 22204 6356 22260 6414
rect 22204 6290 22260 6300
rect 22428 6466 22596 6468
rect 22428 6414 22542 6466
rect 22594 6414 22596 6466
rect 22428 6412 22596 6414
rect 22092 5294 22094 5346
rect 22146 5294 22148 5346
rect 22092 5282 22148 5294
rect 22204 5906 22260 5918
rect 22204 5854 22206 5906
rect 22258 5854 22260 5906
rect 22204 5348 22260 5854
rect 22316 5906 22372 5918
rect 22316 5854 22318 5906
rect 22370 5854 22372 5906
rect 22316 5572 22372 5854
rect 22428 5908 22484 6412
rect 22540 6402 22596 6412
rect 22540 6132 22596 6142
rect 22652 6132 22708 7198
rect 22764 6468 22820 7310
rect 23212 6802 23268 8092
rect 23548 8082 23604 8092
rect 25452 7588 25508 7598
rect 23212 6750 23214 6802
rect 23266 6750 23268 6802
rect 23212 6738 23268 6750
rect 23436 7364 23492 7374
rect 23100 6692 23156 6702
rect 23100 6578 23156 6636
rect 23100 6526 23102 6578
rect 23154 6526 23156 6578
rect 23100 6514 23156 6526
rect 23212 6578 23268 6590
rect 23212 6526 23214 6578
rect 23266 6526 23268 6578
rect 22876 6468 22932 6478
rect 22988 6468 23044 6478
rect 22764 6466 22988 6468
rect 22764 6414 22878 6466
rect 22930 6414 22988 6466
rect 22764 6412 22988 6414
rect 22876 6402 22932 6412
rect 22540 6130 22708 6132
rect 22540 6078 22542 6130
rect 22594 6078 22708 6130
rect 22540 6076 22708 6078
rect 22764 6244 22820 6254
rect 22764 6130 22820 6188
rect 22764 6078 22766 6130
rect 22818 6078 22820 6130
rect 22540 6066 22596 6076
rect 22764 6066 22820 6078
rect 22764 5908 22820 5918
rect 22428 5852 22764 5908
rect 22764 5814 22820 5852
rect 22316 5506 22372 5516
rect 22428 5348 22484 5358
rect 22204 5346 22484 5348
rect 22204 5294 22430 5346
rect 22482 5294 22484 5346
rect 22204 5292 22484 5294
rect 22428 5282 22484 5292
rect 22764 5236 22820 5246
rect 22316 5124 22372 5134
rect 22204 5122 22372 5124
rect 22204 5070 22318 5122
rect 22370 5070 22372 5122
rect 22204 5068 22372 5070
rect 22204 4676 22260 5068
rect 22316 5058 22372 5068
rect 22428 5124 22484 5134
rect 21980 4564 22036 4574
rect 21644 4562 22036 4564
rect 21644 4510 21982 4562
rect 22034 4510 22036 4562
rect 21644 4508 22036 4510
rect 21532 4228 21588 4238
rect 21644 4228 21700 4508
rect 21980 4498 22036 4508
rect 22092 4564 22148 4574
rect 22092 4470 22148 4508
rect 22204 4562 22260 4620
rect 22204 4510 22206 4562
rect 22258 4510 22260 4562
rect 22204 4498 22260 4510
rect 22316 4900 22372 4910
rect 22316 4450 22372 4844
rect 22316 4398 22318 4450
rect 22370 4398 22372 4450
rect 22316 4386 22372 4398
rect 21532 4226 21700 4228
rect 21532 4174 21534 4226
rect 21586 4174 21700 4226
rect 21532 4172 21700 4174
rect 21532 4162 21588 4172
rect 20300 3490 20356 3500
rect 20860 3668 20916 3678
rect 19836 3164 20100 3174
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 19836 3098 20100 3108
rect 20860 800 20916 3612
rect 22092 3668 22148 3678
rect 22092 3574 22148 3612
rect 21084 3556 21140 3566
rect 21084 3462 21140 3500
rect 22428 3388 22484 5068
rect 22764 4676 22820 5180
rect 22876 5122 22932 5134
rect 22876 5070 22878 5122
rect 22930 5070 22932 5122
rect 22876 5012 22932 5070
rect 22876 4946 22932 4956
rect 22764 4620 22932 4676
rect 22764 4452 22820 4462
rect 22764 4338 22820 4396
rect 22764 4286 22766 4338
rect 22818 4286 22820 4338
rect 22764 4274 22820 4286
rect 22876 4340 22932 4620
rect 22988 4564 23044 6412
rect 23100 6020 23156 6030
rect 23100 5926 23156 5964
rect 23100 5572 23156 5582
rect 23212 5572 23268 6526
rect 23324 6020 23380 6030
rect 23324 5684 23380 5964
rect 23324 5618 23380 5628
rect 23436 5906 23492 7308
rect 23548 7362 23604 7374
rect 23548 7310 23550 7362
rect 23602 7310 23604 7362
rect 23548 6020 23604 7310
rect 24444 7364 24500 7374
rect 24444 7270 24500 7308
rect 23660 6690 23716 6702
rect 23660 6638 23662 6690
rect 23714 6638 23716 6690
rect 23660 6580 23716 6638
rect 24780 6690 24836 6702
rect 24780 6638 24782 6690
rect 24834 6638 24836 6690
rect 23660 6514 23716 6524
rect 23996 6578 24052 6590
rect 23996 6526 23998 6578
rect 24050 6526 24052 6578
rect 23996 6468 24052 6526
rect 24332 6580 24388 6590
rect 24332 6486 24388 6524
rect 23996 6402 24052 6412
rect 24108 6466 24164 6478
rect 24108 6414 24110 6466
rect 24162 6414 24164 6466
rect 23884 6020 23940 6030
rect 23548 5964 23716 6020
rect 23436 5854 23438 5906
rect 23490 5854 23492 5906
rect 23156 5516 23268 5572
rect 23100 5010 23156 5516
rect 23436 5124 23492 5854
rect 23436 5058 23492 5068
rect 23548 5796 23604 5806
rect 23548 5122 23604 5740
rect 23548 5070 23550 5122
rect 23602 5070 23604 5122
rect 23548 5058 23604 5070
rect 23100 4958 23102 5010
rect 23154 4958 23156 5010
rect 23100 4946 23156 4958
rect 23436 4564 23492 4574
rect 22988 4562 23492 4564
rect 22988 4510 23438 4562
rect 23490 4510 23492 4562
rect 22988 4508 23492 4510
rect 23436 4498 23492 4508
rect 23660 4452 23716 5964
rect 23884 6018 24052 6020
rect 23884 5966 23886 6018
rect 23938 5966 24052 6018
rect 23884 5964 24052 5966
rect 23884 5954 23940 5964
rect 23772 5906 23828 5918
rect 23772 5854 23774 5906
rect 23826 5854 23828 5906
rect 23772 5348 23828 5854
rect 23772 5282 23828 5292
rect 23884 5682 23940 5694
rect 23884 5630 23886 5682
rect 23938 5630 23940 5682
rect 23772 4452 23828 4462
rect 23660 4450 23828 4452
rect 23660 4398 23774 4450
rect 23826 4398 23828 4450
rect 23660 4396 23828 4398
rect 23100 4340 23156 4350
rect 22876 4338 23156 4340
rect 22876 4286 23102 4338
rect 23154 4286 23156 4338
rect 22876 4284 23156 4286
rect 22204 3332 22484 3388
rect 22204 800 22260 3332
rect 22988 980 23044 4284
rect 23100 4274 23156 4284
rect 23660 3388 23716 4396
rect 23772 4386 23828 4396
rect 23884 4452 23940 5630
rect 23996 4788 24052 5964
rect 23996 4722 24052 4732
rect 24108 4562 24164 6414
rect 24444 5796 24500 5806
rect 24444 5702 24500 5740
rect 24780 5796 24836 6638
rect 25452 6690 25508 7532
rect 25452 6638 25454 6690
rect 25506 6638 25508 6690
rect 25452 6626 25508 6638
rect 25676 6244 25732 8318
rect 27916 8372 27972 8382
rect 27132 8148 27188 8158
rect 27132 8054 27188 8092
rect 27580 8148 27636 8158
rect 27580 8054 27636 8092
rect 27804 8146 27860 8158
rect 27804 8094 27806 8146
rect 27858 8094 27860 8146
rect 26012 8036 26068 8046
rect 26012 7700 26068 7980
rect 27692 8034 27748 8046
rect 27692 7982 27694 8034
rect 27746 7982 27748 8034
rect 26012 7606 26068 7644
rect 27468 7924 27524 7934
rect 26348 7586 26404 7598
rect 26348 7534 26350 7586
rect 26402 7534 26404 7586
rect 26348 6468 26404 7534
rect 27132 7588 27188 7598
rect 27132 7494 27188 7532
rect 26348 6402 26404 6412
rect 26572 7474 26628 7486
rect 26572 7422 26574 7474
rect 26626 7422 26628 7474
rect 24780 5730 24836 5740
rect 25340 5796 25396 5806
rect 25340 5794 25620 5796
rect 25340 5742 25342 5794
rect 25394 5742 25620 5794
rect 25340 5740 25620 5742
rect 25340 5730 25396 5740
rect 24220 5684 24276 5694
rect 24220 5234 24276 5628
rect 25228 5684 25284 5694
rect 25228 5590 25284 5628
rect 25452 5572 25508 5582
rect 24220 5182 24222 5234
rect 24274 5182 24276 5234
rect 24220 5170 24276 5182
rect 24780 5348 24836 5358
rect 24668 5124 24724 5134
rect 24108 4510 24110 4562
rect 24162 4510 24164 4562
rect 24108 4498 24164 4510
rect 24556 4788 24612 4798
rect 24556 4562 24612 4732
rect 24556 4510 24558 4562
rect 24610 4510 24612 4562
rect 24556 4498 24612 4510
rect 23884 4386 23940 4396
rect 24668 4450 24724 5068
rect 24668 4398 24670 4450
rect 24722 4398 24724 4450
rect 24668 4386 24724 4398
rect 24556 4228 24612 4238
rect 24556 4114 24612 4172
rect 24556 4062 24558 4114
rect 24610 4062 24612 4114
rect 24556 4050 24612 4062
rect 24668 3556 24724 3566
rect 24780 3556 24836 5292
rect 24668 3554 24836 3556
rect 24668 3502 24670 3554
rect 24722 3502 24836 3554
rect 24668 3500 24836 3502
rect 24668 3490 24724 3500
rect 22876 924 23044 980
rect 23548 3332 23716 3388
rect 22876 800 22932 924
rect 23548 800 23604 3332
rect 24780 3108 24836 3500
rect 24892 5236 24948 5246
rect 24892 3442 24948 5180
rect 25228 4338 25284 4350
rect 25228 4286 25230 4338
rect 25282 4286 25284 4338
rect 25228 4228 25284 4286
rect 25228 4162 25284 4172
rect 25452 3554 25508 5516
rect 25564 4228 25620 5740
rect 25676 5572 25732 6188
rect 26572 6244 26628 7422
rect 27468 7474 27524 7868
rect 27468 7422 27470 7474
rect 27522 7422 27524 7474
rect 27468 7410 27524 7422
rect 27468 7250 27524 7262
rect 27468 7198 27470 7250
rect 27522 7198 27524 7250
rect 26572 6178 26628 6188
rect 26684 6468 26740 6478
rect 26348 6132 26404 6142
rect 25788 6130 26404 6132
rect 25788 6078 26350 6130
rect 26402 6078 26404 6130
rect 25788 6076 26404 6078
rect 25788 6018 25844 6076
rect 26348 6066 26404 6076
rect 25788 5966 25790 6018
rect 25842 5966 25844 6018
rect 25788 5954 25844 5966
rect 26236 5908 26292 5918
rect 26460 5908 26516 5918
rect 25676 5506 25732 5516
rect 25900 5682 25956 5694
rect 25900 5630 25902 5682
rect 25954 5630 25956 5682
rect 25676 5012 25732 5022
rect 25676 4450 25732 4956
rect 25788 4900 25844 4910
rect 25788 4676 25844 4844
rect 25788 4562 25844 4620
rect 25788 4510 25790 4562
rect 25842 4510 25844 4562
rect 25788 4498 25844 4510
rect 25676 4398 25678 4450
rect 25730 4398 25732 4450
rect 25676 4386 25732 4398
rect 25676 4228 25732 4238
rect 25564 4226 25732 4228
rect 25564 4174 25678 4226
rect 25730 4174 25732 4226
rect 25564 4172 25732 4174
rect 25676 4162 25732 4172
rect 25452 3502 25454 3554
rect 25506 3502 25508 3554
rect 25452 3490 25508 3502
rect 25900 3556 25956 5630
rect 26236 5684 26292 5852
rect 26236 5618 26292 5628
rect 26348 5906 26516 5908
rect 26348 5854 26462 5906
rect 26514 5854 26516 5906
rect 26348 5852 26516 5854
rect 26348 5236 26404 5852
rect 26460 5842 26516 5852
rect 26684 5572 26740 6412
rect 27468 6130 27524 7198
rect 27468 6078 27470 6130
rect 27522 6078 27524 6130
rect 27468 6066 27524 6078
rect 27692 6130 27748 7982
rect 27804 6802 27860 8094
rect 27916 7698 27972 8316
rect 27916 7646 27918 7698
rect 27970 7646 27972 7698
rect 27916 6916 27972 7646
rect 28364 7474 28420 9772
rect 28588 9734 28644 9772
rect 29036 9826 29092 9996
rect 29036 9774 29038 9826
rect 29090 9774 29092 9826
rect 29036 9762 29092 9774
rect 29148 9828 29204 9838
rect 29148 9266 29204 9772
rect 29372 9828 29428 9838
rect 29484 9828 29540 10556
rect 29596 10610 29652 10622
rect 29596 10558 29598 10610
rect 29650 10558 29652 10610
rect 29596 10276 29652 10558
rect 29932 10388 29988 11004
rect 30268 10612 30324 12236
rect 30268 10546 30324 10556
rect 30380 12404 30436 12414
rect 29932 10322 29988 10332
rect 30156 10500 30212 10510
rect 29596 10210 29652 10220
rect 30156 10276 30212 10444
rect 30156 10210 30212 10220
rect 30156 10052 30212 10062
rect 29372 9826 29540 9828
rect 29372 9774 29374 9826
rect 29426 9774 29540 9826
rect 29372 9772 29540 9774
rect 30044 9938 30100 9950
rect 30044 9886 30046 9938
rect 30098 9886 30100 9938
rect 29372 9762 29428 9772
rect 29260 9604 29316 9614
rect 29260 9510 29316 9548
rect 29148 9214 29150 9266
rect 29202 9214 29204 9266
rect 29148 9202 29204 9214
rect 28700 8930 28756 8942
rect 28700 8878 28702 8930
rect 28754 8878 28756 8930
rect 28700 8708 28756 8878
rect 28700 8642 28756 8652
rect 29932 8932 29988 8942
rect 29932 8484 29988 8876
rect 29932 8418 29988 8428
rect 28700 8372 28756 8382
rect 28700 8278 28756 8316
rect 30044 8260 30100 9886
rect 30156 9716 30212 9996
rect 30380 10050 30436 12348
rect 30380 9998 30382 10050
rect 30434 9998 30436 10050
rect 30380 9986 30436 9998
rect 30156 9622 30212 9660
rect 30044 8194 30100 8204
rect 30380 8930 30436 8942
rect 30380 8878 30382 8930
rect 30434 8878 30436 8930
rect 30380 8818 30436 8878
rect 30380 8766 30382 8818
rect 30434 8766 30436 8818
rect 29372 8148 29428 8158
rect 28364 7422 28366 7474
rect 28418 7422 28420 7474
rect 28364 7410 28420 7422
rect 28924 7476 28980 7486
rect 28924 7382 28980 7420
rect 27916 6850 27972 6860
rect 27804 6750 27806 6802
rect 27858 6750 27860 6802
rect 27804 6738 27860 6750
rect 29372 6692 29428 8092
rect 29820 8146 29876 8158
rect 29820 8094 29822 8146
rect 29874 8094 29876 8146
rect 29484 8036 29540 8046
rect 29820 8036 29876 8094
rect 29484 8034 29652 8036
rect 29484 7982 29486 8034
rect 29538 7982 29652 8034
rect 29484 7980 29652 7982
rect 29484 7970 29540 7980
rect 29596 7924 29652 7980
rect 29484 6692 29540 6702
rect 29372 6690 29540 6692
rect 29372 6638 29486 6690
rect 29538 6638 29540 6690
rect 29372 6636 29540 6638
rect 27692 6078 27694 6130
rect 27746 6078 27748 6130
rect 27692 6066 27748 6078
rect 28700 6466 28756 6478
rect 28700 6414 28702 6466
rect 28754 6414 28756 6466
rect 28700 6020 28756 6414
rect 29484 6356 29540 6636
rect 29484 6290 29540 6300
rect 29484 6132 29540 6142
rect 28700 5954 28756 5964
rect 28924 6130 29540 6132
rect 28924 6078 29486 6130
rect 29538 6078 29540 6130
rect 28924 6076 29540 6078
rect 29596 6132 29652 7868
rect 29820 7476 29876 7980
rect 29820 7410 29876 7420
rect 29932 8034 29988 8046
rect 29932 7982 29934 8034
rect 29986 7982 29988 8034
rect 29708 6692 29764 6702
rect 29708 6598 29764 6636
rect 29932 6580 29988 7982
rect 30044 8034 30100 8046
rect 30044 7982 30046 8034
rect 30098 7982 30100 8034
rect 30044 7924 30100 7982
rect 30044 7858 30100 7868
rect 30380 7028 30436 8766
rect 30492 8260 30548 15036
rect 31164 15026 31220 15036
rect 30940 14756 30996 14766
rect 30716 14308 30772 14346
rect 30716 14242 30772 14252
rect 30716 14084 30772 14094
rect 30716 13746 30772 14028
rect 30940 13970 30996 14700
rect 31164 14420 31220 14430
rect 30940 13918 30942 13970
rect 30994 13918 30996 13970
rect 30940 13906 30996 13918
rect 31052 14418 31220 14420
rect 31052 14366 31166 14418
rect 31218 14366 31220 14418
rect 31052 14364 31220 14366
rect 31052 13970 31108 14364
rect 31164 14354 31220 14364
rect 31276 14420 31332 14430
rect 31276 14326 31332 14364
rect 31052 13918 31054 13970
rect 31106 13918 31108 13970
rect 31052 13906 31108 13918
rect 30716 13694 30718 13746
rect 30770 13694 30772 13746
rect 30716 13682 30772 13694
rect 31164 13858 31220 13870
rect 31164 13806 31166 13858
rect 31218 13806 31220 13858
rect 31164 13748 31220 13806
rect 31276 13860 31332 13870
rect 31276 13766 31332 13804
rect 31164 13682 31220 13692
rect 31500 13524 31556 13534
rect 31164 13412 31220 13422
rect 31220 13356 31444 13412
rect 31164 13346 31220 13356
rect 30716 13132 31220 13188
rect 30604 12964 30660 12974
rect 30716 12964 30772 13132
rect 30604 12962 30772 12964
rect 30604 12910 30606 12962
rect 30658 12910 30772 12962
rect 30604 12908 30772 12910
rect 30828 12962 30884 12974
rect 30828 12910 30830 12962
rect 30882 12910 30884 12962
rect 30604 12898 30660 12908
rect 30604 11394 30660 11406
rect 30828 11396 30884 12910
rect 30940 12180 30996 12190
rect 30940 12086 30996 12124
rect 31164 12178 31220 13132
rect 31164 12126 31166 12178
rect 31218 12126 31220 12178
rect 31164 12114 31220 12126
rect 31052 12066 31108 12078
rect 31052 12014 31054 12066
rect 31106 12014 31108 12066
rect 31052 11620 31108 12014
rect 31052 11554 31108 11564
rect 31164 11956 31220 11966
rect 30604 11342 30606 11394
rect 30658 11342 30660 11394
rect 30604 11284 30660 11342
rect 30604 11218 30660 11228
rect 30716 11340 30828 11396
rect 30604 11060 30660 11070
rect 30604 10722 30660 11004
rect 30604 10670 30606 10722
rect 30658 10670 30660 10722
rect 30604 10658 30660 10670
rect 30716 9828 30772 11340
rect 30828 11330 30884 11340
rect 31052 11396 31108 11406
rect 31164 11396 31220 11900
rect 31052 11394 31220 11396
rect 31052 11342 31054 11394
rect 31106 11342 31220 11394
rect 31052 11340 31220 11342
rect 31052 11330 31108 11340
rect 31276 11282 31332 11294
rect 31276 11230 31278 11282
rect 31330 11230 31332 11282
rect 30828 11172 30884 11182
rect 30828 11078 30884 11116
rect 31164 10836 31220 10846
rect 31276 10836 31332 11230
rect 31220 10780 31332 10836
rect 31164 10770 31220 10780
rect 30828 10610 30884 10622
rect 30828 10558 30830 10610
rect 30882 10558 30884 10610
rect 30828 10052 30884 10558
rect 31164 10612 31220 10622
rect 31164 10518 31220 10556
rect 31388 10612 31444 13356
rect 31500 13076 31556 13468
rect 31612 13300 31668 15092
rect 33292 14420 33348 15262
rect 33180 14196 33236 14206
rect 31724 14084 31780 14094
rect 31724 13746 31780 14028
rect 31724 13694 31726 13746
rect 31778 13694 31780 13746
rect 31724 13682 31780 13694
rect 32284 13636 32340 13646
rect 31612 13244 31780 13300
rect 31612 13076 31668 13086
rect 31500 13074 31668 13076
rect 31500 13022 31614 13074
rect 31666 13022 31668 13074
rect 31500 13020 31668 13022
rect 31612 13010 31668 13020
rect 31724 12404 31780 13244
rect 31724 12338 31780 12348
rect 31836 12292 31892 12302
rect 31836 12198 31892 12236
rect 31948 12292 32004 12302
rect 31948 12290 32228 12292
rect 31948 12238 31950 12290
rect 32002 12238 32228 12290
rect 31948 12236 32228 12238
rect 31948 12226 32004 12236
rect 31500 12178 31556 12190
rect 31500 12126 31502 12178
rect 31554 12126 31556 12178
rect 31500 11788 31556 12126
rect 31948 11956 32004 11966
rect 31948 11862 32004 11900
rect 32172 11956 32228 12236
rect 32172 11890 32228 11900
rect 31500 11732 31780 11788
rect 31724 10836 31780 11732
rect 31836 11396 31892 11406
rect 31892 11340 32004 11396
rect 31836 11302 31892 11340
rect 31724 10742 31780 10780
rect 31388 10546 31444 10556
rect 31500 10612 31556 10622
rect 31948 10612 32004 11340
rect 32060 10612 32116 10622
rect 31500 10610 31780 10612
rect 31500 10558 31502 10610
rect 31554 10558 31780 10610
rect 31500 10556 31780 10558
rect 31948 10556 32060 10612
rect 31500 10546 31556 10556
rect 31052 10498 31108 10510
rect 31052 10446 31054 10498
rect 31106 10446 31108 10498
rect 31052 10388 31108 10446
rect 31052 10322 31108 10332
rect 31724 10388 31780 10556
rect 31724 10322 31780 10332
rect 31836 10388 31892 10398
rect 31836 10386 32004 10388
rect 31836 10334 31838 10386
rect 31890 10334 32004 10386
rect 31836 10332 32004 10334
rect 31836 10322 31892 10332
rect 31948 10052 32004 10332
rect 30828 9986 30884 9996
rect 31500 9996 32004 10052
rect 31500 9938 31556 9996
rect 31500 9886 31502 9938
rect 31554 9886 31556 9938
rect 31500 9874 31556 9886
rect 30716 9734 30772 9772
rect 30828 8932 30884 8942
rect 30828 8930 31108 8932
rect 30828 8878 30830 8930
rect 30882 8878 31108 8930
rect 30828 8876 31108 8878
rect 30828 8818 30884 8876
rect 30828 8766 30830 8818
rect 30882 8766 30884 8818
rect 30828 8754 30884 8766
rect 30940 8260 30996 8270
rect 30492 8258 30996 8260
rect 30492 8206 30942 8258
rect 30994 8206 30996 8258
rect 30492 8204 30996 8206
rect 30940 8194 30996 8204
rect 30716 8036 30772 8046
rect 30716 7942 30772 7980
rect 31052 7924 31108 8876
rect 31276 8930 31332 8942
rect 31276 8878 31278 8930
rect 31330 8878 31332 8930
rect 31276 8484 31332 8878
rect 31276 8418 31332 8428
rect 31724 8930 31780 8942
rect 31724 8878 31726 8930
rect 31778 8878 31780 8930
rect 31612 8260 31668 8270
rect 31612 8166 31668 8204
rect 31052 7858 31108 7868
rect 31388 8034 31444 8046
rect 31388 7982 31390 8034
rect 31442 7982 31444 8034
rect 31388 7588 31444 7982
rect 31724 7588 31780 8878
rect 32060 7700 32116 10556
rect 32284 8820 32340 13580
rect 32284 8754 32340 8764
rect 32396 12068 32452 12078
rect 32396 10500 32452 12012
rect 32620 12068 32676 12078
rect 32620 12066 32788 12068
rect 32620 12014 32622 12066
rect 32674 12014 32788 12066
rect 32620 12012 32788 12014
rect 32620 12002 32676 12012
rect 32508 11620 32564 11630
rect 32508 11506 32564 11564
rect 32508 11454 32510 11506
rect 32562 11454 32564 11506
rect 32508 11442 32564 11454
rect 32508 10500 32564 10510
rect 32396 10498 32564 10500
rect 32396 10446 32510 10498
rect 32562 10446 32564 10498
rect 32396 10444 32564 10446
rect 32396 8484 32452 10444
rect 32508 10434 32564 10444
rect 32508 8930 32564 8942
rect 32508 8878 32510 8930
rect 32562 8878 32564 8930
rect 32508 8820 32564 8878
rect 32508 8754 32564 8764
rect 32508 8484 32564 8494
rect 32396 8428 32508 8484
rect 32508 8418 32564 8428
rect 32172 8036 32228 8046
rect 32620 8036 32676 8046
rect 32172 8034 32340 8036
rect 32172 7982 32174 8034
rect 32226 7982 32340 8034
rect 32172 7980 32340 7982
rect 32172 7970 32228 7980
rect 32172 7700 32228 7710
rect 31388 7522 31444 7532
rect 31500 7532 31780 7588
rect 31948 7698 32228 7700
rect 31948 7646 32174 7698
rect 32226 7646 32228 7698
rect 31948 7644 32228 7646
rect 31276 7364 31332 7374
rect 30380 6962 30436 6972
rect 31052 7362 31332 7364
rect 31052 7310 31278 7362
rect 31330 7310 31332 7362
rect 31052 7308 31332 7310
rect 31052 6914 31108 7308
rect 31276 7298 31332 7308
rect 31052 6862 31054 6914
rect 31106 6862 31108 6914
rect 31052 6850 31108 6862
rect 30716 6804 30772 6814
rect 30380 6802 30772 6804
rect 30380 6750 30718 6802
rect 30770 6750 30772 6802
rect 30380 6748 30772 6750
rect 30380 6690 30436 6748
rect 30716 6738 30772 6748
rect 30380 6638 30382 6690
rect 30434 6638 30436 6690
rect 30380 6626 30436 6638
rect 29932 6524 30212 6580
rect 30156 6466 30212 6524
rect 30156 6414 30158 6466
rect 30210 6414 30212 6466
rect 30156 6402 30212 6414
rect 30268 6466 30324 6478
rect 30268 6414 30270 6466
rect 30322 6414 30324 6466
rect 30268 6244 30324 6414
rect 30828 6466 30884 6478
rect 30828 6414 30830 6466
rect 30882 6414 30884 6466
rect 30716 6356 30772 6366
rect 30828 6356 30884 6414
rect 30772 6300 30884 6356
rect 30716 6290 30772 6300
rect 31500 6244 31556 7532
rect 30044 6188 30324 6244
rect 31388 6188 31556 6244
rect 31612 7362 31668 7374
rect 31612 7310 31614 7362
rect 31666 7310 31668 7362
rect 29708 6132 29764 6142
rect 29596 6076 29708 6132
rect 28924 6018 28980 6076
rect 29484 6066 29540 6076
rect 29708 6066 29764 6076
rect 28924 5966 28926 6018
rect 28978 5966 28980 6018
rect 28924 5954 28980 5966
rect 26796 5908 26852 5918
rect 26796 5814 26852 5852
rect 27020 5906 27076 5918
rect 27020 5854 27022 5906
rect 27074 5854 27076 5906
rect 26684 5506 26740 5516
rect 26908 5796 26964 5806
rect 26012 5234 26404 5236
rect 26012 5182 26350 5234
rect 26402 5182 26404 5234
rect 26012 5180 26404 5182
rect 26012 4562 26068 5180
rect 26348 5170 26404 5180
rect 26796 5236 26852 5246
rect 26796 5142 26852 5180
rect 26684 5124 26740 5134
rect 26684 5030 26740 5068
rect 26908 5124 26964 5740
rect 27020 5572 27076 5854
rect 27580 5908 27636 5918
rect 27580 5814 27636 5852
rect 28028 5908 28084 5918
rect 27020 5506 27076 5516
rect 27244 5124 27300 5134
rect 26908 5122 27300 5124
rect 26908 5070 27246 5122
rect 27298 5070 27300 5122
rect 26908 5068 27300 5070
rect 26908 4788 26964 5068
rect 27244 5058 27300 5068
rect 27804 5124 27860 5134
rect 27804 5010 27860 5068
rect 28028 5122 28084 5852
rect 28588 5908 28644 5918
rect 28588 5814 28644 5852
rect 29372 5906 29428 5918
rect 29372 5854 29374 5906
rect 29426 5854 29428 5906
rect 28140 5794 28196 5806
rect 28140 5742 28142 5794
rect 28194 5742 28196 5794
rect 28140 5348 28196 5742
rect 29372 5796 29428 5854
rect 29596 5908 29652 5918
rect 29596 5906 29764 5908
rect 29596 5854 29598 5906
rect 29650 5854 29764 5906
rect 29596 5852 29764 5854
rect 29596 5842 29652 5852
rect 29372 5730 29428 5740
rect 29036 5682 29092 5694
rect 29036 5630 29038 5682
rect 29090 5630 29092 5682
rect 29036 5460 29092 5630
rect 29260 5684 29316 5694
rect 29148 5460 29204 5470
rect 29036 5404 29148 5460
rect 29148 5394 29204 5404
rect 28140 5282 28196 5292
rect 28588 5236 28644 5246
rect 29148 5236 29204 5246
rect 28588 5234 29204 5236
rect 28588 5182 28590 5234
rect 28642 5182 29150 5234
rect 29202 5182 29204 5234
rect 28588 5180 29204 5182
rect 28588 5170 28644 5180
rect 29148 5170 29204 5180
rect 28028 5070 28030 5122
rect 28082 5070 28084 5122
rect 28028 5058 28084 5070
rect 29260 5122 29316 5628
rect 29260 5070 29262 5122
rect 29314 5070 29316 5122
rect 29260 5058 29316 5070
rect 29484 5124 29540 5134
rect 29484 5030 29540 5068
rect 27804 4958 27806 5010
rect 27858 4958 27860 5010
rect 27804 4946 27860 4958
rect 29708 5010 29764 5852
rect 30044 5906 30100 6188
rect 30380 6020 30436 6030
rect 30044 5854 30046 5906
rect 30098 5854 30100 5906
rect 30044 5842 30100 5854
rect 30268 6018 30436 6020
rect 30268 5966 30382 6018
rect 30434 5966 30436 6018
rect 30268 5964 30436 5966
rect 29708 4958 29710 5010
rect 29762 4958 29764 5010
rect 28476 4900 28532 4910
rect 26012 4510 26014 4562
rect 26066 4510 26068 4562
rect 26012 4498 26068 4510
rect 26796 4732 26964 4788
rect 28252 4898 28532 4900
rect 28252 4846 28478 4898
rect 28530 4846 28532 4898
rect 28252 4844 28532 4846
rect 26796 4338 26852 4732
rect 28252 4564 28308 4844
rect 28476 4834 28532 4844
rect 27468 4508 28308 4564
rect 27468 4450 27524 4508
rect 27468 4398 27470 4450
rect 27522 4398 27524 4450
rect 27468 4386 27524 4398
rect 26796 4286 26798 4338
rect 26850 4286 26852 4338
rect 26796 4274 26852 4286
rect 29596 4228 29652 4238
rect 29708 4228 29764 4958
rect 29820 5460 29876 5470
rect 29820 4340 29876 5404
rect 30268 5124 30324 5964
rect 30380 5954 30436 5964
rect 31164 6020 31220 6030
rect 31164 5926 31220 5964
rect 31388 6020 31444 6188
rect 31388 5954 31444 5964
rect 31500 6018 31556 6030
rect 31500 5966 31502 6018
rect 31554 5966 31556 6018
rect 30492 5908 30548 5918
rect 30492 5906 30660 5908
rect 30492 5854 30494 5906
rect 30546 5854 30660 5906
rect 30492 5852 30660 5854
rect 30492 5842 30548 5852
rect 30380 5684 30436 5694
rect 30380 5590 30436 5628
rect 30604 5124 30660 5852
rect 31052 5124 31108 5134
rect 31500 5124 31556 5966
rect 30268 5068 30436 5124
rect 30380 5012 30436 5068
rect 30604 5122 31556 5124
rect 30604 5070 30606 5122
rect 30658 5070 31054 5122
rect 31106 5070 31556 5122
rect 30604 5068 31556 5070
rect 31612 5124 31668 7310
rect 31724 7250 31780 7262
rect 31724 7198 31726 7250
rect 31778 7198 31780 7250
rect 31724 6580 31780 7198
rect 31724 6514 31780 6524
rect 31836 6466 31892 6478
rect 31836 6414 31838 6466
rect 31890 6414 31892 6466
rect 31724 5796 31780 5806
rect 31836 5796 31892 6414
rect 31780 5740 31892 5796
rect 31724 5730 31780 5740
rect 30604 5058 30660 5068
rect 31052 5058 31108 5068
rect 30380 4946 30436 4956
rect 29932 4900 29988 4910
rect 30268 4900 30324 4910
rect 29932 4898 30324 4900
rect 29932 4846 29934 4898
rect 29986 4846 30270 4898
rect 30322 4846 30324 4898
rect 29932 4844 30324 4846
rect 29932 4834 29988 4844
rect 30268 4564 30324 4844
rect 30268 4498 30324 4508
rect 29932 4340 29988 4350
rect 29820 4338 29988 4340
rect 29820 4286 29934 4338
rect 29986 4286 29988 4338
rect 29820 4284 29988 4286
rect 29932 4274 29988 4284
rect 29596 4226 29764 4228
rect 29596 4174 29598 4226
rect 29650 4174 29764 4226
rect 29596 4172 29764 4174
rect 29596 4162 29652 4172
rect 30940 4114 30996 4126
rect 30940 4062 30942 4114
rect 30994 4062 30996 4114
rect 29596 3780 29652 3790
rect 25900 3490 25956 3500
rect 26236 3668 26292 3678
rect 24892 3390 24894 3442
rect 24946 3390 24948 3442
rect 24892 3378 24948 3390
rect 24780 3052 24948 3108
rect 24892 800 24948 3052
rect 26236 800 26292 3612
rect 29372 3668 29428 3678
rect 29372 3574 29428 3612
rect 28588 3556 28644 3566
rect 28588 3462 28644 3500
rect 26908 3442 26964 3454
rect 26908 3390 26910 3442
rect 26962 3390 26964 3442
rect 26908 800 26964 3390
rect 29596 800 29652 3724
rect 30940 3780 30996 4062
rect 30940 3714 30996 3724
rect 30268 3556 30324 3566
rect 31164 3556 31220 5068
rect 31612 5058 31668 5068
rect 31836 5572 31892 5582
rect 31276 4900 31332 4910
rect 31276 4806 31332 4844
rect 31836 4900 31892 5516
rect 31948 5122 32004 7644
rect 32172 7634 32228 7644
rect 32284 7364 32340 7980
rect 32620 7942 32676 7980
rect 32732 7924 32788 12012
rect 33180 10836 33236 14140
rect 33292 12516 33348 14364
rect 33404 13748 33460 13758
rect 33404 13654 33460 13692
rect 33292 12450 33348 12460
rect 33292 12068 33348 12078
rect 33292 11974 33348 12012
rect 33180 10780 33348 10836
rect 33180 10612 33236 10622
rect 33180 10518 33236 10556
rect 33292 9380 33348 10780
rect 33628 10164 33684 17052
rect 33852 16772 33908 17390
rect 33964 16996 34020 18956
rect 34076 18946 34132 18956
rect 34188 19124 34244 19134
rect 33964 16930 34020 16940
rect 34076 18338 34132 18350
rect 34076 18286 34078 18338
rect 34130 18286 34132 18338
rect 33852 16706 33908 16716
rect 33852 16324 33908 16334
rect 33852 16210 33908 16268
rect 33852 16158 33854 16210
rect 33906 16158 33908 16210
rect 33852 15540 33908 16158
rect 33852 15474 33908 15484
rect 34076 15148 34132 18286
rect 34188 17556 34244 19068
rect 34860 19124 34916 19134
rect 34860 19030 34916 19068
rect 34300 19010 34356 19022
rect 34300 18958 34302 19010
rect 34354 18958 34356 19010
rect 34300 18788 34356 18958
rect 34300 18722 34356 18732
rect 35308 18564 35364 19404
rect 35980 19348 36036 19358
rect 36092 19348 36148 19740
rect 35980 19346 36148 19348
rect 35980 19294 35982 19346
rect 36034 19294 36148 19346
rect 35980 19292 36148 19294
rect 35980 19282 36036 19292
rect 35420 19124 35476 19134
rect 35420 19030 35476 19068
rect 36764 19124 36820 21644
rect 37548 21606 37604 21644
rect 36428 19012 36484 19022
rect 36428 19010 36596 19012
rect 36428 18958 36430 19010
rect 36482 18958 36596 19010
rect 36428 18956 36596 18958
rect 36428 18946 36484 18956
rect 36428 18788 36484 18798
rect 35308 18450 35364 18508
rect 36204 18564 36260 18574
rect 36260 18508 36372 18564
rect 36204 18498 36260 18508
rect 35308 18398 35310 18450
rect 35362 18398 35364 18450
rect 35308 18386 35364 18398
rect 36092 18450 36148 18462
rect 36092 18398 36094 18450
rect 36146 18398 36148 18450
rect 36092 18116 36148 18398
rect 36204 18116 36260 18126
rect 35196 18060 35460 18070
rect 34412 18004 34468 18014
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35196 17994 35460 18004
rect 35980 18060 36204 18116
rect 34300 17556 34356 17566
rect 34188 17554 34356 17556
rect 34188 17502 34302 17554
rect 34354 17502 34356 17554
rect 34188 17500 34356 17502
rect 34300 17490 34356 17500
rect 34188 16882 34244 16894
rect 34188 16830 34190 16882
rect 34242 16830 34244 16882
rect 34188 16772 34244 16830
rect 34412 16882 34468 17948
rect 35196 17668 35252 17678
rect 35084 17666 35252 17668
rect 35084 17614 35198 17666
rect 35250 17614 35252 17666
rect 35084 17612 35252 17614
rect 34636 17442 34692 17454
rect 34636 17390 34638 17442
rect 34690 17390 34692 17442
rect 34636 17108 34692 17390
rect 34972 17444 35028 17454
rect 34972 17350 35028 17388
rect 34412 16830 34414 16882
rect 34466 16830 34468 16882
rect 34412 16818 34468 16830
rect 34524 17052 34636 17108
rect 34188 15876 34244 16716
rect 34300 16100 34356 16110
rect 34300 16006 34356 16044
rect 34524 15986 34580 17052
rect 34636 17042 34692 17052
rect 34972 16996 35028 17006
rect 34972 16902 35028 16940
rect 34860 16884 34916 16894
rect 34860 16322 34916 16828
rect 34860 16270 34862 16322
rect 34914 16270 34916 16322
rect 34860 16258 34916 16270
rect 34524 15934 34526 15986
rect 34578 15934 34580 15986
rect 34524 15922 34580 15934
rect 34860 16100 34916 16110
rect 35084 16100 35140 17612
rect 35196 17602 35252 17612
rect 35980 17666 36036 18060
rect 36204 18050 36260 18060
rect 36316 17780 36372 18508
rect 36428 18562 36484 18732
rect 36428 18510 36430 18562
rect 36482 18510 36484 18562
rect 36428 18340 36484 18510
rect 36428 18274 36484 18284
rect 36428 17780 36484 17790
rect 36316 17778 36484 17780
rect 36316 17726 36430 17778
rect 36482 17726 36484 17778
rect 36316 17724 36484 17726
rect 36428 17714 36484 17724
rect 35980 17614 35982 17666
rect 36034 17614 36036 17666
rect 35980 17602 36036 17614
rect 35644 17556 35700 17566
rect 35644 17462 35700 17500
rect 35532 17444 35588 17454
rect 35420 17108 35476 17118
rect 35420 17014 35476 17052
rect 35196 16492 35460 16502
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35196 16426 35460 16436
rect 35196 16100 35252 16110
rect 35084 16044 35196 16100
rect 34188 15810 34244 15820
rect 34412 15652 34468 15662
rect 33964 15092 34132 15148
rect 34300 15314 34356 15326
rect 34300 15262 34302 15314
rect 34354 15262 34356 15314
rect 33964 13972 34020 15092
rect 34300 14756 34356 15262
rect 34300 14690 34356 14700
rect 34412 14754 34468 15596
rect 34524 15540 34580 15550
rect 34524 15446 34580 15484
rect 34860 15538 34916 16044
rect 35196 16006 35252 16044
rect 35532 16098 35588 17388
rect 36540 17220 36596 18956
rect 36540 17154 36596 17164
rect 36652 18452 36708 18462
rect 36540 16996 36596 17006
rect 36540 16902 36596 16940
rect 36204 16884 36260 16894
rect 35644 16882 36260 16884
rect 35644 16830 36206 16882
rect 36258 16830 36260 16882
rect 35644 16828 36260 16830
rect 35644 16210 35700 16828
rect 36204 16818 36260 16828
rect 35644 16158 35646 16210
rect 35698 16158 35700 16210
rect 35644 16146 35700 16158
rect 35532 16046 35534 16098
rect 35586 16046 35588 16098
rect 35532 16034 35588 16046
rect 36204 16098 36260 16110
rect 36204 16046 36206 16098
rect 36258 16046 36260 16098
rect 34972 15874 35028 15886
rect 34972 15822 34974 15874
rect 35026 15822 35028 15874
rect 34972 15652 35028 15822
rect 34972 15586 35028 15596
rect 35756 15874 35812 15886
rect 35756 15822 35758 15874
rect 35810 15822 35812 15874
rect 35756 15652 35812 15822
rect 35756 15586 35812 15596
rect 35868 15876 35924 15886
rect 34860 15486 34862 15538
rect 34914 15486 34916 15538
rect 34860 15474 34916 15486
rect 35868 15538 35924 15820
rect 35868 15486 35870 15538
rect 35922 15486 35924 15538
rect 35868 15474 35924 15486
rect 36204 15428 36260 16046
rect 36652 15538 36708 18396
rect 36652 15486 36654 15538
rect 36706 15486 36708 15538
rect 36652 15474 36708 15486
rect 36316 15428 36372 15438
rect 36204 15426 36372 15428
rect 36204 15374 36318 15426
rect 36370 15374 36372 15426
rect 36204 15372 36372 15374
rect 34412 14702 34414 14754
rect 34466 14702 34468 14754
rect 34412 14690 34468 14702
rect 35084 15314 35140 15326
rect 35084 15262 35086 15314
rect 35138 15262 35140 15314
rect 35084 14756 35140 15262
rect 35532 15314 35588 15326
rect 35532 15262 35534 15314
rect 35586 15262 35588 15314
rect 35532 15148 35588 15262
rect 36092 15316 36148 15326
rect 36092 15148 36148 15260
rect 35532 15092 35924 15148
rect 36092 15092 36260 15148
rect 35196 14924 35460 14934
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35196 14858 35460 14868
rect 35644 14868 35700 14878
rect 35084 14700 35364 14756
rect 35308 14642 35364 14700
rect 35308 14590 35310 14642
rect 35362 14590 35364 14642
rect 34300 14418 34356 14430
rect 34300 14366 34302 14418
rect 34354 14366 34356 14418
rect 34300 13972 34356 14366
rect 34636 14308 34692 14318
rect 33964 13916 34244 13972
rect 33964 13748 34020 13758
rect 33740 13692 33964 13748
rect 33740 13074 33796 13692
rect 33964 13654 34020 13692
rect 33740 13022 33742 13074
rect 33794 13022 33796 13074
rect 33740 13010 33796 13022
rect 34188 13074 34244 13916
rect 34300 13916 34580 13972
rect 34300 13748 34356 13916
rect 34300 13682 34356 13692
rect 34412 13746 34468 13758
rect 34412 13694 34414 13746
rect 34466 13694 34468 13746
rect 34188 13022 34190 13074
rect 34242 13022 34244 13074
rect 33740 12068 33796 12078
rect 33740 11974 33796 12012
rect 34188 11956 34244 13022
rect 34412 12852 34468 13694
rect 34524 13074 34580 13916
rect 34524 13022 34526 13074
rect 34578 13022 34580 13074
rect 34524 13010 34580 13022
rect 34636 13524 34692 14252
rect 34860 13748 34916 13758
rect 35308 13748 35364 14590
rect 35644 14530 35700 14812
rect 35644 14478 35646 14530
rect 35698 14478 35700 14530
rect 35644 13972 35700 14478
rect 35644 13906 35700 13916
rect 35756 14756 35812 14766
rect 35420 13748 35476 13758
rect 34860 13746 35700 13748
rect 34860 13694 34862 13746
rect 34914 13694 35422 13746
rect 35474 13694 35700 13746
rect 34860 13692 35700 13694
rect 34860 13682 34916 13692
rect 35420 13682 35476 13692
rect 34468 12796 34580 12852
rect 34412 12786 34468 12796
rect 34076 11954 34244 11956
rect 34076 11902 34190 11954
rect 34242 11902 34244 11954
rect 34076 11900 34244 11902
rect 33852 11172 33908 11182
rect 33852 10722 33908 11116
rect 33852 10670 33854 10722
rect 33906 10670 33908 10722
rect 33852 10658 33908 10670
rect 33292 9266 33348 9324
rect 33292 9214 33294 9266
rect 33346 9214 33348 9266
rect 33292 9202 33348 9214
rect 33516 10108 33684 10164
rect 34076 10612 34132 11900
rect 34188 11890 34244 11900
rect 34300 12066 34356 12078
rect 34300 12014 34302 12066
rect 34354 12014 34356 12066
rect 33516 9154 33572 10108
rect 33740 10052 33796 10062
rect 33628 9996 33740 10052
rect 33628 9938 33684 9996
rect 33740 9986 33796 9996
rect 33628 9886 33630 9938
rect 33682 9886 33684 9938
rect 33628 9874 33684 9886
rect 34076 9940 34132 10556
rect 34300 10052 34356 12014
rect 34524 11508 34580 12796
rect 34636 12402 34692 13468
rect 35196 13356 35460 13366
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35196 13290 35460 13300
rect 35420 13188 35476 13198
rect 35420 13094 35476 13132
rect 34636 12350 34638 12402
rect 34690 12350 34692 12402
rect 34636 12338 34692 12350
rect 34748 12962 34804 12974
rect 34748 12910 34750 12962
rect 34802 12910 34804 12962
rect 34748 12180 34804 12910
rect 34972 12962 35028 12974
rect 34972 12910 34974 12962
rect 35026 12910 35028 12962
rect 34972 12852 35028 12910
rect 35644 12962 35700 13692
rect 35756 13524 35812 14700
rect 35868 14306 35924 15092
rect 35868 14254 35870 14306
rect 35922 14254 35924 14306
rect 35868 13746 35924 14254
rect 35868 13694 35870 13746
rect 35922 13694 35924 13746
rect 35868 13682 35924 13694
rect 35980 14530 36036 14542
rect 35980 14478 35982 14530
rect 36034 14478 36036 14530
rect 35868 13524 35924 13534
rect 35756 13468 35868 13524
rect 35868 13430 35924 13468
rect 35644 12910 35646 12962
rect 35698 12910 35700 12962
rect 35644 12898 35700 12910
rect 35980 13412 36036 14478
rect 34972 12786 35028 12796
rect 35980 12290 36036 13356
rect 36092 13972 36148 13982
rect 36092 12962 36148 13916
rect 36092 12910 36094 12962
rect 36146 12910 36148 12962
rect 36092 12898 36148 12910
rect 35980 12238 35982 12290
rect 36034 12238 36036 12290
rect 35980 12226 36036 12238
rect 34748 12114 34804 12124
rect 35532 12180 35588 12190
rect 35084 12068 35140 12078
rect 35084 11974 35140 12012
rect 34972 11954 35028 11966
rect 34972 11902 34974 11954
rect 35026 11902 35028 11954
rect 34972 11788 35028 11902
rect 35196 11788 35460 11798
rect 34972 11732 35140 11788
rect 34636 11508 34692 11518
rect 34524 11506 34692 11508
rect 34524 11454 34638 11506
rect 34690 11454 34692 11506
rect 34524 11452 34692 11454
rect 34636 11442 34692 11452
rect 35084 11508 35140 11732
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35196 11722 35460 11732
rect 35084 11414 35140 11452
rect 35532 11172 35588 12124
rect 35532 11106 35588 11116
rect 35644 11956 35700 11966
rect 35196 10220 35460 10230
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35196 10154 35460 10164
rect 35532 10052 35588 10062
rect 35644 10052 35700 11900
rect 36204 11732 36260 15092
rect 36316 14532 36372 15372
rect 36540 15314 36596 15326
rect 36540 15262 36542 15314
rect 36594 15262 36596 15314
rect 36540 14868 36596 15262
rect 36540 14802 36596 14812
rect 36316 14466 36372 14476
rect 36428 13748 36484 13758
rect 36428 13074 36484 13692
rect 36428 13022 36430 13074
rect 36482 13022 36484 13074
rect 36204 11666 36260 11676
rect 36316 12068 36372 12078
rect 36204 11508 36260 11518
rect 36204 11414 36260 11452
rect 35868 11170 35924 11182
rect 35868 11118 35870 11170
rect 35922 11118 35924 11170
rect 35868 10276 35924 11118
rect 35980 11172 36036 11182
rect 35980 10498 36036 11116
rect 36316 10610 36372 12012
rect 36316 10558 36318 10610
rect 36370 10558 36372 10610
rect 36316 10546 36372 10558
rect 35980 10446 35982 10498
rect 36034 10446 36036 10498
rect 35980 10434 36036 10446
rect 35868 10210 35924 10220
rect 34300 9996 34580 10052
rect 34076 9938 34468 9940
rect 34076 9886 34078 9938
rect 34130 9886 34468 9938
rect 34076 9884 34468 9886
rect 34076 9874 34132 9884
rect 34300 9268 34356 9278
rect 34300 9174 34356 9212
rect 33516 9102 33518 9154
rect 33570 9102 33572 9154
rect 33516 9090 33572 9102
rect 33180 8818 33236 8830
rect 33180 8766 33182 8818
rect 33234 8766 33236 8818
rect 33180 8258 33236 8766
rect 33964 8372 34020 8382
rect 33964 8278 34020 8316
rect 34412 8370 34468 9884
rect 34412 8318 34414 8370
rect 34466 8318 34468 8370
rect 34412 8306 34468 8318
rect 34524 8932 34580 9996
rect 35532 10050 35700 10052
rect 35532 9998 35534 10050
rect 35586 9998 35700 10050
rect 35532 9996 35700 9998
rect 36092 10052 36148 10062
rect 35532 9986 35588 9996
rect 34636 9716 34692 9726
rect 34636 9266 34692 9660
rect 36092 9716 36148 9996
rect 36316 9828 36372 9838
rect 36428 9828 36484 13022
rect 36764 13076 36820 19068
rect 36876 21476 36932 21486
rect 36876 16994 36932 21420
rect 36988 21474 37044 21486
rect 36988 21422 36990 21474
rect 37042 21422 37044 21474
rect 36988 20692 37044 21422
rect 37660 21476 37716 23548
rect 38444 23492 38500 23502
rect 37884 23380 37940 23390
rect 37884 22372 37940 23324
rect 38444 23154 38500 23436
rect 38892 23380 38948 23548
rect 39004 23380 39060 23390
rect 38892 23378 39060 23380
rect 38892 23326 39006 23378
rect 39058 23326 39060 23378
rect 38892 23324 39060 23326
rect 39004 23314 39060 23324
rect 39340 23380 39396 24220
rect 39676 23940 39732 24446
rect 39900 23940 39956 23950
rect 39676 23938 39956 23940
rect 39676 23886 39902 23938
rect 39954 23886 39956 23938
rect 39676 23884 39956 23886
rect 39340 23378 39732 23380
rect 39340 23326 39342 23378
rect 39394 23326 39732 23378
rect 39340 23324 39732 23326
rect 39340 23314 39396 23324
rect 38444 23102 38446 23154
rect 38498 23102 38500 23154
rect 38444 23090 38500 23102
rect 38668 23266 38724 23278
rect 38668 23214 38670 23266
rect 38722 23214 38724 23266
rect 37996 23044 38052 23054
rect 37996 22950 38052 22988
rect 37884 21586 37940 22316
rect 38108 22148 38164 22158
rect 38108 22054 38164 22092
rect 38444 22148 38500 22158
rect 38668 22148 38724 23214
rect 39676 23266 39732 23324
rect 39676 23214 39678 23266
rect 39730 23214 39732 23266
rect 39676 22932 39732 23214
rect 39676 22866 39732 22876
rect 39788 23042 39844 23054
rect 39788 22990 39790 23042
rect 39842 22990 39844 23042
rect 39788 22596 39844 22990
rect 39900 23044 39956 23884
rect 40012 23828 40068 24556
rect 40236 24610 40292 24622
rect 40236 24558 40238 24610
rect 40290 24558 40292 24610
rect 40236 24498 40292 24558
rect 40236 24446 40238 24498
rect 40290 24446 40292 24498
rect 40236 24434 40292 24446
rect 40348 24500 40404 24510
rect 40012 23734 40068 23772
rect 39900 22978 39956 22988
rect 40012 23380 40068 23390
rect 40012 23154 40068 23324
rect 40012 23102 40014 23154
rect 40066 23102 40068 23154
rect 39340 22540 39844 22596
rect 38780 22428 39284 22484
rect 38780 22370 38836 22428
rect 38780 22318 38782 22370
rect 38834 22318 38836 22370
rect 38780 22306 38836 22318
rect 38892 22316 39172 22372
rect 38892 22148 38948 22316
rect 39116 22258 39172 22316
rect 39116 22206 39118 22258
rect 39170 22206 39172 22258
rect 39116 22194 39172 22206
rect 38668 22092 38948 22148
rect 38444 22054 38500 22092
rect 38892 22036 38948 22092
rect 38892 21970 38948 21980
rect 39004 22146 39060 22158
rect 39004 22094 39006 22146
rect 39058 22094 39060 22146
rect 39004 21924 39060 22094
rect 39004 21868 39172 21924
rect 39004 21700 39060 21710
rect 39004 21606 39060 21644
rect 37884 21534 37886 21586
rect 37938 21534 37940 21586
rect 37884 21522 37940 21534
rect 37660 21410 37716 21420
rect 37212 21362 37268 21374
rect 37212 21310 37214 21362
rect 37266 21310 37268 21362
rect 37212 21028 37268 21310
rect 37212 20962 37268 20972
rect 38332 21364 38388 21374
rect 37660 20916 37716 20926
rect 37660 20822 37716 20860
rect 38332 20802 38388 21308
rect 38332 20750 38334 20802
rect 38386 20750 38388 20802
rect 38332 20738 38388 20750
rect 38444 21028 38500 21038
rect 37212 20692 37268 20702
rect 36988 20690 37492 20692
rect 36988 20638 37214 20690
rect 37266 20638 37492 20690
rect 36988 20636 37492 20638
rect 37212 20626 37268 20636
rect 37436 19906 37492 20636
rect 37436 19854 37438 19906
rect 37490 19854 37492 19906
rect 37436 19842 37492 19854
rect 37772 20018 37828 20030
rect 37772 19966 37774 20018
rect 37826 19966 37828 20018
rect 37548 19236 37604 19246
rect 37772 19236 37828 19966
rect 37548 19234 37828 19236
rect 37548 19182 37550 19234
rect 37602 19182 37828 19234
rect 37548 19180 37828 19182
rect 37212 19012 37268 19022
rect 37548 19012 37604 19180
rect 37212 19010 37604 19012
rect 37212 18958 37214 19010
rect 37266 18958 37604 19010
rect 37212 18956 37604 18958
rect 37212 18564 37268 18956
rect 37212 18498 37268 18508
rect 37660 18900 37716 18910
rect 37100 18452 37156 18490
rect 37100 18386 37156 18396
rect 37548 18340 37604 18350
rect 37660 18340 37716 18844
rect 37548 18338 37716 18340
rect 37548 18286 37550 18338
rect 37602 18286 37716 18338
rect 37548 18284 37716 18286
rect 37548 18274 37604 18284
rect 37100 18226 37156 18238
rect 37100 18174 37102 18226
rect 37154 18174 37156 18226
rect 37100 17666 37156 18174
rect 37100 17614 37102 17666
rect 37154 17614 37156 17666
rect 37100 17602 37156 17614
rect 37324 18116 37380 18126
rect 36876 16942 36878 16994
rect 36930 16942 36932 16994
rect 36876 16930 36932 16942
rect 37212 16882 37268 16894
rect 37212 16830 37214 16882
rect 37266 16830 37268 16882
rect 37212 16324 37268 16830
rect 37212 16258 37268 16268
rect 37212 16100 37268 16110
rect 37212 16006 37268 16044
rect 37324 15540 37380 18060
rect 37324 15474 37380 15484
rect 37548 17220 37604 17230
rect 37548 16548 37604 17164
rect 37548 15426 37604 16492
rect 37660 16322 37716 18284
rect 37884 18450 37940 18462
rect 37884 18398 37886 18450
rect 37938 18398 37940 18450
rect 37884 17220 37940 18398
rect 38444 18450 38500 20972
rect 39116 20914 39172 21868
rect 39228 21810 39284 22428
rect 39340 22370 39396 22540
rect 39340 22318 39342 22370
rect 39394 22318 39396 22370
rect 39340 22306 39396 22318
rect 39900 22370 39956 22382
rect 39900 22318 39902 22370
rect 39954 22318 39956 22370
rect 39564 22260 39620 22270
rect 39564 22036 39620 22204
rect 39788 22260 39844 22270
rect 39788 22166 39844 22204
rect 39900 22036 39956 22318
rect 40012 22372 40068 23102
rect 40012 22306 40068 22316
rect 40124 23268 40180 23278
rect 39564 21980 39956 22036
rect 39228 21758 39230 21810
rect 39282 21758 39284 21810
rect 39228 21746 39284 21758
rect 39116 20862 39118 20914
rect 39170 20862 39172 20914
rect 39116 20850 39172 20862
rect 39228 21586 39284 21598
rect 39228 21534 39230 21586
rect 39282 21534 39284 21586
rect 38444 18398 38446 18450
rect 38498 18398 38500 18450
rect 38444 18228 38500 18398
rect 38444 18162 38500 18172
rect 38668 20468 38724 20478
rect 38668 17890 38724 20412
rect 39004 20132 39060 20142
rect 39004 18674 39060 20076
rect 39228 19908 39284 21534
rect 39228 19842 39284 19852
rect 39900 21586 39956 21980
rect 39900 21534 39902 21586
rect 39954 21534 39956 21586
rect 39900 19796 39956 21534
rect 40012 21924 40068 21934
rect 40012 21698 40068 21868
rect 40012 21646 40014 21698
rect 40066 21646 40068 21698
rect 40012 20804 40068 21646
rect 40012 20738 40068 20748
rect 39900 19730 39956 19740
rect 40012 20020 40068 20030
rect 39900 19348 39956 19358
rect 39900 19254 39956 19292
rect 39004 18622 39006 18674
rect 39058 18622 39060 18674
rect 39004 18610 39060 18622
rect 38668 17838 38670 17890
rect 38722 17838 38724 17890
rect 38668 17826 38724 17838
rect 39452 18450 39508 18462
rect 39676 18452 39732 18462
rect 39452 18398 39454 18450
rect 39506 18398 39508 18450
rect 37884 17154 37940 17164
rect 38220 17666 38276 17678
rect 38220 17614 38222 17666
rect 38274 17614 38276 17666
rect 38220 16996 38276 17614
rect 39228 17666 39284 17678
rect 39228 17614 39230 17666
rect 39282 17614 39284 17666
rect 39228 17556 39284 17614
rect 39228 17490 39284 17500
rect 38220 16930 38276 16940
rect 38444 17444 38500 17454
rect 37660 16270 37662 16322
rect 37714 16270 37716 16322
rect 37660 16258 37716 16270
rect 37772 16882 37828 16894
rect 37772 16830 37774 16882
rect 37826 16830 37828 16882
rect 37772 16772 37828 16830
rect 38108 16772 38164 16782
rect 37772 16770 38164 16772
rect 37772 16718 38110 16770
rect 38162 16718 38164 16770
rect 37772 16716 38164 16718
rect 37660 16100 37716 16110
rect 37772 16100 37828 16716
rect 38108 16706 38164 16716
rect 38220 16770 38276 16782
rect 38220 16718 38222 16770
rect 38274 16718 38276 16770
rect 38108 16324 38164 16334
rect 37660 16098 37828 16100
rect 37660 16046 37662 16098
rect 37714 16046 37828 16098
rect 37660 16044 37828 16046
rect 37996 16268 38108 16324
rect 37996 16098 38052 16268
rect 38108 16258 38164 16268
rect 38220 16100 38276 16718
rect 37996 16046 37998 16098
rect 38050 16046 38052 16098
rect 37660 16034 37716 16044
rect 37996 16034 38052 16046
rect 38108 16044 38276 16100
rect 37996 15652 38052 15662
rect 37772 15540 37828 15550
rect 37772 15446 37828 15484
rect 37996 15538 38052 15596
rect 37996 15486 37998 15538
rect 38050 15486 38052 15538
rect 37996 15474 38052 15486
rect 37548 15374 37550 15426
rect 37602 15374 37604 15426
rect 37548 15362 37604 15374
rect 36876 15316 36932 15326
rect 38108 15316 38164 16044
rect 38332 15986 38388 15998
rect 38332 15934 38334 15986
rect 38386 15934 38388 15986
rect 38220 15876 38276 15886
rect 38220 15782 38276 15820
rect 38332 15540 38388 15934
rect 38444 15876 38500 17388
rect 38668 17332 38724 17342
rect 38668 17106 38724 17276
rect 38668 17054 38670 17106
rect 38722 17054 38724 17106
rect 38668 17042 38724 17054
rect 39004 16996 39060 17006
rect 38668 16324 38724 16334
rect 39004 16324 39060 16940
rect 39452 16996 39508 18398
rect 39564 18450 39732 18452
rect 39564 18398 39678 18450
rect 39730 18398 39732 18450
rect 39564 18396 39732 18398
rect 39564 17556 39620 18396
rect 39676 18386 39732 18396
rect 39900 18452 39956 18462
rect 40012 18452 40068 19964
rect 40124 19906 40180 23212
rect 40124 19854 40126 19906
rect 40178 19854 40180 19906
rect 40124 19842 40180 19854
rect 40348 18676 40404 24444
rect 40460 23938 40516 25452
rect 40460 23886 40462 23938
rect 40514 23886 40516 23938
rect 40460 23156 40516 23886
rect 40572 25396 40628 25406
rect 40572 23714 40628 25340
rect 40684 25394 40740 26852
rect 40908 26180 40964 26190
rect 40908 26086 40964 26124
rect 41132 26066 41188 26078
rect 41132 26014 41134 26066
rect 41186 26014 41188 26066
rect 40684 25342 40686 25394
rect 40738 25342 40740 25394
rect 40684 24724 40740 25342
rect 40796 25506 40852 25518
rect 40796 25454 40798 25506
rect 40850 25454 40852 25506
rect 40796 25284 40852 25454
rect 40796 25218 40852 25228
rect 41132 24724 41188 26014
rect 41244 25508 41300 27806
rect 42700 27858 42756 29372
rect 43484 29988 43540 29998
rect 43484 28980 43540 29932
rect 43372 28644 43428 28654
rect 43260 28530 43316 28542
rect 43260 28478 43262 28530
rect 43314 28478 43316 28530
rect 43260 28308 43316 28478
rect 43260 28242 43316 28252
rect 43372 27970 43428 28588
rect 43484 28530 43540 28924
rect 43484 28478 43486 28530
rect 43538 28478 43540 28530
rect 43484 28466 43540 28478
rect 43372 27918 43374 27970
rect 43426 27918 43428 27970
rect 43372 27906 43428 27918
rect 42700 27806 42702 27858
rect 42754 27806 42756 27858
rect 42700 27794 42756 27806
rect 43372 26852 43428 26862
rect 43260 26796 43372 26852
rect 41916 26180 41972 26190
rect 41916 26086 41972 26124
rect 43260 26180 43316 26796
rect 43372 26786 43428 26796
rect 41468 26068 41524 26078
rect 41244 25442 41300 25452
rect 41356 26066 41524 26068
rect 41356 26014 41470 26066
rect 41522 26014 41524 26066
rect 41356 26012 41524 26014
rect 41356 25394 41412 26012
rect 41468 26002 41524 26012
rect 41356 25342 41358 25394
rect 41410 25342 41412 25394
rect 41356 25330 41412 25342
rect 41692 25508 41748 25518
rect 40684 24668 40852 24724
rect 40684 24500 40740 24510
rect 40684 23826 40740 24444
rect 40684 23774 40686 23826
rect 40738 23774 40740 23826
rect 40684 23762 40740 23774
rect 40572 23662 40574 23714
rect 40626 23662 40628 23714
rect 40572 23650 40628 23662
rect 40796 23380 40852 24668
rect 41132 24658 41188 24668
rect 41020 24612 41076 24622
rect 41020 24518 41076 24556
rect 40796 23314 40852 23324
rect 41692 23938 41748 25452
rect 41804 25506 41860 25518
rect 41804 25454 41806 25506
rect 41858 25454 41860 25506
rect 41804 24836 41860 25454
rect 42364 25508 42420 25518
rect 42364 25414 42420 25452
rect 43036 25506 43092 25518
rect 43036 25454 43038 25506
rect 43090 25454 43092 25506
rect 43036 25396 43092 25454
rect 43036 25330 43092 25340
rect 43148 25284 43204 25294
rect 41804 24770 41860 24780
rect 42700 24836 42756 24846
rect 42476 24724 42532 24734
rect 42140 24500 42196 24510
rect 42140 24406 42196 24444
rect 41692 23886 41694 23938
rect 41746 23886 41748 23938
rect 41244 23156 41300 23166
rect 40460 23154 41412 23156
rect 40460 23102 41246 23154
rect 41298 23102 41412 23154
rect 40460 23100 41412 23102
rect 41244 23090 41300 23100
rect 40908 22932 40964 22942
rect 40908 22838 40964 22876
rect 41244 22932 41300 22942
rect 41244 22838 41300 22876
rect 40572 22372 40628 22382
rect 40628 22316 40740 22372
rect 40572 22278 40628 22316
rect 40684 22036 40740 22316
rect 40796 22260 40852 22270
rect 40796 22166 40852 22204
rect 40684 21980 40964 22036
rect 40908 21586 40964 21980
rect 41356 21812 41412 23100
rect 41692 22372 41748 23886
rect 41916 23828 41972 23838
rect 41804 23492 41860 23502
rect 41804 23378 41860 23436
rect 41804 23326 41806 23378
rect 41858 23326 41860 23378
rect 41804 23314 41860 23326
rect 41804 22372 41860 22382
rect 41692 22370 41860 22372
rect 41692 22318 41806 22370
rect 41858 22318 41860 22370
rect 41692 22316 41860 22318
rect 41804 22036 41860 22316
rect 41916 22148 41972 23772
rect 42364 23492 42420 23502
rect 42028 23266 42084 23278
rect 42028 23214 42030 23266
rect 42082 23214 42084 23266
rect 42028 23156 42084 23214
rect 42364 23266 42420 23436
rect 42364 23214 42366 23266
rect 42418 23214 42420 23266
rect 42364 23202 42420 23214
rect 42028 23090 42084 23100
rect 42476 22372 42532 24668
rect 42700 24722 42756 24780
rect 43148 24724 43204 25228
rect 43260 24946 43316 26124
rect 43596 25732 43652 30156
rect 43820 29314 43876 29326
rect 43820 29262 43822 29314
rect 43874 29262 43876 29314
rect 43820 28868 43876 29262
rect 43820 28774 43876 28812
rect 43932 27972 43988 34188
rect 44156 34150 44212 34188
rect 44268 34020 44324 35196
rect 45052 35028 45108 35644
rect 45836 35252 45892 37214
rect 47068 35700 47124 38670
rect 47852 37268 47908 38894
rect 48076 38668 48132 44156
rect 48188 43092 48244 45166
rect 48300 43764 48356 45612
rect 48300 43698 48356 43708
rect 48188 43026 48244 43036
rect 48188 42756 48244 42766
rect 48244 42700 48356 42756
rect 48188 42662 48244 42700
rect 48188 42420 48244 42430
rect 48188 42194 48244 42364
rect 48188 42142 48190 42194
rect 48242 42142 48244 42194
rect 48188 42130 48244 42142
rect 48188 39732 48244 39742
rect 48300 39732 48356 42700
rect 48188 39730 48356 39732
rect 48188 39678 48190 39730
rect 48242 39678 48356 39730
rect 48188 39676 48356 39678
rect 48188 39666 48244 39676
rect 48076 38612 48356 38668
rect 48188 38164 48244 38174
rect 48300 38164 48356 38612
rect 48188 38162 48356 38164
rect 48188 38110 48190 38162
rect 48242 38110 48356 38162
rect 48188 38108 48356 38110
rect 48188 38052 48244 38108
rect 48188 37986 48244 37996
rect 47852 37212 48132 37268
rect 47964 37042 48020 37054
rect 47964 36990 47966 37042
rect 48018 36990 48020 37042
rect 47068 35634 47124 35644
rect 47404 36370 47460 36382
rect 47404 36318 47406 36370
rect 47458 36318 47460 36370
rect 45836 35186 45892 35196
rect 44940 34804 44996 34814
rect 44940 34710 44996 34748
rect 44604 34692 44660 34702
rect 44604 34130 44660 34636
rect 44604 34078 44606 34130
rect 44658 34078 44660 34130
rect 44604 34066 44660 34078
rect 44268 33954 44324 33964
rect 45052 33458 45108 34972
rect 45836 34916 45892 34926
rect 45724 34914 45892 34916
rect 45724 34862 45838 34914
rect 45890 34862 45892 34914
rect 45724 34860 45892 34862
rect 45164 34692 45220 34702
rect 45164 34354 45220 34636
rect 45164 34302 45166 34354
rect 45218 34302 45220 34354
rect 45164 34290 45220 34302
rect 45276 34690 45332 34702
rect 45276 34638 45278 34690
rect 45330 34638 45332 34690
rect 45052 33406 45054 33458
rect 45106 33406 45108 33458
rect 45052 33394 45108 33406
rect 45276 33460 45332 34638
rect 45276 33394 45332 33404
rect 45388 33346 45444 33358
rect 45388 33294 45390 33346
rect 45442 33294 45444 33346
rect 45052 32338 45108 32350
rect 45052 32286 45054 32338
rect 45106 32286 45108 32338
rect 45052 31948 45108 32286
rect 45388 31948 45444 33294
rect 45612 32564 45668 32574
rect 45612 32470 45668 32508
rect 45724 31948 45780 34860
rect 45836 34850 45892 34860
rect 47180 34802 47236 34814
rect 47180 34750 47182 34802
rect 47234 34750 47236 34802
rect 46284 33906 46340 33918
rect 46284 33854 46286 33906
rect 46338 33854 46340 33906
rect 46060 33460 46116 33470
rect 46060 33366 46116 33404
rect 45052 31892 45332 31948
rect 45388 31892 45556 31948
rect 45724 31892 45892 31948
rect 44156 31668 44212 31678
rect 44828 31668 44884 31678
rect 44156 31666 44884 31668
rect 44156 31614 44158 31666
rect 44210 31614 44830 31666
rect 44882 31614 44884 31666
rect 44156 31612 44884 31614
rect 44156 31602 44212 31612
rect 44828 31602 44884 31612
rect 45164 31556 45220 31566
rect 44940 31554 45220 31556
rect 44940 31502 45166 31554
rect 45218 31502 45220 31554
rect 44940 31500 45220 31502
rect 44940 31106 44996 31500
rect 45164 31490 45220 31500
rect 44940 31054 44942 31106
rect 44994 31054 44996 31106
rect 44940 31042 44996 31054
rect 45276 30996 45332 31892
rect 45500 30996 45556 31892
rect 45724 31778 45780 31790
rect 45724 31726 45726 31778
rect 45778 31726 45780 31778
rect 45612 30996 45668 31006
rect 45500 30994 45668 30996
rect 45500 30942 45614 30994
rect 45666 30942 45668 30994
rect 45500 30940 45668 30942
rect 45276 30930 45332 30940
rect 45388 30212 45444 30222
rect 45612 30212 45668 30940
rect 45444 30156 45668 30212
rect 45388 30118 45444 30156
rect 44044 29988 44100 29998
rect 44044 28532 44100 29932
rect 44940 29988 44996 29998
rect 44940 29894 44996 29932
rect 45724 29652 45780 31726
rect 45836 31780 45892 31892
rect 45836 31714 45892 31724
rect 46060 31106 46116 31118
rect 46060 31054 46062 31106
rect 46114 31054 46116 31106
rect 46060 30322 46116 31054
rect 46060 30270 46062 30322
rect 46114 30270 46116 30322
rect 46060 30258 46116 30270
rect 46284 30324 46340 33854
rect 47068 32338 47124 32350
rect 47068 32286 47070 32338
rect 47122 32286 47124 32338
rect 46396 30996 46452 31006
rect 46844 30996 46900 31006
rect 46396 30994 46900 30996
rect 46396 30942 46398 30994
rect 46450 30942 46846 30994
rect 46898 30942 46900 30994
rect 46396 30940 46900 30942
rect 46396 30930 46452 30940
rect 46844 30930 46900 30940
rect 46284 30258 46340 30268
rect 45500 29596 45780 29652
rect 46060 29764 46116 29774
rect 45276 29538 45332 29550
rect 45276 29486 45278 29538
rect 45330 29486 45332 29538
rect 45052 29428 45108 29438
rect 45052 29426 45220 29428
rect 45052 29374 45054 29426
rect 45106 29374 45220 29426
rect 45052 29372 45220 29374
rect 45052 29362 45108 29372
rect 44156 28756 44212 28766
rect 44156 28754 45108 28756
rect 44156 28702 44158 28754
rect 44210 28702 45108 28754
rect 44156 28700 45108 28702
rect 44156 28690 44212 28700
rect 45052 28642 45108 28700
rect 45052 28590 45054 28642
rect 45106 28590 45108 28642
rect 45052 28578 45108 28590
rect 44044 28476 44212 28532
rect 43932 26962 43988 27916
rect 43932 26910 43934 26962
rect 43986 26910 43988 26962
rect 43932 26898 43988 26910
rect 44044 26178 44100 26190
rect 44044 26126 44046 26178
rect 44098 26126 44100 26178
rect 43596 25676 43764 25732
rect 43372 25620 43428 25630
rect 43372 25282 43428 25564
rect 43596 25506 43652 25518
rect 43596 25454 43598 25506
rect 43650 25454 43652 25506
rect 43372 25230 43374 25282
rect 43426 25230 43428 25282
rect 43372 25218 43428 25230
rect 43484 25394 43540 25406
rect 43484 25342 43486 25394
rect 43538 25342 43540 25394
rect 43484 25284 43540 25342
rect 43484 25218 43540 25228
rect 43596 25060 43652 25454
rect 43260 24894 43262 24946
rect 43314 24894 43316 24946
rect 43260 24882 43316 24894
rect 43372 25004 43652 25060
rect 43708 25060 43764 25676
rect 44044 25620 44100 26126
rect 44044 25554 44100 25564
rect 42700 24670 42702 24722
rect 42754 24670 42756 24722
rect 42700 24658 42756 24670
rect 42924 24668 43204 24724
rect 42588 23938 42644 23950
rect 42924 23940 42980 24668
rect 43372 24610 43428 25004
rect 43708 24994 43764 25004
rect 43372 24558 43374 24610
rect 43426 24558 43428 24610
rect 43372 24546 43428 24558
rect 43820 24836 43876 24846
rect 43036 24498 43092 24510
rect 43036 24446 43038 24498
rect 43090 24446 43092 24498
rect 43036 24388 43092 24446
rect 43092 24332 43204 24388
rect 43036 24322 43092 24332
rect 42588 23886 42590 23938
rect 42642 23886 42644 23938
rect 42588 23828 42644 23886
rect 42588 23762 42644 23772
rect 42812 23938 42980 23940
rect 42812 23886 42926 23938
rect 42978 23886 42980 23938
rect 42812 23884 42980 23886
rect 42812 23156 42868 23884
rect 42924 23874 42980 23884
rect 43148 23828 43204 24332
rect 43708 24052 43764 24062
rect 43260 24050 43764 24052
rect 43260 23998 43710 24050
rect 43762 23998 43764 24050
rect 43260 23996 43764 23998
rect 43260 23938 43316 23996
rect 43708 23986 43764 23996
rect 43260 23886 43262 23938
rect 43314 23886 43316 23938
rect 43260 23874 43316 23886
rect 43148 23762 43204 23772
rect 43596 23828 43652 23838
rect 43596 23734 43652 23772
rect 43820 23826 43876 24780
rect 43820 23774 43822 23826
rect 43874 23774 43876 23826
rect 43820 23762 43876 23774
rect 44044 24276 44100 24286
rect 42924 23714 42980 23726
rect 42924 23662 42926 23714
rect 42978 23662 42980 23714
rect 42924 23492 42980 23662
rect 44044 23492 44100 24220
rect 42924 23436 43652 23492
rect 42812 23090 42868 23100
rect 42924 23268 42980 23278
rect 42924 23154 42980 23212
rect 43596 23266 43652 23436
rect 44044 23426 44100 23436
rect 43596 23214 43598 23266
rect 43650 23214 43652 23266
rect 43596 23202 43652 23214
rect 42924 23102 42926 23154
rect 42978 23102 42980 23154
rect 42924 23090 42980 23102
rect 43484 23156 43540 23166
rect 43148 22932 43204 22942
rect 42588 22372 42644 22382
rect 42476 22370 42644 22372
rect 42476 22318 42590 22370
rect 42642 22318 42644 22370
rect 42476 22316 42644 22318
rect 42252 22260 42308 22270
rect 42252 22166 42308 22204
rect 42028 22148 42084 22158
rect 41916 22146 42084 22148
rect 41916 22094 42030 22146
rect 42082 22094 42084 22146
rect 41916 22092 42084 22094
rect 42028 22082 42084 22092
rect 41804 21980 41972 22036
rect 41804 21812 41860 21822
rect 41356 21810 41860 21812
rect 41356 21758 41806 21810
rect 41858 21758 41860 21810
rect 41356 21756 41860 21758
rect 41804 21746 41860 21756
rect 40908 21534 40910 21586
rect 40962 21534 40964 21586
rect 40908 21522 40964 21534
rect 41356 21586 41412 21598
rect 41356 21534 41358 21586
rect 41410 21534 41412 21586
rect 41244 20916 41300 20926
rect 41356 20916 41412 21534
rect 41916 21252 41972 21980
rect 42140 21812 42196 21822
rect 42140 21718 42196 21756
rect 42476 21700 42532 22316
rect 42588 22306 42644 22316
rect 42812 22370 42868 22382
rect 42812 22318 42814 22370
rect 42866 22318 42868 22370
rect 42812 21812 42868 22318
rect 43148 22370 43204 22876
rect 43148 22318 43150 22370
rect 43202 22318 43204 22370
rect 43148 22306 43204 22318
rect 43484 22370 43540 23100
rect 43484 22318 43486 22370
rect 43538 22318 43540 22370
rect 43484 22036 43540 22318
rect 43708 22258 43764 22270
rect 43708 22206 43710 22258
rect 43762 22206 43764 22258
rect 43484 21970 43540 21980
rect 43596 22146 43652 22158
rect 43596 22094 43598 22146
rect 43650 22094 43652 22146
rect 42812 21746 42868 21756
rect 43260 21812 43316 21822
rect 41916 21186 41972 21196
rect 42364 21698 42532 21700
rect 42364 21646 42478 21698
rect 42530 21646 42532 21698
rect 42364 21644 42532 21646
rect 41244 20914 41412 20916
rect 41244 20862 41246 20914
rect 41298 20862 41412 20914
rect 41244 20860 41412 20862
rect 41244 20850 41300 20860
rect 41244 20132 41300 20142
rect 40908 20018 40964 20030
rect 40908 19966 40910 20018
rect 40962 19966 40964 20018
rect 40460 19012 40516 19022
rect 40460 19010 40628 19012
rect 40460 18958 40462 19010
rect 40514 18958 40628 19010
rect 40460 18956 40628 18958
rect 40460 18946 40516 18956
rect 39956 18396 40068 18452
rect 40236 18620 40404 18676
rect 40460 18676 40516 18686
rect 39900 18358 39956 18396
rect 40124 18338 40180 18350
rect 40124 18286 40126 18338
rect 40178 18286 40180 18338
rect 39564 17500 39732 17556
rect 39452 16930 39508 16940
rect 39116 16884 39172 16894
rect 39116 16770 39172 16828
rect 39228 16884 39284 16894
rect 39228 16882 39396 16884
rect 39228 16830 39230 16882
rect 39282 16830 39396 16882
rect 39228 16828 39396 16830
rect 39228 16818 39284 16828
rect 39116 16718 39118 16770
rect 39170 16718 39172 16770
rect 39116 16706 39172 16718
rect 39228 16324 39284 16334
rect 38668 16230 38724 16268
rect 38780 16322 39284 16324
rect 38780 16270 39230 16322
rect 39282 16270 39284 16322
rect 38780 16268 39284 16270
rect 38444 15810 38500 15820
rect 38332 15474 38388 15484
rect 36876 15222 36932 15260
rect 37996 15260 38164 15316
rect 37548 14532 37604 14542
rect 37212 14418 37268 14430
rect 37212 14366 37214 14418
rect 37266 14366 37268 14418
rect 37212 13858 37268 14366
rect 37548 14418 37604 14476
rect 37548 14366 37550 14418
rect 37602 14366 37604 14418
rect 37548 14354 37604 14366
rect 37884 14530 37940 14542
rect 37884 14478 37886 14530
rect 37938 14478 37940 14530
rect 37884 14420 37940 14478
rect 37884 14354 37940 14364
rect 37884 13972 37940 13982
rect 37996 13972 38052 15260
rect 38780 15202 38836 16268
rect 39228 16258 39284 16268
rect 38780 15150 38782 15202
rect 38834 15150 38836 15202
rect 38780 15138 38836 15150
rect 38892 15986 38948 15998
rect 38892 15934 38894 15986
rect 38946 15934 38948 15986
rect 38108 15090 38164 15102
rect 38108 15038 38110 15090
rect 38162 15038 38164 15090
rect 38108 14754 38164 15038
rect 38108 14702 38110 14754
rect 38162 14702 38164 14754
rect 38108 14690 38164 14702
rect 38444 14308 38500 14318
rect 38444 14214 38500 14252
rect 38780 14308 38836 14318
rect 38892 14308 38948 15934
rect 39116 15314 39172 15326
rect 39116 15262 39118 15314
rect 39170 15262 39172 15314
rect 39116 14980 39172 15262
rect 39004 14532 39060 14542
rect 39004 14438 39060 14476
rect 38780 14306 38948 14308
rect 38780 14254 38782 14306
rect 38834 14254 38948 14306
rect 38780 14252 38948 14254
rect 37940 13916 38052 13972
rect 37884 13878 37940 13916
rect 37212 13806 37214 13858
rect 37266 13806 37268 13858
rect 36876 13748 36932 13758
rect 36876 13654 36932 13692
rect 37212 13412 37268 13806
rect 38556 13748 38612 13758
rect 38556 13654 38612 13692
rect 37212 13346 37268 13356
rect 37660 13412 37716 13422
rect 36764 13010 36820 13020
rect 37660 12962 37716 13356
rect 37660 12910 37662 12962
rect 37714 12910 37716 12962
rect 37660 12898 37716 12910
rect 38780 12852 38836 14252
rect 39116 13972 39172 14924
rect 39340 14532 39396 16828
rect 39564 16882 39620 16894
rect 39564 16830 39566 16882
rect 39618 16830 39620 16882
rect 39564 16436 39620 16830
rect 39564 16370 39620 16380
rect 39452 16098 39508 16110
rect 39452 16046 39454 16098
rect 39506 16046 39508 16098
rect 39452 15428 39508 16046
rect 39564 15876 39620 15886
rect 39676 15876 39732 17500
rect 39900 16996 39956 17006
rect 39900 16660 39956 16940
rect 39900 16594 39956 16604
rect 40124 16212 40180 18286
rect 40236 17892 40292 18620
rect 40460 18582 40516 18620
rect 40348 18452 40404 18462
rect 40348 18358 40404 18396
rect 40572 18116 40628 18956
rect 40572 18050 40628 18060
rect 40236 17826 40292 17836
rect 40460 17778 40516 17790
rect 40460 17726 40462 17778
rect 40514 17726 40516 17778
rect 40348 17668 40404 17678
rect 40348 17574 40404 17612
rect 40460 17332 40516 17726
rect 40460 17266 40516 17276
rect 40572 17556 40628 17566
rect 40236 17220 40292 17230
rect 40236 17106 40292 17164
rect 40236 17054 40238 17106
rect 40290 17054 40292 17106
rect 40236 17042 40292 17054
rect 40124 16146 40180 16156
rect 40348 16324 40404 16334
rect 40348 16098 40404 16268
rect 40572 16212 40628 17500
rect 40908 17444 40964 19966
rect 41020 19908 41076 19918
rect 41020 19346 41076 19852
rect 41244 19684 41300 20076
rect 41356 20020 41412 20860
rect 42028 20916 42084 20926
rect 42028 20802 42084 20860
rect 42028 20750 42030 20802
rect 42082 20750 42084 20802
rect 42028 20738 42084 20750
rect 42140 20692 42196 20702
rect 42140 20242 42196 20636
rect 42140 20190 42142 20242
rect 42194 20190 42196 20242
rect 42140 20178 42196 20190
rect 41580 20020 41636 20030
rect 41356 20018 41636 20020
rect 41356 19966 41582 20018
rect 41634 19966 41636 20018
rect 41356 19964 41636 19966
rect 41580 19954 41636 19964
rect 41804 20020 41860 20030
rect 42364 20020 42420 21644
rect 42476 21634 42532 21644
rect 42812 21588 42868 21598
rect 42700 21586 42868 21588
rect 42700 21534 42814 21586
rect 42866 21534 42868 21586
rect 42700 21532 42868 21534
rect 41804 20018 42420 20020
rect 41804 19966 41806 20018
rect 41858 19966 42420 20018
rect 41804 19964 42420 19966
rect 42476 20020 42532 20030
rect 41804 19954 41860 19964
rect 42476 19926 42532 19964
rect 41244 19618 41300 19628
rect 42700 19684 42756 21532
rect 42812 21522 42868 21532
rect 43260 21474 43316 21756
rect 43596 21812 43652 22094
rect 43596 21746 43652 21756
rect 43708 21588 43764 22206
rect 43260 21422 43262 21474
rect 43314 21422 43316 21474
rect 43260 21410 43316 21422
rect 43596 21532 43764 21588
rect 44156 21588 44212 28476
rect 44828 28420 44884 28430
rect 44828 28326 44884 28364
rect 45164 28084 45220 29372
rect 45164 28018 45220 28028
rect 45276 27188 45332 29486
rect 45500 28308 45556 29596
rect 45612 29426 45668 29438
rect 45612 29374 45614 29426
rect 45666 29374 45668 29426
rect 45612 28868 45668 29374
rect 45612 28802 45668 28812
rect 45500 27746 45556 28252
rect 45500 27694 45502 27746
rect 45554 27694 45556 27746
rect 45500 27682 45556 27694
rect 45612 28642 45668 28654
rect 45612 28590 45614 28642
rect 45666 28590 45668 28642
rect 45612 27300 45668 28590
rect 46060 28084 46116 29708
rect 47068 29652 47124 32286
rect 47180 32004 47236 34750
rect 47404 33684 47460 36318
rect 47852 35700 47908 35710
rect 47852 35586 47908 35644
rect 47852 35534 47854 35586
rect 47906 35534 47908 35586
rect 47852 35522 47908 35534
rect 47964 34356 48020 36990
rect 47964 34290 48020 34300
rect 47404 33618 47460 33628
rect 47964 34130 48020 34142
rect 47964 34078 47966 34130
rect 48018 34078 48020 34130
rect 47180 31938 47236 31948
rect 47740 31890 47796 31902
rect 47740 31838 47742 31890
rect 47794 31838 47796 31890
rect 47404 31106 47460 31118
rect 47404 31054 47406 31106
rect 47458 31054 47460 31106
rect 47180 30772 47236 30782
rect 47180 30770 47348 30772
rect 47180 30718 47182 30770
rect 47234 30718 47348 30770
rect 47180 30716 47348 30718
rect 47180 30706 47236 30716
rect 47068 29586 47124 29596
rect 46060 28082 46564 28084
rect 46060 28030 46062 28082
rect 46114 28030 46564 28082
rect 46060 28028 46564 28030
rect 46060 28018 46116 28028
rect 45612 27234 45668 27244
rect 46508 27858 46564 28028
rect 46620 27972 46676 27982
rect 46620 27878 46676 27916
rect 46508 27806 46510 27858
rect 46562 27806 46564 27858
rect 45276 27122 45332 27132
rect 46060 27188 46116 27198
rect 46060 27094 46116 27132
rect 45388 27074 45444 27086
rect 45388 27022 45390 27074
rect 45442 27022 45444 27074
rect 44268 26852 44324 26862
rect 44268 26758 44324 26796
rect 44716 26292 44772 26302
rect 44716 26198 44772 26236
rect 45388 26292 45444 27022
rect 46508 26908 46564 27806
rect 47292 27860 47348 30716
rect 47404 29988 47460 31054
rect 47404 29922 47460 29932
rect 47740 28980 47796 31838
rect 47964 31106 48020 34078
rect 48076 33460 48132 37212
rect 48188 33460 48244 33470
rect 48076 33458 48244 33460
rect 48076 33406 48190 33458
rect 48242 33406 48244 33458
rect 48076 33404 48244 33406
rect 48188 32340 48244 33404
rect 48188 32274 48244 32284
rect 47964 31054 47966 31106
rect 48018 31054 48020 31106
rect 47964 30324 48020 31054
rect 48188 30324 48244 30334
rect 47964 30322 48244 30324
rect 47964 30270 48190 30322
rect 48242 30270 48244 30322
rect 47964 30268 48244 30270
rect 48188 30258 48244 30268
rect 47740 28914 47796 28924
rect 47964 29202 48020 29214
rect 47964 29150 47966 29202
rect 48018 29150 48020 29202
rect 47852 28754 47908 28766
rect 47852 28702 47854 28754
rect 47906 28702 47908 28754
rect 47628 28084 47684 28094
rect 47628 27990 47684 28028
rect 47852 28084 47908 28702
rect 47964 28308 48020 29150
rect 47964 28242 48020 28252
rect 47852 28018 47908 28028
rect 47292 27858 48244 27860
rect 47292 27806 47294 27858
rect 47346 27806 48244 27858
rect 47292 27804 48244 27806
rect 47292 27794 47348 27804
rect 48188 27186 48244 27804
rect 48188 27134 48190 27186
rect 48242 27134 48244 27186
rect 48188 27122 48244 27134
rect 46284 26852 46564 26908
rect 45388 25506 45444 26236
rect 45612 26290 45668 26302
rect 45612 26238 45614 26290
rect 45666 26238 45668 26290
rect 45612 25956 45668 26238
rect 45612 25890 45668 25900
rect 45388 25454 45390 25506
rect 45442 25454 45444 25506
rect 44604 25396 44660 25406
rect 44604 24946 44660 25340
rect 45276 25060 45332 25070
rect 44604 24894 44606 24946
rect 44658 24894 44660 24946
rect 44604 24882 44660 24894
rect 45164 24948 45220 24958
rect 44940 24836 44996 24846
rect 44940 24742 44996 24780
rect 44380 24722 44436 24734
rect 44380 24670 44382 24722
rect 44434 24670 44436 24722
rect 44380 23380 44436 24670
rect 44940 24052 44996 24062
rect 44940 23826 44996 23996
rect 45164 23940 45220 24892
rect 45276 24946 45332 25004
rect 45276 24894 45278 24946
rect 45330 24894 45332 24946
rect 45276 24882 45332 24894
rect 44940 23774 44942 23826
rect 44994 23774 44996 23826
rect 44940 23762 44996 23774
rect 45052 23938 45220 23940
rect 45052 23886 45166 23938
rect 45218 23886 45220 23938
rect 45052 23884 45220 23886
rect 44380 23314 44436 23324
rect 44380 22484 44436 22494
rect 44380 22390 44436 22428
rect 45052 22482 45108 23884
rect 45164 23874 45220 23884
rect 45052 22430 45054 22482
rect 45106 22430 45108 22482
rect 45052 22418 45108 22430
rect 45388 23268 45444 25454
rect 46060 25396 46116 25406
rect 46060 25302 46116 25340
rect 45724 24836 45780 24846
rect 45612 23940 45668 23950
rect 45612 23846 45668 23884
rect 45388 22370 45444 23212
rect 45724 23042 45780 24780
rect 45724 22990 45726 23042
rect 45778 22990 45780 23042
rect 45724 22978 45780 22990
rect 46284 22484 46340 26852
rect 47964 26066 48020 26078
rect 47964 26014 47966 26066
rect 48018 26014 48020 26066
rect 47964 25620 48020 26014
rect 47964 25554 48020 25564
rect 48188 25618 48244 25630
rect 48188 25566 48190 25618
rect 48242 25566 48244 25618
rect 47404 25060 47460 25070
rect 46956 24610 47012 24622
rect 46956 24558 46958 24610
rect 47010 24558 47012 24610
rect 46508 23380 46564 23390
rect 46508 23286 46564 23324
rect 46844 23268 46900 23278
rect 46844 23154 46900 23212
rect 46844 23102 46846 23154
rect 46898 23102 46900 23154
rect 46844 23090 46900 23102
rect 46956 22932 47012 24558
rect 47404 23716 47460 25004
rect 48076 24722 48132 24734
rect 48076 24670 48078 24722
rect 48130 24670 48132 24722
rect 46956 22866 47012 22876
rect 47068 23266 47124 23278
rect 47068 23214 47070 23266
rect 47122 23214 47124 23266
rect 46284 22418 46340 22428
rect 47068 22484 47124 23214
rect 47068 22418 47124 22428
rect 47180 23268 47236 23278
rect 45388 22318 45390 22370
rect 45442 22318 45444 22370
rect 43260 21252 43316 21262
rect 43148 20916 43204 20926
rect 42700 19618 42756 19628
rect 42812 20802 42868 20814
rect 42812 20750 42814 20802
rect 42866 20750 42868 20802
rect 42364 19460 42420 19470
rect 41020 19294 41022 19346
rect 41074 19294 41076 19346
rect 41020 19236 41076 19294
rect 42140 19458 42420 19460
rect 42140 19406 42366 19458
rect 42418 19406 42420 19458
rect 42140 19404 42420 19406
rect 41020 19170 41076 19180
rect 41692 19236 41748 19274
rect 41692 19170 41748 19180
rect 42028 19236 42084 19246
rect 42140 19236 42196 19404
rect 42364 19394 42420 19404
rect 42028 19234 42196 19236
rect 42028 19182 42030 19234
rect 42082 19182 42196 19234
rect 42028 19180 42196 19182
rect 42028 19170 42084 19180
rect 41356 19122 41412 19134
rect 41356 19070 41358 19122
rect 41410 19070 41412 19122
rect 41356 18676 41412 19070
rect 41692 19012 41748 19022
rect 41356 18610 41412 18620
rect 41468 19010 41748 19012
rect 41468 18958 41694 19010
rect 41746 18958 41748 19010
rect 41468 18956 41748 18958
rect 40908 17378 40964 17388
rect 41132 17220 41188 17230
rect 40796 16996 40852 17006
rect 40796 16772 40852 16940
rect 40908 16884 40964 16894
rect 40908 16790 40964 16828
rect 41132 16884 41188 17164
rect 41356 17108 41412 17118
rect 41356 17014 41412 17052
rect 41468 16884 41524 18956
rect 41692 18946 41748 18956
rect 41804 18452 41860 18462
rect 41804 18450 42084 18452
rect 41804 18398 41806 18450
rect 41858 18398 42084 18450
rect 41804 18396 42084 18398
rect 41804 18386 41860 18396
rect 42028 17780 42084 18396
rect 42140 18450 42196 19180
rect 42588 19236 42644 19246
rect 42812 19236 42868 20750
rect 42924 20692 42980 20702
rect 42924 20598 42980 20636
rect 43148 20244 43204 20860
rect 42924 20188 43204 20244
rect 42924 19346 42980 20188
rect 43036 20020 43092 20030
rect 43260 20020 43316 21196
rect 43596 20914 43652 21532
rect 43596 20862 43598 20914
rect 43650 20862 43652 20914
rect 43596 20850 43652 20862
rect 43708 20802 43764 20814
rect 43708 20750 43710 20802
rect 43762 20750 43764 20802
rect 43708 20356 43764 20750
rect 43596 20300 43764 20356
rect 43820 20690 43876 20702
rect 43820 20638 43822 20690
rect 43874 20638 43876 20690
rect 43596 20244 43652 20300
rect 43036 20018 43316 20020
rect 43036 19966 43038 20018
rect 43090 19966 43316 20018
rect 43036 19964 43316 19966
rect 43372 20188 43652 20244
rect 43036 19954 43092 19964
rect 42924 19294 42926 19346
rect 42978 19294 42980 19346
rect 42924 19282 42980 19294
rect 43372 19796 43428 20188
rect 43708 20132 43764 20142
rect 43708 20038 43764 20076
rect 43372 19346 43428 19740
rect 43372 19294 43374 19346
rect 43426 19294 43428 19346
rect 43372 19282 43428 19294
rect 43484 20018 43540 20030
rect 43484 19966 43486 20018
rect 43538 19966 43540 20018
rect 43484 19908 43540 19966
rect 43820 19908 43876 20638
rect 44156 20244 44212 21532
rect 45276 22260 45332 22270
rect 45052 21364 45108 21374
rect 45052 20802 45108 21308
rect 45052 20750 45054 20802
rect 45106 20750 45108 20802
rect 45052 20738 45108 20750
rect 45276 20690 45332 22204
rect 45388 22036 45444 22318
rect 46060 22260 46116 22298
rect 46060 22194 46116 22204
rect 45612 22148 45668 22158
rect 45444 21980 45556 22036
rect 45388 21970 45444 21980
rect 45388 21812 45444 21822
rect 45388 21698 45444 21756
rect 45388 21646 45390 21698
rect 45442 21646 45444 21698
rect 45388 21634 45444 21646
rect 45276 20638 45278 20690
rect 45330 20638 45332 20690
rect 45276 20626 45332 20638
rect 44156 20178 44212 20188
rect 45052 20244 45108 20254
rect 44380 20132 44436 20142
rect 44380 20130 44548 20132
rect 44380 20078 44382 20130
rect 44434 20078 44548 20130
rect 44380 20076 44548 20078
rect 44380 20066 44436 20076
rect 43484 19852 43876 19908
rect 44044 20018 44100 20030
rect 44044 19966 44046 20018
rect 44098 19966 44100 20018
rect 42644 19180 42868 19236
rect 42588 19170 42644 19180
rect 42252 19122 42308 19134
rect 42252 19070 42254 19122
rect 42306 19070 42308 19122
rect 42252 18564 42308 19070
rect 42364 19012 42420 19022
rect 42364 19010 42532 19012
rect 42364 18958 42366 19010
rect 42418 18958 42532 19010
rect 42364 18956 42532 18958
rect 42364 18946 42420 18956
rect 42476 18676 42532 18956
rect 42476 18610 42532 18620
rect 42700 18674 42756 19180
rect 42700 18622 42702 18674
rect 42754 18622 42756 18674
rect 42700 18610 42756 18622
rect 43484 18676 43540 19852
rect 43484 18610 43540 18620
rect 43708 19684 43764 19694
rect 44044 19684 44100 19966
rect 43764 19628 44100 19684
rect 43708 18674 43764 19628
rect 43708 18622 43710 18674
rect 43762 18622 43764 18674
rect 43708 18610 43764 18622
rect 43820 19346 43876 19358
rect 43820 19294 43822 19346
rect 43874 19294 43876 19346
rect 42252 18498 42308 18508
rect 42140 18398 42142 18450
rect 42194 18398 42196 18450
rect 42140 18386 42196 18398
rect 42588 18450 42644 18462
rect 42588 18398 42590 18450
rect 42642 18398 42644 18450
rect 42252 18340 42308 18350
rect 42588 18340 42644 18398
rect 43260 18452 43316 18462
rect 43484 18452 43540 18462
rect 43260 18358 43316 18396
rect 43372 18450 43540 18452
rect 43372 18398 43486 18450
rect 43538 18398 43540 18450
rect 43372 18396 43540 18398
rect 42252 18338 42644 18340
rect 42252 18286 42254 18338
rect 42306 18286 42644 18338
rect 42252 18284 42644 18286
rect 42252 18274 42308 18284
rect 41132 16790 41188 16828
rect 41244 16828 41524 16884
rect 41916 17666 41972 17678
rect 41916 17614 41918 17666
rect 41970 17614 41972 17666
rect 41916 16884 41972 17614
rect 42028 17666 42084 17724
rect 42028 17614 42030 17666
rect 42082 17614 42084 17666
rect 42028 17602 42084 17614
rect 42140 18228 42196 18238
rect 42140 17442 42196 18172
rect 42700 18228 42756 18238
rect 42700 18134 42756 18172
rect 42700 17780 42756 17790
rect 42700 17686 42756 17724
rect 42364 17556 42420 17566
rect 42364 17462 42420 17500
rect 42700 17556 42756 17566
rect 42140 17390 42142 17442
rect 42194 17390 42196 17442
rect 42140 17378 42196 17390
rect 40796 16706 40852 16716
rect 41020 16770 41076 16782
rect 41020 16718 41022 16770
rect 41074 16718 41076 16770
rect 40684 16660 40740 16670
rect 40684 16322 40740 16604
rect 40684 16270 40686 16322
rect 40738 16270 40740 16322
rect 40684 16258 40740 16270
rect 41020 16324 41076 16718
rect 41020 16258 41076 16268
rect 41244 16212 41300 16828
rect 41916 16818 41972 16828
rect 42700 16996 42756 17500
rect 42812 17554 42868 17566
rect 42812 17502 42814 17554
rect 42866 17502 42868 17554
rect 42812 17220 42868 17502
rect 42812 17154 42868 17164
rect 43260 17108 43316 17118
rect 43372 17108 43428 18396
rect 43484 18386 43540 18396
rect 43484 18228 43540 18238
rect 43484 17778 43540 18172
rect 43708 17892 43764 17902
rect 43484 17726 43486 17778
rect 43538 17726 43540 17778
rect 43484 17714 43540 17726
rect 43596 17836 43708 17892
rect 43596 17666 43652 17836
rect 43708 17826 43764 17836
rect 43596 17614 43598 17666
rect 43650 17614 43652 17666
rect 43596 17602 43652 17614
rect 43708 17668 43764 17678
rect 43316 17052 43428 17108
rect 43708 17108 43764 17612
rect 43820 17444 43876 19294
rect 44268 19012 44324 19022
rect 44268 18918 44324 18956
rect 43932 18450 43988 18462
rect 43932 18398 43934 18450
rect 43986 18398 43988 18450
rect 43932 17780 43988 18398
rect 44044 18340 44100 18350
rect 44380 18340 44436 18350
rect 44044 18338 44436 18340
rect 44044 18286 44046 18338
rect 44098 18286 44382 18338
rect 44434 18286 44436 18338
rect 44044 18284 44436 18286
rect 44044 18274 44100 18284
rect 44380 18274 44436 18284
rect 44380 18004 44436 18014
rect 44492 18004 44548 20076
rect 45052 20130 45108 20188
rect 45052 20078 45054 20130
rect 45106 20078 45108 20130
rect 45052 20066 45108 20078
rect 45388 20020 45444 20030
rect 45500 20020 45556 21980
rect 45612 20802 45668 22092
rect 46060 22036 46116 22046
rect 46060 21586 46116 21980
rect 46060 21534 46062 21586
rect 46114 21534 46116 21586
rect 46060 21522 46116 21534
rect 47180 21588 47236 23212
rect 47404 23266 47460 23660
rect 47964 24050 48020 24062
rect 47964 23998 47966 24050
rect 48018 23998 48020 24050
rect 47964 23604 48020 23998
rect 47964 23538 48020 23548
rect 47404 23214 47406 23266
rect 47458 23214 47460 23266
rect 47404 23202 47460 23214
rect 48076 22484 48132 24670
rect 48188 23268 48244 25566
rect 48188 23202 48244 23212
rect 48300 23716 48356 23726
rect 48188 23044 48244 23054
rect 48300 23044 48356 23660
rect 48188 23042 48356 23044
rect 48188 22990 48190 23042
rect 48242 22990 48356 23042
rect 48188 22988 48356 22990
rect 48188 22978 48244 22988
rect 48188 22484 48244 22494
rect 48076 22482 48244 22484
rect 48076 22430 48190 22482
rect 48242 22430 48244 22482
rect 48076 22428 48244 22430
rect 47964 22260 48020 22270
rect 47516 21698 47572 21710
rect 47516 21646 47518 21698
rect 47570 21646 47572 21698
rect 47292 21588 47348 21598
rect 47180 21586 47348 21588
rect 47180 21534 47294 21586
rect 47346 21534 47348 21586
rect 47180 21532 47348 21534
rect 47292 21522 47348 21532
rect 47516 21588 47572 21646
rect 47516 21522 47572 21532
rect 46956 21364 47012 21374
rect 46956 21270 47012 21308
rect 47964 21026 48020 22204
rect 48076 21698 48132 22428
rect 48188 22418 48244 22428
rect 48076 21646 48078 21698
rect 48130 21646 48132 21698
rect 48076 21634 48132 21646
rect 47964 20974 47966 21026
rect 48018 20974 48020 21026
rect 47964 20962 48020 20974
rect 48300 21588 48356 21598
rect 47516 20916 47572 20926
rect 45612 20750 45614 20802
rect 45666 20750 45668 20802
rect 45612 20738 45668 20750
rect 46620 20804 46676 20814
rect 45388 20018 45556 20020
rect 45388 19966 45390 20018
rect 45442 19966 45556 20018
rect 45388 19964 45556 19966
rect 45388 19954 45444 19964
rect 44940 19346 44996 19358
rect 44940 19294 44942 19346
rect 44994 19294 44996 19346
rect 44436 17948 44548 18004
rect 44716 19234 44772 19246
rect 44716 19182 44718 19234
rect 44770 19182 44772 19234
rect 44716 18452 44772 19182
rect 44380 17938 44436 17948
rect 44044 17780 44100 17790
rect 43932 17724 44044 17780
rect 44044 17714 44100 17724
rect 44156 17780 44212 17790
rect 44716 17780 44772 18396
rect 44156 17778 44772 17780
rect 44156 17726 44158 17778
rect 44210 17726 44772 17778
rect 44156 17724 44772 17726
rect 44828 18450 44884 18462
rect 44828 18398 44830 18450
rect 44882 18398 44884 18450
rect 44156 17714 44212 17724
rect 44044 17444 44100 17454
rect 44268 17444 44324 17454
rect 43820 17442 44100 17444
rect 43820 17390 44046 17442
rect 44098 17390 44100 17442
rect 43820 17388 44100 17390
rect 44044 17220 44100 17388
rect 44044 17154 44100 17164
rect 44156 17442 44324 17444
rect 44156 17390 44270 17442
rect 44322 17390 44324 17442
rect 44156 17388 44324 17390
rect 42700 16882 42756 16940
rect 42700 16830 42702 16882
rect 42754 16830 42756 16882
rect 41804 16772 41860 16782
rect 40348 16046 40350 16098
rect 40402 16046 40404 16098
rect 40348 16034 40404 16046
rect 40460 16156 40628 16212
rect 41132 16156 41300 16212
rect 41356 16770 41860 16772
rect 41356 16718 41806 16770
rect 41858 16718 41860 16770
rect 41356 16716 41860 16718
rect 40012 15988 40068 15998
rect 40012 15894 40068 15932
rect 39564 15874 39732 15876
rect 39564 15822 39566 15874
rect 39618 15822 39732 15874
rect 39564 15820 39732 15822
rect 39788 15876 39844 15886
rect 39564 15810 39620 15820
rect 39676 15428 39732 15438
rect 39452 15426 39732 15428
rect 39452 15374 39678 15426
rect 39730 15374 39732 15426
rect 39452 15372 39732 15374
rect 39676 15316 39732 15372
rect 39788 15426 39844 15820
rect 40236 15876 40292 15886
rect 40236 15782 40292 15820
rect 40012 15540 40068 15550
rect 40012 15446 40068 15484
rect 39788 15374 39790 15426
rect 39842 15374 39844 15426
rect 39788 15362 39844 15374
rect 40236 15426 40292 15438
rect 40236 15374 40238 15426
rect 40290 15374 40292 15426
rect 39676 15250 39732 15260
rect 39676 15090 39732 15102
rect 39676 15038 39678 15090
rect 39730 15038 39732 15090
rect 39340 14466 39396 14476
rect 39564 14644 39620 14654
rect 38556 12796 38836 12852
rect 38892 13916 39172 13972
rect 39452 14306 39508 14318
rect 39452 14254 39454 14306
rect 39506 14254 39508 14306
rect 38892 12962 38948 13916
rect 38892 12910 38894 12962
rect 38946 12910 38948 12962
rect 37772 12740 37828 12750
rect 38556 12740 38612 12796
rect 37100 12292 37156 12302
rect 36652 12066 36708 12078
rect 36652 12014 36654 12066
rect 36706 12014 36708 12066
rect 36316 9826 36484 9828
rect 36316 9774 36318 9826
rect 36370 9774 36484 9826
rect 36316 9772 36484 9774
rect 36540 11732 36596 11742
rect 36316 9762 36372 9772
rect 36092 9714 36260 9716
rect 36092 9662 36094 9714
rect 36146 9662 36260 9714
rect 36092 9660 36260 9662
rect 36092 9650 36148 9660
rect 34636 9214 34638 9266
rect 34690 9214 34692 9266
rect 34636 9202 34692 9214
rect 34860 9602 34916 9614
rect 35196 9604 35252 9614
rect 34860 9550 34862 9602
rect 34914 9550 34916 9602
rect 33180 8206 33182 8258
rect 33234 8206 33236 8258
rect 33180 8194 33236 8206
rect 34524 8260 34580 8876
rect 34524 8194 34580 8204
rect 32732 7858 32788 7868
rect 33404 8034 33460 8046
rect 33404 7982 33406 8034
rect 33458 7982 33460 8034
rect 33404 7476 33460 7982
rect 32060 7308 32340 7364
rect 33068 7362 33124 7374
rect 33068 7310 33070 7362
rect 33122 7310 33124 7362
rect 32060 6466 32116 7308
rect 32284 6916 32340 6926
rect 32172 6804 32228 6814
rect 32172 6710 32228 6748
rect 32284 6690 32340 6860
rect 33068 6916 33124 7310
rect 33068 6850 33124 6860
rect 32956 6804 33012 6814
rect 32956 6710 33012 6748
rect 32284 6638 32286 6690
rect 32338 6638 32340 6690
rect 32284 6626 32340 6638
rect 33292 6690 33348 6702
rect 33292 6638 33294 6690
rect 33346 6638 33348 6690
rect 32060 6414 32062 6466
rect 32114 6414 32116 6466
rect 32060 6356 32116 6414
rect 32060 6290 32116 6300
rect 33068 6578 33124 6590
rect 33068 6526 33070 6578
rect 33122 6526 33124 6578
rect 32060 6020 32116 6030
rect 32060 5926 32116 5964
rect 32396 6018 32452 6030
rect 32396 5966 32398 6018
rect 32450 5966 32452 6018
rect 31948 5070 31950 5122
rect 32002 5070 32004 5122
rect 31948 5058 32004 5070
rect 31836 4834 31892 4844
rect 31500 4788 31556 4798
rect 31276 3556 31332 3566
rect 31164 3554 31332 3556
rect 31164 3502 31278 3554
rect 31330 3502 31332 3554
rect 31164 3500 31332 3502
rect 30268 800 30324 3500
rect 31276 3490 31332 3500
rect 30940 3444 30996 3454
rect 31500 3444 31556 4732
rect 31724 4788 31780 4798
rect 31612 3444 31668 3454
rect 31500 3442 31668 3444
rect 31500 3390 31614 3442
rect 31666 3390 31668 3442
rect 31500 3388 31668 3390
rect 30940 800 30996 3388
rect 31612 3378 31668 3388
rect 31724 1764 31780 4732
rect 32396 4452 32452 5966
rect 32620 5684 32676 5694
rect 32620 5234 32676 5628
rect 32620 5182 32622 5234
rect 32674 5182 32676 5234
rect 32620 5170 32676 5182
rect 33068 5236 33124 6526
rect 33180 6132 33236 6142
rect 33180 6038 33236 6076
rect 33292 6130 33348 6638
rect 33292 6078 33294 6130
rect 33346 6078 33348 6130
rect 33292 6066 33348 6078
rect 33404 6018 33460 7420
rect 34076 6692 34132 6702
rect 34300 6692 34356 6702
rect 34076 6690 34356 6692
rect 34076 6638 34078 6690
rect 34130 6638 34302 6690
rect 34354 6638 34356 6690
rect 34076 6636 34356 6638
rect 34076 6626 34132 6636
rect 34300 6626 34356 6636
rect 34636 6692 34692 6702
rect 34636 6598 34692 6636
rect 33404 5966 33406 6018
rect 33458 5966 33460 6018
rect 33404 5954 33460 5966
rect 33740 6580 33796 6590
rect 33740 6018 33796 6524
rect 34524 6466 34580 6478
rect 34524 6414 34526 6466
rect 34578 6414 34580 6466
rect 34524 6132 34580 6414
rect 34860 6468 34916 9550
rect 35084 9602 35252 9604
rect 35084 9550 35198 9602
rect 35250 9550 35252 9602
rect 35084 9548 35252 9550
rect 36204 9604 36260 9660
rect 36204 9548 36484 9604
rect 35084 8372 35140 9548
rect 35196 9538 35252 9548
rect 35196 9380 35252 9390
rect 35196 9042 35252 9324
rect 35196 8990 35198 9042
rect 35250 8990 35252 9042
rect 35196 8820 35252 8990
rect 36428 9042 36484 9548
rect 36428 8990 36430 9042
rect 36482 8990 36484 9042
rect 36428 8978 36484 8990
rect 35196 8754 35252 8764
rect 35756 8930 35812 8942
rect 35756 8878 35758 8930
rect 35810 8878 35812 8930
rect 35644 8708 35700 8718
rect 35196 8652 35460 8662
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35196 8586 35460 8596
rect 35308 8372 35364 8382
rect 35084 8370 35364 8372
rect 35084 8318 35310 8370
rect 35362 8318 35364 8370
rect 35084 8316 35364 8318
rect 35308 8306 35364 8316
rect 35644 8258 35700 8652
rect 35644 8206 35646 8258
rect 35698 8206 35700 8258
rect 35644 8194 35700 8206
rect 34972 8036 35028 8046
rect 34972 8034 35140 8036
rect 34972 7982 34974 8034
rect 35026 7982 35140 8034
rect 34972 7980 35140 7982
rect 34972 7970 35028 7980
rect 34860 6402 34916 6412
rect 34524 6076 34692 6132
rect 33740 5966 33742 6018
rect 33794 5966 33796 6018
rect 33740 5954 33796 5966
rect 33852 6018 33908 6030
rect 33852 5966 33854 6018
rect 33906 5966 33908 6018
rect 33852 5908 33908 5966
rect 34412 6018 34468 6030
rect 34412 5966 34414 6018
rect 34466 5966 34468 6018
rect 34188 5908 34244 5918
rect 33852 5842 33908 5852
rect 33964 5906 34244 5908
rect 33964 5854 34190 5906
rect 34242 5854 34244 5906
rect 33964 5852 34244 5854
rect 33852 5682 33908 5694
rect 33852 5630 33854 5682
rect 33906 5630 33908 5682
rect 33852 5348 33908 5630
rect 33852 5282 33908 5292
rect 33068 5180 33348 5236
rect 33068 5012 33124 5022
rect 33068 4562 33124 4956
rect 33068 4510 33070 4562
rect 33122 4510 33124 4562
rect 33068 4498 33124 4510
rect 32396 4386 32452 4396
rect 33180 4226 33236 4238
rect 33180 4174 33182 4226
rect 33234 4174 33236 4226
rect 33180 3892 33236 4174
rect 32508 3836 33236 3892
rect 32284 3556 32340 3566
rect 32284 3462 32340 3500
rect 32508 3442 32564 3836
rect 32508 3390 32510 3442
rect 32562 3390 32564 3442
rect 32508 3378 32564 3390
rect 32956 3668 33012 3678
rect 31612 1708 31780 1764
rect 31612 800 31668 1708
rect 32956 800 33012 3612
rect 33292 3554 33348 5180
rect 33964 5012 34020 5852
rect 34188 5842 34244 5852
rect 33852 4956 34020 5012
rect 33852 4450 33908 4956
rect 34412 4788 34468 5966
rect 34524 5908 34580 5918
rect 34524 5814 34580 5852
rect 34636 5236 34692 6076
rect 34972 5794 35028 5806
rect 34972 5742 34974 5794
rect 35026 5742 35028 5794
rect 34860 5684 34916 5694
rect 34860 5590 34916 5628
rect 34748 5236 34804 5246
rect 34188 4732 34468 4788
rect 34524 5234 34804 5236
rect 34524 5182 34750 5234
rect 34802 5182 34804 5234
rect 34524 5180 34804 5182
rect 34188 4676 34244 4732
rect 34188 4610 34244 4620
rect 34076 4564 34132 4574
rect 34076 4470 34132 4508
rect 34300 4564 34356 4574
rect 34524 4564 34580 5180
rect 34748 5170 34804 5180
rect 34300 4562 34580 4564
rect 34300 4510 34302 4562
rect 34354 4510 34580 4562
rect 34300 4508 34580 4510
rect 34636 5012 34692 5022
rect 34972 5012 35028 5742
rect 34636 4562 34692 4956
rect 34636 4510 34638 4562
rect 34690 4510 34692 4562
rect 34300 4498 34356 4508
rect 34636 4498 34692 4510
rect 34860 4956 35028 5012
rect 33852 4398 33854 4450
rect 33906 4398 33908 4450
rect 33852 4386 33908 4398
rect 33964 4452 34020 4462
rect 33964 4358 34020 4396
rect 34188 4228 34244 4238
rect 34860 4228 34916 4956
rect 34972 4788 35028 4798
rect 34972 4450 35028 4732
rect 34972 4398 34974 4450
rect 35026 4398 35028 4450
rect 34972 4386 35028 4398
rect 34188 4226 34916 4228
rect 34188 4174 34190 4226
rect 34242 4174 34916 4226
rect 34188 4172 34916 4174
rect 34188 4162 34244 4172
rect 33852 3668 33908 3678
rect 33852 3574 33908 3612
rect 33292 3502 33294 3554
rect 33346 3502 33348 3554
rect 33292 3490 33348 3502
rect 33628 3556 33684 3566
rect 33628 800 33684 3500
rect 35084 3556 35140 7980
rect 35420 7476 35476 7486
rect 35420 7382 35476 7420
rect 35196 7084 35460 7094
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35196 7018 35460 7028
rect 35308 6916 35364 6926
rect 35308 6822 35364 6860
rect 35756 6804 35812 8878
rect 36204 8932 36260 8942
rect 36204 8930 36372 8932
rect 36204 8878 36206 8930
rect 36258 8878 36372 8930
rect 36204 8876 36372 8878
rect 36204 8866 36260 8876
rect 36316 8820 36372 8876
rect 36540 8820 36596 11676
rect 36652 10500 36708 12014
rect 36988 11620 37044 11630
rect 36988 11506 37044 11564
rect 37100 11618 37156 12236
rect 37324 12180 37380 12190
rect 37324 12086 37380 12124
rect 37772 12178 37828 12684
rect 38332 12684 38612 12740
rect 37772 12126 37774 12178
rect 37826 12126 37828 12178
rect 37772 12068 37828 12126
rect 37996 12628 38052 12638
rect 37996 12178 38052 12572
rect 37996 12126 37998 12178
rect 38050 12126 38052 12178
rect 37828 12012 37940 12068
rect 37772 12002 37828 12012
rect 37100 11566 37102 11618
rect 37154 11566 37156 11618
rect 37100 11554 37156 11566
rect 37436 11844 37492 11854
rect 36988 11454 36990 11506
rect 37042 11454 37044 11506
rect 36988 11284 37044 11454
rect 36988 11218 37044 11228
rect 37100 10724 37156 10734
rect 37100 10630 37156 10668
rect 36652 10434 36708 10444
rect 37436 9938 37492 11788
rect 37548 11284 37604 11294
rect 37548 11190 37604 11228
rect 37436 9886 37438 9938
rect 37490 9886 37492 9938
rect 37436 9874 37492 9886
rect 37884 9938 37940 12012
rect 37996 11844 38052 12126
rect 37996 11778 38052 11788
rect 38220 11954 38276 11966
rect 38220 11902 38222 11954
rect 38274 11902 38276 11954
rect 37996 11506 38052 11518
rect 37996 11454 37998 11506
rect 38050 11454 38052 11506
rect 37996 10724 38052 11454
rect 38220 11396 38276 11902
rect 38220 11330 38276 11340
rect 38332 11956 38388 12684
rect 38780 12292 38836 12302
rect 38780 12178 38836 12236
rect 38780 12126 38782 12178
rect 38834 12126 38836 12178
rect 38780 12114 38836 12126
rect 38332 11060 38388 11900
rect 38444 12066 38500 12078
rect 38444 12014 38446 12066
rect 38498 12014 38500 12066
rect 38444 11508 38500 12014
rect 38892 12068 38948 12910
rect 38892 12002 38948 12012
rect 39004 13748 39060 13758
rect 39004 11508 39060 13692
rect 39452 13076 39508 14254
rect 39452 13010 39508 13020
rect 39340 12180 39396 12190
rect 39340 12086 39396 12124
rect 39452 12068 39508 12078
rect 39564 12068 39620 14588
rect 39676 14308 39732 15038
rect 40012 14980 40068 14990
rect 40236 14980 40292 15374
rect 40348 15428 40404 15438
rect 40348 15334 40404 15372
rect 40460 15148 40516 16156
rect 40796 16098 40852 16110
rect 41132 16100 41188 16156
rect 40796 16046 40798 16098
rect 40850 16046 40852 16098
rect 40796 15540 40852 16046
rect 41020 16044 41188 16100
rect 41356 16098 41412 16716
rect 41804 16706 41860 16716
rect 41916 16660 41972 16670
rect 41356 16046 41358 16098
rect 41410 16046 41412 16098
rect 40796 15474 40852 15484
rect 40908 15764 40964 15774
rect 40068 14924 40292 14980
rect 40348 15092 40516 15148
rect 40012 14914 40068 14924
rect 40124 14756 40180 14766
rect 40012 14532 40068 14542
rect 39676 14242 39732 14252
rect 39788 14306 39844 14318
rect 39788 14254 39790 14306
rect 39842 14254 39844 14306
rect 39788 14084 39844 14254
rect 39788 14018 39844 14028
rect 40012 13972 40068 14476
rect 40012 13906 40068 13916
rect 40012 13748 40068 13758
rect 40124 13748 40180 14700
rect 40012 13746 40180 13748
rect 40012 13694 40014 13746
rect 40066 13694 40180 13746
rect 40012 13692 40180 13694
rect 40012 13682 40068 13692
rect 39676 13636 39732 13646
rect 39676 13074 39732 13580
rect 40348 13186 40404 15092
rect 40572 14644 40628 14654
rect 40572 14550 40628 14588
rect 40684 14532 40740 14542
rect 40908 14532 40964 15708
rect 41020 15652 41076 16044
rect 41356 16034 41412 16046
rect 41580 16436 41636 16446
rect 41580 16098 41636 16380
rect 41580 16046 41582 16098
rect 41634 16046 41636 16098
rect 41580 16034 41636 16046
rect 41244 15988 41300 15998
rect 41132 15932 41244 15988
rect 41132 15874 41188 15932
rect 41244 15922 41300 15932
rect 41468 15988 41524 15998
rect 41468 15894 41524 15932
rect 41132 15822 41134 15874
rect 41186 15822 41188 15874
rect 41132 15810 41188 15822
rect 41916 15652 41972 16604
rect 42140 16658 42196 16670
rect 42140 16606 42142 16658
rect 42194 16606 42196 16658
rect 42028 16212 42084 16222
rect 42140 16212 42196 16606
rect 42252 16658 42308 16670
rect 42252 16606 42254 16658
rect 42306 16606 42308 16658
rect 42252 16548 42308 16606
rect 42700 16548 42756 16830
rect 42812 16994 42868 17006
rect 42812 16942 42814 16994
rect 42866 16942 42868 16994
rect 42812 16884 42868 16942
rect 43260 16994 43316 17052
rect 43708 17014 43764 17052
rect 43260 16942 43262 16994
rect 43314 16942 43316 16994
rect 43260 16930 43316 16942
rect 43484 16884 43540 16894
rect 43820 16884 43876 16894
rect 42812 16828 43204 16884
rect 42812 16660 42868 16670
rect 42812 16658 42980 16660
rect 42812 16606 42814 16658
rect 42866 16606 42980 16658
rect 42812 16604 42980 16606
rect 42812 16594 42868 16604
rect 42252 16492 42756 16548
rect 42924 16548 42980 16604
rect 42140 16156 42532 16212
rect 42028 16100 42084 16156
rect 42028 16044 42196 16100
rect 42140 15986 42196 16044
rect 42140 15934 42142 15986
rect 42194 15934 42196 15986
rect 42140 15922 42196 15934
rect 42476 15986 42532 16156
rect 42476 15934 42478 15986
rect 42530 15934 42532 15986
rect 41020 15596 41524 15652
rect 41132 15484 41300 15540
rect 40684 14530 40964 14532
rect 40684 14478 40686 14530
rect 40738 14478 40964 14530
rect 40684 14476 40964 14478
rect 41020 15204 41076 15214
rect 41020 14530 41076 15148
rect 41020 14478 41022 14530
rect 41074 14478 41076 14530
rect 40684 14466 40740 14476
rect 41020 14466 41076 14478
rect 41132 14532 41188 15484
rect 41244 15426 41300 15484
rect 41468 15538 41524 15596
rect 41468 15486 41470 15538
rect 41522 15486 41524 15538
rect 41468 15474 41524 15486
rect 41692 15596 41972 15652
rect 42028 15874 42084 15886
rect 42028 15822 42030 15874
rect 42082 15822 42084 15874
rect 41692 15538 41748 15596
rect 41692 15486 41694 15538
rect 41746 15486 41748 15538
rect 41692 15474 41748 15486
rect 42028 15540 42084 15822
rect 42252 15876 42308 15886
rect 42140 15540 42196 15550
rect 42028 15484 42140 15540
rect 42140 15474 42196 15484
rect 41244 15374 41246 15426
rect 41298 15374 41300 15426
rect 41244 15362 41300 15374
rect 41580 15316 41636 15326
rect 41580 15222 41636 15260
rect 41916 15314 41972 15326
rect 41916 15262 41918 15314
rect 41970 15262 41972 15314
rect 41916 15092 41972 15262
rect 42252 15148 42308 15820
rect 41804 15036 41972 15092
rect 42140 15092 42308 15148
rect 42364 15204 42420 15242
rect 42364 15138 42420 15148
rect 41580 14754 41636 14766
rect 41580 14702 41582 14754
rect 41634 14702 41636 14754
rect 41132 14466 41188 14476
rect 41468 14532 41524 14542
rect 41468 14438 41524 14476
rect 40460 14308 40516 14318
rect 40460 13748 40516 14252
rect 40796 14308 40852 14318
rect 40460 13682 40516 13692
rect 40684 14196 40740 14206
rect 40348 13134 40350 13186
rect 40402 13134 40404 13186
rect 40348 13122 40404 13134
rect 40684 13186 40740 14140
rect 40796 13746 40852 14252
rect 41244 14306 41300 14318
rect 41244 14254 41246 14306
rect 41298 14254 41300 14306
rect 41244 14196 41300 14254
rect 40796 13694 40798 13746
rect 40850 13694 40852 13746
rect 40796 13682 40852 13694
rect 41020 14084 41076 14094
rect 40684 13134 40686 13186
rect 40738 13134 40740 13186
rect 40684 13122 40740 13134
rect 40908 13412 40964 13422
rect 39676 13022 39678 13074
rect 39730 13022 39732 13074
rect 39676 13010 39732 13022
rect 40012 12962 40068 12974
rect 40012 12910 40014 12962
rect 40066 12910 40068 12962
rect 40012 12852 40068 12910
rect 39452 12066 39620 12068
rect 39452 12014 39454 12066
rect 39506 12014 39620 12066
rect 39452 12012 39620 12014
rect 39900 12290 39956 12302
rect 39900 12238 39902 12290
rect 39954 12238 39956 12290
rect 39452 12002 39508 12012
rect 39900 11618 39956 12238
rect 40012 12292 40068 12796
rect 40908 12962 40964 13356
rect 40908 12910 40910 12962
rect 40962 12910 40964 12962
rect 40348 12292 40404 12302
rect 40012 12290 40404 12292
rect 40012 12238 40350 12290
rect 40402 12238 40404 12290
rect 40012 12236 40404 12238
rect 40348 12226 40404 12236
rect 40236 11954 40292 11966
rect 40236 11902 40238 11954
rect 40290 11902 40292 11954
rect 40236 11732 40292 11902
rect 40236 11666 40292 11676
rect 39900 11566 39902 11618
rect 39954 11566 39956 11618
rect 39900 11554 39956 11566
rect 40908 11620 40964 12910
rect 41020 12066 41076 14028
rect 41020 12014 41022 12066
rect 41074 12014 41076 12066
rect 41020 12002 41076 12014
rect 41132 13076 41188 13086
rect 40908 11554 40964 11564
rect 38444 11442 38500 11452
rect 38892 11452 39060 11508
rect 39788 11508 39844 11518
rect 38332 11004 38612 11060
rect 37996 10658 38052 10668
rect 37884 9886 37886 9938
rect 37938 9886 37940 9938
rect 37884 9874 37940 9886
rect 38108 10052 38164 10062
rect 38108 9826 38164 9996
rect 38108 9774 38110 9826
rect 38162 9774 38164 9826
rect 36876 9716 36932 9726
rect 36876 9042 36932 9660
rect 38108 9268 38164 9774
rect 38220 9268 38276 9278
rect 38108 9266 38276 9268
rect 38108 9214 38222 9266
rect 38274 9214 38276 9266
rect 38108 9212 38276 9214
rect 37324 9156 37380 9166
rect 37324 9062 37380 9100
rect 36876 8990 36878 9042
rect 36930 8990 36932 9042
rect 36876 8978 36932 8990
rect 37884 8932 37940 8942
rect 37884 8930 38052 8932
rect 37884 8878 37886 8930
rect 37938 8878 38052 8930
rect 37884 8876 38052 8878
rect 37884 8866 37940 8876
rect 36316 8764 36596 8820
rect 36652 8818 36708 8830
rect 36652 8766 36654 8818
rect 36706 8766 36708 8818
rect 35980 8372 36036 8382
rect 35868 8258 35924 8270
rect 35868 8206 35870 8258
rect 35922 8206 35924 8258
rect 35868 8148 35924 8206
rect 35868 8082 35924 8092
rect 35980 7700 36036 8316
rect 36540 8372 36596 8382
rect 36540 8258 36596 8316
rect 36540 8206 36542 8258
rect 36594 8206 36596 8258
rect 36540 8194 36596 8206
rect 35980 7476 36036 7644
rect 36652 7812 36708 8766
rect 37324 8148 37380 8158
rect 37324 8054 37380 8092
rect 36988 8034 37044 8046
rect 36988 7982 36990 8034
rect 37042 7982 37044 8034
rect 36988 7812 37044 7982
rect 36652 7756 37044 7812
rect 37772 8034 37828 8046
rect 37772 7982 37774 8034
rect 37826 7982 37828 8034
rect 35756 6738 35812 6748
rect 35868 7474 36036 7476
rect 35868 7422 35982 7474
rect 36034 7422 36036 7474
rect 35868 7420 36036 7422
rect 35196 6578 35252 6590
rect 35196 6526 35198 6578
rect 35250 6526 35252 6578
rect 35196 6244 35252 6526
rect 35196 6178 35252 6188
rect 35756 6466 35812 6478
rect 35756 6414 35758 6466
rect 35810 6414 35812 6466
rect 35756 6132 35812 6414
rect 35756 6066 35812 6076
rect 35308 5908 35364 5918
rect 35308 5814 35364 5852
rect 35868 5906 35924 7420
rect 35980 7410 36036 7420
rect 36428 7476 36484 7486
rect 36652 7476 36708 7756
rect 37212 7700 37268 7710
rect 37212 7606 37268 7644
rect 36428 7474 36708 7476
rect 36428 7422 36430 7474
rect 36482 7422 36708 7474
rect 36428 7420 36708 7422
rect 36764 7586 36820 7598
rect 36764 7534 36766 7586
rect 36818 7534 36820 7586
rect 36428 6916 36484 7420
rect 36428 6850 36484 6860
rect 36652 6692 36708 6702
rect 36764 6692 36820 7534
rect 37660 7362 37716 7374
rect 37660 7310 37662 7362
rect 37714 7310 37716 7362
rect 37660 6804 37716 7310
rect 37660 6738 37716 6748
rect 36708 6636 36820 6692
rect 36652 6626 36708 6636
rect 35868 5854 35870 5906
rect 35922 5854 35924 5906
rect 35868 5842 35924 5854
rect 36316 6578 36372 6590
rect 36316 6526 36318 6578
rect 36370 6526 36372 6578
rect 35420 5796 35476 5806
rect 35420 5794 35812 5796
rect 35420 5742 35422 5794
rect 35474 5742 35812 5794
rect 35420 5740 35812 5742
rect 35420 5730 35476 5740
rect 35196 5516 35460 5526
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35196 5450 35460 5460
rect 35196 5346 35252 5358
rect 35196 5294 35198 5346
rect 35250 5294 35252 5346
rect 35196 5236 35252 5294
rect 35644 5348 35700 5358
rect 35196 5180 35476 5236
rect 35308 5012 35364 5022
rect 35308 4918 35364 4956
rect 35196 4898 35252 4910
rect 35196 4846 35198 4898
rect 35250 4846 35252 4898
rect 35196 4676 35252 4846
rect 35196 4610 35252 4620
rect 35420 4340 35476 5180
rect 35644 5122 35700 5292
rect 35644 5070 35646 5122
rect 35698 5070 35700 5122
rect 35644 5058 35700 5070
rect 35532 4340 35588 4350
rect 35420 4338 35588 4340
rect 35420 4286 35534 4338
rect 35586 4286 35588 4338
rect 35420 4284 35588 4286
rect 35532 4274 35588 4284
rect 35756 4004 35812 5740
rect 36092 5572 36148 5582
rect 35868 5124 35924 5134
rect 35868 4228 35924 5068
rect 36092 5012 36148 5516
rect 36316 5234 36372 6526
rect 36428 6466 36484 6478
rect 36428 6414 36430 6466
rect 36482 6414 36484 6466
rect 36428 6020 36484 6414
rect 36652 6468 36708 6478
rect 36540 6020 36596 6030
rect 36428 6018 36596 6020
rect 36428 5966 36542 6018
rect 36594 5966 36596 6018
rect 36428 5964 36596 5966
rect 36540 5954 36596 5964
rect 36652 5796 36708 6412
rect 36764 6132 36820 6636
rect 36764 6066 36820 6076
rect 37100 6580 37156 6590
rect 36316 5182 36318 5234
rect 36370 5182 36372 5234
rect 36316 5170 36372 5182
rect 36428 5740 36708 5796
rect 36428 5122 36484 5740
rect 36652 5684 36708 5740
rect 36652 5618 36708 5628
rect 36428 5070 36430 5122
rect 36482 5070 36484 5122
rect 36428 5058 36484 5070
rect 36540 5348 36596 5358
rect 35980 5010 36148 5012
rect 35980 4958 36094 5010
rect 36146 4958 36148 5010
rect 35980 4956 36148 4958
rect 35980 4452 36036 4956
rect 36092 4946 36148 4956
rect 36204 4898 36260 4910
rect 36204 4846 36206 4898
rect 36258 4846 36260 4898
rect 36092 4564 36148 4574
rect 36204 4564 36260 4846
rect 36148 4508 36260 4564
rect 36316 4564 36372 4574
rect 36540 4564 36596 5292
rect 37100 5124 37156 6524
rect 37324 6578 37380 6590
rect 37324 6526 37326 6578
rect 37378 6526 37380 6578
rect 37324 6132 37380 6526
rect 37772 6580 37828 7982
rect 37884 6804 37940 6814
rect 37884 6690 37940 6748
rect 37884 6638 37886 6690
rect 37938 6638 37940 6690
rect 37884 6626 37940 6638
rect 37996 6692 38052 8876
rect 38108 8372 38164 9212
rect 38220 9202 38276 9212
rect 38556 9266 38612 11004
rect 38892 9940 38948 11452
rect 39228 11396 39284 11406
rect 39004 11284 39060 11294
rect 39004 11190 39060 11228
rect 39228 10498 39284 11340
rect 39676 11396 39732 11406
rect 39676 11302 39732 11340
rect 39676 10724 39732 10734
rect 39788 10724 39844 11452
rect 40236 11508 40292 11518
rect 40236 11282 40292 11452
rect 40684 11508 40740 11518
rect 40684 11414 40740 11452
rect 40236 11230 40238 11282
rect 40290 11230 40292 11282
rect 40236 11218 40292 11230
rect 40012 11172 40068 11182
rect 40012 11170 40180 11172
rect 40012 11118 40014 11170
rect 40066 11118 40180 11170
rect 40012 11116 40180 11118
rect 40012 11106 40068 11116
rect 40124 10836 40180 11116
rect 40236 10836 40292 10846
rect 40124 10834 40292 10836
rect 40124 10782 40238 10834
rect 40290 10782 40292 10834
rect 40124 10780 40292 10782
rect 40236 10770 40292 10780
rect 41132 10834 41188 13020
rect 41244 12962 41300 14140
rect 41580 13972 41636 14702
rect 41804 14644 41860 15036
rect 42140 14980 42196 15092
rect 41804 14578 41860 14588
rect 41916 14924 42196 14980
rect 41692 14532 41748 14542
rect 41692 14438 41748 14476
rect 41580 13916 41748 13972
rect 41468 13860 41524 13870
rect 41244 12910 41246 12962
rect 41298 12910 41300 12962
rect 41244 12898 41300 12910
rect 41356 13804 41468 13860
rect 41356 12516 41412 13804
rect 41468 13794 41524 13804
rect 41580 13748 41636 13758
rect 41580 13654 41636 13692
rect 41692 13524 41748 13916
rect 41580 13468 41748 13524
rect 41468 13074 41524 13086
rect 41468 13022 41470 13074
rect 41522 13022 41524 13074
rect 41468 12964 41524 13022
rect 41468 12898 41524 12908
rect 41580 12850 41636 13468
rect 41580 12798 41582 12850
rect 41634 12798 41636 12850
rect 41580 12786 41636 12798
rect 41692 13076 41748 13086
rect 41692 12850 41748 13020
rect 41916 12964 41972 14924
rect 42140 14420 42196 14430
rect 42028 14308 42084 14318
rect 42028 13524 42084 14252
rect 42140 13746 42196 14364
rect 42364 14306 42420 14318
rect 42364 14254 42366 14306
rect 42418 14254 42420 14306
rect 42364 14196 42420 14254
rect 42364 14130 42420 14140
rect 42252 13860 42308 13870
rect 42252 13766 42308 13804
rect 42140 13694 42142 13746
rect 42194 13694 42196 13746
rect 42140 13682 42196 13694
rect 42476 13636 42532 15934
rect 42588 15428 42644 16492
rect 42924 16482 42980 16492
rect 42812 16436 42868 16446
rect 42588 15362 42644 15372
rect 42700 16380 42812 16436
rect 43148 16436 43204 16828
rect 43148 16380 43428 16436
rect 42700 14308 42756 16380
rect 42812 16370 42868 16380
rect 43372 16322 43428 16380
rect 43372 16270 43374 16322
rect 43426 16270 43428 16322
rect 43372 16258 43428 16270
rect 43036 16212 43092 16222
rect 43092 16156 43204 16212
rect 43036 16118 43092 16156
rect 43036 15652 43092 15662
rect 42700 14242 42756 14252
rect 42812 15202 42868 15214
rect 42812 15150 42814 15202
rect 42866 15150 42868 15202
rect 42812 13860 42868 15150
rect 43036 14530 43092 15596
rect 43148 14868 43204 16156
rect 43484 15874 43540 16828
rect 43484 15822 43486 15874
rect 43538 15822 43540 15874
rect 43484 15538 43540 15822
rect 43484 15486 43486 15538
rect 43538 15486 43540 15538
rect 43484 15474 43540 15486
rect 43596 16828 43820 16884
rect 43148 14802 43204 14812
rect 43596 14756 43652 16828
rect 43820 16790 43876 16828
rect 44156 16884 44212 17388
rect 44268 17378 44324 17388
rect 44604 17444 44660 17454
rect 44380 17332 44436 17342
rect 44268 16996 44324 17006
rect 44268 16902 44324 16940
rect 44156 16818 44212 16828
rect 44380 16210 44436 17276
rect 44380 16158 44382 16210
rect 44434 16158 44436 16210
rect 44380 16146 44436 16158
rect 44492 17108 44548 17118
rect 43708 15986 43764 15998
rect 43708 15934 43710 15986
rect 43762 15934 43764 15986
rect 43708 15540 43764 15934
rect 43708 15484 44212 15540
rect 43820 15316 43876 15326
rect 43596 14690 43652 14700
rect 43708 15260 43820 15316
rect 43484 14644 43540 14654
rect 43484 14550 43540 14588
rect 43708 14532 43764 15260
rect 43820 15222 43876 15260
rect 43036 14478 43038 14530
rect 43090 14478 43092 14530
rect 43036 14466 43092 14478
rect 43596 14476 43764 14532
rect 44156 15092 44212 15484
rect 43484 14420 43540 14430
rect 43484 14326 43540 14364
rect 42812 13794 42868 13804
rect 43596 13860 43652 14476
rect 43820 14418 43876 14430
rect 43820 14366 43822 14418
rect 43874 14366 43876 14418
rect 43708 13860 43764 13870
rect 43596 13858 43764 13860
rect 43596 13806 43710 13858
rect 43762 13806 43764 13858
rect 43596 13804 43764 13806
rect 43372 13746 43428 13758
rect 43372 13694 43374 13746
rect 43426 13694 43428 13746
rect 42476 13570 42532 13580
rect 42700 13634 42756 13646
rect 42700 13582 42702 13634
rect 42754 13582 42756 13634
rect 42028 13468 42308 13524
rect 42140 13188 42196 13198
rect 41916 12908 42084 12964
rect 41692 12798 41694 12850
rect 41746 12798 41748 12850
rect 41692 12786 41748 12798
rect 41468 12740 41524 12750
rect 41468 12646 41524 12684
rect 41356 12460 41636 12516
rect 41132 10782 41134 10834
rect 41186 10782 41188 10834
rect 39676 10722 39844 10724
rect 39676 10670 39678 10722
rect 39730 10670 39844 10722
rect 39676 10668 39844 10670
rect 39676 10658 39732 10668
rect 39228 10446 39230 10498
rect 39282 10446 39284 10498
rect 39228 10434 39284 10446
rect 40348 10500 40404 10510
rect 40348 10498 40852 10500
rect 40348 10446 40350 10498
rect 40402 10446 40852 10498
rect 40348 10444 40852 10446
rect 40348 10434 40404 10444
rect 39564 10388 39620 10398
rect 38892 9874 38948 9884
rect 39340 10386 39620 10388
rect 39340 10334 39566 10386
rect 39618 10334 39620 10386
rect 39340 10332 39620 10334
rect 38892 9714 38948 9726
rect 39340 9716 39396 10332
rect 39564 10322 39620 10332
rect 38892 9662 38894 9714
rect 38946 9662 38948 9714
rect 38556 9214 38558 9266
rect 38610 9214 38612 9266
rect 38556 9202 38612 9214
rect 38780 9268 38836 9278
rect 38780 9174 38836 9212
rect 38892 8930 38948 9662
rect 39116 9660 39396 9716
rect 39900 10164 39956 10174
rect 39116 9042 39172 9660
rect 39116 8990 39118 9042
rect 39170 8990 39172 9042
rect 39116 8978 39172 8990
rect 38892 8878 38894 8930
rect 38946 8878 38948 8930
rect 38892 8866 38948 8878
rect 39004 8932 39060 8942
rect 39004 8820 39060 8876
rect 39452 8930 39508 8942
rect 39452 8878 39454 8930
rect 39506 8878 39508 8930
rect 39004 8764 39172 8820
rect 38444 8596 38500 8606
rect 38332 8372 38388 8382
rect 38108 8370 38388 8372
rect 38108 8318 38334 8370
rect 38386 8318 38388 8370
rect 38108 8316 38388 8318
rect 38108 8036 38164 8316
rect 38332 8306 38388 8316
rect 38108 7700 38164 7980
rect 38108 7634 38164 7644
rect 38220 8148 38276 8158
rect 38220 8036 38276 8092
rect 38444 8036 38500 8540
rect 38220 7980 38500 8036
rect 38780 8258 38836 8270
rect 38780 8206 38782 8258
rect 38834 8206 38836 8258
rect 38220 7698 38276 7980
rect 38220 7646 38222 7698
rect 38274 7646 38276 7698
rect 38220 7634 38276 7646
rect 38780 7588 38836 8206
rect 38780 7522 38836 7532
rect 39004 8034 39060 8046
rect 39004 7982 39006 8034
rect 39058 7982 39060 8034
rect 38444 7476 38500 7486
rect 38332 7474 38500 7476
rect 38332 7422 38446 7474
rect 38498 7422 38500 7474
rect 38332 7420 38500 7422
rect 37996 6626 38052 6636
rect 38220 6692 38276 6702
rect 38332 6692 38388 7420
rect 38444 7410 38500 7420
rect 39004 7140 39060 7982
rect 39004 7074 39060 7084
rect 38780 6802 38836 6814
rect 38780 6750 38782 6802
rect 38834 6750 38836 6802
rect 38220 6690 38388 6692
rect 38220 6638 38222 6690
rect 38274 6638 38388 6690
rect 38220 6636 38388 6638
rect 38444 6690 38500 6702
rect 38444 6638 38446 6690
rect 38498 6638 38500 6690
rect 38220 6626 38276 6636
rect 37772 6514 37828 6524
rect 37324 6066 37380 6076
rect 37436 6466 37492 6478
rect 37436 6414 37438 6466
rect 37490 6414 37492 6466
rect 37436 5348 37492 6414
rect 37660 6466 37716 6478
rect 37660 6414 37662 6466
rect 37714 6414 37716 6466
rect 37660 6356 37716 6414
rect 37996 6468 38052 6478
rect 37996 6374 38052 6412
rect 37660 6300 37940 6356
rect 37884 6244 37940 6300
rect 38444 6244 38500 6638
rect 37884 6188 38500 6244
rect 38556 6692 38612 6702
rect 38556 5796 38612 6636
rect 38780 6244 38836 6750
rect 39116 6690 39172 8764
rect 39452 8818 39508 8878
rect 39900 8932 39956 10108
rect 40684 9940 40740 9950
rect 40796 9940 40852 10444
rect 41020 9940 41076 9950
rect 40796 9938 41076 9940
rect 40796 9886 41022 9938
rect 41074 9886 41076 9938
rect 40796 9884 41076 9886
rect 39900 8866 39956 8876
rect 40012 8930 40068 8942
rect 40012 8878 40014 8930
rect 40066 8878 40068 8930
rect 39452 8766 39454 8818
rect 39506 8766 39508 8818
rect 39340 8146 39396 8158
rect 39340 8094 39342 8146
rect 39394 8094 39396 8146
rect 39340 7588 39396 8094
rect 39116 6638 39118 6690
rect 39170 6638 39172 6690
rect 39116 6626 39172 6638
rect 39228 7532 39396 7588
rect 39452 8036 39508 8766
rect 39228 6244 39284 7532
rect 39340 7362 39396 7374
rect 39340 7310 39342 7362
rect 39394 7310 39396 7362
rect 39340 6804 39396 7310
rect 39452 6804 39508 7980
rect 39564 8820 39620 8830
rect 39564 7474 39620 8764
rect 40012 8708 40068 8878
rect 40348 8932 40404 8942
rect 40348 8818 40404 8876
rect 40348 8766 40350 8818
rect 40402 8766 40404 8818
rect 40348 8754 40404 8766
rect 40012 8642 40068 8652
rect 40460 8372 40516 8382
rect 40012 8260 40068 8270
rect 39676 8204 39956 8260
rect 39676 8146 39732 8204
rect 39676 8094 39678 8146
rect 39730 8094 39732 8146
rect 39676 8082 39732 8094
rect 39900 7924 39956 8204
rect 40012 8258 40292 8260
rect 40012 8206 40014 8258
rect 40066 8206 40292 8258
rect 40012 8204 40292 8206
rect 40012 8194 40068 8204
rect 40124 8034 40180 8046
rect 40124 7982 40126 8034
rect 40178 7982 40180 8034
rect 39900 7868 40068 7924
rect 39564 7422 39566 7474
rect 39618 7422 39620 7474
rect 39564 7410 39620 7422
rect 39900 7588 39956 7598
rect 39900 6916 39956 7532
rect 39900 6850 39956 6860
rect 39564 6804 39620 6814
rect 39452 6748 39564 6804
rect 39340 6710 39396 6748
rect 38780 6188 39284 6244
rect 39452 6580 39508 6590
rect 38892 6020 38948 6030
rect 38556 5730 38612 5740
rect 38668 5794 38724 5806
rect 38668 5742 38670 5794
rect 38722 5742 38724 5794
rect 38668 5684 38724 5742
rect 38668 5618 38724 5628
rect 37436 5282 37492 5292
rect 37660 5348 37716 5358
rect 37660 5254 37716 5292
rect 38892 5346 38948 5964
rect 39004 5684 39060 6188
rect 39452 6130 39508 6524
rect 39452 6078 39454 6130
rect 39506 6078 39508 6130
rect 39452 6066 39508 6078
rect 39116 5908 39172 5918
rect 39340 5908 39396 5918
rect 39116 5906 39340 5908
rect 39116 5854 39118 5906
rect 39170 5854 39340 5906
rect 39116 5852 39340 5854
rect 39116 5842 39172 5852
rect 39340 5842 39396 5852
rect 39004 5628 39172 5684
rect 38892 5294 38894 5346
rect 38946 5294 38948 5346
rect 38892 5282 38948 5294
rect 37772 5124 37828 5134
rect 36764 5122 37156 5124
rect 36764 5070 37102 5122
rect 37154 5070 37156 5122
rect 36764 5068 37156 5070
rect 36316 4562 36708 4564
rect 36316 4510 36318 4562
rect 36370 4510 36708 4562
rect 36316 4508 36708 4510
rect 36092 4470 36148 4508
rect 36316 4498 36372 4508
rect 35980 4386 36036 4396
rect 35980 4228 36036 4238
rect 35868 4226 36036 4228
rect 35868 4174 35982 4226
rect 36034 4174 36036 4226
rect 35868 4172 36036 4174
rect 35980 4162 36036 4172
rect 36652 4226 36708 4508
rect 36652 4174 36654 4226
rect 36706 4174 36708 4226
rect 36652 4162 36708 4174
rect 35196 3948 35460 3958
rect 35756 3948 36036 4004
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35196 3882 35460 3892
rect 35084 3490 35140 3500
rect 35980 3442 36036 3948
rect 36204 3556 36260 3566
rect 36204 3462 36260 3500
rect 35980 3390 35982 3442
rect 36034 3390 36036 3442
rect 35980 3378 36036 3390
rect 36764 3388 36820 5068
rect 37100 5058 37156 5068
rect 37324 5122 37828 5124
rect 37324 5070 37774 5122
rect 37826 5070 37828 5122
rect 37324 5068 37828 5070
rect 37324 5010 37380 5068
rect 37772 5058 37828 5068
rect 38108 5124 38164 5134
rect 38108 5030 38164 5068
rect 37324 4958 37326 5010
rect 37378 4958 37380 5010
rect 37324 4946 37380 4958
rect 38780 5012 38836 5022
rect 38780 4918 38836 4956
rect 38220 4900 38276 4910
rect 38220 4898 38724 4900
rect 38220 4846 38222 4898
rect 38274 4846 38724 4898
rect 38220 4844 38724 4846
rect 38220 4834 38276 4844
rect 38668 4452 38724 4844
rect 38892 4898 38948 4910
rect 38892 4846 38894 4898
rect 38946 4846 38948 4898
rect 38780 4452 38836 4462
rect 38668 4450 38836 4452
rect 38668 4398 38782 4450
rect 38834 4398 38836 4450
rect 38668 4396 38836 4398
rect 38780 4386 38836 4396
rect 38332 4228 38388 4238
rect 36428 3332 36820 3388
rect 36988 3666 37044 3678
rect 36988 3614 36990 3666
rect 37042 3614 37044 3666
rect 35644 924 36036 980
rect 35644 800 35700 924
rect 0 0 112 800
rect 672 0 784 800
rect 1344 0 1456 800
rect 2016 0 2128 800
rect 2688 0 2800 800
rect 3360 0 3472 800
rect 4032 0 4144 800
rect 4704 0 4816 800
rect 5376 0 5488 800
rect 6048 0 6160 800
rect 6720 0 6832 800
rect 7392 0 7504 800
rect 8064 0 8176 800
rect 8736 0 8848 800
rect 9408 0 9520 800
rect 10080 0 10192 800
rect 10752 0 10864 800
rect 11424 0 11536 800
rect 12096 0 12208 800
rect 12768 0 12880 800
rect 13440 0 13552 800
rect 14112 0 14224 800
rect 14784 0 14896 800
rect 15456 0 15568 800
rect 16128 0 16240 800
rect 16800 0 16912 800
rect 17472 0 17584 800
rect 18144 0 18256 800
rect 18816 0 18928 800
rect 19488 0 19600 800
rect 20160 0 20272 800
rect 20832 0 20944 800
rect 22176 0 22288 800
rect 22848 0 22960 800
rect 23520 0 23632 800
rect 24864 0 24976 800
rect 26208 0 26320 800
rect 26880 0 26992 800
rect 29568 0 29680 800
rect 30240 0 30352 800
rect 30912 0 31024 800
rect 31584 0 31696 800
rect 32928 0 33040 800
rect 33600 0 33712 800
rect 35616 0 35728 800
rect 35980 756 36036 924
rect 36428 756 36484 3332
rect 36988 800 37044 3614
rect 37660 3668 37716 3678
rect 37660 800 37716 3612
rect 38332 800 38388 4172
rect 38892 3332 38948 4846
rect 39116 3554 39172 5628
rect 39452 5124 39508 5134
rect 39564 5124 39620 6748
rect 39788 6356 39844 6366
rect 39788 6132 39844 6300
rect 39788 6018 39844 6076
rect 39788 5966 39790 6018
rect 39842 5966 39844 6018
rect 39788 5954 39844 5966
rect 39900 5908 39956 5918
rect 39900 5814 39956 5852
rect 39452 5122 39620 5124
rect 39452 5070 39454 5122
rect 39506 5070 39620 5122
rect 39452 5068 39620 5070
rect 39452 5058 39508 5068
rect 39564 4338 39620 5068
rect 39564 4286 39566 4338
rect 39618 4286 39620 4338
rect 39564 4274 39620 4286
rect 39900 5348 39956 5358
rect 39116 3502 39118 3554
rect 39170 3502 39172 3554
rect 39116 3490 39172 3502
rect 38892 3266 38948 3276
rect 39004 3444 39060 3454
rect 39004 800 39060 3388
rect 39900 2884 39956 5292
rect 40012 3554 40068 7868
rect 40124 6804 40180 7982
rect 40236 7476 40292 8204
rect 40236 7410 40292 7420
rect 40460 8258 40516 8316
rect 40460 8206 40462 8258
rect 40514 8206 40516 8258
rect 40348 7364 40404 7374
rect 40348 7270 40404 7308
rect 40236 7250 40292 7262
rect 40236 7198 40238 7250
rect 40290 7198 40292 7250
rect 40236 7028 40292 7198
rect 40236 6962 40292 6972
rect 40124 6748 40292 6804
rect 40236 6692 40292 6748
rect 40236 6636 40404 6692
rect 40124 6580 40180 6590
rect 40124 6486 40180 6524
rect 40236 6468 40292 6478
rect 40236 6374 40292 6412
rect 40348 6244 40404 6636
rect 40236 6188 40404 6244
rect 40124 5908 40180 5918
rect 40124 5814 40180 5852
rect 40124 5684 40180 5694
rect 40124 5234 40180 5628
rect 40124 5182 40126 5234
rect 40178 5182 40180 5234
rect 40124 5170 40180 5182
rect 40236 5012 40292 6188
rect 40460 6132 40516 8206
rect 40684 8146 40740 9884
rect 41020 9874 41076 9884
rect 41132 9268 41188 10782
rect 41356 12292 41412 12302
rect 41356 11844 41412 12236
rect 41356 10834 41412 11788
rect 41468 12178 41524 12190
rect 41468 12126 41470 12178
rect 41522 12126 41524 12178
rect 41468 11620 41524 12126
rect 41468 11554 41524 11564
rect 41580 11956 41636 12460
rect 41916 12292 41972 12302
rect 41916 12198 41972 12236
rect 42028 12068 42084 12908
rect 41356 10782 41358 10834
rect 41410 10782 41412 10834
rect 41356 10770 41412 10782
rect 41468 11284 41524 11294
rect 41468 10834 41524 11228
rect 41468 10782 41470 10834
rect 41522 10782 41524 10834
rect 41468 10770 41524 10782
rect 41580 10834 41636 11900
rect 41580 10782 41582 10834
rect 41634 10782 41636 10834
rect 41580 10770 41636 10782
rect 41916 12012 42084 12068
rect 41916 10834 41972 12012
rect 41916 10782 41918 10834
rect 41970 10782 41972 10834
rect 41916 9940 41972 10782
rect 42140 10610 42196 13132
rect 42252 12740 42308 13468
rect 42700 13412 42756 13582
rect 43372 13636 43428 13694
rect 43372 13570 43428 13580
rect 42700 13346 42756 13356
rect 43148 13524 43204 13534
rect 42700 13188 42756 13198
rect 42700 13094 42756 13132
rect 42252 12674 42308 12684
rect 42588 12850 42644 12862
rect 42588 12798 42590 12850
rect 42642 12798 42644 12850
rect 42588 12180 42644 12798
rect 42812 12180 42868 12190
rect 42588 12124 42812 12180
rect 42812 12086 42868 12124
rect 43148 12178 43204 13468
rect 43596 12962 43652 13804
rect 43708 13794 43764 13804
rect 43596 12910 43598 12962
rect 43650 12910 43652 12962
rect 43596 12898 43652 12910
rect 43820 13412 43876 14366
rect 44156 14196 44212 15036
rect 44268 14532 44324 14542
rect 44268 14438 44324 14476
rect 44156 14130 44212 14140
rect 43260 12292 43316 12302
rect 43260 12198 43316 12236
rect 43148 12126 43150 12178
rect 43202 12126 43204 12178
rect 43148 12114 43204 12126
rect 43820 12180 43876 13356
rect 43932 13634 43988 13646
rect 43932 13582 43934 13634
rect 43986 13582 43988 13634
rect 43932 12740 43988 13582
rect 44380 13524 44436 13534
rect 44156 13186 44212 13198
rect 44156 13134 44158 13186
rect 44210 13134 44212 13186
rect 43932 12684 44100 12740
rect 43932 12180 43988 12190
rect 43820 12124 43932 12180
rect 43932 12114 43988 12124
rect 44044 12178 44100 12684
rect 44156 12516 44212 13134
rect 44380 12962 44436 13468
rect 44380 12910 44382 12962
rect 44434 12910 44436 12962
rect 44380 12898 44436 12910
rect 44156 12460 44436 12516
rect 44044 12126 44046 12178
rect 44098 12126 44100 12178
rect 44044 12114 44100 12126
rect 44380 12180 44436 12460
rect 44492 12404 44548 17052
rect 44604 15988 44660 17388
rect 44828 17220 44884 18398
rect 44940 18116 44996 19294
rect 45052 19010 45108 19022
rect 45052 18958 45054 19010
rect 45106 18958 45108 19010
rect 45052 18900 45108 18958
rect 45052 18834 45108 18844
rect 45276 19010 45332 19022
rect 45276 18958 45278 19010
rect 45330 18958 45332 19010
rect 45276 18564 45332 18958
rect 45500 18788 45556 19964
rect 45612 20132 45668 20142
rect 45612 19234 45668 20076
rect 46060 19908 46116 19918
rect 46060 19906 46564 19908
rect 46060 19854 46062 19906
rect 46114 19854 46564 19906
rect 46060 19852 46564 19854
rect 46060 19842 46116 19852
rect 45612 19182 45614 19234
rect 45666 19182 45668 19234
rect 45612 19170 45668 19182
rect 44940 18050 44996 18060
rect 45052 18508 45332 18564
rect 45388 18732 45556 18788
rect 45612 18900 45668 18910
rect 44940 17892 44996 17902
rect 44940 17778 44996 17836
rect 44940 17726 44942 17778
rect 44994 17726 44996 17778
rect 44940 17714 44996 17726
rect 45052 17444 45108 18508
rect 45276 18340 45332 18350
rect 45276 18246 45332 18284
rect 45388 17666 45444 18732
rect 45612 18674 45668 18844
rect 45612 18622 45614 18674
rect 45666 18622 45668 18674
rect 45612 18610 45668 18622
rect 46508 18674 46564 19852
rect 46508 18622 46510 18674
rect 46562 18622 46564 18674
rect 46508 18610 46564 18622
rect 45836 18564 45892 18574
rect 45836 18470 45892 18508
rect 46060 18452 46116 18462
rect 46060 18358 46116 18396
rect 46620 18452 46676 20748
rect 47180 18676 47236 18686
rect 47180 18582 47236 18620
rect 46620 18386 46676 18396
rect 46732 18450 46788 18462
rect 46732 18398 46734 18450
rect 46786 18398 46788 18450
rect 45388 17614 45390 17666
rect 45442 17614 45444 17666
rect 45388 17602 45444 17614
rect 45724 18338 45780 18350
rect 45724 18286 45726 18338
rect 45778 18286 45780 18338
rect 45052 17378 45108 17388
rect 44828 16882 44884 17164
rect 44828 16830 44830 16882
rect 44882 16830 44884 16882
rect 44716 16770 44772 16782
rect 44716 16718 44718 16770
rect 44770 16718 44772 16770
rect 44716 16212 44772 16718
rect 44716 16146 44772 16156
rect 44604 15932 44772 15988
rect 44604 15202 44660 15214
rect 44604 15150 44606 15202
rect 44658 15150 44660 15202
rect 44604 14756 44660 15150
rect 44604 14690 44660 14700
rect 44492 12348 44660 12404
rect 44492 12180 44548 12190
rect 44380 12178 44548 12180
rect 44380 12126 44494 12178
rect 44546 12126 44548 12178
rect 44380 12124 44548 12126
rect 44492 12114 44548 12124
rect 42140 10558 42142 10610
rect 42194 10558 42196 10610
rect 42140 10546 42196 10558
rect 42252 12066 42308 12078
rect 42252 12014 42254 12066
rect 42306 12014 42308 12066
rect 42252 10164 42308 12014
rect 42700 11620 42756 11630
rect 42700 10834 42756 11564
rect 43596 11396 43652 11406
rect 42812 11284 42868 11294
rect 42812 11190 42868 11228
rect 42700 10782 42702 10834
rect 42754 10782 42756 10834
rect 42700 10770 42756 10782
rect 43372 10724 43428 10734
rect 43372 10630 43428 10668
rect 43484 10612 43540 10622
rect 43484 10518 43540 10556
rect 42252 10098 42308 10108
rect 42700 10276 42756 10286
rect 41916 9874 41972 9884
rect 41132 9202 41188 9212
rect 41356 9826 41412 9838
rect 41356 9774 41358 9826
rect 41410 9774 41412 9826
rect 41132 8932 41188 8942
rect 41356 8932 41412 9774
rect 42140 9716 42196 9726
rect 41580 9714 42196 9716
rect 41580 9662 42142 9714
rect 42194 9662 42196 9714
rect 41580 9660 42196 9662
rect 41580 9266 41636 9660
rect 42140 9650 42196 9660
rect 41580 9214 41582 9266
rect 41634 9214 41636 9266
rect 41580 9202 41636 9214
rect 41916 9268 41972 9278
rect 41916 9174 41972 9212
rect 42476 9154 42532 9166
rect 42476 9102 42478 9154
rect 42530 9102 42532 9154
rect 41468 9044 41524 9054
rect 41468 8950 41524 8988
rect 41692 9042 41748 9054
rect 41692 8990 41694 9042
rect 41746 8990 41748 9042
rect 41132 8930 41300 8932
rect 41132 8878 41134 8930
rect 41186 8878 41300 8930
rect 41132 8876 41300 8878
rect 41132 8866 41188 8876
rect 41244 8484 41300 8876
rect 41356 8866 41412 8876
rect 41692 8820 41748 8990
rect 41692 8754 41748 8764
rect 42476 8484 42532 9102
rect 41244 8428 41860 8484
rect 40684 8094 40686 8146
rect 40738 8094 40740 8146
rect 40684 8082 40740 8094
rect 41356 8258 41412 8270
rect 41356 8206 41358 8258
rect 41410 8206 41412 8258
rect 40796 8036 40852 8046
rect 40796 8034 40964 8036
rect 40796 7982 40798 8034
rect 40850 7982 40964 8034
rect 40796 7980 40964 7982
rect 40796 7970 40852 7980
rect 40908 7586 40964 7980
rect 40908 7534 40910 7586
rect 40962 7534 40964 7586
rect 40572 6690 40628 6702
rect 40572 6638 40574 6690
rect 40626 6638 40628 6690
rect 40572 6580 40628 6638
rect 40572 6514 40628 6524
rect 40348 6076 40516 6132
rect 40348 6018 40404 6076
rect 40348 5966 40350 6018
rect 40402 5966 40404 6018
rect 40348 5954 40404 5966
rect 40908 5906 40964 7534
rect 41020 7252 41076 7262
rect 41020 7158 41076 7196
rect 41244 7140 41300 7150
rect 40908 5854 40910 5906
rect 40962 5854 40964 5906
rect 40908 5842 40964 5854
rect 41132 6916 41188 6926
rect 41020 5684 41076 5694
rect 40460 5236 40516 5246
rect 40124 4956 40292 5012
rect 40348 5124 40404 5134
rect 40124 4450 40180 4956
rect 40236 4564 40292 4574
rect 40236 4470 40292 4508
rect 40124 4398 40126 4450
rect 40178 4398 40180 4450
rect 40124 4386 40180 4398
rect 40012 3502 40014 3554
rect 40066 3502 40068 3554
rect 40012 3490 40068 3502
rect 39676 2828 39956 2884
rect 39676 800 39732 2828
rect 40348 800 40404 5068
rect 40460 4562 40516 5180
rect 40460 4510 40462 4562
rect 40514 4510 40516 4562
rect 40460 4498 40516 4510
rect 40796 3668 40852 3678
rect 40796 3574 40852 3612
rect 41020 800 41076 5628
rect 41132 4338 41188 6860
rect 41132 4286 41134 4338
rect 41186 4286 41188 4338
rect 41132 4274 41188 4286
rect 41244 3556 41300 7084
rect 41356 6356 41412 8206
rect 41468 7474 41524 7486
rect 41468 7422 41470 7474
rect 41522 7422 41524 7474
rect 41468 6804 41524 7422
rect 41468 6738 41524 6748
rect 41356 6290 41412 6300
rect 41580 6466 41636 6478
rect 41580 6414 41582 6466
rect 41634 6414 41636 6466
rect 41580 5124 41636 6414
rect 41580 5058 41636 5068
rect 41244 3490 41300 3500
rect 41692 4900 41748 4910
rect 41692 800 41748 4844
rect 41804 4340 41860 8428
rect 42476 8418 42532 8428
rect 42028 8204 42420 8260
rect 41916 8148 41972 8158
rect 41916 8054 41972 8092
rect 41916 7924 41972 7934
rect 42028 7924 42084 8204
rect 42364 8146 42420 8204
rect 42364 8094 42366 8146
rect 42418 8094 42420 8146
rect 42364 8082 42420 8094
rect 42476 8146 42532 8158
rect 42476 8094 42478 8146
rect 42530 8094 42532 8146
rect 41972 7868 42084 7924
rect 41916 7858 41972 7868
rect 42028 6020 42084 7868
rect 42140 8034 42196 8046
rect 42140 7982 42142 8034
rect 42194 7982 42196 8034
rect 42140 7924 42196 7982
rect 42140 7858 42196 7868
rect 42364 7700 42420 7710
rect 42140 7644 42364 7700
rect 42140 7586 42196 7644
rect 42364 7634 42420 7644
rect 42140 7534 42142 7586
rect 42194 7534 42196 7586
rect 42140 7522 42196 7534
rect 42476 6356 42532 8094
rect 42700 7588 42756 10220
rect 43484 10052 43540 10062
rect 43596 10052 43652 11340
rect 44268 11172 44324 11182
rect 44156 11170 44324 11172
rect 44156 11118 44270 11170
rect 44322 11118 44324 11170
rect 44156 11116 44324 11118
rect 43932 10836 43988 10846
rect 43932 10722 43988 10780
rect 43932 10670 43934 10722
rect 43986 10670 43988 10722
rect 43932 10658 43988 10670
rect 43540 9996 43652 10052
rect 43708 10610 43764 10622
rect 43708 10558 43710 10610
rect 43762 10558 43764 10610
rect 43484 9986 43540 9996
rect 42812 8932 42868 8942
rect 42812 8838 42868 8876
rect 43260 8930 43316 8942
rect 43260 8878 43262 8930
rect 43314 8878 43316 8930
rect 42924 8820 42980 8830
rect 42924 8818 43092 8820
rect 42924 8766 42926 8818
rect 42978 8766 43092 8818
rect 42924 8764 43092 8766
rect 42924 8754 42980 8764
rect 42924 8146 42980 8158
rect 42924 8094 42926 8146
rect 42978 8094 42980 8146
rect 42812 8034 42868 8046
rect 42812 7982 42814 8034
rect 42866 7982 42868 8034
rect 42812 7700 42868 7982
rect 42812 7634 42868 7644
rect 42700 7522 42756 7532
rect 42476 6290 42532 6300
rect 42700 7364 42756 7374
rect 42028 5964 42196 6020
rect 41804 4274 41860 4284
rect 41916 5796 41972 5806
rect 41916 3388 41972 5740
rect 42028 5794 42084 5806
rect 42028 5742 42030 5794
rect 42082 5742 42084 5794
rect 42028 5348 42084 5742
rect 42028 5282 42084 5292
rect 42140 4564 42196 5964
rect 42252 5908 42308 5918
rect 42252 5236 42308 5852
rect 42252 5234 42644 5236
rect 42252 5182 42254 5234
rect 42306 5182 42644 5234
rect 42252 5180 42644 5182
rect 42252 5170 42308 5180
rect 42588 5122 42644 5180
rect 42700 5234 42756 7308
rect 42924 7364 42980 8094
rect 42924 7298 42980 7308
rect 42700 5182 42702 5234
rect 42754 5182 42756 5234
rect 42700 5170 42756 5182
rect 42812 5796 42868 5806
rect 42588 5070 42590 5122
rect 42642 5070 42644 5122
rect 42588 5058 42644 5070
rect 42140 4498 42196 4508
rect 42700 5012 42756 5022
rect 42028 4228 42084 4238
rect 42028 4134 42084 4172
rect 42364 3668 42420 3678
rect 42364 3388 42420 3612
rect 42700 3554 42756 4956
rect 42700 3502 42702 3554
rect 42754 3502 42756 3554
rect 42700 3490 42756 3502
rect 42812 4898 42868 5740
rect 42924 5124 42980 5134
rect 42924 5010 42980 5068
rect 42924 4958 42926 5010
rect 42978 4958 42980 5010
rect 42924 4946 42980 4958
rect 42812 4846 42814 4898
rect 42866 4846 42868 4898
rect 42812 3444 42868 4846
rect 43036 4452 43092 8764
rect 43036 4386 43092 4396
rect 43148 8708 43204 8718
rect 43148 3780 43204 8652
rect 43260 8372 43316 8878
rect 43372 8820 43428 8830
rect 43708 8820 43764 10558
rect 44156 10164 44212 11116
rect 44268 11106 44324 11116
rect 44604 10948 44660 12348
rect 44268 10892 44660 10948
rect 44268 10724 44324 10892
rect 44268 10630 44324 10668
rect 44716 10836 44772 15932
rect 44828 15426 44884 16830
rect 45500 16996 45556 17006
rect 45500 16772 45556 16940
rect 45724 16882 45780 18286
rect 46396 18340 46452 18350
rect 46396 18246 46452 18284
rect 46060 17780 46116 17790
rect 45724 16830 45726 16882
rect 45778 16830 45780 16882
rect 45724 16818 45780 16830
rect 45948 17724 46060 17780
rect 45388 16770 45556 16772
rect 45388 16718 45502 16770
rect 45554 16718 45556 16770
rect 45388 16716 45556 16718
rect 44940 16322 44996 16334
rect 44940 16270 44942 16322
rect 44994 16270 44996 16322
rect 44940 15764 44996 16270
rect 44940 15698 44996 15708
rect 45164 16098 45220 16110
rect 45164 16046 45166 16098
rect 45218 16046 45220 16098
rect 44828 15374 44830 15426
rect 44882 15374 44884 15426
rect 44828 15362 44884 15374
rect 45164 15148 45220 16046
rect 44828 15092 45220 15148
rect 44828 13412 44884 15092
rect 44940 14868 44996 14878
rect 44940 14644 44996 14812
rect 44940 14642 45332 14644
rect 44940 14590 44942 14642
rect 44994 14590 45332 14642
rect 44940 14588 45332 14590
rect 44940 14578 44996 14588
rect 44828 13346 44884 13356
rect 45276 14530 45332 14588
rect 45276 14478 45278 14530
rect 45330 14478 45332 14530
rect 45164 13300 45220 13310
rect 44828 12964 44884 12974
rect 44828 12870 44884 12908
rect 44940 12852 44996 12862
rect 44940 12758 44996 12796
rect 44828 11396 44884 11406
rect 44828 11302 44884 11340
rect 45164 11060 45220 13244
rect 45276 12962 45332 14478
rect 45388 13300 45444 16716
rect 45500 16706 45556 16716
rect 45612 16212 45668 16222
rect 45612 16098 45668 16156
rect 45948 16100 46004 17724
rect 46060 17714 46116 17724
rect 46060 17554 46116 17566
rect 46060 17502 46062 17554
rect 46114 17502 46116 17554
rect 46060 17106 46116 17502
rect 46060 17054 46062 17106
rect 46114 17054 46116 17106
rect 46060 17042 46116 17054
rect 46284 16996 46340 17006
rect 46732 16996 46788 18398
rect 47516 18450 47572 20860
rect 47964 20132 48020 20142
rect 47964 19458 48020 20076
rect 48188 19908 48244 19918
rect 47964 19406 47966 19458
rect 48018 19406 48020 19458
rect 47964 19394 48020 19406
rect 48076 19906 48244 19908
rect 48076 19854 48190 19906
rect 48242 19854 48244 19906
rect 48076 19852 48244 19854
rect 48076 19012 48132 19852
rect 48188 19842 48244 19852
rect 47516 18398 47518 18450
rect 47570 18398 47572 18450
rect 47516 18228 47572 18398
rect 47852 18562 47908 18574
rect 47852 18510 47854 18562
rect 47906 18510 47908 18562
rect 47852 18452 47908 18510
rect 47852 18386 47908 18396
rect 47516 18162 47572 18172
rect 47628 18116 47684 18126
rect 46956 16996 47012 17006
rect 46732 16940 46956 16996
rect 46172 16884 46228 16894
rect 46172 16790 46228 16828
rect 46284 16882 46340 16940
rect 46284 16830 46286 16882
rect 46338 16830 46340 16882
rect 46284 16818 46340 16830
rect 45612 16046 45614 16098
rect 45666 16046 45668 16098
rect 45612 16034 45668 16046
rect 45836 16098 46004 16100
rect 45836 16046 45950 16098
rect 46002 16046 46004 16098
rect 45836 16044 46004 16046
rect 45836 14532 45892 16044
rect 45948 16034 46004 16044
rect 46060 16772 46116 16782
rect 45948 15316 46004 15326
rect 45948 15222 46004 15260
rect 46060 14642 46116 16716
rect 46844 16772 46900 16782
rect 46844 16678 46900 16716
rect 46732 16658 46788 16670
rect 46732 16606 46734 16658
rect 46786 16606 46788 16658
rect 46396 16212 46452 16222
rect 46396 15314 46452 16156
rect 46732 15428 46788 16606
rect 46956 16210 47012 16940
rect 47516 16994 47572 17006
rect 47516 16942 47518 16994
rect 47570 16942 47572 16994
rect 47292 16884 47348 16894
rect 47292 16790 47348 16828
rect 46956 16158 46958 16210
rect 47010 16158 47012 16210
rect 46956 16146 47012 16158
rect 47516 16212 47572 16942
rect 47628 16994 47684 18060
rect 48076 17556 48132 18956
rect 48188 18452 48244 18462
rect 48300 18452 48356 21532
rect 48188 18450 48356 18452
rect 48188 18398 48190 18450
rect 48242 18398 48356 18450
rect 48188 18396 48356 18398
rect 48188 18386 48244 18396
rect 48188 17780 48244 17790
rect 48188 17686 48244 17724
rect 48076 17500 48244 17556
rect 48188 17108 48244 17500
rect 48300 17332 48356 18396
rect 48300 17266 48356 17276
rect 48188 17052 48356 17108
rect 47628 16942 47630 16994
rect 47682 16942 47684 16994
rect 47628 16930 47684 16942
rect 48076 16996 48132 17006
rect 48076 16902 48132 16940
rect 47516 16146 47572 16156
rect 46732 15362 46788 15372
rect 47292 15986 47348 15998
rect 47292 15934 47294 15986
rect 47346 15934 47348 15986
rect 46396 15262 46398 15314
rect 46450 15262 46452 15314
rect 46396 15250 46452 15262
rect 47292 15316 47348 15934
rect 47852 15874 47908 15886
rect 47852 15822 47854 15874
rect 47906 15822 47908 15874
rect 47292 15250 47348 15260
rect 47404 15426 47460 15438
rect 47404 15374 47406 15426
rect 47458 15374 47460 15426
rect 47404 15092 47460 15374
rect 47852 15148 47908 15822
rect 46060 14590 46062 14642
rect 46114 14590 46116 14642
rect 46060 14578 46116 14590
rect 47068 14644 47124 14654
rect 45836 13748 45892 14476
rect 47068 13970 47124 14588
rect 47068 13918 47070 13970
rect 47122 13918 47124 13970
rect 47068 13906 47124 13918
rect 46284 13748 46340 13758
rect 45836 13746 46340 13748
rect 45836 13694 46286 13746
rect 46338 13694 46340 13746
rect 45836 13692 46340 13694
rect 46284 13682 46340 13692
rect 46732 13748 46788 13758
rect 46732 13654 46788 13692
rect 47404 13748 47460 15036
rect 45388 13234 45444 13244
rect 45276 12910 45278 12962
rect 45330 12910 45332 12962
rect 45276 11396 45332 12910
rect 46060 12852 46116 12862
rect 46060 12758 46116 12796
rect 47404 12290 47460 13692
rect 47740 15092 47908 15148
rect 47740 14644 47796 15092
rect 48188 14644 48244 14654
rect 47740 14642 48244 14644
rect 47740 14590 48190 14642
rect 48242 14590 48244 14642
rect 47740 14588 48244 14590
rect 47740 13746 47796 14588
rect 48188 14578 48244 14588
rect 47740 13694 47742 13746
rect 47794 13694 47796 13746
rect 47740 13682 47796 13694
rect 47964 13636 48020 13646
rect 48300 13636 48356 17052
rect 47964 13634 48356 13636
rect 47964 13582 47966 13634
rect 48018 13582 48356 13634
rect 47964 13580 48356 13582
rect 47516 13524 47572 13534
rect 47964 13524 48020 13580
rect 47516 13522 47908 13524
rect 47516 13470 47518 13522
rect 47570 13470 47908 13522
rect 47516 13468 47908 13470
rect 47516 13458 47572 13468
rect 47852 13188 47908 13468
rect 47964 13458 48020 13468
rect 47852 13132 48244 13188
rect 47964 12402 48020 13132
rect 48188 13074 48244 13132
rect 48188 13022 48190 13074
rect 48242 13022 48244 13074
rect 48188 13010 48244 13022
rect 47964 12350 47966 12402
rect 48018 12350 48020 12402
rect 47964 12338 48020 12350
rect 47404 12238 47406 12290
rect 47458 12238 47460 12290
rect 47404 12226 47460 12238
rect 46508 12180 46564 12190
rect 45948 12066 46004 12078
rect 45948 12014 45950 12066
rect 46002 12014 46004 12066
rect 45836 11956 45892 11966
rect 45276 11330 45332 11340
rect 45724 11954 45892 11956
rect 45724 11902 45838 11954
rect 45890 11902 45892 11954
rect 45724 11900 45892 11902
rect 44604 10612 44660 10622
rect 44716 10612 44772 10780
rect 44940 11004 45220 11060
rect 45612 11282 45668 11294
rect 45612 11230 45614 11282
rect 45666 11230 45668 11282
rect 44604 10610 44772 10612
rect 44604 10558 44606 10610
rect 44658 10558 44772 10610
rect 44604 10556 44772 10558
rect 44828 10612 44884 10622
rect 44604 10546 44660 10556
rect 44828 10518 44884 10556
rect 44828 10388 44884 10398
rect 44940 10388 44996 11004
rect 45052 10836 45108 10846
rect 45612 10836 45668 11230
rect 45052 10834 45668 10836
rect 45052 10782 45054 10834
rect 45106 10782 45668 10834
rect 45052 10780 45668 10782
rect 45052 10770 45108 10780
rect 44828 10386 44996 10388
rect 44828 10334 44830 10386
rect 44882 10334 44996 10386
rect 44828 10332 44996 10334
rect 45388 10498 45444 10510
rect 45388 10446 45390 10498
rect 45442 10446 45444 10498
rect 44828 10322 44884 10332
rect 44156 10108 44436 10164
rect 44268 9940 44324 9950
rect 43820 9938 44324 9940
rect 43820 9886 44270 9938
rect 44322 9886 44324 9938
rect 43820 9884 44324 9886
rect 43820 9154 43876 9884
rect 44268 9874 44324 9884
rect 43820 9102 43822 9154
rect 43874 9102 43876 9154
rect 43820 9090 43876 9102
rect 44156 9268 44212 9278
rect 43372 8818 43652 8820
rect 43372 8766 43374 8818
rect 43426 8766 43652 8818
rect 43372 8764 43652 8766
rect 43372 8754 43428 8764
rect 43260 8306 43316 8316
rect 43484 7364 43540 7374
rect 43484 6802 43540 7308
rect 43484 6750 43486 6802
rect 43538 6750 43540 6802
rect 43484 6738 43540 6750
rect 43596 6356 43652 8764
rect 43708 8726 43764 8764
rect 44156 9042 44212 9212
rect 44156 8990 44158 9042
rect 44210 8990 44212 9042
rect 44156 8596 44212 8990
rect 44156 8530 44212 8540
rect 44268 9154 44324 9166
rect 44268 9102 44270 9154
rect 44322 9102 44324 9154
rect 44156 8372 44212 8382
rect 44156 8278 44212 8316
rect 43820 8146 43876 8158
rect 43820 8094 43822 8146
rect 43874 8094 43876 8146
rect 43708 7924 43764 7934
rect 43708 6578 43764 7868
rect 43820 6916 43876 8094
rect 43820 6850 43876 6860
rect 43932 8146 43988 8158
rect 43932 8094 43934 8146
rect 43986 8094 43988 8146
rect 43932 8036 43988 8094
rect 44156 8148 44212 8158
rect 43708 6526 43710 6578
rect 43762 6526 43764 6578
rect 43708 6514 43764 6526
rect 43932 6578 43988 7980
rect 43932 6526 43934 6578
rect 43986 6526 43988 6578
rect 43820 6468 43876 6478
rect 43596 6300 43764 6356
rect 43708 5684 43764 6300
rect 43820 5906 43876 6412
rect 43820 5854 43822 5906
rect 43874 5854 43876 5906
rect 43820 5842 43876 5854
rect 43708 5628 43876 5684
rect 43260 5236 43316 5246
rect 43260 5122 43316 5180
rect 43260 5070 43262 5122
rect 43314 5070 43316 5122
rect 43260 5058 43316 5070
rect 43708 5122 43764 5134
rect 43708 5070 43710 5122
rect 43762 5070 43764 5122
rect 43708 4564 43764 5070
rect 43708 4498 43764 4508
rect 43820 4450 43876 5628
rect 43932 5124 43988 6526
rect 44044 8034 44100 8046
rect 44044 7982 44046 8034
rect 44098 7982 44100 8034
rect 44044 6466 44100 7982
rect 44156 7364 44212 8092
rect 44268 8036 44324 9102
rect 44268 7942 44324 7980
rect 44268 7364 44324 7374
rect 44156 7362 44324 7364
rect 44156 7310 44270 7362
rect 44322 7310 44324 7362
rect 44156 7308 44324 7310
rect 44380 7364 44436 10108
rect 44940 9714 44996 9726
rect 44940 9662 44942 9714
rect 44994 9662 44996 9714
rect 44940 9268 44996 9662
rect 45052 9604 45108 9614
rect 45276 9604 45332 9614
rect 45052 9510 45108 9548
rect 45164 9602 45332 9604
rect 45164 9550 45278 9602
rect 45330 9550 45332 9602
rect 45164 9548 45332 9550
rect 44940 9202 44996 9212
rect 44716 9156 44772 9166
rect 44492 9044 44548 9054
rect 44716 9044 44772 9100
rect 44940 9044 44996 9054
rect 45164 9044 45220 9548
rect 45276 9538 45332 9548
rect 45388 9268 45444 10446
rect 45500 10388 45556 10398
rect 45500 10386 45668 10388
rect 45500 10334 45502 10386
rect 45554 10334 45668 10386
rect 45500 10332 45668 10334
rect 45500 10322 45556 10332
rect 45388 9212 45556 9268
rect 44492 9042 44660 9044
rect 44492 8990 44494 9042
rect 44546 8990 44660 9042
rect 44492 8988 44660 8990
rect 44492 8978 44548 8988
rect 44604 7476 44660 8988
rect 44716 9042 44884 9044
rect 44716 8990 44718 9042
rect 44770 8990 44884 9042
rect 44716 8988 44884 8990
rect 44716 8978 44772 8988
rect 44716 7476 44772 7486
rect 44604 7474 44772 7476
rect 44604 7422 44718 7474
rect 44770 7422 44772 7474
rect 44604 7420 44772 7422
rect 44828 7476 44884 8988
rect 44940 9042 45220 9044
rect 44940 8990 44942 9042
rect 44994 8990 45220 9042
rect 44940 8988 45220 8990
rect 45388 9044 45444 9054
rect 44940 8978 44996 8988
rect 45276 8820 45332 8830
rect 45052 8818 45332 8820
rect 45052 8766 45278 8818
rect 45330 8766 45332 8818
rect 45052 8764 45332 8766
rect 44940 8484 44996 8494
rect 44940 8036 44996 8428
rect 45052 8258 45108 8764
rect 45276 8754 45332 8764
rect 45052 8206 45054 8258
rect 45106 8206 45108 8258
rect 45052 8194 45108 8206
rect 45164 8596 45220 8606
rect 45388 8596 45444 8988
rect 44940 7980 45108 8036
rect 45052 7588 45108 7980
rect 45164 7700 45220 8540
rect 45276 8540 45444 8596
rect 45276 8146 45332 8540
rect 45388 8372 45444 8382
rect 45500 8372 45556 9212
rect 45444 8316 45556 8372
rect 45388 8306 45444 8316
rect 45276 8094 45278 8146
rect 45330 8094 45332 8146
rect 45276 8082 45332 8094
rect 45276 7700 45332 7710
rect 45164 7698 45332 7700
rect 45164 7646 45278 7698
rect 45330 7646 45332 7698
rect 45164 7644 45332 7646
rect 45276 7634 45332 7644
rect 45052 7532 45220 7588
rect 44940 7476 44996 7486
rect 44828 7474 44996 7476
rect 44828 7422 44942 7474
rect 44994 7422 44996 7474
rect 44828 7420 44996 7422
rect 44716 7410 44772 7420
rect 44940 7410 44996 7420
rect 44380 7308 44660 7364
rect 44044 6414 44046 6466
rect 44098 6414 44100 6466
rect 44044 5796 44100 6414
rect 44044 5730 44100 5740
rect 44156 6916 44212 6926
rect 43932 5058 43988 5068
rect 43932 4564 43988 4574
rect 43932 4470 43988 4508
rect 44156 4562 44212 6860
rect 44268 6578 44324 7308
rect 44268 6526 44270 6578
rect 44322 6526 44324 6578
rect 44268 6514 44324 6526
rect 44492 6580 44548 6590
rect 44268 5236 44324 5246
rect 44268 5122 44324 5180
rect 44268 5070 44270 5122
rect 44322 5070 44324 5122
rect 44268 5012 44324 5070
rect 44268 4946 44324 4956
rect 44156 4510 44158 4562
rect 44210 4510 44212 4562
rect 44156 4498 44212 4510
rect 43820 4398 43822 4450
rect 43874 4398 43876 4450
rect 43820 4386 43876 4398
rect 43036 3444 43092 3454
rect 42812 3442 43092 3444
rect 42812 3390 43038 3442
rect 43090 3390 43092 3442
rect 42812 3388 43092 3390
rect 41916 3332 42420 3388
rect 43036 3378 43092 3388
rect 42364 800 42420 3332
rect 43148 3220 43204 3724
rect 43932 4340 43988 4350
rect 43708 3556 43764 3566
rect 43708 3462 43764 3500
rect 43036 3164 43204 3220
rect 43036 800 43092 3164
rect 43932 2996 43988 4284
rect 44492 4338 44548 6524
rect 44604 4788 44660 7308
rect 45052 7252 45108 7262
rect 44940 6578 44996 6590
rect 44940 6526 44942 6578
rect 44994 6526 44996 6578
rect 44828 6466 44884 6478
rect 44828 6414 44830 6466
rect 44882 6414 44884 6466
rect 44828 6356 44884 6414
rect 44828 6290 44884 6300
rect 44604 4722 44660 4732
rect 44716 6244 44772 6254
rect 44716 5348 44772 6188
rect 44828 5684 44884 5694
rect 44828 5590 44884 5628
rect 44492 4286 44494 4338
rect 44546 4286 44548 4338
rect 44492 4274 44548 4286
rect 44716 4116 44772 5292
rect 43708 2940 43988 2996
rect 44380 4060 44772 4116
rect 44828 5460 44884 5470
rect 43708 800 43764 2940
rect 44380 800 44436 4060
rect 44604 3666 44660 3678
rect 44604 3614 44606 3666
rect 44658 3614 44660 3666
rect 44604 3444 44660 3614
rect 44604 3378 44660 3388
rect 44828 3388 44884 5404
rect 44940 5124 44996 6526
rect 44940 5058 44996 5068
rect 45052 5122 45108 7196
rect 45164 6244 45220 7532
rect 45388 6690 45444 6702
rect 45388 6638 45390 6690
rect 45442 6638 45444 6690
rect 45276 6580 45332 6590
rect 45388 6580 45444 6638
rect 45612 6692 45668 10332
rect 45724 7474 45780 11900
rect 45836 11890 45892 11900
rect 45836 10836 45892 10846
rect 45836 10742 45892 10780
rect 45948 10500 46004 12014
rect 46284 12068 46340 12078
rect 46172 10836 46228 10846
rect 46284 10836 46340 12012
rect 46172 10834 46340 10836
rect 46172 10782 46174 10834
rect 46226 10782 46340 10834
rect 46172 10780 46340 10782
rect 46172 10770 46228 10780
rect 46508 10722 46564 12124
rect 46508 10670 46510 10722
rect 46562 10670 46564 10722
rect 46508 10658 46564 10670
rect 46844 12178 46900 12190
rect 46844 12126 46846 12178
rect 46898 12126 46900 12178
rect 46844 11508 46900 12126
rect 46844 10722 46900 11452
rect 47740 11508 47796 11518
rect 47740 11414 47796 11452
rect 48188 11170 48244 11182
rect 48188 11118 48190 11170
rect 48242 11118 48244 11170
rect 46844 10670 46846 10722
rect 46898 10670 46900 10722
rect 46844 10658 46900 10670
rect 47180 10722 47236 10734
rect 47180 10670 47182 10722
rect 47234 10670 47236 10722
rect 45948 10444 46228 10500
rect 46172 10276 46228 10444
rect 46172 10210 46228 10220
rect 47180 10276 47236 10670
rect 47180 10210 47236 10220
rect 47404 10610 47460 10622
rect 47404 10558 47406 10610
rect 47458 10558 47460 10610
rect 45948 10164 46004 10174
rect 45836 9044 45892 9054
rect 45836 8950 45892 8988
rect 45948 8258 46004 10108
rect 46844 10164 46900 10174
rect 45948 8206 45950 8258
rect 46002 8206 46004 8258
rect 45948 8194 46004 8206
rect 46620 8260 46676 8270
rect 45724 7422 45726 7474
rect 45778 7422 45780 7474
rect 45724 7410 45780 7422
rect 46396 7476 46452 7486
rect 46060 6692 46116 6702
rect 45612 6690 46116 6692
rect 45612 6638 46062 6690
rect 46114 6638 46116 6690
rect 45612 6636 46116 6638
rect 46060 6626 46116 6636
rect 45332 6524 45444 6580
rect 45276 6514 45332 6524
rect 45164 6188 45332 6244
rect 45052 5070 45054 5122
rect 45106 5070 45108 5122
rect 45052 5058 45108 5070
rect 45164 4452 45220 4462
rect 45164 4358 45220 4396
rect 45276 3556 45332 6188
rect 46396 5012 46452 7420
rect 46396 4946 46452 4956
rect 46508 5124 46564 5134
rect 45836 4900 45892 4910
rect 45836 4806 45892 4844
rect 45276 3490 45332 3500
rect 46508 3442 46564 5068
rect 46620 4564 46676 8204
rect 46732 5906 46788 5918
rect 46732 5854 46734 5906
rect 46786 5854 46788 5906
rect 46732 5796 46788 5854
rect 46732 5730 46788 5740
rect 46620 4498 46676 4508
rect 46844 4116 46900 10108
rect 46956 9604 47012 9614
rect 46956 6130 47012 9548
rect 47180 9604 47236 9614
rect 47180 9510 47236 9548
rect 46956 6078 46958 6130
rect 47010 6078 47012 6130
rect 46956 5012 47012 6078
rect 47068 8932 47124 8942
rect 47068 5794 47124 8876
rect 47404 8596 47460 10558
rect 47964 10498 48020 10510
rect 47964 10446 47966 10498
rect 48018 10446 48020 10498
rect 47852 10386 47908 10398
rect 47852 10334 47854 10386
rect 47906 10334 47908 10386
rect 47852 9826 47908 10334
rect 47852 9774 47854 9826
rect 47906 9774 47908 9826
rect 47852 9762 47908 9774
rect 47964 9044 48020 10446
rect 48188 10164 48244 11118
rect 48188 10098 48244 10108
rect 47964 8978 48020 8988
rect 47964 8820 48020 8830
rect 47964 8726 48020 8764
rect 47404 8530 47460 8540
rect 47964 8370 48020 8382
rect 47964 8318 47966 8370
rect 48018 8318 48020 8370
rect 47964 8148 48020 8318
rect 47964 8082 48020 8092
rect 48188 8036 48244 8046
rect 47964 7476 48020 7486
rect 47964 7362 48020 7420
rect 47964 7310 47966 7362
rect 48018 7310 48020 7362
rect 47964 7298 48020 7310
rect 48188 6802 48244 7980
rect 48188 6750 48190 6802
rect 48242 6750 48244 6802
rect 48188 6738 48244 6750
rect 47292 6020 47348 6030
rect 47292 5926 47348 5964
rect 48188 6018 48244 6030
rect 48188 5966 48190 6018
rect 48242 5966 48244 6018
rect 47068 5742 47070 5794
rect 47122 5742 47124 5794
rect 47068 5730 47124 5742
rect 47180 5906 47236 5918
rect 47180 5854 47182 5906
rect 47234 5854 47236 5906
rect 47068 5572 47124 5582
rect 47180 5572 47236 5854
rect 47124 5516 47236 5572
rect 47852 5906 47908 5918
rect 47852 5854 47854 5906
rect 47906 5854 47908 5906
rect 47068 5506 47124 5516
rect 47852 5460 47908 5854
rect 47852 5394 47908 5404
rect 47964 5348 48020 5358
rect 47740 5236 47796 5246
rect 47404 5012 47460 5022
rect 46956 4956 47348 5012
rect 47292 4226 47348 4956
rect 47292 4174 47294 4226
rect 47346 4174 47348 4226
rect 47292 4162 47348 4174
rect 46956 4116 47012 4126
rect 46844 4060 46956 4116
rect 46956 4050 47012 4060
rect 46732 3668 46788 3678
rect 46732 3554 46788 3612
rect 46732 3502 46734 3554
rect 46786 3502 46788 3554
rect 46732 3490 46788 3502
rect 46508 3390 46510 3442
rect 46562 3390 46564 3442
rect 44828 3332 45108 3388
rect 46508 3378 46564 3390
rect 47404 3442 47460 4956
rect 47740 5010 47796 5180
rect 47964 5122 48020 5292
rect 47964 5070 47966 5122
rect 48018 5070 48020 5122
rect 47964 5058 48020 5070
rect 47740 4958 47742 5010
rect 47794 4958 47796 5010
rect 47740 4946 47796 4958
rect 47628 4564 47684 4574
rect 47628 4470 47684 4508
rect 47852 4340 47908 4350
rect 47852 4246 47908 4284
rect 47628 3780 47684 3790
rect 47628 3554 47684 3724
rect 48188 3666 48244 5966
rect 48188 3614 48190 3666
rect 48242 3614 48244 3666
rect 48188 3602 48244 3614
rect 47628 3502 47630 3554
rect 47682 3502 47684 3554
rect 47628 3490 47684 3502
rect 47404 3390 47406 3442
rect 47458 3390 47460 3442
rect 47404 3378 47460 3390
rect 48076 3444 48132 3482
rect 48076 3378 48132 3388
rect 45052 800 45108 3332
rect 35980 700 36484 756
rect 36960 0 37072 800
rect 37632 0 37744 800
rect 38304 0 38416 800
rect 38976 0 39088 800
rect 39648 0 39760 800
rect 40320 0 40432 800
rect 40992 0 41104 800
rect 41664 0 41776 800
rect 42336 0 42448 800
rect 43008 0 43120 800
rect 43680 0 43792 800
rect 44352 0 44464 800
rect 45024 0 45136 800
<< via2 >>
rect 4476 46282 4532 46284
rect 4476 46230 4478 46282
rect 4478 46230 4530 46282
rect 4530 46230 4532 46282
rect 4476 46228 4532 46230
rect 4580 46282 4636 46284
rect 4580 46230 4582 46282
rect 4582 46230 4634 46282
rect 4634 46230 4636 46282
rect 4580 46228 4636 46230
rect 4684 46282 4740 46284
rect 4684 46230 4686 46282
rect 4686 46230 4738 46282
rect 4738 46230 4740 46282
rect 4684 46228 4740 46230
rect 10668 46002 10724 46004
rect 10668 45950 10670 46002
rect 10670 45950 10722 46002
rect 10722 45950 10724 46002
rect 10668 45948 10724 45950
rect 13916 45948 13972 46004
rect 15260 45890 15316 45892
rect 15260 45838 15262 45890
rect 15262 45838 15314 45890
rect 15314 45838 15316 45890
rect 15260 45836 15316 45838
rect 16268 45890 16324 45892
rect 16268 45838 16270 45890
rect 16270 45838 16322 45890
rect 16322 45838 16324 45890
rect 16268 45836 16324 45838
rect 1708 45388 1764 45444
rect 7420 45612 7476 45668
rect 6188 44940 6244 44996
rect 4476 44714 4532 44716
rect 4476 44662 4478 44714
rect 4478 44662 4530 44714
rect 4530 44662 4532 44714
rect 4476 44660 4532 44662
rect 4580 44714 4636 44716
rect 4580 44662 4582 44714
rect 4582 44662 4634 44714
rect 4634 44662 4636 44714
rect 4580 44660 4636 44662
rect 4684 44714 4740 44716
rect 4684 44662 4686 44714
rect 4686 44662 4738 44714
rect 4738 44662 4740 44714
rect 4684 44660 4740 44662
rect 1484 44044 1540 44100
rect 1372 39116 1428 39172
rect 3948 43596 4004 43652
rect 1708 41970 1764 41972
rect 1708 41918 1710 41970
rect 1710 41918 1762 41970
rect 1762 41918 1764 41970
rect 1708 41916 1764 41918
rect 1596 40348 1652 40404
rect 1708 38332 1764 38388
rect 1820 40962 1876 40964
rect 1820 40910 1822 40962
rect 1822 40910 1874 40962
rect 1874 40910 1876 40962
rect 1820 40908 1876 40910
rect 1708 38050 1764 38052
rect 1708 37998 1710 38050
rect 1710 37998 1762 38050
rect 1762 37998 1764 38050
rect 1708 37996 1764 37998
rect 1708 36876 1764 36932
rect 2156 42476 2212 42532
rect 4844 43596 4900 43652
rect 5628 43596 5684 43652
rect 2268 42028 2324 42084
rect 2268 41356 2324 41412
rect 2156 40908 2212 40964
rect 2268 39788 2324 39844
rect 2492 40290 2548 40292
rect 2492 40238 2494 40290
rect 2494 40238 2546 40290
rect 2546 40238 2548 40290
rect 2492 40236 2548 40238
rect 2604 39676 2660 39732
rect 2940 40124 2996 40180
rect 2940 39506 2996 39508
rect 2940 39454 2942 39506
rect 2942 39454 2994 39506
rect 2994 39454 2996 39506
rect 2940 39452 2996 39454
rect 2044 36988 2100 37044
rect 1708 35644 1764 35700
rect 1820 35196 1876 35252
rect 1708 34860 1764 34916
rect 1820 34524 1876 34580
rect 1372 33180 1428 33236
rect 1708 33852 1764 33908
rect 1484 32284 1540 32340
rect 2268 38162 2324 38164
rect 2268 38110 2270 38162
rect 2270 38110 2322 38162
rect 2322 38110 2324 38162
rect 2268 38108 2324 38110
rect 2828 37884 2884 37940
rect 2828 37436 2884 37492
rect 2268 36204 2324 36260
rect 2156 35196 2212 35252
rect 2268 35084 2324 35140
rect 2604 34524 2660 34580
rect 2716 35196 2772 35252
rect 2604 34354 2660 34356
rect 2604 34302 2606 34354
rect 2606 34302 2658 34354
rect 2658 34302 2660 34354
rect 2604 34300 2660 34302
rect 2044 33852 2100 33908
rect 2156 33292 2212 33348
rect 1820 31612 1876 31668
rect 1708 30940 1764 30996
rect 3388 40124 3444 40180
rect 3164 39788 3220 39844
rect 3164 38892 3220 38948
rect 3276 39676 3332 39732
rect 3500 40012 3556 40068
rect 3500 39564 3556 39620
rect 3500 39394 3556 39396
rect 3500 39342 3502 39394
rect 3502 39342 3554 39394
rect 3554 39342 3556 39394
rect 3500 39340 3556 39342
rect 3948 42530 4004 42532
rect 3948 42478 3950 42530
rect 3950 42478 4002 42530
rect 4002 42478 4004 42530
rect 3948 42476 4004 42478
rect 3836 41970 3892 41972
rect 3836 41918 3838 41970
rect 3838 41918 3890 41970
rect 3890 41918 3892 41970
rect 3836 41916 3892 41918
rect 3052 37548 3108 37604
rect 3724 40236 3780 40292
rect 3052 37378 3108 37380
rect 3052 37326 3054 37378
rect 3054 37326 3106 37378
rect 3106 37326 3108 37378
rect 3052 37324 3108 37326
rect 2940 36876 2996 36932
rect 3164 36204 3220 36260
rect 4844 43426 4900 43428
rect 4844 43374 4846 43426
rect 4846 43374 4898 43426
rect 4898 43374 4900 43426
rect 4844 43372 4900 43374
rect 4476 43146 4532 43148
rect 4476 43094 4478 43146
rect 4478 43094 4530 43146
rect 4530 43094 4532 43146
rect 4476 43092 4532 43094
rect 4580 43146 4636 43148
rect 4580 43094 4582 43146
rect 4582 43094 4634 43146
rect 4634 43094 4636 43146
rect 4580 43092 4636 43094
rect 4684 43146 4740 43148
rect 4684 43094 4686 43146
rect 4686 43094 4738 43146
rect 4738 43094 4740 43146
rect 4684 43092 4740 43094
rect 4060 40012 4116 40068
rect 3948 39788 4004 39844
rect 3388 37996 3444 38052
rect 3500 38108 3556 38164
rect 4284 42028 4340 42084
rect 8092 45666 8148 45668
rect 8092 45614 8094 45666
rect 8094 45614 8146 45666
rect 8146 45614 8148 45666
rect 8092 45612 8148 45614
rect 7980 44994 8036 44996
rect 7980 44942 7982 44994
rect 7982 44942 8034 44994
rect 8034 44942 8036 44994
rect 7980 44940 8036 44942
rect 8428 44994 8484 44996
rect 8428 44942 8430 44994
rect 8430 44942 8482 44994
rect 8482 44942 8484 44994
rect 8428 44940 8484 44942
rect 6076 43596 6132 43652
rect 5740 43372 5796 43428
rect 6636 42924 6692 42980
rect 6412 42642 6468 42644
rect 6412 42590 6414 42642
rect 6414 42590 6466 42642
rect 6466 42590 6468 42642
rect 6412 42588 6468 42590
rect 6300 42252 6356 42308
rect 5404 41916 5460 41972
rect 4956 41804 5012 41860
rect 4476 41578 4532 41580
rect 4476 41526 4478 41578
rect 4478 41526 4530 41578
rect 4530 41526 4532 41578
rect 4476 41524 4532 41526
rect 4580 41578 4636 41580
rect 4580 41526 4582 41578
rect 4582 41526 4634 41578
rect 4634 41526 4636 41578
rect 4580 41524 4636 41526
rect 4684 41578 4740 41580
rect 4684 41526 4686 41578
rect 4686 41526 4738 41578
rect 4738 41526 4740 41578
rect 4684 41524 4740 41526
rect 5852 41298 5908 41300
rect 5852 41246 5854 41298
rect 5854 41246 5906 41298
rect 5906 41246 5908 41298
rect 5852 41244 5908 41246
rect 5068 41020 5124 41076
rect 5740 41132 5796 41188
rect 4476 40010 4532 40012
rect 4476 39958 4478 40010
rect 4478 39958 4530 40010
rect 4530 39958 4532 40010
rect 4476 39956 4532 39958
rect 4580 40010 4636 40012
rect 4580 39958 4582 40010
rect 4582 39958 4634 40010
rect 4634 39958 4636 40010
rect 4580 39956 4636 39958
rect 4684 40010 4740 40012
rect 4684 39958 4686 40010
rect 4686 39958 4738 40010
rect 4738 39958 4740 40010
rect 4684 39956 4740 39958
rect 4396 39116 4452 39172
rect 4284 39004 4340 39060
rect 3612 37826 3668 37828
rect 3612 37774 3614 37826
rect 3614 37774 3666 37826
rect 3666 37774 3668 37826
rect 3612 37772 3668 37774
rect 3836 37660 3892 37716
rect 3612 37490 3668 37492
rect 3612 37438 3614 37490
rect 3614 37438 3666 37490
rect 3666 37438 3668 37490
rect 3612 37436 3668 37438
rect 3948 37436 4004 37492
rect 3500 37154 3556 37156
rect 3500 37102 3502 37154
rect 3502 37102 3554 37154
rect 3554 37102 3556 37154
rect 3500 37100 3556 37102
rect 3724 36988 3780 37044
rect 3276 35644 3332 35700
rect 2940 34860 2996 34916
rect 2940 34690 2996 34692
rect 2940 34638 2942 34690
rect 2942 34638 2994 34690
rect 2994 34638 2996 34690
rect 2940 34636 2996 34638
rect 2940 34354 2996 34356
rect 2940 34302 2942 34354
rect 2942 34302 2994 34354
rect 2994 34302 2996 34354
rect 2940 34300 2996 34302
rect 2828 34188 2884 34244
rect 2604 33628 2660 33684
rect 2268 32844 2324 32900
rect 2828 33516 2884 33572
rect 3612 34972 3668 35028
rect 3948 37100 4004 37156
rect 5292 39004 5348 39060
rect 5404 39452 5460 39508
rect 4732 38780 4788 38836
rect 4620 38556 4676 38612
rect 4476 38442 4532 38444
rect 4476 38390 4478 38442
rect 4478 38390 4530 38442
rect 4530 38390 4532 38442
rect 4476 38388 4532 38390
rect 4580 38442 4636 38444
rect 4580 38390 4582 38442
rect 4582 38390 4634 38442
rect 4634 38390 4636 38442
rect 4580 38388 4636 38390
rect 4684 38442 4740 38444
rect 4684 38390 4686 38442
rect 4686 38390 4738 38442
rect 4738 38390 4740 38442
rect 4684 38388 4740 38390
rect 4172 38108 4228 38164
rect 4396 37996 4452 38052
rect 4956 37996 5012 38052
rect 4508 37938 4564 37940
rect 4508 37886 4510 37938
rect 4510 37886 4562 37938
rect 4562 37886 4564 37938
rect 4508 37884 4564 37886
rect 4172 37660 4228 37716
rect 4172 37212 4228 37268
rect 5180 37884 5236 37940
rect 4732 37212 4788 37268
rect 4732 36988 4788 37044
rect 4060 35196 4116 35252
rect 4172 36540 4228 36596
rect 3836 34972 3892 35028
rect 5068 37548 5124 37604
rect 4476 36874 4532 36876
rect 4476 36822 4478 36874
rect 4478 36822 4530 36874
rect 4530 36822 4532 36874
rect 4476 36820 4532 36822
rect 4580 36874 4636 36876
rect 4580 36822 4582 36874
rect 4582 36822 4634 36874
rect 4634 36822 4636 36874
rect 4580 36820 4636 36822
rect 4684 36874 4740 36876
rect 4684 36822 4686 36874
rect 4686 36822 4738 36874
rect 4738 36822 4740 36874
rect 4684 36820 4740 36822
rect 4732 36540 4788 36596
rect 4956 37436 5012 37492
rect 3388 34802 3444 34804
rect 3388 34750 3390 34802
rect 3390 34750 3442 34802
rect 3442 34750 3444 34802
rect 3388 34748 3444 34750
rect 3500 34860 3556 34916
rect 4476 35306 4532 35308
rect 4476 35254 4478 35306
rect 4478 35254 4530 35306
rect 4530 35254 4532 35306
rect 4476 35252 4532 35254
rect 4580 35306 4636 35308
rect 4580 35254 4582 35306
rect 4582 35254 4634 35306
rect 4634 35254 4636 35306
rect 4580 35252 4636 35254
rect 4684 35306 4740 35308
rect 4684 35254 4686 35306
rect 4686 35254 4738 35306
rect 4738 35254 4740 35306
rect 4684 35252 4740 35254
rect 3724 34860 3780 34916
rect 3612 34690 3668 34692
rect 3612 34638 3614 34690
rect 3614 34638 3666 34690
rect 3666 34638 3668 34690
rect 3612 34636 3668 34638
rect 3612 34412 3668 34468
rect 3836 34300 3892 34356
rect 3276 33516 3332 33572
rect 3388 33852 3444 33908
rect 3836 33570 3892 33572
rect 3836 33518 3838 33570
rect 3838 33518 3890 33570
rect 3890 33518 3892 33570
rect 3836 33516 3892 33518
rect 3612 33458 3668 33460
rect 3612 33406 3614 33458
rect 3614 33406 3666 33458
rect 3666 33406 3668 33458
rect 3612 33404 3668 33406
rect 3052 32732 3108 32788
rect 2940 32674 2996 32676
rect 2940 32622 2942 32674
rect 2942 32622 2994 32674
rect 2994 32622 2996 32674
rect 2940 32620 2996 32622
rect 2268 32450 2324 32452
rect 2268 32398 2270 32450
rect 2270 32398 2322 32450
rect 2322 32398 2324 32450
rect 2268 32396 2324 32398
rect 3836 33068 3892 33124
rect 3612 32732 3668 32788
rect 3948 32674 4004 32676
rect 3948 32622 3950 32674
rect 3950 32622 4002 32674
rect 4002 32622 4004 32674
rect 3948 32620 4004 32622
rect 3164 31724 3220 31780
rect 3276 31666 3332 31668
rect 3276 31614 3278 31666
rect 3278 31614 3330 31666
rect 3330 31614 3332 31666
rect 3276 31612 3332 31614
rect 2380 30940 2436 30996
rect 1820 30268 1876 30324
rect 1708 30156 1764 30212
rect 1820 29148 1876 29204
rect 2492 29596 2548 29652
rect 1708 28252 1764 28308
rect 2716 29538 2772 29540
rect 2716 29486 2718 29538
rect 2718 29486 2770 29538
rect 2770 29486 2772 29538
rect 2716 29484 2772 29486
rect 2492 29426 2548 29428
rect 2492 29374 2494 29426
rect 2494 29374 2546 29426
rect 2546 29374 2548 29426
rect 2492 29372 2548 29374
rect 2828 29372 2884 29428
rect 3164 29426 3220 29428
rect 3164 29374 3166 29426
rect 3166 29374 3218 29426
rect 3218 29374 3220 29426
rect 3164 29372 3220 29374
rect 4396 34748 4452 34804
rect 4732 34354 4788 34356
rect 4732 34302 4734 34354
rect 4734 34302 4786 34354
rect 4786 34302 4788 34354
rect 4732 34300 4788 34302
rect 4172 33458 4228 33460
rect 4172 33406 4174 33458
rect 4174 33406 4226 33458
rect 4226 33406 4228 33458
rect 4172 33404 4228 33406
rect 4396 34076 4452 34132
rect 4476 33738 4532 33740
rect 4476 33686 4478 33738
rect 4478 33686 4530 33738
rect 4530 33686 4532 33738
rect 4476 33684 4532 33686
rect 4580 33738 4636 33740
rect 4580 33686 4582 33738
rect 4582 33686 4634 33738
rect 4634 33686 4636 33738
rect 4580 33684 4636 33686
rect 4684 33738 4740 33740
rect 4684 33686 4686 33738
rect 4686 33686 4738 33738
rect 4738 33686 4740 33738
rect 4684 33684 4740 33686
rect 4844 33516 4900 33572
rect 5068 35756 5124 35812
rect 5068 35026 5124 35028
rect 5068 34974 5070 35026
rect 5070 34974 5122 35026
rect 5122 34974 5124 35026
rect 5068 34972 5124 34974
rect 5180 34300 5236 34356
rect 6300 40460 6356 40516
rect 6188 40348 6244 40404
rect 5964 39676 6020 39732
rect 5852 39564 5908 39620
rect 6188 39506 6244 39508
rect 6188 39454 6190 39506
rect 6190 39454 6242 39506
rect 6242 39454 6244 39506
rect 6188 39452 6244 39454
rect 6636 42252 6692 42308
rect 7196 44098 7252 44100
rect 7196 44046 7198 44098
rect 7198 44046 7250 44098
rect 7250 44046 7252 44098
rect 7196 44044 7252 44046
rect 8764 44828 8820 44884
rect 8428 44210 8484 44212
rect 8428 44158 8430 44210
rect 8430 44158 8482 44210
rect 8482 44158 8484 44210
rect 8428 44156 8484 44158
rect 8316 44098 8372 44100
rect 8316 44046 8318 44098
rect 8318 44046 8370 44098
rect 8370 44046 8372 44098
rect 8316 44044 8372 44046
rect 8988 44044 9044 44100
rect 8652 42530 8708 42532
rect 8652 42478 8654 42530
rect 8654 42478 8706 42530
rect 8706 42478 8708 42530
rect 8652 42476 8708 42478
rect 7980 42194 8036 42196
rect 7980 42142 7982 42194
rect 7982 42142 8034 42194
rect 8034 42142 8036 42194
rect 7980 42140 8036 42142
rect 7420 41970 7476 41972
rect 7420 41918 7422 41970
rect 7422 41918 7474 41970
rect 7474 41918 7476 41970
rect 7420 41916 7476 41918
rect 6748 41804 6804 41860
rect 6636 40124 6692 40180
rect 6748 39564 6804 39620
rect 6972 41244 7028 41300
rect 7084 41074 7140 41076
rect 7084 41022 7086 41074
rect 7086 41022 7138 41074
rect 7138 41022 7140 41074
rect 7084 41020 7140 41022
rect 7420 41020 7476 41076
rect 7980 40572 8036 40628
rect 8092 40684 8148 40740
rect 7532 40236 7588 40292
rect 6524 39228 6580 39284
rect 5740 38834 5796 38836
rect 5740 38782 5742 38834
rect 5742 38782 5794 38834
rect 5794 38782 5796 38834
rect 5740 38780 5796 38782
rect 5852 39004 5908 39060
rect 6636 39340 6692 39396
rect 6300 38892 6356 38948
rect 6860 39228 6916 39284
rect 6748 39058 6804 39060
rect 6748 39006 6750 39058
rect 6750 39006 6802 39058
rect 6802 39006 6804 39058
rect 6748 39004 6804 39006
rect 5964 38556 6020 38612
rect 6188 37884 6244 37940
rect 6076 37772 6132 37828
rect 5964 36988 6020 37044
rect 5852 35980 5908 36036
rect 5628 35922 5684 35924
rect 5628 35870 5630 35922
rect 5630 35870 5682 35922
rect 5682 35870 5684 35922
rect 5628 35868 5684 35870
rect 7084 38892 7140 38948
rect 8316 39788 8372 39844
rect 6188 36370 6244 36372
rect 6188 36318 6190 36370
rect 6190 36318 6242 36370
rect 6242 36318 6244 36370
rect 6188 36316 6244 36318
rect 6860 38108 6916 38164
rect 6860 37660 6916 37716
rect 6636 35868 6692 35924
rect 5740 35698 5796 35700
rect 5740 35646 5742 35698
rect 5742 35646 5794 35698
rect 5794 35646 5796 35698
rect 5740 35644 5796 35646
rect 4508 33122 4564 33124
rect 4508 33070 4510 33122
rect 4510 33070 4562 33122
rect 4562 33070 4564 33122
rect 4508 33068 4564 33070
rect 4508 32786 4564 32788
rect 4508 32734 4510 32786
rect 4510 32734 4562 32786
rect 4562 32734 4564 32786
rect 4508 32732 4564 32734
rect 5180 33516 5236 33572
rect 4844 32956 4900 33012
rect 4844 32732 4900 32788
rect 4284 32284 4340 32340
rect 4172 31836 4228 31892
rect 4060 31778 4116 31780
rect 4060 31726 4062 31778
rect 4062 31726 4114 31778
rect 4114 31726 4116 31778
rect 4060 31724 4116 31726
rect 4060 31500 4116 31556
rect 3724 30940 3780 30996
rect 3948 30882 4004 30884
rect 3948 30830 3950 30882
rect 3950 30830 4002 30882
rect 4002 30830 4004 30882
rect 3948 30828 4004 30830
rect 4476 32170 4532 32172
rect 4476 32118 4478 32170
rect 4478 32118 4530 32170
rect 4530 32118 4532 32170
rect 4476 32116 4532 32118
rect 4580 32170 4636 32172
rect 4580 32118 4582 32170
rect 4582 32118 4634 32170
rect 4634 32118 4636 32170
rect 4580 32116 4636 32118
rect 4684 32170 4740 32172
rect 4684 32118 4686 32170
rect 4686 32118 4738 32170
rect 4738 32118 4740 32170
rect 4684 32116 4740 32118
rect 4508 31948 4564 32004
rect 5404 32508 5460 32564
rect 5964 35196 6020 35252
rect 5964 34972 6020 35028
rect 7756 38332 7812 38388
rect 7644 38162 7700 38164
rect 7644 38110 7646 38162
rect 7646 38110 7698 38162
rect 7698 38110 7700 38162
rect 7644 38108 7700 38110
rect 8316 38556 8372 38612
rect 8316 38162 8372 38164
rect 8316 38110 8318 38162
rect 8318 38110 8370 38162
rect 8370 38110 8372 38162
rect 8316 38108 8372 38110
rect 8204 37378 8260 37380
rect 8204 37326 8206 37378
rect 8206 37326 8258 37378
rect 8258 37326 8260 37378
rect 8204 37324 8260 37326
rect 8092 37266 8148 37268
rect 8092 37214 8094 37266
rect 8094 37214 8146 37266
rect 8146 37214 8148 37266
rect 8092 37212 8148 37214
rect 6860 35756 6916 35812
rect 7084 36092 7140 36148
rect 6300 34972 6356 35028
rect 6636 34972 6692 35028
rect 5180 32284 5236 32340
rect 5068 31836 5124 31892
rect 4844 31052 4900 31108
rect 4956 30940 5012 30996
rect 4476 30602 4532 30604
rect 4476 30550 4478 30602
rect 4478 30550 4530 30602
rect 4530 30550 4532 30602
rect 4476 30548 4532 30550
rect 4580 30602 4636 30604
rect 4580 30550 4582 30602
rect 4582 30550 4634 30602
rect 4634 30550 4636 30602
rect 4580 30548 4636 30550
rect 4684 30602 4740 30604
rect 4684 30550 4686 30602
rect 4686 30550 4738 30602
rect 4738 30550 4740 30602
rect 4684 30548 4740 30550
rect 4172 30156 4228 30212
rect 4284 30044 4340 30100
rect 4284 29596 4340 29652
rect 2604 28700 2660 28756
rect 2716 29260 2772 29316
rect 3500 29148 3556 29204
rect 3052 28924 3108 28980
rect 2268 28252 2324 28308
rect 2268 28028 2324 28084
rect 1372 27916 1428 27972
rect 1708 26236 1764 26292
rect 1708 25788 1764 25844
rect 1708 25564 1764 25620
rect 2492 27746 2548 27748
rect 2492 27694 2494 27746
rect 2494 27694 2546 27746
rect 2546 27694 2548 27746
rect 2492 27692 2548 27694
rect 2380 26796 2436 26852
rect 2156 26572 2212 26628
rect 2716 26796 2772 26852
rect 2492 26684 2548 26740
rect 2492 25228 2548 25284
rect 2380 24722 2436 24724
rect 2380 24670 2382 24722
rect 2382 24670 2434 24722
rect 2434 24670 2436 24722
rect 2380 24668 2436 24670
rect 2044 24108 2100 24164
rect 2156 24556 2212 24612
rect 1708 23548 1764 23604
rect 1820 22988 1876 23044
rect 2044 22876 2100 22932
rect 1708 20076 1764 20132
rect 2156 19346 2212 19348
rect 2156 19294 2158 19346
rect 2158 19294 2210 19346
rect 2210 19294 2212 19346
rect 2156 19292 2212 19294
rect 3164 28588 3220 28644
rect 5404 30828 5460 30884
rect 4956 30268 5012 30324
rect 5068 30380 5124 30436
rect 4396 29260 4452 29316
rect 4956 29260 5012 29316
rect 4476 29034 4532 29036
rect 4476 28982 4478 29034
rect 4478 28982 4530 29034
rect 4530 28982 4532 29034
rect 4476 28980 4532 28982
rect 4580 29034 4636 29036
rect 4580 28982 4582 29034
rect 4582 28982 4634 29034
rect 4634 28982 4636 29034
rect 4580 28980 4636 28982
rect 4684 29034 4740 29036
rect 4684 28982 4686 29034
rect 4686 28982 4738 29034
rect 4738 28982 4740 29034
rect 4684 28980 4740 28982
rect 4844 28924 4900 28980
rect 4396 28700 4452 28756
rect 4620 28588 4676 28644
rect 5180 28812 5236 28868
rect 3164 27132 3220 27188
rect 3388 27580 3444 27636
rect 2940 26460 2996 26516
rect 2940 26178 2996 26180
rect 2940 26126 2942 26178
rect 2942 26126 2994 26178
rect 2994 26126 2996 26178
rect 2940 26124 2996 26126
rect 3052 25788 3108 25844
rect 2716 25564 2772 25620
rect 2940 25116 2996 25172
rect 2492 22540 2548 22596
rect 3724 27580 3780 27636
rect 4476 27466 4532 27468
rect 4476 27414 4478 27466
rect 4478 27414 4530 27466
rect 4530 27414 4532 27466
rect 4476 27412 4532 27414
rect 4580 27466 4636 27468
rect 4580 27414 4582 27466
rect 4582 27414 4634 27466
rect 4634 27414 4636 27466
rect 4580 27412 4636 27414
rect 4684 27466 4740 27468
rect 4684 27414 4686 27466
rect 4686 27414 4738 27466
rect 4738 27414 4740 27466
rect 4684 27412 4740 27414
rect 3612 26850 3668 26852
rect 3612 26798 3614 26850
rect 3614 26798 3666 26850
rect 3666 26798 3668 26850
rect 3612 26796 3668 26798
rect 3500 26572 3556 26628
rect 3276 25228 3332 25284
rect 4060 27244 4116 27300
rect 5068 27746 5124 27748
rect 5068 27694 5070 27746
rect 5070 27694 5122 27746
rect 5122 27694 5124 27746
rect 5068 27692 5124 27694
rect 5964 33068 6020 33124
rect 6188 34300 6244 34356
rect 6412 34354 6468 34356
rect 6412 34302 6414 34354
rect 6414 34302 6466 34354
rect 6466 34302 6468 34354
rect 6412 34300 6468 34302
rect 6412 33628 6468 33684
rect 6300 33180 6356 33236
rect 6748 34354 6804 34356
rect 6748 34302 6750 34354
rect 6750 34302 6802 34354
rect 6802 34302 6804 34354
rect 6748 34300 6804 34302
rect 6860 34242 6916 34244
rect 6860 34190 6862 34242
rect 6862 34190 6914 34242
rect 6914 34190 6916 34242
rect 6860 34188 6916 34190
rect 6636 33964 6692 34020
rect 6972 33628 7028 33684
rect 6636 33346 6692 33348
rect 6636 33294 6638 33346
rect 6638 33294 6690 33346
rect 6690 33294 6692 33346
rect 6636 33292 6692 33294
rect 5628 32450 5684 32452
rect 5628 32398 5630 32450
rect 5630 32398 5682 32450
rect 5682 32398 5684 32450
rect 5628 32396 5684 32398
rect 5740 31948 5796 32004
rect 6300 32508 6356 32564
rect 5852 31778 5908 31780
rect 5852 31726 5854 31778
rect 5854 31726 5906 31778
rect 5906 31726 5908 31778
rect 5852 31724 5908 31726
rect 6636 32396 6692 32452
rect 6748 32060 6804 32116
rect 6636 31890 6692 31892
rect 6636 31838 6638 31890
rect 6638 31838 6690 31890
rect 6690 31838 6692 31890
rect 6636 31836 6692 31838
rect 6412 31500 6468 31556
rect 6636 31276 6692 31332
rect 5740 28866 5796 28868
rect 5740 28814 5742 28866
rect 5742 28814 5794 28866
rect 5794 28814 5796 28866
rect 5740 28812 5796 28814
rect 6188 30828 6244 30884
rect 5628 28642 5684 28644
rect 5628 28590 5630 28642
rect 5630 28590 5682 28642
rect 5682 28590 5684 28642
rect 5628 28588 5684 28590
rect 5852 28364 5908 28420
rect 5740 28028 5796 28084
rect 4732 26962 4788 26964
rect 4732 26910 4734 26962
rect 4734 26910 4786 26962
rect 4786 26910 4788 26962
rect 4732 26908 4788 26910
rect 4396 26460 4452 26516
rect 4620 26684 4676 26740
rect 4844 26572 4900 26628
rect 3836 25788 3892 25844
rect 3388 24556 3444 24612
rect 4476 25898 4532 25900
rect 4476 25846 4478 25898
rect 4478 25846 4530 25898
rect 4530 25846 4532 25898
rect 4476 25844 4532 25846
rect 4580 25898 4636 25900
rect 4580 25846 4582 25898
rect 4582 25846 4634 25898
rect 4634 25846 4636 25898
rect 4580 25844 4636 25846
rect 4684 25898 4740 25900
rect 4684 25846 4686 25898
rect 4686 25846 4738 25898
rect 4738 25846 4740 25898
rect 4684 25844 4740 25846
rect 4620 25618 4676 25620
rect 4620 25566 4622 25618
rect 4622 25566 4674 25618
rect 4674 25566 4676 25618
rect 4620 25564 4676 25566
rect 4956 27132 5012 27188
rect 5628 26850 5684 26852
rect 5628 26798 5630 26850
rect 5630 26798 5682 26850
rect 5682 26798 5684 26850
rect 5628 26796 5684 26798
rect 5068 26572 5124 26628
rect 5180 26684 5236 26740
rect 5068 26402 5124 26404
rect 5068 26350 5070 26402
rect 5070 26350 5122 26402
rect 5122 26350 5124 26402
rect 5068 26348 5124 26350
rect 5516 26514 5572 26516
rect 5516 26462 5518 26514
rect 5518 26462 5570 26514
rect 5570 26462 5572 26514
rect 5516 26460 5572 26462
rect 5964 27244 6020 27300
rect 5740 26684 5796 26740
rect 5964 26684 6020 26740
rect 5404 26124 5460 26180
rect 5180 25116 5236 25172
rect 4476 24330 4532 24332
rect 4476 24278 4478 24330
rect 4478 24278 4530 24330
rect 4530 24278 4532 24330
rect 4476 24276 4532 24278
rect 4580 24330 4636 24332
rect 4580 24278 4582 24330
rect 4582 24278 4634 24330
rect 4634 24278 4636 24330
rect 4580 24276 4636 24278
rect 4684 24330 4740 24332
rect 4684 24278 4686 24330
rect 4686 24278 4738 24330
rect 4738 24278 4740 24330
rect 4684 24276 4740 24278
rect 4620 24050 4676 24052
rect 4620 23998 4622 24050
rect 4622 23998 4674 24050
rect 4674 23998 4676 24050
rect 4620 23996 4676 23998
rect 3948 23042 4004 23044
rect 3948 22990 3950 23042
rect 3950 22990 4002 23042
rect 4002 22990 4004 23042
rect 3948 22988 4004 22990
rect 5068 24332 5124 24388
rect 4844 22988 4900 23044
rect 4476 22762 4532 22764
rect 4476 22710 4478 22762
rect 4478 22710 4530 22762
rect 4530 22710 4532 22762
rect 4476 22708 4532 22710
rect 4580 22762 4636 22764
rect 4580 22710 4582 22762
rect 4582 22710 4634 22762
rect 4634 22710 4636 22762
rect 4580 22708 4636 22710
rect 4684 22762 4740 22764
rect 4684 22710 4686 22762
rect 4686 22710 4738 22762
rect 4738 22710 4740 22762
rect 4684 22708 4740 22710
rect 4620 22482 4676 22484
rect 4620 22430 4622 22482
rect 4622 22430 4674 22482
rect 4674 22430 4676 22482
rect 4620 22428 4676 22430
rect 6524 30940 6580 30996
rect 6412 30716 6468 30772
rect 6300 30380 6356 30436
rect 6412 29708 6468 29764
rect 8204 37100 8260 37156
rect 7420 37042 7476 37044
rect 7420 36990 7422 37042
rect 7422 36990 7474 37042
rect 7474 36990 7476 37042
rect 7420 36988 7476 36990
rect 7420 36594 7476 36596
rect 7420 36542 7422 36594
rect 7422 36542 7474 36594
rect 7474 36542 7476 36594
rect 7420 36540 7476 36542
rect 7308 36428 7364 36484
rect 7532 36482 7588 36484
rect 7532 36430 7534 36482
rect 7534 36430 7586 36482
rect 7586 36430 7588 36482
rect 7532 36428 7588 36430
rect 7756 36428 7812 36484
rect 7644 36092 7700 36148
rect 7196 34972 7252 35028
rect 7420 35196 7476 35252
rect 8876 42082 8932 42084
rect 8876 42030 8878 42082
rect 8878 42030 8930 42082
rect 8930 42030 8932 42082
rect 8876 42028 8932 42030
rect 8764 41356 8820 41412
rect 8764 41186 8820 41188
rect 8764 41134 8766 41186
rect 8766 41134 8818 41186
rect 8818 41134 8820 41186
rect 8764 41132 8820 41134
rect 8540 40178 8596 40180
rect 8540 40126 8542 40178
rect 8542 40126 8594 40178
rect 8594 40126 8596 40178
rect 8540 40124 8596 40126
rect 8540 39340 8596 39396
rect 8652 39116 8708 39172
rect 8540 39058 8596 39060
rect 8540 39006 8542 39058
rect 8542 39006 8594 39058
rect 8594 39006 8596 39058
rect 8540 39004 8596 39006
rect 8540 38444 8596 38500
rect 11116 45388 11172 45444
rect 11564 45612 11620 45668
rect 10108 45052 10164 45108
rect 9660 44994 9716 44996
rect 9660 44942 9662 44994
rect 9662 44942 9714 44994
rect 9714 44942 9716 44994
rect 9660 44940 9716 44942
rect 9548 44828 9604 44884
rect 10108 44828 10164 44884
rect 9548 43596 9604 43652
rect 9212 42642 9268 42644
rect 9212 42590 9214 42642
rect 9214 42590 9266 42642
rect 9266 42590 9268 42642
rect 9212 42588 9268 42590
rect 9100 41804 9156 41860
rect 9996 42140 10052 42196
rect 10108 42866 10164 42868
rect 10108 42814 10110 42866
rect 10110 42814 10162 42866
rect 10162 42814 10164 42866
rect 10108 42812 10164 42814
rect 10220 42476 10276 42532
rect 11004 43708 11060 43764
rect 10892 42812 10948 42868
rect 10556 42700 10612 42756
rect 11452 43650 11508 43652
rect 11452 43598 11454 43650
rect 11454 43598 11506 43650
rect 11506 43598 11508 43650
rect 11452 43596 11508 43598
rect 11788 44940 11844 44996
rect 12236 45388 12292 45444
rect 11676 43708 11732 43764
rect 11900 43708 11956 43764
rect 11564 43538 11620 43540
rect 11564 43486 11566 43538
rect 11566 43486 11618 43538
rect 11618 43486 11620 43538
rect 11564 43484 11620 43486
rect 11676 43036 11732 43092
rect 11340 42754 11396 42756
rect 11340 42702 11342 42754
rect 11342 42702 11394 42754
rect 11394 42702 11396 42754
rect 11340 42700 11396 42702
rect 11452 42642 11508 42644
rect 11452 42590 11454 42642
rect 11454 42590 11506 42642
rect 11506 42590 11508 42642
rect 11452 42588 11508 42590
rect 10108 42028 10164 42084
rect 9436 41916 9492 41972
rect 9884 41916 9940 41972
rect 8876 39004 8932 39060
rect 8988 37996 9044 38052
rect 8540 36092 8596 36148
rect 8092 35810 8148 35812
rect 8092 35758 8094 35810
rect 8094 35758 8146 35810
rect 8146 35758 8148 35810
rect 8092 35756 8148 35758
rect 7868 35698 7924 35700
rect 7868 35646 7870 35698
rect 7870 35646 7922 35698
rect 7922 35646 7924 35698
rect 7868 35644 7924 35646
rect 8204 35644 8260 35700
rect 8428 35698 8484 35700
rect 8428 35646 8430 35698
rect 8430 35646 8482 35698
rect 8482 35646 8484 35698
rect 8428 35644 8484 35646
rect 8428 35084 8484 35140
rect 7532 34802 7588 34804
rect 7532 34750 7534 34802
rect 7534 34750 7586 34802
rect 7586 34750 7588 34802
rect 7532 34748 7588 34750
rect 7308 34018 7364 34020
rect 7308 33966 7310 34018
rect 7310 33966 7362 34018
rect 7362 33966 7364 34018
rect 7308 33964 7364 33966
rect 7420 33628 7476 33684
rect 7308 32450 7364 32452
rect 7308 32398 7310 32450
rect 7310 32398 7362 32450
rect 7362 32398 7364 32450
rect 7308 32396 7364 32398
rect 6972 31778 7028 31780
rect 6972 31726 6974 31778
rect 6974 31726 7026 31778
rect 7026 31726 7028 31778
rect 6972 31724 7028 31726
rect 6748 29426 6804 29428
rect 6748 29374 6750 29426
rect 6750 29374 6802 29426
rect 6802 29374 6804 29426
rect 6748 29372 6804 29374
rect 7084 30828 7140 30884
rect 6972 30770 7028 30772
rect 6972 30718 6974 30770
rect 6974 30718 7026 30770
rect 7026 30718 7028 30770
rect 6972 30716 7028 30718
rect 6972 29314 7028 29316
rect 6972 29262 6974 29314
rect 6974 29262 7026 29314
rect 7026 29262 7028 29314
rect 6972 29260 7028 29262
rect 6860 28812 6916 28868
rect 6412 28364 6468 28420
rect 6300 28028 6356 28084
rect 7196 28588 7252 28644
rect 6412 27356 6468 27412
rect 6524 27244 6580 27300
rect 6524 26908 6580 26964
rect 5628 24722 5684 24724
rect 5628 24670 5630 24722
rect 5630 24670 5682 24722
rect 5682 24670 5684 24722
rect 5628 24668 5684 24670
rect 6300 26066 6356 26068
rect 6300 26014 6302 26066
rect 6302 26014 6354 26066
rect 6354 26014 6356 26066
rect 6300 26012 6356 26014
rect 6860 27356 6916 27412
rect 6972 26962 7028 26964
rect 6972 26910 6974 26962
rect 6974 26910 7026 26962
rect 7026 26910 7028 26962
rect 6972 26908 7028 26910
rect 6636 26684 6692 26740
rect 6636 26460 6692 26516
rect 6748 26572 6804 26628
rect 6748 26236 6804 26292
rect 7196 27858 7252 27860
rect 7196 27806 7198 27858
rect 7198 27806 7250 27858
rect 7250 27806 7252 27858
rect 7196 27804 7252 27806
rect 7196 27020 7252 27076
rect 6860 26012 6916 26068
rect 8204 34412 8260 34468
rect 7756 33740 7812 33796
rect 7868 32562 7924 32564
rect 7868 32510 7870 32562
rect 7870 32510 7922 32562
rect 7922 32510 7924 32562
rect 7868 32508 7924 32510
rect 7532 31948 7588 32004
rect 7532 31666 7588 31668
rect 7532 31614 7534 31666
rect 7534 31614 7586 31666
rect 7586 31614 7588 31666
rect 7532 31612 7588 31614
rect 8540 34748 8596 34804
rect 9548 40236 9604 40292
rect 9324 38332 9380 38388
rect 9772 40684 9828 40740
rect 9660 38444 9716 38500
rect 9772 40460 9828 40516
rect 9436 37996 9492 38052
rect 9100 36204 9156 36260
rect 9324 37212 9380 37268
rect 8988 35756 9044 35812
rect 8876 34972 8932 35028
rect 8764 34300 8820 34356
rect 8876 34242 8932 34244
rect 8876 34190 8878 34242
rect 8878 34190 8930 34242
rect 8930 34190 8932 34242
rect 8876 34188 8932 34190
rect 8540 33628 8596 33684
rect 8652 33852 8708 33908
rect 8428 33180 8484 33236
rect 9436 36092 9492 36148
rect 9660 37436 9716 37492
rect 9660 36988 9716 37044
rect 10108 41804 10164 41860
rect 11116 42028 11172 42084
rect 10220 40684 10276 40740
rect 10108 40290 10164 40292
rect 10108 40238 10110 40290
rect 10110 40238 10162 40290
rect 10162 40238 10164 40290
rect 10108 40236 10164 40238
rect 9996 39564 10052 39620
rect 9884 38892 9940 38948
rect 10668 41970 10724 41972
rect 10668 41918 10670 41970
rect 10670 41918 10722 41970
rect 10722 41918 10724 41970
rect 10668 41916 10724 41918
rect 11004 41020 11060 41076
rect 10332 39452 10388 39508
rect 11228 40684 11284 40740
rect 10220 37548 10276 37604
rect 9996 37324 10052 37380
rect 9884 37266 9940 37268
rect 9884 37214 9886 37266
rect 9886 37214 9938 37266
rect 9938 37214 9940 37266
rect 9884 37212 9940 37214
rect 10108 37100 10164 37156
rect 9772 36204 9828 36260
rect 10332 37324 10388 37380
rect 9996 36764 10052 36820
rect 9884 35756 9940 35812
rect 9660 35698 9716 35700
rect 9660 35646 9662 35698
rect 9662 35646 9714 35698
rect 9714 35646 9716 35698
rect 9660 35644 9716 35646
rect 9548 35196 9604 35252
rect 9436 35084 9492 35140
rect 9436 34914 9492 34916
rect 9436 34862 9438 34914
rect 9438 34862 9490 34914
rect 9490 34862 9492 34914
rect 9436 34860 9492 34862
rect 10668 37212 10724 37268
rect 10892 39676 10948 39732
rect 10892 37772 10948 37828
rect 11452 40460 11508 40516
rect 11340 40402 11396 40404
rect 11340 40350 11342 40402
rect 11342 40350 11394 40402
rect 11394 40350 11396 40402
rect 11340 40348 11396 40350
rect 11900 41132 11956 41188
rect 13692 45106 13748 45108
rect 13692 45054 13694 45106
rect 13694 45054 13746 45106
rect 13746 45054 13748 45106
rect 13692 45052 13748 45054
rect 12572 43708 12628 43764
rect 12348 43596 12404 43652
rect 12908 44210 12964 44212
rect 12908 44158 12910 44210
rect 12910 44158 12962 44210
rect 12962 44158 12964 44210
rect 12908 44156 12964 44158
rect 12908 43708 12964 43764
rect 12796 43596 12852 43652
rect 12684 43484 12740 43540
rect 13132 43426 13188 43428
rect 13132 43374 13134 43426
rect 13134 43374 13186 43426
rect 13186 43374 13188 43426
rect 13132 43372 13188 43374
rect 13692 43820 13748 43876
rect 12460 42700 12516 42756
rect 12348 42028 12404 42084
rect 12908 41858 12964 41860
rect 12908 41806 12910 41858
rect 12910 41806 12962 41858
rect 12962 41806 12964 41858
rect 12908 41804 12964 41806
rect 12572 41692 12628 41748
rect 11788 40124 11844 40180
rect 11564 39788 11620 39844
rect 11788 39004 11844 39060
rect 12684 41580 12740 41636
rect 12908 41468 12964 41524
rect 12572 40796 12628 40852
rect 12348 39788 12404 39844
rect 12124 39004 12180 39060
rect 12236 39340 12292 39396
rect 11340 38780 11396 38836
rect 11340 38332 11396 38388
rect 11116 38050 11172 38052
rect 11116 37998 11118 38050
rect 11118 37998 11170 38050
rect 11170 37998 11172 38050
rect 11116 37996 11172 37998
rect 11228 37938 11284 37940
rect 11228 37886 11230 37938
rect 11230 37886 11282 37938
rect 11282 37886 11284 37938
rect 11228 37884 11284 37886
rect 10444 36764 10500 36820
rect 9884 34748 9940 34804
rect 10108 34972 10164 35028
rect 10108 34748 10164 34804
rect 9212 34188 9268 34244
rect 9436 34300 9492 34356
rect 9324 33964 9380 34020
rect 9660 33852 9716 33908
rect 9100 33516 9156 33572
rect 9212 33628 9268 33684
rect 8764 33122 8820 33124
rect 8764 33070 8766 33122
rect 8766 33070 8818 33122
rect 8818 33070 8820 33122
rect 8764 33068 8820 33070
rect 8876 32956 8932 33012
rect 8316 32508 8372 32564
rect 7756 30770 7812 30772
rect 7756 30718 7758 30770
rect 7758 30718 7810 30770
rect 7810 30718 7812 30770
rect 7756 30716 7812 30718
rect 7868 30210 7924 30212
rect 7868 30158 7870 30210
rect 7870 30158 7922 30210
rect 7922 30158 7924 30210
rect 7868 30156 7924 30158
rect 8204 31778 8260 31780
rect 8204 31726 8206 31778
rect 8206 31726 8258 31778
rect 8258 31726 8260 31778
rect 8204 31724 8260 31726
rect 8540 31666 8596 31668
rect 8540 31614 8542 31666
rect 8542 31614 8594 31666
rect 8594 31614 8596 31666
rect 8540 31612 8596 31614
rect 8988 32450 9044 32452
rect 8988 32398 8990 32450
rect 8990 32398 9042 32450
rect 9042 32398 9044 32450
rect 8988 32396 9044 32398
rect 9100 31948 9156 32004
rect 8764 31724 8820 31780
rect 8764 31388 8820 31444
rect 8204 30882 8260 30884
rect 8204 30830 8206 30882
rect 8206 30830 8258 30882
rect 8258 30830 8260 30882
rect 8204 30828 8260 30830
rect 7644 29596 7700 29652
rect 8204 30268 8260 30324
rect 8428 30156 8484 30212
rect 8764 31164 8820 31220
rect 8988 30940 9044 30996
rect 8316 29538 8372 29540
rect 8316 29486 8318 29538
rect 8318 29486 8370 29538
rect 8370 29486 8372 29538
rect 8316 29484 8372 29486
rect 8092 28642 8148 28644
rect 8092 28590 8094 28642
rect 8094 28590 8146 28642
rect 8146 28590 8148 28642
rect 8092 28588 8148 28590
rect 9996 33628 10052 33684
rect 11116 37100 11172 37156
rect 11004 36988 11060 37044
rect 11116 36764 11172 36820
rect 10892 35810 10948 35812
rect 10892 35758 10894 35810
rect 10894 35758 10946 35810
rect 10946 35758 10948 35810
rect 10892 35756 10948 35758
rect 10556 34860 10612 34916
rect 10444 34748 10500 34804
rect 10556 34300 10612 34356
rect 10332 34188 10388 34244
rect 10220 34130 10276 34132
rect 10220 34078 10222 34130
rect 10222 34078 10274 34130
rect 10274 34078 10276 34130
rect 10220 34076 10276 34078
rect 10444 33964 10500 34020
rect 10108 33404 10164 33460
rect 9884 33292 9940 33348
rect 9548 33234 9604 33236
rect 9548 33182 9550 33234
rect 9550 33182 9602 33234
rect 9602 33182 9604 33234
rect 9548 33180 9604 33182
rect 9324 32844 9380 32900
rect 9548 32620 9604 32676
rect 9324 31388 9380 31444
rect 8764 28812 8820 28868
rect 8540 28588 8596 28644
rect 8428 28476 8484 28532
rect 8204 27916 8260 27972
rect 6972 25564 7028 25620
rect 6748 25452 6804 25508
rect 6972 25116 7028 25172
rect 6076 23714 6132 23716
rect 6076 23662 6078 23714
rect 6078 23662 6130 23714
rect 6130 23662 6132 23714
rect 6076 23660 6132 23662
rect 6300 23772 6356 23828
rect 6412 24444 6468 24500
rect 6524 23884 6580 23940
rect 6300 23548 6356 23604
rect 6748 24610 6804 24612
rect 6748 24558 6750 24610
rect 6750 24558 6802 24610
rect 6802 24558 6804 24610
rect 6748 24556 6804 24558
rect 7868 27692 7924 27748
rect 8092 27020 8148 27076
rect 7196 26236 7252 26292
rect 7644 26124 7700 26180
rect 7756 26012 7812 26068
rect 6748 23938 6804 23940
rect 6748 23886 6750 23938
rect 6750 23886 6802 23938
rect 6802 23886 6804 23938
rect 6748 23884 6804 23886
rect 7868 25900 7924 25956
rect 8092 26290 8148 26292
rect 8092 26238 8094 26290
rect 8094 26238 8146 26290
rect 8146 26238 8148 26290
rect 8092 26236 8148 26238
rect 8204 25788 8260 25844
rect 8764 27132 8820 27188
rect 8652 27074 8708 27076
rect 8652 27022 8654 27074
rect 8654 27022 8706 27074
rect 8706 27022 8708 27074
rect 8652 27020 8708 27022
rect 10332 33852 10388 33908
rect 9996 32562 10052 32564
rect 9996 32510 9998 32562
rect 9998 32510 10050 32562
rect 10050 32510 10052 32562
rect 9996 32508 10052 32510
rect 9660 32450 9716 32452
rect 9660 32398 9662 32450
rect 9662 32398 9714 32450
rect 9714 32398 9716 32450
rect 9660 32396 9716 32398
rect 9772 32172 9828 32228
rect 9660 31948 9716 32004
rect 9548 31218 9604 31220
rect 9548 31166 9550 31218
rect 9550 31166 9602 31218
rect 9602 31166 9604 31218
rect 9548 31164 9604 31166
rect 9436 31052 9492 31108
rect 9548 30994 9604 30996
rect 9548 30942 9550 30994
rect 9550 30942 9602 30994
rect 9602 30942 9604 30994
rect 9548 30940 9604 30942
rect 10332 32844 10388 32900
rect 9772 31388 9828 31444
rect 10108 31612 10164 31668
rect 9660 30716 9716 30772
rect 9772 31106 9828 31108
rect 9772 31054 9774 31106
rect 9774 31054 9826 31106
rect 9826 31054 9828 31106
rect 9772 31052 9828 31054
rect 9660 29650 9716 29652
rect 9660 29598 9662 29650
rect 9662 29598 9714 29650
rect 9714 29598 9716 29650
rect 9660 29596 9716 29598
rect 10108 30994 10164 30996
rect 10108 30942 10110 30994
rect 10110 30942 10162 30994
rect 10162 30942 10164 30994
rect 10108 30940 10164 30942
rect 8988 27580 9044 27636
rect 8316 26796 8372 26852
rect 8092 25506 8148 25508
rect 8092 25454 8094 25506
rect 8094 25454 8146 25506
rect 8146 25454 8148 25506
rect 8092 25452 8148 25454
rect 7196 23884 7252 23940
rect 6860 23826 6916 23828
rect 6860 23774 6862 23826
rect 6862 23774 6914 23826
rect 6914 23774 6916 23826
rect 6860 23772 6916 23774
rect 6636 23324 6692 23380
rect 6524 23212 6580 23268
rect 5852 22764 5908 22820
rect 7196 22764 7252 22820
rect 7420 23100 7476 23156
rect 7308 22482 7364 22484
rect 7308 22430 7310 22482
rect 7310 22430 7362 22482
rect 7362 22430 7364 22482
rect 7308 22428 7364 22430
rect 6748 22204 6804 22260
rect 6076 22092 6132 22148
rect 5628 21810 5684 21812
rect 5628 21758 5630 21810
rect 5630 21758 5682 21810
rect 5682 21758 5684 21810
rect 5628 21756 5684 21758
rect 5068 21532 5124 21588
rect 4620 21308 4676 21364
rect 4476 21194 4532 21196
rect 4476 21142 4478 21194
rect 4478 21142 4530 21194
rect 4530 21142 4532 21194
rect 4476 21140 4532 21142
rect 4580 21194 4636 21196
rect 4580 21142 4582 21194
rect 4582 21142 4634 21194
rect 4634 21142 4636 21194
rect 4580 21140 4636 21142
rect 4684 21194 4740 21196
rect 4684 21142 4686 21194
rect 4686 21142 4738 21194
rect 4738 21142 4740 21194
rect 4684 21140 4740 21142
rect 5180 21474 5236 21476
rect 5180 21422 5182 21474
rect 5182 21422 5234 21474
rect 5234 21422 5236 21474
rect 5180 21420 5236 21422
rect 3612 20130 3668 20132
rect 3612 20078 3614 20130
rect 3614 20078 3666 20130
rect 3666 20078 3668 20130
rect 3612 20076 3668 20078
rect 2492 19852 2548 19908
rect 3500 19964 3556 20020
rect 1820 18450 1876 18452
rect 1820 18398 1822 18450
rect 1822 18398 1874 18450
rect 1874 18398 1876 18450
rect 1820 18396 1876 18398
rect 1708 16716 1764 16772
rect 2492 18338 2548 18340
rect 2492 18286 2494 18338
rect 2494 18286 2546 18338
rect 2546 18286 2548 18338
rect 2492 18284 2548 18286
rect 1932 17778 1988 17780
rect 1932 17726 1934 17778
rect 1934 17726 1986 17778
rect 1986 17726 1988 17778
rect 1932 17724 1988 17726
rect 3276 17106 3332 17108
rect 3276 17054 3278 17106
rect 3278 17054 3330 17106
rect 3330 17054 3332 17106
rect 3276 17052 3332 17054
rect 2828 16882 2884 16884
rect 2828 16830 2830 16882
rect 2830 16830 2882 16882
rect 2882 16830 2884 16882
rect 2828 16828 2884 16830
rect 3164 16770 3220 16772
rect 3164 16718 3166 16770
rect 3166 16718 3218 16770
rect 3218 16718 3220 16770
rect 3164 16716 3220 16718
rect 3500 19346 3556 19348
rect 3500 19294 3502 19346
rect 3502 19294 3554 19346
rect 3554 19294 3556 19346
rect 3500 19292 3556 19294
rect 3612 19180 3668 19236
rect 4172 20130 4228 20132
rect 4172 20078 4174 20130
rect 4174 20078 4226 20130
rect 4226 20078 4228 20130
rect 4172 20076 4228 20078
rect 4060 19906 4116 19908
rect 4060 19854 4062 19906
rect 4062 19854 4114 19906
rect 4114 19854 4116 19906
rect 4060 19852 4116 19854
rect 5740 20188 5796 20244
rect 5852 21532 5908 21588
rect 4396 20018 4452 20020
rect 4396 19966 4398 20018
rect 4398 19966 4450 20018
rect 4450 19966 4452 20018
rect 4396 19964 4452 19966
rect 5628 20076 5684 20132
rect 4956 19906 5012 19908
rect 4956 19854 4958 19906
rect 4958 19854 5010 19906
rect 5010 19854 5012 19906
rect 4956 19852 5012 19854
rect 4732 19740 4788 19796
rect 4476 19626 4532 19628
rect 4476 19574 4478 19626
rect 4478 19574 4530 19626
rect 4530 19574 4532 19626
rect 4476 19572 4532 19574
rect 4580 19626 4636 19628
rect 4580 19574 4582 19626
rect 4582 19574 4634 19626
rect 4634 19574 4636 19626
rect 4580 19572 4636 19574
rect 4684 19626 4740 19628
rect 4684 19574 4686 19626
rect 4686 19574 4738 19626
rect 4738 19574 4740 19626
rect 4684 19572 4740 19574
rect 3948 19234 4004 19236
rect 3948 19182 3950 19234
rect 3950 19182 4002 19234
rect 4002 19182 4004 19234
rect 3948 19180 4004 19182
rect 4844 19458 4900 19460
rect 4844 19406 4846 19458
rect 4846 19406 4898 19458
rect 4898 19406 4900 19458
rect 4844 19404 4900 19406
rect 3836 18956 3892 19012
rect 4060 18396 4116 18452
rect 3948 17836 4004 17892
rect 3836 17276 3892 17332
rect 3388 16716 3444 16772
rect 3500 16828 3556 16884
rect 2492 15148 2548 15204
rect 4284 19010 4340 19012
rect 4284 18958 4286 19010
rect 4286 18958 4338 19010
rect 4338 18958 4340 19010
rect 4284 18956 4340 18958
rect 5068 19180 5124 19236
rect 5180 19404 5236 19460
rect 4620 18396 4676 18452
rect 4844 18508 4900 18564
rect 4172 18172 4228 18228
rect 4476 18058 4532 18060
rect 4476 18006 4478 18058
rect 4478 18006 4530 18058
rect 4530 18006 4532 18058
rect 4476 18004 4532 18006
rect 4580 18058 4636 18060
rect 4580 18006 4582 18058
rect 4582 18006 4634 18058
rect 4634 18006 4636 18058
rect 4580 18004 4636 18006
rect 4684 18058 4740 18060
rect 4684 18006 4686 18058
rect 4686 18006 4738 18058
rect 4738 18006 4740 18058
rect 4684 18004 4740 18006
rect 4172 17052 4228 17108
rect 4508 16604 4564 16660
rect 4476 16490 4532 16492
rect 4476 16438 4478 16490
rect 4478 16438 4530 16490
rect 4530 16438 4532 16490
rect 4476 16436 4532 16438
rect 4580 16490 4636 16492
rect 4580 16438 4582 16490
rect 4582 16438 4634 16490
rect 4634 16438 4636 16490
rect 4580 16436 4636 16438
rect 4684 16490 4740 16492
rect 4684 16438 4686 16490
rect 4686 16438 4738 16490
rect 4738 16438 4740 16490
rect 4684 16436 4740 16438
rect 3612 16268 3668 16324
rect 4620 16156 4676 16212
rect 5292 19292 5348 19348
rect 5292 18956 5348 19012
rect 5740 19906 5796 19908
rect 5740 19854 5742 19906
rect 5742 19854 5794 19906
rect 5794 19854 5796 19906
rect 5740 19852 5796 19854
rect 5404 19180 5460 19236
rect 5068 18562 5124 18564
rect 5068 18510 5070 18562
rect 5070 18510 5122 18562
rect 5122 18510 5124 18562
rect 5068 18508 5124 18510
rect 5180 18338 5236 18340
rect 5180 18286 5182 18338
rect 5182 18286 5234 18338
rect 5234 18286 5236 18338
rect 5180 18284 5236 18286
rect 5180 17948 5236 18004
rect 5068 17442 5124 17444
rect 5068 17390 5070 17442
rect 5070 17390 5122 17442
rect 5122 17390 5124 17442
rect 5068 17388 5124 17390
rect 5068 17106 5124 17108
rect 5068 17054 5070 17106
rect 5070 17054 5122 17106
rect 5122 17054 5124 17106
rect 5068 17052 5124 17054
rect 5292 16994 5348 16996
rect 5292 16942 5294 16994
rect 5294 16942 5346 16994
rect 5346 16942 5348 16994
rect 5292 16940 5348 16942
rect 5292 16716 5348 16772
rect 4956 16604 5012 16660
rect 5180 16492 5236 16548
rect 5068 16210 5124 16212
rect 5068 16158 5070 16210
rect 5070 16158 5122 16210
rect 5122 16158 5124 16210
rect 5068 16156 5124 16158
rect 4956 15260 5012 15316
rect 2492 13580 2548 13636
rect 3164 12402 3220 12404
rect 3164 12350 3166 12402
rect 3166 12350 3218 12402
rect 3218 12350 3220 12402
rect 3164 12348 3220 12350
rect 3612 12236 3668 12292
rect 2492 12012 2548 12068
rect 3276 12066 3332 12068
rect 3276 12014 3278 12066
rect 3278 12014 3330 12066
rect 3330 12014 3332 12066
rect 3276 12012 3332 12014
rect 3388 11564 3444 11620
rect 1708 9938 1764 9940
rect 1708 9886 1710 9938
rect 1710 9886 1762 9938
rect 1762 9886 1764 9938
rect 1708 9884 1764 9886
rect 2492 9212 2548 9268
rect 1820 8258 1876 8260
rect 1820 8206 1822 8258
rect 1822 8206 1874 8258
rect 1874 8206 1876 8258
rect 1820 8204 1876 8206
rect 3276 8204 3332 8260
rect 4844 15202 4900 15204
rect 4844 15150 4846 15202
rect 4846 15150 4898 15202
rect 4898 15150 4900 15202
rect 4844 15148 4900 15150
rect 4476 14922 4532 14924
rect 4476 14870 4478 14922
rect 4478 14870 4530 14922
rect 4530 14870 4532 14922
rect 4476 14868 4532 14870
rect 4580 14922 4636 14924
rect 4580 14870 4582 14922
rect 4582 14870 4634 14922
rect 4634 14870 4636 14922
rect 4580 14868 4636 14870
rect 4684 14922 4740 14924
rect 4684 14870 4686 14922
rect 4686 14870 4738 14922
rect 4738 14870 4740 14922
rect 4684 14868 4740 14870
rect 4620 14642 4676 14644
rect 4620 14590 4622 14642
rect 4622 14590 4674 14642
rect 4674 14590 4676 14642
rect 4620 14588 4676 14590
rect 5068 14028 5124 14084
rect 4732 13634 4788 13636
rect 4732 13582 4734 13634
rect 4734 13582 4786 13634
rect 4786 13582 4788 13634
rect 4732 13580 4788 13582
rect 4476 13354 4532 13356
rect 4476 13302 4478 13354
rect 4478 13302 4530 13354
rect 4530 13302 4532 13354
rect 4476 13300 4532 13302
rect 4580 13354 4636 13356
rect 4580 13302 4582 13354
rect 4582 13302 4634 13354
rect 4634 13302 4636 13354
rect 4580 13300 4636 13302
rect 4684 13354 4740 13356
rect 4684 13302 4686 13354
rect 4686 13302 4738 13354
rect 4738 13302 4740 13354
rect 4684 13300 4740 13302
rect 5292 15260 5348 15316
rect 6748 21644 6804 21700
rect 5964 20076 6020 20132
rect 6076 19964 6132 20020
rect 6524 20802 6580 20804
rect 6524 20750 6526 20802
rect 6526 20750 6578 20802
rect 6578 20750 6580 20802
rect 6524 20748 6580 20750
rect 6412 19906 6468 19908
rect 6412 19854 6414 19906
rect 6414 19854 6466 19906
rect 6466 19854 6468 19906
rect 6412 19852 6468 19854
rect 6524 20188 6580 20244
rect 6076 18956 6132 19012
rect 5740 17948 5796 18004
rect 5852 17724 5908 17780
rect 5628 17666 5684 17668
rect 5628 17614 5630 17666
rect 5630 17614 5682 17666
rect 5682 17614 5684 17666
rect 5628 17612 5684 17614
rect 5964 17554 6020 17556
rect 5964 17502 5966 17554
rect 5966 17502 6018 17554
rect 6018 17502 6020 17554
rect 5964 17500 6020 17502
rect 5740 17442 5796 17444
rect 5740 17390 5742 17442
rect 5742 17390 5794 17442
rect 5794 17390 5796 17442
rect 5740 17388 5796 17390
rect 5628 16604 5684 16660
rect 6076 16716 6132 16772
rect 5852 16268 5908 16324
rect 6972 21810 7028 21812
rect 6972 21758 6974 21810
rect 6974 21758 7026 21810
rect 7026 21758 7028 21810
rect 6972 21756 7028 21758
rect 7420 21420 7476 21476
rect 6524 18060 6580 18116
rect 6860 20018 6916 20020
rect 6860 19966 6862 20018
rect 6862 19966 6914 20018
rect 6914 19966 6916 20018
rect 6860 19964 6916 19966
rect 6300 17612 6356 17668
rect 6636 17500 6692 17556
rect 7420 20300 7476 20356
rect 8988 27244 9044 27300
rect 9100 27132 9156 27188
rect 8204 23996 8260 24052
rect 8652 25788 8708 25844
rect 7644 23042 7700 23044
rect 7644 22990 7646 23042
rect 7646 22990 7698 23042
rect 7698 22990 7700 23042
rect 7644 22988 7700 22990
rect 8092 22652 8148 22708
rect 7756 22146 7812 22148
rect 7756 22094 7758 22146
rect 7758 22094 7810 22146
rect 7810 22094 7812 22146
rect 7756 22092 7812 22094
rect 7868 21756 7924 21812
rect 8652 23660 8708 23716
rect 8988 26514 9044 26516
rect 8988 26462 8990 26514
rect 8990 26462 9042 26514
rect 9042 26462 9044 26514
rect 8988 26460 9044 26462
rect 8876 24556 8932 24612
rect 9436 28812 9492 28868
rect 9772 29148 9828 29204
rect 10108 29036 10164 29092
rect 9772 28642 9828 28644
rect 9772 28590 9774 28642
rect 9774 28590 9826 28642
rect 9826 28590 9828 28642
rect 9772 28588 9828 28590
rect 9772 27746 9828 27748
rect 9772 27694 9774 27746
rect 9774 27694 9826 27746
rect 9826 27694 9828 27746
rect 9772 27692 9828 27694
rect 9548 27580 9604 27636
rect 10108 27858 10164 27860
rect 10108 27806 10110 27858
rect 10110 27806 10162 27858
rect 10162 27806 10164 27858
rect 10108 27804 10164 27806
rect 9996 27580 10052 27636
rect 10108 27468 10164 27524
rect 11676 37378 11732 37380
rect 11676 37326 11678 37378
rect 11678 37326 11730 37378
rect 11730 37326 11732 37378
rect 11676 37324 11732 37326
rect 11564 37266 11620 37268
rect 11564 37214 11566 37266
rect 11566 37214 11618 37266
rect 11618 37214 11620 37266
rect 11564 37212 11620 37214
rect 11452 36764 11508 36820
rect 11340 35810 11396 35812
rect 11340 35758 11342 35810
rect 11342 35758 11394 35810
rect 11394 35758 11396 35810
rect 11340 35756 11396 35758
rect 11116 35196 11172 35252
rect 10892 35084 10948 35140
rect 10556 33628 10612 33684
rect 10668 33180 10724 33236
rect 10668 31948 10724 32004
rect 10668 31500 10724 31556
rect 10780 31612 10836 31668
rect 10556 30492 10612 30548
rect 11340 35084 11396 35140
rect 11116 34748 11172 34804
rect 11564 36706 11620 36708
rect 11564 36654 11566 36706
rect 11566 36654 11618 36706
rect 11618 36654 11620 36706
rect 11564 36652 11620 36654
rect 11676 36540 11732 36596
rect 11340 34300 11396 34356
rect 11452 34636 11508 34692
rect 11452 33740 11508 33796
rect 11116 33404 11172 33460
rect 11116 32060 11172 32116
rect 11340 31948 11396 32004
rect 11004 31778 11060 31780
rect 11004 31726 11006 31778
rect 11006 31726 11058 31778
rect 11058 31726 11060 31778
rect 11004 31724 11060 31726
rect 10668 30380 10724 30436
rect 11116 31388 11172 31444
rect 10444 29932 10500 29988
rect 11116 30604 11172 30660
rect 11228 30380 11284 30436
rect 10892 30156 10948 30212
rect 10556 29596 10612 29652
rect 10668 29484 10724 29540
rect 10332 29202 10388 29204
rect 10332 29150 10334 29202
rect 10334 29150 10386 29202
rect 10386 29150 10388 29202
rect 10332 29148 10388 29150
rect 10556 29202 10612 29204
rect 10556 29150 10558 29202
rect 10558 29150 10610 29202
rect 10610 29150 10612 29202
rect 10556 29148 10612 29150
rect 10444 29036 10500 29092
rect 10444 28700 10500 28756
rect 10332 27804 10388 27860
rect 9324 27020 9380 27076
rect 10332 26796 10388 26852
rect 9996 26290 10052 26292
rect 9996 26238 9998 26290
rect 9998 26238 10050 26290
rect 10050 26238 10052 26290
rect 9996 26236 10052 26238
rect 10556 26908 10612 26964
rect 11116 29538 11172 29540
rect 11116 29486 11118 29538
rect 11118 29486 11170 29538
rect 11170 29486 11172 29538
rect 11116 29484 11172 29486
rect 11004 29036 11060 29092
rect 10780 27804 10836 27860
rect 10892 28588 10948 28644
rect 10668 26796 10724 26852
rect 10780 27020 10836 27076
rect 11228 28642 11284 28644
rect 11228 28590 11230 28642
rect 11230 28590 11282 28642
rect 11282 28590 11284 28642
rect 11228 28588 11284 28590
rect 11228 27692 11284 27748
rect 11676 34802 11732 34804
rect 11676 34750 11678 34802
rect 11678 34750 11730 34802
rect 11730 34750 11732 34802
rect 11676 34748 11732 34750
rect 12348 38050 12404 38052
rect 12348 37998 12350 38050
rect 12350 37998 12402 38050
rect 12402 37998 12404 38050
rect 12348 37996 12404 37998
rect 12460 37938 12516 37940
rect 12460 37886 12462 37938
rect 12462 37886 12514 37938
rect 12514 37886 12516 37938
rect 12460 37884 12516 37886
rect 12460 37660 12516 37716
rect 12348 36258 12404 36260
rect 12348 36206 12350 36258
rect 12350 36206 12402 36258
rect 12402 36206 12404 36258
rect 12348 36204 12404 36206
rect 12348 35420 12404 35476
rect 12236 35196 12292 35252
rect 12124 33516 12180 33572
rect 12012 33404 12068 33460
rect 13020 40514 13076 40516
rect 13020 40462 13022 40514
rect 13022 40462 13074 40514
rect 13074 40462 13076 40514
rect 13020 40460 13076 40462
rect 12908 39788 12964 39844
rect 12684 39340 12740 39396
rect 12796 37212 12852 37268
rect 12796 36764 12852 36820
rect 12908 36540 12964 36596
rect 13020 36204 13076 36260
rect 12908 34914 12964 34916
rect 12908 34862 12910 34914
rect 12910 34862 12962 34914
rect 12962 34862 12964 34914
rect 12908 34860 12964 34862
rect 12572 34412 12628 34468
rect 12460 34242 12516 34244
rect 12460 34190 12462 34242
rect 12462 34190 12514 34242
rect 12514 34190 12516 34242
rect 12460 34188 12516 34190
rect 12684 34188 12740 34244
rect 12348 33404 12404 33460
rect 11676 33122 11732 33124
rect 11676 33070 11678 33122
rect 11678 33070 11730 33122
rect 11730 33070 11732 33122
rect 11676 33068 11732 33070
rect 11788 32562 11844 32564
rect 11788 32510 11790 32562
rect 11790 32510 11842 32562
rect 11842 32510 11844 32562
rect 11788 32508 11844 32510
rect 12012 32396 12068 32452
rect 11564 31778 11620 31780
rect 11564 31726 11566 31778
rect 11566 31726 11618 31778
rect 11618 31726 11620 31778
rect 11564 31724 11620 31726
rect 11452 31666 11508 31668
rect 11452 31614 11454 31666
rect 11454 31614 11506 31666
rect 11506 31614 11508 31666
rect 11452 31612 11508 31614
rect 11564 30994 11620 30996
rect 11564 30942 11566 30994
rect 11566 30942 11618 30994
rect 11618 30942 11620 30994
rect 11564 30940 11620 30942
rect 12236 32396 12292 32452
rect 12348 32956 12404 33012
rect 12124 31778 12180 31780
rect 12124 31726 12126 31778
rect 12126 31726 12178 31778
rect 12178 31726 12180 31778
rect 12124 31724 12180 31726
rect 11788 29314 11844 29316
rect 11788 29262 11790 29314
rect 11790 29262 11842 29314
rect 11842 29262 11844 29314
rect 11788 29260 11844 29262
rect 11340 27356 11396 27412
rect 11116 27186 11172 27188
rect 11116 27134 11118 27186
rect 11118 27134 11170 27186
rect 11170 27134 11172 27186
rect 11116 27132 11172 27134
rect 10892 26460 10948 26516
rect 10108 26124 10164 26180
rect 9884 25900 9940 25956
rect 9548 25788 9604 25844
rect 10108 25788 10164 25844
rect 9324 25564 9380 25620
rect 10444 25506 10500 25508
rect 10444 25454 10446 25506
rect 10446 25454 10498 25506
rect 10498 25454 10500 25506
rect 10444 25452 10500 25454
rect 9212 23772 9268 23828
rect 8988 23660 9044 23716
rect 9212 23548 9268 23604
rect 8652 23266 8708 23268
rect 8652 23214 8654 23266
rect 8654 23214 8706 23266
rect 8706 23214 8708 23266
rect 8652 23212 8708 23214
rect 8428 22652 8484 22708
rect 8764 22764 8820 22820
rect 8876 22258 8932 22260
rect 8876 22206 8878 22258
rect 8878 22206 8930 22258
rect 8930 22206 8932 22258
rect 8876 22204 8932 22206
rect 7644 21698 7700 21700
rect 7644 21646 7646 21698
rect 7646 21646 7698 21698
rect 7698 21646 7700 21698
rect 7644 21644 7700 21646
rect 7532 20188 7588 20244
rect 7420 19906 7476 19908
rect 7420 19854 7422 19906
rect 7422 19854 7474 19906
rect 7474 19854 7476 19906
rect 7420 19852 7476 19854
rect 7420 19010 7476 19012
rect 7420 18958 7422 19010
rect 7422 18958 7474 19010
rect 7474 18958 7476 19010
rect 7420 18956 7476 18958
rect 8092 21644 8148 21700
rect 8764 21868 8820 21924
rect 8652 21810 8708 21812
rect 8652 21758 8654 21810
rect 8654 21758 8706 21810
rect 8706 21758 8708 21810
rect 8652 21756 8708 21758
rect 8428 21196 8484 21252
rect 8988 21420 9044 21476
rect 7868 20802 7924 20804
rect 7868 20750 7870 20802
rect 7870 20750 7922 20802
rect 7922 20750 7924 20802
rect 7868 20748 7924 20750
rect 8876 20802 8932 20804
rect 8876 20750 8878 20802
rect 8878 20750 8930 20802
rect 8930 20750 8932 20802
rect 8876 20748 8932 20750
rect 8204 20188 8260 20244
rect 8652 20076 8708 20132
rect 9212 22428 9268 22484
rect 9996 25116 10052 25172
rect 9548 24722 9604 24724
rect 9548 24670 9550 24722
rect 9550 24670 9602 24722
rect 9602 24670 9604 24722
rect 9548 24668 9604 24670
rect 9996 23660 10052 23716
rect 10780 24834 10836 24836
rect 10780 24782 10782 24834
rect 10782 24782 10834 24834
rect 10834 24782 10836 24834
rect 10780 24780 10836 24782
rect 10556 23660 10612 23716
rect 10108 23548 10164 23604
rect 9436 23324 9492 23380
rect 10108 23212 10164 23268
rect 9660 23154 9716 23156
rect 9660 23102 9662 23154
rect 9662 23102 9714 23154
rect 9714 23102 9716 23154
rect 9660 23100 9716 23102
rect 9436 22876 9492 22932
rect 9772 22428 9828 22484
rect 9884 22876 9940 22932
rect 9324 22258 9380 22260
rect 9324 22206 9326 22258
rect 9326 22206 9378 22258
rect 9378 22206 9380 22258
rect 9324 22204 9380 22206
rect 9100 20300 9156 20356
rect 8540 20018 8596 20020
rect 8540 19966 8542 20018
rect 8542 19966 8594 20018
rect 8594 19966 8596 20018
rect 8540 19964 8596 19966
rect 8764 19740 8820 19796
rect 8428 19234 8484 19236
rect 8428 19182 8430 19234
rect 8430 19182 8482 19234
rect 8482 19182 8484 19234
rect 8428 19180 8484 19182
rect 8204 18956 8260 19012
rect 7084 18172 7140 18228
rect 7308 18172 7364 18228
rect 6972 17948 7028 18004
rect 7084 17778 7140 17780
rect 7084 17726 7086 17778
rect 7086 17726 7138 17778
rect 7138 17726 7140 17778
rect 7084 17724 7140 17726
rect 7196 17612 7252 17668
rect 6748 17276 6804 17332
rect 6636 16380 6692 16436
rect 6188 16210 6244 16212
rect 6188 16158 6190 16210
rect 6190 16158 6242 16210
rect 6242 16158 6244 16210
rect 6188 16156 6244 16158
rect 7868 18060 7924 18116
rect 8204 17948 8260 18004
rect 7980 17388 8036 17444
rect 7420 16492 7476 16548
rect 7084 15426 7140 15428
rect 7084 15374 7086 15426
rect 7086 15374 7138 15426
rect 7138 15374 7140 15426
rect 7084 15372 7140 15374
rect 6860 15314 6916 15316
rect 6860 15262 6862 15314
rect 6862 15262 6914 15314
rect 6914 15262 6916 15314
rect 6860 15260 6916 15262
rect 7420 16098 7476 16100
rect 7420 16046 7422 16098
rect 7422 16046 7474 16098
rect 7474 16046 7476 16098
rect 7420 16044 7476 16046
rect 9548 20018 9604 20020
rect 9548 19966 9550 20018
rect 9550 19966 9602 20018
rect 9602 19966 9604 20018
rect 9548 19964 9604 19966
rect 9436 19852 9492 19908
rect 10556 23154 10612 23156
rect 10556 23102 10558 23154
rect 10558 23102 10610 23154
rect 10610 23102 10612 23154
rect 10556 23100 10612 23102
rect 10332 22764 10388 22820
rect 10444 22370 10500 22372
rect 10444 22318 10446 22370
rect 10446 22318 10498 22370
rect 10498 22318 10500 22370
rect 10444 22316 10500 22318
rect 9996 22258 10052 22260
rect 9996 22206 9998 22258
rect 9998 22206 10050 22258
rect 10050 22206 10052 22258
rect 9996 22204 10052 22206
rect 10892 24722 10948 24724
rect 10892 24670 10894 24722
rect 10894 24670 10946 24722
rect 10946 24670 10948 24722
rect 10892 24668 10948 24670
rect 10780 23548 10836 23604
rect 10892 23772 10948 23828
rect 10332 21308 10388 21364
rect 9772 20076 9828 20132
rect 9772 19852 9828 19908
rect 9324 19122 9380 19124
rect 9324 19070 9326 19122
rect 9326 19070 9378 19122
rect 9378 19070 9380 19122
rect 9324 19068 9380 19070
rect 9100 18732 9156 18788
rect 8988 18508 9044 18564
rect 8652 17500 8708 17556
rect 8540 17388 8596 17444
rect 8428 17276 8484 17332
rect 9100 17500 9156 17556
rect 8092 16882 8148 16884
rect 8092 16830 8094 16882
rect 8094 16830 8146 16882
rect 8146 16830 8148 16882
rect 8092 16828 8148 16830
rect 8540 16828 8596 16884
rect 7644 16210 7700 16212
rect 7644 16158 7646 16210
rect 7646 16158 7698 16210
rect 7698 16158 7700 16210
rect 7644 16156 7700 16158
rect 8428 16156 8484 16212
rect 8092 16098 8148 16100
rect 8092 16046 8094 16098
rect 8094 16046 8146 16098
rect 8146 16046 8148 16098
rect 8092 16044 8148 16046
rect 6076 14588 6132 14644
rect 5852 14028 5908 14084
rect 4732 13132 4788 13188
rect 4620 12796 4676 12852
rect 4284 12402 4340 12404
rect 4284 12350 4286 12402
rect 4286 12350 4338 12402
rect 4338 12350 4340 12402
rect 4284 12348 4340 12350
rect 5404 13916 5460 13972
rect 5180 13132 5236 13188
rect 4732 12236 4788 12292
rect 3836 12178 3892 12180
rect 3836 12126 3838 12178
rect 3838 12126 3890 12178
rect 3890 12126 3892 12178
rect 3836 12124 3892 12126
rect 4508 12178 4564 12180
rect 4508 12126 4510 12178
rect 4510 12126 4562 12178
rect 4562 12126 4564 12178
rect 4508 12124 4564 12126
rect 5292 13020 5348 13076
rect 5068 12850 5124 12852
rect 5068 12798 5070 12850
rect 5070 12798 5122 12850
rect 5122 12798 5124 12850
rect 5068 12796 5124 12798
rect 4476 11786 4532 11788
rect 4476 11734 4478 11786
rect 4478 11734 4530 11786
rect 4530 11734 4532 11786
rect 4476 11732 4532 11734
rect 4580 11786 4636 11788
rect 4580 11734 4582 11786
rect 4582 11734 4634 11786
rect 4634 11734 4636 11786
rect 4580 11732 4636 11734
rect 4684 11786 4740 11788
rect 4684 11734 4686 11786
rect 4686 11734 4738 11786
rect 4738 11734 4740 11786
rect 4684 11732 4740 11734
rect 5292 12178 5348 12180
rect 5292 12126 5294 12178
rect 5294 12126 5346 12178
rect 5346 12126 5348 12178
rect 5292 12124 5348 12126
rect 4732 11564 4788 11620
rect 4620 11506 4676 11508
rect 4620 11454 4622 11506
rect 4622 11454 4674 11506
rect 4674 11454 4676 11506
rect 4620 11452 4676 11454
rect 5068 11282 5124 11284
rect 5068 11230 5070 11282
rect 5070 11230 5122 11282
rect 5122 11230 5124 11282
rect 5068 11228 5124 11230
rect 4956 10610 5012 10612
rect 4956 10558 4958 10610
rect 4958 10558 5010 10610
rect 5010 10558 5012 10610
rect 4956 10556 5012 10558
rect 5292 10556 5348 10612
rect 3836 9266 3892 9268
rect 3836 9214 3838 9266
rect 3838 9214 3890 9266
rect 3890 9214 3892 9266
rect 3836 9212 3892 9214
rect 4060 9212 4116 9268
rect 3948 9042 4004 9044
rect 3948 8990 3950 9042
rect 3950 8990 4002 9042
rect 4002 8990 4004 9042
rect 3948 8988 4004 8990
rect 4476 10218 4532 10220
rect 4476 10166 4478 10218
rect 4478 10166 4530 10218
rect 4530 10166 4532 10218
rect 4476 10164 4532 10166
rect 4580 10218 4636 10220
rect 4580 10166 4582 10218
rect 4582 10166 4634 10218
rect 4634 10166 4636 10218
rect 4580 10164 4636 10166
rect 4684 10218 4740 10220
rect 4684 10166 4686 10218
rect 4686 10166 4738 10218
rect 4738 10166 4740 10218
rect 4684 10164 4740 10166
rect 5292 9996 5348 10052
rect 6636 14028 6692 14084
rect 7196 14028 7252 14084
rect 7868 15260 7924 15316
rect 5852 12796 5908 12852
rect 5740 12738 5796 12740
rect 5740 12686 5742 12738
rect 5742 12686 5794 12738
rect 5794 12686 5796 12738
rect 5740 12684 5796 12686
rect 5628 11452 5684 11508
rect 9548 18396 9604 18452
rect 9884 19068 9940 19124
rect 10892 21868 10948 21924
rect 10668 20860 10724 20916
rect 10556 20690 10612 20692
rect 10556 20638 10558 20690
rect 10558 20638 10610 20690
rect 10610 20638 10612 20690
rect 10556 20636 10612 20638
rect 10892 20748 10948 20804
rect 11340 26796 11396 26852
rect 11564 28082 11620 28084
rect 11564 28030 11566 28082
rect 11566 28030 11618 28082
rect 11618 28030 11620 28082
rect 11564 28028 11620 28030
rect 11788 28252 11844 28308
rect 11788 28028 11844 28084
rect 11900 27692 11956 27748
rect 12012 27468 12068 27524
rect 12124 28812 12180 28868
rect 11900 27244 11956 27300
rect 11564 27132 11620 27188
rect 11788 27132 11844 27188
rect 11900 27074 11956 27076
rect 11900 27022 11902 27074
rect 11902 27022 11954 27074
rect 11954 27022 11956 27074
rect 11900 27020 11956 27022
rect 11564 26850 11620 26852
rect 11564 26798 11566 26850
rect 11566 26798 11618 26850
rect 11618 26798 11620 26850
rect 11564 26796 11620 26798
rect 11452 26460 11508 26516
rect 12236 28588 12292 28644
rect 12460 32508 12516 32564
rect 12796 34130 12852 34132
rect 12796 34078 12798 34130
rect 12798 34078 12850 34130
rect 12850 34078 12852 34130
rect 12796 34076 12852 34078
rect 13020 34130 13076 34132
rect 13020 34078 13022 34130
rect 13022 34078 13074 34130
rect 13074 34078 13076 34130
rect 13020 34076 13076 34078
rect 13356 41692 13412 41748
rect 13244 40124 13300 40180
rect 13916 43484 13972 43540
rect 13692 43372 13748 43428
rect 13804 43260 13860 43316
rect 13580 41804 13636 41860
rect 13580 41132 13636 41188
rect 13580 40962 13636 40964
rect 13580 40910 13582 40962
rect 13582 40910 13634 40962
rect 13634 40910 13636 40962
rect 13580 40908 13636 40910
rect 13804 42364 13860 42420
rect 14028 43036 14084 43092
rect 14028 42812 14084 42868
rect 14028 42476 14084 42532
rect 14140 43820 14196 43876
rect 14028 41970 14084 41972
rect 14028 41918 14030 41970
rect 14030 41918 14082 41970
rect 14082 41918 14084 41970
rect 14028 41916 14084 41918
rect 13804 41244 13860 41300
rect 13916 41132 13972 41188
rect 13468 39842 13524 39844
rect 13468 39790 13470 39842
rect 13470 39790 13522 39842
rect 13522 39790 13524 39842
rect 13468 39788 13524 39790
rect 13692 40402 13748 40404
rect 13692 40350 13694 40402
rect 13694 40350 13746 40402
rect 13746 40350 13748 40402
rect 13692 40348 13748 40350
rect 14252 43260 14308 43316
rect 14476 43596 14532 43652
rect 14700 43708 14756 43764
rect 14364 42476 14420 42532
rect 14700 42476 14756 42532
rect 14700 42252 14756 42308
rect 14028 40796 14084 40852
rect 14252 40348 14308 40404
rect 14252 39618 14308 39620
rect 14252 39566 14254 39618
rect 14254 39566 14306 39618
rect 14306 39566 14308 39618
rect 14252 39564 14308 39566
rect 15260 42588 15316 42644
rect 15036 42530 15092 42532
rect 15036 42478 15038 42530
rect 15038 42478 15090 42530
rect 15090 42478 15092 42530
rect 15036 42476 15092 42478
rect 14924 41580 14980 41636
rect 14924 41356 14980 41412
rect 15596 43596 15652 43652
rect 18172 45666 18228 45668
rect 18172 45614 18174 45666
rect 18174 45614 18226 45666
rect 18226 45614 18228 45666
rect 18172 45612 18228 45614
rect 17612 45388 17668 45444
rect 17164 45052 17220 45108
rect 15708 43538 15764 43540
rect 15708 43486 15710 43538
rect 15710 43486 15762 43538
rect 15762 43486 15764 43538
rect 15708 43484 15764 43486
rect 15596 42194 15652 42196
rect 15596 42142 15598 42194
rect 15598 42142 15650 42194
rect 15650 42142 15652 42194
rect 15596 42140 15652 42142
rect 15036 41298 15092 41300
rect 15036 41246 15038 41298
rect 15038 41246 15090 41298
rect 15090 41246 15092 41298
rect 15036 41244 15092 41246
rect 15260 41692 15316 41748
rect 15260 41244 15316 41300
rect 15372 41580 15428 41636
rect 14588 39394 14644 39396
rect 14588 39342 14590 39394
rect 14590 39342 14642 39394
rect 14642 39342 14644 39394
rect 14588 39340 14644 39342
rect 14700 39116 14756 39172
rect 14476 39004 14532 39060
rect 15260 39394 15316 39396
rect 15260 39342 15262 39394
rect 15262 39342 15314 39394
rect 15314 39342 15316 39394
rect 15260 39340 15316 39342
rect 14924 39004 14980 39060
rect 13804 37996 13860 38052
rect 13916 38108 13972 38164
rect 13244 37436 13300 37492
rect 13580 37266 13636 37268
rect 13580 37214 13582 37266
rect 13582 37214 13634 37266
rect 13634 37214 13636 37266
rect 13580 37212 13636 37214
rect 14364 37938 14420 37940
rect 14364 37886 14366 37938
rect 14366 37886 14418 37938
rect 14418 37886 14420 37938
rect 14364 37884 14420 37886
rect 13804 37826 13860 37828
rect 13804 37774 13806 37826
rect 13806 37774 13858 37826
rect 13858 37774 13860 37826
rect 13804 37772 13860 37774
rect 14028 37826 14084 37828
rect 14028 37774 14030 37826
rect 14030 37774 14082 37826
rect 14082 37774 14084 37826
rect 14028 37772 14084 37774
rect 14140 36652 14196 36708
rect 13692 36594 13748 36596
rect 13692 36542 13694 36594
rect 13694 36542 13746 36594
rect 13746 36542 13748 36594
rect 13692 36540 13748 36542
rect 13356 36316 13412 36372
rect 13804 36258 13860 36260
rect 13804 36206 13806 36258
rect 13806 36206 13858 36258
rect 13858 36206 13860 36258
rect 13804 36204 13860 36206
rect 13580 35980 13636 36036
rect 13244 35308 13300 35364
rect 13580 35196 13636 35252
rect 13580 34412 13636 34468
rect 13468 33740 13524 33796
rect 13132 33628 13188 33684
rect 12908 33234 12964 33236
rect 12908 33182 12910 33234
rect 12910 33182 12962 33234
rect 12962 33182 12964 33234
rect 12908 33180 12964 33182
rect 12796 32620 12852 32676
rect 12572 31612 12628 31668
rect 12796 31612 12852 31668
rect 13020 31500 13076 31556
rect 12460 30492 12516 30548
rect 12572 30434 12628 30436
rect 12572 30382 12574 30434
rect 12574 30382 12626 30434
rect 12626 30382 12628 30434
rect 12572 30380 12628 30382
rect 12908 30322 12964 30324
rect 12908 30270 12910 30322
rect 12910 30270 12962 30322
rect 12962 30270 12964 30322
rect 12908 30268 12964 30270
rect 12572 29820 12628 29876
rect 12684 28924 12740 28980
rect 12796 29986 12852 29988
rect 12796 29934 12798 29986
rect 12798 29934 12850 29986
rect 12850 29934 12852 29986
rect 12796 29932 12852 29934
rect 13020 29538 13076 29540
rect 13020 29486 13022 29538
rect 13022 29486 13074 29538
rect 13074 29486 13076 29538
rect 13020 29484 13076 29486
rect 12908 28700 12964 28756
rect 12684 28028 12740 28084
rect 12460 27858 12516 27860
rect 12460 27806 12462 27858
rect 12462 27806 12514 27858
rect 12514 27806 12516 27858
rect 12460 27804 12516 27806
rect 12572 27468 12628 27524
rect 12236 27298 12292 27300
rect 12236 27246 12238 27298
rect 12238 27246 12290 27298
rect 12290 27246 12292 27298
rect 12236 27244 12292 27246
rect 12124 26796 12180 26852
rect 11676 26348 11732 26404
rect 11116 25116 11172 25172
rect 11340 26124 11396 26180
rect 11340 25340 11396 25396
rect 11452 25116 11508 25172
rect 11228 24668 11284 24724
rect 11564 24668 11620 24724
rect 11676 25004 11732 25060
rect 11340 24444 11396 24500
rect 11340 24220 11396 24276
rect 11900 26124 11956 26180
rect 11900 24780 11956 24836
rect 12012 24668 12068 24724
rect 11788 23996 11844 24052
rect 11900 23884 11956 23940
rect 11340 22652 11396 22708
rect 11676 23714 11732 23716
rect 11676 23662 11678 23714
rect 11678 23662 11730 23714
rect 11730 23662 11732 23714
rect 11676 23660 11732 23662
rect 11564 23436 11620 23492
rect 11788 23324 11844 23380
rect 11452 21644 11508 21700
rect 11228 21420 11284 21476
rect 10108 19906 10164 19908
rect 10108 19854 10110 19906
rect 10110 19854 10162 19906
rect 10162 19854 10164 19906
rect 10108 19852 10164 19854
rect 10220 19740 10276 19796
rect 10220 19068 10276 19124
rect 10556 20076 10612 20132
rect 10332 18284 10388 18340
rect 10444 19068 10500 19124
rect 9772 16716 9828 16772
rect 9548 15426 9604 15428
rect 9548 15374 9550 15426
rect 9550 15374 9602 15426
rect 9602 15374 9604 15426
rect 9548 15372 9604 15374
rect 8652 14476 8708 14532
rect 8876 12684 8932 12740
rect 8540 12124 8596 12180
rect 8876 12460 8932 12516
rect 5964 11282 6020 11284
rect 5964 11230 5966 11282
rect 5966 11230 6018 11282
rect 6018 11230 6020 11282
rect 5964 11228 6020 11230
rect 7756 11676 7812 11732
rect 8316 11452 8372 11508
rect 6188 9996 6244 10052
rect 6524 11228 6580 11284
rect 5404 9884 5460 9940
rect 6076 9884 6132 9940
rect 4956 9266 5012 9268
rect 4956 9214 4958 9266
rect 4958 9214 5010 9266
rect 5010 9214 5012 9266
rect 4956 9212 5012 9214
rect 4620 9154 4676 9156
rect 4620 9102 4622 9154
rect 4622 9102 4674 9154
rect 4674 9102 4676 9154
rect 4620 9100 4676 9102
rect 4956 9042 5012 9044
rect 4956 8990 4958 9042
rect 4958 8990 5010 9042
rect 5010 8990 5012 9042
rect 4956 8988 5012 8990
rect 4396 8764 4452 8820
rect 5180 9100 5236 9156
rect 5516 9548 5572 9604
rect 5740 9154 5796 9156
rect 5740 9102 5742 9154
rect 5742 9102 5794 9154
rect 5794 9102 5796 9154
rect 5740 9100 5796 9102
rect 6636 11116 6692 11172
rect 7868 11170 7924 11172
rect 7868 11118 7870 11170
rect 7870 11118 7922 11170
rect 7922 11118 7924 11170
rect 7868 11116 7924 11118
rect 8204 11170 8260 11172
rect 8204 11118 8206 11170
rect 8206 11118 8258 11170
rect 8258 11118 8260 11170
rect 8204 11116 8260 11118
rect 8204 10834 8260 10836
rect 8204 10782 8206 10834
rect 8206 10782 8258 10834
rect 8258 10782 8260 10834
rect 8204 10780 8260 10782
rect 8764 11676 8820 11732
rect 8988 12236 9044 12292
rect 9212 13580 9268 13636
rect 9660 14476 9716 14532
rect 9660 14028 9716 14084
rect 9436 13468 9492 13524
rect 9884 15986 9940 15988
rect 9884 15934 9886 15986
rect 9886 15934 9938 15986
rect 9938 15934 9940 15986
rect 9884 15932 9940 15934
rect 9884 15484 9940 15540
rect 9996 14642 10052 14644
rect 9996 14590 9998 14642
rect 9998 14590 10050 14642
rect 10050 14590 10052 14642
rect 9996 14588 10052 14590
rect 9884 13804 9940 13860
rect 10332 15932 10388 15988
rect 10332 15148 10388 15204
rect 10892 20578 10948 20580
rect 10892 20526 10894 20578
rect 10894 20526 10946 20578
rect 10946 20526 10948 20578
rect 10892 20524 10948 20526
rect 10892 20300 10948 20356
rect 11340 20914 11396 20916
rect 11340 20862 11342 20914
rect 11342 20862 11394 20914
rect 11394 20862 11396 20914
rect 11340 20860 11396 20862
rect 11564 20802 11620 20804
rect 11564 20750 11566 20802
rect 11566 20750 11618 20802
rect 11618 20750 11620 20802
rect 11564 20748 11620 20750
rect 11116 20076 11172 20132
rect 11004 19740 11060 19796
rect 11564 19964 11620 20020
rect 10668 19180 10724 19236
rect 10556 18620 10612 18676
rect 10780 18060 10836 18116
rect 10892 18172 10948 18228
rect 10668 16828 10724 16884
rect 10556 16156 10612 16212
rect 10780 16716 10836 16772
rect 10780 14642 10836 14644
rect 10780 14590 10782 14642
rect 10782 14590 10834 14642
rect 10834 14590 10836 14642
rect 10780 14588 10836 14590
rect 10220 14028 10276 14084
rect 10444 13916 10500 13972
rect 10668 14530 10724 14532
rect 10668 14478 10670 14530
rect 10670 14478 10722 14530
rect 10722 14478 10724 14530
rect 10668 14476 10724 14478
rect 10444 13580 10500 13636
rect 10220 13468 10276 13524
rect 11116 19068 11172 19124
rect 11564 18338 11620 18340
rect 11564 18286 11566 18338
rect 11566 18286 11618 18338
rect 11618 18286 11620 18338
rect 11564 18284 11620 18286
rect 11788 21474 11844 21476
rect 11788 21422 11790 21474
rect 11790 21422 11842 21474
rect 11842 21422 11844 21474
rect 11788 21420 11844 21422
rect 11788 20524 11844 20580
rect 11900 18450 11956 18452
rect 11900 18398 11902 18450
rect 11902 18398 11954 18450
rect 11954 18398 11956 18450
rect 11900 18396 11956 18398
rect 11788 18060 11844 18116
rect 11116 17724 11172 17780
rect 11452 17724 11508 17780
rect 11340 17164 11396 17220
rect 11004 16044 11060 16100
rect 11004 15538 11060 15540
rect 11004 15486 11006 15538
rect 11006 15486 11058 15538
rect 11058 15486 11060 15538
rect 11004 15484 11060 15486
rect 11340 15372 11396 15428
rect 11116 15260 11172 15316
rect 9324 11564 9380 11620
rect 8988 10780 9044 10836
rect 6972 9996 7028 10052
rect 8876 10444 8932 10500
rect 9996 12460 10052 12516
rect 11900 17276 11956 17332
rect 12348 26908 12404 26964
rect 12460 26348 12516 26404
rect 12684 25452 12740 25508
rect 12460 25394 12516 25396
rect 12460 25342 12462 25394
rect 12462 25342 12514 25394
rect 12514 25342 12516 25394
rect 12460 25340 12516 25342
rect 12236 23772 12292 23828
rect 12348 24444 12404 24500
rect 13020 28588 13076 28644
rect 12908 27580 12964 27636
rect 14252 35026 14308 35028
rect 14252 34974 14254 35026
rect 14254 34974 14306 35026
rect 14306 34974 14308 35026
rect 14252 34972 14308 34974
rect 14028 34914 14084 34916
rect 14028 34862 14030 34914
rect 14030 34862 14082 34914
rect 14082 34862 14084 34914
rect 14028 34860 14084 34862
rect 15148 39228 15204 39284
rect 15036 37548 15092 37604
rect 15260 39116 15316 39172
rect 15820 41468 15876 41524
rect 15708 41356 15764 41412
rect 15932 41074 15988 41076
rect 15932 41022 15934 41074
rect 15934 41022 15986 41074
rect 15986 41022 15988 41074
rect 15932 41020 15988 41022
rect 15596 40908 15652 40964
rect 15484 40572 15540 40628
rect 16268 43260 16324 43316
rect 16044 40684 16100 40740
rect 16156 41858 16212 41860
rect 16156 41806 16158 41858
rect 16158 41806 16210 41858
rect 16210 41806 16212 41858
rect 16156 41804 16212 41806
rect 17052 44098 17108 44100
rect 17052 44046 17054 44098
rect 17054 44046 17106 44098
rect 17106 44046 17108 44098
rect 17052 44044 17108 44046
rect 16492 41804 16548 41860
rect 16604 42140 16660 42196
rect 16268 41580 16324 41636
rect 16156 40572 16212 40628
rect 16604 41356 16660 41412
rect 16268 41244 16324 41300
rect 16268 40460 16324 40516
rect 16044 40290 16100 40292
rect 16044 40238 16046 40290
rect 16046 40238 16098 40290
rect 16098 40238 16100 40290
rect 16044 40236 16100 40238
rect 16268 40178 16324 40180
rect 16268 40126 16270 40178
rect 16270 40126 16322 40178
rect 16322 40126 16324 40178
rect 16268 40124 16324 40126
rect 16716 40402 16772 40404
rect 16716 40350 16718 40402
rect 16718 40350 16770 40402
rect 16770 40350 16772 40402
rect 16716 40348 16772 40350
rect 16044 39676 16100 39732
rect 15596 39340 15652 39396
rect 15820 39618 15876 39620
rect 15820 39566 15822 39618
rect 15822 39566 15874 39618
rect 15874 39566 15876 39618
rect 15820 39564 15876 39566
rect 15820 39116 15876 39172
rect 15708 39004 15764 39060
rect 15484 38668 15540 38724
rect 15372 38556 15428 38612
rect 15148 37436 15204 37492
rect 15372 37996 15428 38052
rect 14812 37324 14868 37380
rect 14588 36594 14644 36596
rect 14588 36542 14590 36594
rect 14590 36542 14642 36594
rect 14642 36542 14644 36594
rect 14588 36540 14644 36542
rect 14588 36204 14644 36260
rect 14924 36370 14980 36372
rect 14924 36318 14926 36370
rect 14926 36318 14978 36370
rect 14978 36318 14980 36370
rect 14924 36316 14980 36318
rect 14700 35868 14756 35924
rect 14588 35420 14644 35476
rect 15036 36204 15092 36260
rect 14924 35026 14980 35028
rect 14924 34974 14926 35026
rect 14926 34974 14978 35026
rect 14978 34974 14980 35026
rect 14924 34972 14980 34974
rect 14476 34860 14532 34916
rect 15036 34860 15092 34916
rect 15260 34972 15316 35028
rect 13804 33516 13860 33572
rect 14140 34748 14196 34804
rect 13244 33180 13300 33236
rect 14588 34636 14644 34692
rect 14364 34412 14420 34468
rect 13804 32956 13860 33012
rect 13580 31948 13636 32004
rect 13916 32284 13972 32340
rect 13244 31276 13300 31332
rect 13356 30940 13412 30996
rect 14028 31164 14084 31220
rect 13692 30770 13748 30772
rect 13692 30718 13694 30770
rect 13694 30718 13746 30770
rect 13746 30718 13748 30770
rect 13692 30716 13748 30718
rect 13916 29932 13972 29988
rect 13804 29820 13860 29876
rect 13804 29260 13860 29316
rect 13468 28700 13524 28756
rect 13244 27468 13300 27524
rect 13356 28364 13412 28420
rect 12684 25228 12740 25284
rect 12460 23884 12516 23940
rect 12572 23378 12628 23380
rect 12572 23326 12574 23378
rect 12574 23326 12626 23378
rect 12626 23326 12628 23378
rect 12572 23324 12628 23326
rect 12124 21980 12180 22036
rect 12124 21644 12180 21700
rect 12236 21586 12292 21588
rect 12236 21534 12238 21586
rect 12238 21534 12290 21586
rect 12290 21534 12292 21586
rect 12236 21532 12292 21534
rect 13356 27132 13412 27188
rect 12796 22652 12852 22708
rect 13692 28754 13748 28756
rect 13692 28702 13694 28754
rect 13694 28702 13746 28754
rect 13746 28702 13748 28754
rect 13692 28700 13748 28702
rect 14028 28588 14084 28644
rect 14588 34076 14644 34132
rect 15260 33852 15316 33908
rect 14700 32284 14756 32340
rect 14476 30828 14532 30884
rect 16044 39340 16100 39396
rect 15932 38668 15988 38724
rect 15932 37996 15988 38052
rect 15708 37548 15764 37604
rect 15820 37490 15876 37492
rect 15820 37438 15822 37490
rect 15822 37438 15874 37490
rect 15874 37438 15876 37490
rect 15820 37436 15876 37438
rect 16044 37772 16100 37828
rect 16492 39004 16548 39060
rect 16380 38668 16436 38724
rect 16268 38050 16324 38052
rect 16268 37998 16270 38050
rect 16270 37998 16322 38050
rect 16322 37998 16324 38050
rect 16268 37996 16324 37998
rect 15932 36652 15988 36708
rect 17948 42588 18004 42644
rect 17500 42028 17556 42084
rect 17388 41916 17444 41972
rect 18060 41804 18116 41860
rect 17388 41020 17444 41076
rect 17276 40684 17332 40740
rect 17164 39452 17220 39508
rect 16828 38722 16884 38724
rect 16828 38670 16830 38722
rect 16830 38670 16882 38722
rect 16882 38670 16884 38722
rect 16828 38668 16884 38670
rect 16380 37212 16436 37268
rect 16604 37266 16660 37268
rect 16604 37214 16606 37266
rect 16606 37214 16658 37266
rect 16658 37214 16660 37266
rect 16604 37212 16660 37214
rect 16604 36370 16660 36372
rect 16604 36318 16606 36370
rect 16606 36318 16658 36370
rect 16658 36318 16660 36370
rect 16604 36316 16660 36318
rect 16268 36092 16324 36148
rect 16044 35810 16100 35812
rect 16044 35758 16046 35810
rect 16046 35758 16098 35810
rect 16098 35758 16100 35810
rect 16044 35756 16100 35758
rect 15484 34860 15540 34916
rect 15708 35420 15764 35476
rect 15596 34412 15652 34468
rect 15596 34242 15652 34244
rect 15596 34190 15598 34242
rect 15598 34190 15650 34242
rect 15650 34190 15652 34242
rect 15596 34188 15652 34190
rect 15708 33740 15764 33796
rect 15596 33234 15652 33236
rect 15596 33182 15598 33234
rect 15598 33182 15650 33234
rect 15650 33182 15652 33234
rect 15596 33180 15652 33182
rect 15820 33180 15876 33236
rect 15372 32732 15428 32788
rect 15708 32786 15764 32788
rect 15708 32734 15710 32786
rect 15710 32734 15762 32786
rect 15762 32734 15764 32786
rect 15708 32732 15764 32734
rect 15036 32620 15092 32676
rect 16828 36540 16884 36596
rect 16156 35532 16212 35588
rect 16380 35420 16436 35476
rect 16268 35308 16324 35364
rect 16380 34690 16436 34692
rect 16380 34638 16382 34690
rect 16382 34638 16434 34690
rect 16434 34638 16436 34690
rect 16380 34636 16436 34638
rect 16044 32956 16100 33012
rect 16268 34300 16324 34356
rect 15932 32620 15988 32676
rect 15484 32562 15540 32564
rect 15484 32510 15486 32562
rect 15486 32510 15538 32562
rect 15538 32510 15540 32562
rect 15484 32508 15540 32510
rect 16268 32732 16324 32788
rect 15148 32450 15204 32452
rect 15148 32398 15150 32450
rect 15150 32398 15202 32450
rect 15202 32398 15204 32450
rect 15148 32396 15204 32398
rect 15036 32060 15092 32116
rect 16156 32060 16212 32116
rect 14252 30380 14308 30436
rect 14476 30268 14532 30324
rect 14588 30156 14644 30212
rect 15036 30492 15092 30548
rect 15036 30268 15092 30324
rect 14588 29820 14644 29876
rect 15484 31612 15540 31668
rect 16156 31500 16212 31556
rect 15372 30716 15428 30772
rect 15260 30268 15316 30324
rect 15372 29986 15428 29988
rect 15372 29934 15374 29986
rect 15374 29934 15426 29986
rect 15426 29934 15428 29986
rect 15372 29932 15428 29934
rect 15372 29484 15428 29540
rect 14252 28700 14308 28756
rect 15260 28476 15316 28532
rect 13916 28252 13972 28308
rect 14252 27692 14308 27748
rect 13804 26684 13860 26740
rect 13916 26908 13972 26964
rect 13692 26178 13748 26180
rect 13692 26126 13694 26178
rect 13694 26126 13746 26178
rect 13746 26126 13748 26178
rect 13692 26124 13748 26126
rect 13468 25900 13524 25956
rect 13580 25618 13636 25620
rect 13580 25566 13582 25618
rect 13582 25566 13634 25618
rect 13634 25566 13636 25618
rect 13580 25564 13636 25566
rect 13356 25452 13412 25508
rect 13020 24722 13076 24724
rect 13020 24670 13022 24722
rect 13022 24670 13074 24722
rect 13074 24670 13076 24722
rect 13020 24668 13076 24670
rect 13244 23154 13300 23156
rect 13244 23102 13246 23154
rect 13246 23102 13298 23154
rect 13298 23102 13300 23154
rect 13244 23100 13300 23102
rect 12908 22146 12964 22148
rect 12908 22094 12910 22146
rect 12910 22094 12962 22146
rect 12962 22094 12964 22146
rect 12908 22092 12964 22094
rect 12908 21698 12964 21700
rect 12908 21646 12910 21698
rect 12910 21646 12962 21698
rect 12962 21646 12964 21698
rect 12908 21644 12964 21646
rect 12684 20524 12740 20580
rect 12124 20300 12180 20356
rect 12236 20412 12292 20468
rect 12236 19234 12292 19236
rect 12236 19182 12238 19234
rect 12238 19182 12290 19234
rect 12290 19182 12292 19234
rect 12236 19180 12292 19182
rect 12124 18956 12180 19012
rect 12236 18226 12292 18228
rect 12236 18174 12238 18226
rect 12238 18174 12290 18226
rect 12290 18174 12292 18226
rect 12236 18172 12292 18174
rect 12236 16940 12292 16996
rect 12124 16882 12180 16884
rect 12124 16830 12126 16882
rect 12126 16830 12178 16882
rect 12178 16830 12180 16882
rect 12124 16828 12180 16830
rect 12012 15986 12068 15988
rect 12012 15934 12014 15986
rect 12014 15934 12066 15986
rect 12066 15934 12068 15986
rect 12012 15932 12068 15934
rect 11900 15484 11956 15540
rect 11788 15314 11844 15316
rect 11788 15262 11790 15314
rect 11790 15262 11842 15314
rect 11842 15262 11844 15314
rect 11788 15260 11844 15262
rect 11564 14588 11620 14644
rect 12012 14642 12068 14644
rect 12012 14590 12014 14642
rect 12014 14590 12066 14642
rect 12066 14590 12068 14642
rect 12012 14588 12068 14590
rect 11340 13692 11396 13748
rect 10444 13074 10500 13076
rect 10444 13022 10446 13074
rect 10446 13022 10498 13074
rect 10498 13022 10500 13074
rect 10444 13020 10500 13022
rect 10444 12348 10500 12404
rect 9884 11676 9940 11732
rect 9996 12236 10052 12292
rect 11116 12402 11172 12404
rect 11116 12350 11118 12402
rect 11118 12350 11170 12402
rect 11170 12350 11172 12402
rect 11116 12348 11172 12350
rect 11228 12290 11284 12292
rect 11228 12238 11230 12290
rect 11230 12238 11282 12290
rect 11282 12238 11284 12290
rect 11228 12236 11284 12238
rect 10108 12012 10164 12068
rect 9660 11116 9716 11172
rect 9884 11340 9940 11396
rect 10668 11452 10724 11508
rect 10220 11394 10276 11396
rect 10220 11342 10222 11394
rect 10222 11342 10274 11394
rect 10274 11342 10276 11394
rect 10220 11340 10276 11342
rect 9772 10556 9828 10612
rect 6524 9602 6580 9604
rect 6524 9550 6526 9602
rect 6526 9550 6578 9602
rect 6578 9550 6580 9602
rect 6524 9548 6580 9550
rect 7084 9602 7140 9604
rect 7084 9550 7086 9602
rect 7086 9550 7138 9602
rect 7138 9550 7140 9602
rect 7084 9548 7140 9550
rect 7756 9548 7812 9604
rect 4476 8650 4532 8652
rect 4476 8598 4478 8650
rect 4478 8598 4530 8650
rect 4530 8598 4532 8650
rect 4476 8596 4532 8598
rect 4580 8650 4636 8652
rect 4580 8598 4582 8650
rect 4582 8598 4634 8650
rect 4634 8598 4636 8650
rect 4580 8596 4636 8598
rect 4684 8650 4740 8652
rect 4684 8598 4686 8650
rect 4686 8598 4738 8650
rect 4738 8598 4740 8650
rect 4684 8596 4740 8598
rect 5180 8540 5236 8596
rect 1708 5404 1764 5460
rect 9996 9826 10052 9828
rect 9996 9774 9998 9826
rect 9998 9774 10050 9826
rect 10050 9774 10052 9826
rect 9996 9772 10052 9774
rect 7980 8988 8036 9044
rect 8988 9548 9044 9604
rect 9996 8930 10052 8932
rect 9996 8878 9998 8930
rect 9998 8878 10050 8930
rect 10050 8878 10052 8930
rect 9996 8876 10052 8878
rect 8988 8652 9044 8708
rect 5852 8316 5908 8372
rect 7084 8316 7140 8372
rect 5516 8092 5572 8148
rect 6636 8092 6692 8148
rect 9436 8258 9492 8260
rect 9436 8206 9438 8258
rect 9438 8206 9490 8258
rect 9490 8206 9492 8258
rect 9436 8204 9492 8206
rect 8988 7980 9044 8036
rect 4476 7082 4532 7084
rect 4476 7030 4478 7082
rect 4478 7030 4530 7082
rect 4530 7030 4532 7082
rect 4476 7028 4532 7030
rect 4580 7082 4636 7084
rect 4580 7030 4582 7082
rect 4582 7030 4634 7082
rect 4634 7030 4636 7082
rect 4580 7028 4636 7030
rect 4684 7082 4740 7084
rect 4684 7030 4686 7082
rect 4686 7030 4738 7082
rect 4738 7030 4740 7082
rect 5292 7084 5348 7140
rect 6524 7084 6580 7140
rect 4684 7028 4740 7030
rect 6524 6188 6580 6244
rect 6300 6130 6356 6132
rect 6300 6078 6302 6130
rect 6302 6078 6354 6130
rect 6354 6078 6356 6130
rect 6300 6076 6356 6078
rect 4476 5514 4532 5516
rect 4476 5462 4478 5514
rect 4478 5462 4530 5514
rect 4530 5462 4532 5514
rect 4476 5460 4532 5462
rect 4580 5514 4636 5516
rect 4580 5462 4582 5514
rect 4582 5462 4634 5514
rect 4634 5462 4636 5514
rect 4580 5460 4636 5462
rect 4684 5514 4740 5516
rect 4684 5462 4686 5514
rect 4686 5462 4738 5514
rect 4738 5462 4740 5514
rect 4684 5460 4740 5462
rect 4060 4956 4116 5012
rect 1708 4898 1764 4900
rect 1708 4846 1710 4898
rect 1710 4846 1762 4898
rect 1762 4846 1764 4898
rect 1708 4844 1764 4846
rect 5068 5010 5124 5012
rect 5068 4958 5070 5010
rect 5070 4958 5122 5010
rect 5122 4958 5124 5010
rect 5068 4956 5124 4958
rect 1708 4060 1764 4116
rect 7420 6130 7476 6132
rect 7420 6078 7422 6130
rect 7422 6078 7474 6130
rect 7474 6078 7476 6130
rect 7420 6076 7476 6078
rect 8092 6524 8148 6580
rect 7644 6188 7700 6244
rect 7084 5906 7140 5908
rect 7084 5854 7086 5906
rect 7086 5854 7138 5906
rect 7138 5854 7140 5906
rect 7084 5852 7140 5854
rect 6748 5740 6804 5796
rect 6748 5292 6804 5348
rect 6748 5068 6804 5124
rect 6300 4898 6356 4900
rect 6300 4846 6302 4898
rect 6302 4846 6354 4898
rect 6354 4846 6356 4898
rect 6300 4844 6356 4846
rect 6524 4396 6580 4452
rect 5516 4060 5572 4116
rect 5852 4284 5908 4340
rect 4476 3946 4532 3948
rect 4476 3894 4478 3946
rect 4478 3894 4530 3946
rect 4530 3894 4532 3946
rect 4476 3892 4532 3894
rect 4580 3946 4636 3948
rect 4580 3894 4582 3946
rect 4582 3894 4634 3946
rect 4634 3894 4636 3946
rect 4580 3892 4636 3894
rect 4684 3946 4740 3948
rect 4684 3894 4686 3946
rect 4686 3894 4738 3946
rect 4738 3894 4740 3946
rect 4684 3892 4740 3894
rect 5068 3836 5124 3892
rect 4620 3666 4676 3668
rect 4620 3614 4622 3666
rect 4622 3614 4674 3666
rect 4674 3614 4676 3666
rect 4620 3612 4676 3614
rect 6188 4172 6244 4228
rect 6748 4060 6804 4116
rect 7420 5740 7476 5796
rect 7756 5292 7812 5348
rect 7532 4562 7588 4564
rect 7532 4510 7534 4562
rect 7534 4510 7586 4562
rect 7586 4510 7588 4562
rect 7532 4508 7588 4510
rect 8652 6300 8708 6356
rect 8540 5906 8596 5908
rect 8540 5854 8542 5906
rect 8542 5854 8594 5906
rect 8594 5854 8596 5906
rect 8540 5852 8596 5854
rect 8764 5852 8820 5908
rect 8540 5180 8596 5236
rect 8204 5122 8260 5124
rect 8204 5070 8206 5122
rect 8206 5070 8258 5122
rect 8258 5070 8260 5122
rect 8204 5068 8260 5070
rect 8428 5068 8484 5124
rect 7084 4338 7140 4340
rect 7084 4286 7086 4338
rect 7086 4286 7138 4338
rect 7138 4286 7140 4338
rect 7084 4284 7140 4286
rect 7420 4338 7476 4340
rect 7420 4286 7422 4338
rect 7422 4286 7474 4338
rect 7474 4286 7476 4338
rect 7420 4284 7476 4286
rect 4172 3554 4228 3556
rect 4172 3502 4174 3554
rect 4174 3502 4226 3554
rect 4226 3502 4228 3554
rect 4172 3500 4228 3502
rect 1708 3388 1764 3444
rect 6076 3442 6132 3444
rect 6076 3390 6078 3442
rect 6078 3390 6130 3442
rect 6130 3390 6132 3442
rect 6076 3388 6132 3390
rect 2156 2716 2212 2772
rect 7420 3500 7476 3556
rect 6972 3442 7028 3444
rect 6972 3390 6974 3442
rect 6974 3390 7026 3442
rect 7026 3390 7028 3442
rect 6972 3388 7028 3390
rect 7980 3724 8036 3780
rect 8428 3612 8484 3668
rect 7868 3554 7924 3556
rect 7868 3502 7870 3554
rect 7870 3502 7922 3554
rect 7922 3502 7924 3554
rect 7868 3500 7924 3502
rect 9772 8034 9828 8036
rect 9772 7982 9774 8034
rect 9774 7982 9826 8034
rect 9826 7982 9828 8034
rect 9772 7980 9828 7982
rect 8988 7084 9044 7140
rect 9100 6972 9156 7028
rect 9772 6860 9828 6916
rect 8876 5740 8932 5796
rect 8876 4844 8932 4900
rect 9884 6748 9940 6804
rect 10556 10780 10612 10836
rect 12236 15260 12292 15316
rect 12908 19852 12964 19908
rect 13020 20076 13076 20132
rect 13132 22204 13188 22260
rect 12908 19180 12964 19236
rect 12796 18620 12852 18676
rect 13244 21868 13300 21924
rect 13692 24892 13748 24948
rect 14028 26460 14084 26516
rect 13580 23826 13636 23828
rect 13580 23774 13582 23826
rect 13582 23774 13634 23826
rect 13634 23774 13636 23826
rect 13580 23772 13636 23774
rect 13916 24444 13972 24500
rect 13916 24220 13972 24276
rect 13468 22258 13524 22260
rect 13468 22206 13470 22258
rect 13470 22206 13522 22258
rect 13522 22206 13524 22258
rect 13468 22204 13524 22206
rect 14476 28252 14532 28308
rect 15036 28082 15092 28084
rect 15036 28030 15038 28082
rect 15038 28030 15090 28082
rect 15090 28030 15092 28082
rect 15036 28028 15092 28030
rect 14812 27468 14868 27524
rect 15036 27356 15092 27412
rect 15260 27804 15316 27860
rect 14924 27244 14980 27300
rect 15708 30604 15764 30660
rect 16604 35756 16660 35812
rect 16828 35644 16884 35700
rect 16716 34524 16772 34580
rect 18060 40572 18116 40628
rect 17724 39564 17780 39620
rect 17612 39228 17668 39284
rect 17388 38668 17444 38724
rect 18284 42082 18340 42084
rect 18284 42030 18286 42082
rect 18286 42030 18338 42082
rect 18338 42030 18340 42082
rect 18284 42028 18340 42030
rect 19292 45388 19348 45444
rect 18732 44492 18788 44548
rect 19292 44940 19348 44996
rect 18620 43708 18676 43764
rect 19068 43820 19124 43876
rect 19292 43708 19348 43764
rect 18956 43538 19012 43540
rect 18956 43486 18958 43538
rect 18958 43486 19010 43538
rect 19010 43486 19012 43538
rect 18956 43484 19012 43486
rect 18620 42588 18676 42644
rect 19516 42588 19572 42644
rect 18508 41970 18564 41972
rect 18508 41918 18510 41970
rect 18510 41918 18562 41970
rect 18562 41918 18564 41970
rect 18508 41916 18564 41918
rect 19068 42476 19124 42532
rect 19180 42364 19236 42420
rect 18284 41074 18340 41076
rect 18284 41022 18286 41074
rect 18286 41022 18338 41074
rect 18338 41022 18340 41074
rect 18284 41020 18340 41022
rect 18284 40626 18340 40628
rect 18284 40574 18286 40626
rect 18286 40574 18338 40626
rect 18338 40574 18340 40626
rect 18284 40572 18340 40574
rect 18508 40348 18564 40404
rect 18620 40460 18676 40516
rect 18172 40124 18228 40180
rect 18060 38780 18116 38836
rect 18620 39004 18676 39060
rect 18844 40796 18900 40852
rect 19180 40402 19236 40404
rect 19180 40350 19182 40402
rect 19182 40350 19234 40402
rect 19234 40350 19236 40402
rect 19180 40348 19236 40350
rect 19292 40124 19348 40180
rect 20076 45612 20132 45668
rect 19836 45498 19892 45500
rect 19836 45446 19838 45498
rect 19838 45446 19890 45498
rect 19890 45446 19892 45498
rect 19836 45444 19892 45446
rect 19940 45498 19996 45500
rect 19940 45446 19942 45498
rect 19942 45446 19994 45498
rect 19994 45446 19996 45498
rect 19940 45444 19996 45446
rect 20044 45498 20100 45500
rect 20044 45446 20046 45498
rect 20046 45446 20098 45498
rect 20098 45446 20100 45498
rect 20044 45444 20100 45446
rect 22988 45276 23044 45332
rect 22876 45052 22932 45108
rect 20412 44994 20468 44996
rect 20412 44942 20414 44994
rect 20414 44942 20466 44994
rect 20466 44942 20468 44994
rect 20412 44940 20468 44942
rect 19836 43930 19892 43932
rect 19836 43878 19838 43930
rect 19838 43878 19890 43930
rect 19890 43878 19892 43930
rect 19836 43876 19892 43878
rect 19940 43930 19996 43932
rect 19940 43878 19942 43930
rect 19942 43878 19994 43930
rect 19994 43878 19996 43930
rect 19940 43876 19996 43878
rect 20044 43930 20100 43932
rect 20044 43878 20046 43930
rect 20046 43878 20098 43930
rect 20098 43878 20100 43930
rect 20044 43876 20100 43878
rect 19740 42700 19796 42756
rect 19964 42476 20020 42532
rect 19836 42362 19892 42364
rect 19836 42310 19838 42362
rect 19838 42310 19890 42362
rect 19890 42310 19892 42362
rect 19836 42308 19892 42310
rect 19940 42362 19996 42364
rect 19940 42310 19942 42362
rect 19942 42310 19994 42362
rect 19994 42310 19996 42362
rect 19940 42308 19996 42310
rect 20044 42362 20100 42364
rect 20044 42310 20046 42362
rect 20046 42310 20098 42362
rect 20098 42310 20100 42362
rect 20044 42308 20100 42310
rect 19852 42028 19908 42084
rect 19964 41916 20020 41972
rect 20412 43708 20468 43764
rect 23100 45164 23156 45220
rect 22652 44940 22708 44996
rect 21980 44380 22036 44436
rect 21868 44322 21924 44324
rect 21868 44270 21870 44322
rect 21870 44270 21922 44322
rect 21922 44270 21924 44322
rect 21868 44268 21924 44270
rect 21084 43426 21140 43428
rect 21084 43374 21086 43426
rect 21086 43374 21138 43426
rect 21138 43374 21140 43426
rect 21084 43372 21140 43374
rect 20636 42588 20692 42644
rect 20412 42140 20468 42196
rect 23660 44994 23716 44996
rect 23660 44942 23662 44994
rect 23662 44942 23714 44994
rect 23714 44942 23716 44994
rect 23660 44940 23716 44942
rect 22092 43372 22148 43428
rect 22428 43484 22484 43540
rect 21980 41916 22036 41972
rect 20860 41692 20916 41748
rect 20636 40908 20692 40964
rect 19836 40794 19892 40796
rect 19836 40742 19838 40794
rect 19838 40742 19890 40794
rect 19890 40742 19892 40794
rect 19836 40740 19892 40742
rect 19940 40794 19996 40796
rect 19940 40742 19942 40794
rect 19942 40742 19994 40794
rect 19994 40742 19996 40794
rect 19940 40740 19996 40742
rect 20044 40794 20100 40796
rect 20044 40742 20046 40794
rect 20046 40742 20098 40794
rect 20098 40742 20100 40794
rect 20044 40740 20100 40742
rect 18844 39506 18900 39508
rect 18844 39454 18846 39506
rect 18846 39454 18898 39506
rect 18898 39454 18900 39506
rect 18844 39452 18900 39454
rect 19068 39506 19124 39508
rect 19068 39454 19070 39506
rect 19070 39454 19122 39506
rect 19122 39454 19124 39506
rect 19068 39452 19124 39454
rect 17164 37996 17220 38052
rect 17500 37938 17556 37940
rect 17500 37886 17502 37938
rect 17502 37886 17554 37938
rect 17554 37886 17556 37938
rect 17500 37884 17556 37886
rect 18508 38220 18564 38276
rect 18060 37938 18116 37940
rect 18060 37886 18062 37938
rect 18062 37886 18114 37938
rect 18114 37886 18116 37938
rect 18060 37884 18116 37886
rect 17724 37826 17780 37828
rect 17724 37774 17726 37826
rect 17726 37774 17778 37826
rect 17778 37774 17780 37826
rect 17724 37772 17780 37774
rect 17276 37436 17332 37492
rect 17052 36370 17108 36372
rect 17052 36318 17054 36370
rect 17054 36318 17106 36370
rect 17106 36318 17108 36370
rect 17052 36316 17108 36318
rect 17164 36258 17220 36260
rect 17164 36206 17166 36258
rect 17166 36206 17218 36258
rect 17218 36206 17220 36258
rect 17164 36204 17220 36206
rect 17388 37266 17444 37268
rect 17388 37214 17390 37266
rect 17390 37214 17442 37266
rect 17442 37214 17444 37266
rect 17388 37212 17444 37214
rect 16940 34300 16996 34356
rect 17724 37378 17780 37380
rect 17724 37326 17726 37378
rect 17726 37326 17778 37378
rect 17778 37326 17780 37378
rect 17724 37324 17780 37326
rect 18284 36540 18340 36596
rect 18732 38444 18788 38500
rect 18508 37938 18564 37940
rect 18508 37886 18510 37938
rect 18510 37886 18562 37938
rect 18562 37886 18564 37938
rect 18508 37884 18564 37886
rect 18732 37548 18788 37604
rect 18732 37100 18788 37156
rect 17612 35980 17668 36036
rect 16828 33180 16884 33236
rect 16828 32732 16884 32788
rect 16268 30210 16324 30212
rect 16268 30158 16270 30210
rect 16270 30158 16322 30210
rect 16322 30158 16324 30210
rect 16268 30156 16324 30158
rect 16604 30156 16660 30212
rect 16492 29708 16548 29764
rect 16380 29596 16436 29652
rect 16044 29538 16100 29540
rect 16044 29486 16046 29538
rect 16046 29486 16098 29538
rect 16098 29486 16100 29538
rect 16044 29484 16100 29486
rect 15596 28812 15652 28868
rect 16268 29260 16324 29316
rect 16044 28476 16100 28532
rect 15820 28028 15876 28084
rect 16044 27746 16100 27748
rect 16044 27694 16046 27746
rect 16046 27694 16098 27746
rect 16098 27694 16100 27746
rect 16044 27692 16100 27694
rect 15708 27132 15764 27188
rect 15372 27074 15428 27076
rect 15372 27022 15374 27074
rect 15374 27022 15426 27074
rect 15426 27022 15428 27074
rect 15372 27020 15428 27022
rect 15820 27074 15876 27076
rect 15820 27022 15822 27074
rect 15822 27022 15874 27074
rect 15874 27022 15876 27074
rect 15820 27020 15876 27022
rect 14476 25228 14532 25284
rect 14588 26684 14644 26740
rect 14252 23548 14308 23604
rect 14028 22988 14084 23044
rect 14140 22652 14196 22708
rect 14028 22370 14084 22372
rect 14028 22318 14030 22370
rect 14030 22318 14082 22370
rect 14082 22318 14084 22370
rect 14028 22316 14084 22318
rect 13692 22092 13748 22148
rect 13804 21644 13860 21700
rect 13580 21196 13636 21252
rect 13916 20802 13972 20804
rect 13916 20750 13918 20802
rect 13918 20750 13970 20802
rect 13970 20750 13972 20802
rect 13916 20748 13972 20750
rect 13580 20076 13636 20132
rect 14140 20524 14196 20580
rect 14476 23660 14532 23716
rect 14476 22764 14532 22820
rect 14812 26684 14868 26740
rect 15708 26684 15764 26740
rect 15372 26572 15428 26628
rect 15260 25564 15316 25620
rect 15596 26124 15652 26180
rect 16156 27634 16212 27636
rect 16156 27582 16158 27634
rect 16158 27582 16210 27634
rect 16210 27582 16212 27634
rect 16156 27580 16212 27582
rect 16940 32620 16996 32676
rect 16604 29260 16660 29316
rect 16716 29202 16772 29204
rect 16716 29150 16718 29202
rect 16718 29150 16770 29202
rect 16770 29150 16772 29202
rect 16716 29148 16772 29150
rect 18284 35980 18340 36036
rect 17724 35810 17780 35812
rect 17724 35758 17726 35810
rect 17726 35758 17778 35810
rect 17778 35758 17780 35810
rect 17724 35756 17780 35758
rect 18060 35756 18116 35812
rect 17836 35644 17892 35700
rect 17724 35026 17780 35028
rect 17724 34974 17726 35026
rect 17726 34974 17778 35026
rect 17778 34974 17780 35026
rect 17724 34972 17780 34974
rect 17612 34860 17668 34916
rect 17388 34018 17444 34020
rect 17388 33966 17390 34018
rect 17390 33966 17442 34018
rect 17442 33966 17444 34018
rect 17388 33964 17444 33966
rect 17388 33628 17444 33684
rect 17500 33740 17556 33796
rect 17164 32396 17220 32452
rect 17388 32338 17444 32340
rect 17388 32286 17390 32338
rect 17390 32286 17442 32338
rect 17442 32286 17444 32338
rect 17388 32284 17444 32286
rect 17500 32060 17556 32116
rect 17164 30210 17220 30212
rect 17164 30158 17166 30210
rect 17166 30158 17218 30210
rect 17218 30158 17220 30210
rect 17164 30156 17220 30158
rect 16940 28812 16996 28868
rect 17052 29596 17108 29652
rect 17276 29484 17332 29540
rect 16492 28140 16548 28196
rect 17276 28028 17332 28084
rect 16828 27804 16884 27860
rect 16044 26908 16100 26964
rect 16716 27468 16772 27524
rect 16156 26290 16212 26292
rect 16156 26238 16158 26290
rect 16158 26238 16210 26290
rect 16210 26238 16212 26290
rect 16156 26236 16212 26238
rect 16492 26684 16548 26740
rect 16492 26460 16548 26516
rect 17164 26684 17220 26740
rect 16716 26236 16772 26292
rect 16380 25618 16436 25620
rect 16380 25566 16382 25618
rect 16382 25566 16434 25618
rect 16434 25566 16436 25618
rect 16380 25564 16436 25566
rect 15708 25452 15764 25508
rect 15708 24780 15764 24836
rect 14924 24220 14980 24276
rect 15372 24220 15428 24276
rect 15372 23772 15428 23828
rect 15820 25340 15876 25396
rect 15036 23212 15092 23268
rect 14924 23154 14980 23156
rect 14924 23102 14926 23154
rect 14926 23102 14978 23154
rect 14978 23102 14980 23154
rect 14924 23100 14980 23102
rect 15708 23772 15764 23828
rect 15148 22764 15204 22820
rect 14476 21868 14532 21924
rect 14812 21532 14868 21588
rect 14700 21420 14756 21476
rect 15372 22540 15428 22596
rect 15596 22092 15652 22148
rect 15484 21586 15540 21588
rect 15484 21534 15486 21586
rect 15486 21534 15538 21586
rect 15538 21534 15540 21586
rect 15484 21532 15540 21534
rect 14700 20636 14756 20692
rect 14588 20524 14644 20580
rect 13356 19794 13412 19796
rect 13356 19742 13358 19794
rect 13358 19742 13410 19794
rect 13410 19742 13412 19794
rect 13356 19740 13412 19742
rect 13916 20018 13972 20020
rect 13916 19966 13918 20018
rect 13918 19966 13970 20018
rect 13970 19966 13972 20018
rect 13916 19964 13972 19966
rect 14028 19852 14084 19908
rect 13692 19180 13748 19236
rect 13468 18956 13524 19012
rect 14252 19628 14308 19684
rect 14476 19404 14532 19460
rect 15484 20412 15540 20468
rect 15372 19906 15428 19908
rect 15372 19854 15374 19906
rect 15374 19854 15426 19906
rect 15426 19854 15428 19906
rect 15372 19852 15428 19854
rect 13244 18562 13300 18564
rect 13244 18510 13246 18562
rect 13246 18510 13298 18562
rect 13298 18510 13300 18562
rect 13244 18508 13300 18510
rect 12572 18450 12628 18452
rect 12572 18398 12574 18450
rect 12574 18398 12626 18450
rect 12626 18398 12628 18450
rect 12572 18396 12628 18398
rect 12572 17836 12628 17892
rect 12684 17948 12740 18004
rect 12572 16268 12628 16324
rect 12684 17276 12740 17332
rect 12796 16380 12852 16436
rect 12572 15874 12628 15876
rect 12572 15822 12574 15874
rect 12574 15822 12626 15874
rect 12626 15822 12628 15874
rect 12572 15820 12628 15822
rect 14924 19234 14980 19236
rect 14924 19182 14926 19234
rect 14926 19182 14978 19234
rect 14978 19182 14980 19234
rect 14924 19180 14980 19182
rect 13580 17948 13636 18004
rect 13468 16828 13524 16884
rect 13804 18172 13860 18228
rect 14028 17666 14084 17668
rect 14028 17614 14030 17666
rect 14030 17614 14082 17666
rect 14082 17614 14084 17666
rect 14028 17612 14084 17614
rect 14588 18396 14644 18452
rect 14812 18226 14868 18228
rect 14812 18174 14814 18226
rect 14814 18174 14866 18226
rect 14866 18174 14868 18226
rect 14812 18172 14868 18174
rect 14476 17276 14532 17332
rect 14588 17612 14644 17668
rect 14476 17106 14532 17108
rect 14476 17054 14478 17106
rect 14478 17054 14530 17106
rect 14530 17054 14532 17106
rect 14476 17052 14532 17054
rect 13804 16828 13860 16884
rect 14140 16604 14196 16660
rect 14476 16268 14532 16324
rect 12236 13804 12292 13860
rect 12012 13020 12068 13076
rect 11004 11618 11060 11620
rect 11004 11566 11006 11618
rect 11006 11566 11058 11618
rect 11058 11566 11060 11618
rect 11004 11564 11060 11566
rect 10780 10668 10836 10724
rect 10892 10610 10948 10612
rect 10892 10558 10894 10610
rect 10894 10558 10946 10610
rect 10946 10558 10948 10610
rect 10892 10556 10948 10558
rect 10780 10498 10836 10500
rect 10780 10446 10782 10498
rect 10782 10446 10834 10498
rect 10834 10446 10836 10498
rect 10780 10444 10836 10446
rect 10556 10332 10612 10388
rect 10444 8876 10500 8932
rect 10332 6860 10388 6916
rect 9772 6300 9828 6356
rect 10108 6076 10164 6132
rect 9996 5906 10052 5908
rect 9996 5854 9998 5906
rect 9998 5854 10050 5906
rect 10050 5854 10052 5906
rect 9996 5852 10052 5854
rect 10444 5906 10500 5908
rect 10444 5854 10446 5906
rect 10446 5854 10498 5906
rect 10498 5854 10500 5906
rect 10444 5852 10500 5854
rect 11676 11564 11732 11620
rect 11228 11394 11284 11396
rect 11228 11342 11230 11394
rect 11230 11342 11282 11394
rect 11282 11342 11284 11394
rect 11228 11340 11284 11342
rect 12236 11394 12292 11396
rect 12236 11342 12238 11394
rect 12238 11342 12290 11394
rect 12290 11342 12292 11394
rect 12236 11340 12292 11342
rect 12012 11170 12068 11172
rect 12012 11118 12014 11170
rect 12014 11118 12066 11170
rect 12066 11118 12068 11170
rect 12012 11116 12068 11118
rect 11116 10332 11172 10388
rect 11900 9884 11956 9940
rect 10668 9826 10724 9828
rect 10668 9774 10670 9826
rect 10670 9774 10722 9826
rect 10722 9774 10724 9826
rect 10668 9772 10724 9774
rect 10668 8988 10724 9044
rect 11452 9772 11508 9828
rect 11676 9714 11732 9716
rect 11676 9662 11678 9714
rect 11678 9662 11730 9714
rect 11730 9662 11732 9714
rect 11676 9660 11732 9662
rect 10892 8988 10948 9044
rect 10780 8482 10836 8484
rect 10780 8430 10782 8482
rect 10782 8430 10834 8482
rect 10834 8430 10836 8482
rect 10780 8428 10836 8430
rect 12236 9436 12292 9492
rect 10780 8258 10836 8260
rect 10780 8206 10782 8258
rect 10782 8206 10834 8258
rect 10834 8206 10836 8258
rect 10780 8204 10836 8206
rect 11452 7644 11508 7700
rect 12684 15148 12740 15204
rect 12908 14588 12964 14644
rect 12460 11452 12516 11508
rect 12460 11170 12516 11172
rect 12460 11118 12462 11170
rect 12462 11118 12514 11170
rect 12514 11118 12516 11170
rect 12460 11116 12516 11118
rect 12796 14306 12852 14308
rect 12796 14254 12798 14306
rect 12798 14254 12850 14306
rect 12850 14254 12852 14306
rect 12796 14252 12852 14254
rect 12796 13970 12852 13972
rect 12796 13918 12798 13970
rect 12798 13918 12850 13970
rect 12850 13918 12852 13970
rect 12796 13916 12852 13918
rect 13692 15932 13748 15988
rect 13244 15820 13300 15876
rect 14028 15820 14084 15876
rect 12684 13746 12740 13748
rect 12684 13694 12686 13746
rect 12686 13694 12738 13746
rect 12738 13694 12740 13746
rect 12684 13692 12740 13694
rect 13132 13244 13188 13300
rect 12796 11340 12852 11396
rect 13468 14588 13524 14644
rect 14924 16994 14980 16996
rect 14924 16942 14926 16994
rect 14926 16942 14978 16994
rect 14978 16942 14980 16994
rect 14924 16940 14980 16942
rect 14588 15148 14644 15204
rect 13468 13074 13524 13076
rect 13468 13022 13470 13074
rect 13470 13022 13522 13074
rect 13522 13022 13524 13074
rect 13468 13020 13524 13022
rect 13020 11452 13076 11508
rect 12684 11282 12740 11284
rect 12684 11230 12686 11282
rect 12686 11230 12738 11282
rect 12738 11230 12740 11282
rect 12684 11228 12740 11230
rect 11900 8876 11956 8932
rect 12684 9602 12740 9604
rect 12684 9550 12686 9602
rect 12686 9550 12738 9602
rect 12738 9550 12740 9602
rect 12684 9548 12740 9550
rect 12572 9436 12628 9492
rect 12572 8764 12628 8820
rect 11900 7980 11956 8036
rect 11564 7532 11620 7588
rect 11676 6860 11732 6916
rect 10668 6748 10724 6804
rect 11452 6748 11508 6804
rect 11004 6578 11060 6580
rect 11004 6526 11006 6578
rect 11006 6526 11058 6578
rect 11058 6526 11060 6578
rect 11004 6524 11060 6526
rect 10780 6018 10836 6020
rect 10780 5966 10782 6018
rect 10782 5966 10834 6018
rect 10834 5966 10836 6018
rect 10780 5964 10836 5966
rect 11228 5964 11284 6020
rect 11116 5906 11172 5908
rect 11116 5854 11118 5906
rect 11118 5854 11170 5906
rect 11170 5854 11172 5906
rect 11116 5852 11172 5854
rect 11004 5292 11060 5348
rect 9772 4508 9828 4564
rect 8988 4226 9044 4228
rect 8988 4174 8990 4226
rect 8990 4174 9042 4226
rect 9042 4174 9044 4226
rect 8988 4172 9044 4174
rect 9436 4060 9492 4116
rect 9324 3724 9380 3780
rect 9548 3836 9604 3892
rect 10108 3612 10164 3668
rect 11452 6188 11508 6244
rect 10892 5010 10948 5012
rect 10892 4958 10894 5010
rect 10894 4958 10946 5010
rect 10946 4958 10948 5010
rect 10892 4956 10948 4958
rect 12124 6860 12180 6916
rect 12908 9884 12964 9940
rect 13468 11394 13524 11396
rect 13468 11342 13470 11394
rect 13470 11342 13522 11394
rect 13522 11342 13524 11394
rect 13468 11340 13524 11342
rect 14028 12738 14084 12740
rect 14028 12686 14030 12738
rect 14030 12686 14082 12738
rect 14082 12686 14084 12738
rect 14028 12684 14084 12686
rect 14476 12850 14532 12852
rect 14476 12798 14478 12850
rect 14478 12798 14530 12850
rect 14530 12798 14532 12850
rect 14476 12796 14532 12798
rect 17276 26012 17332 26068
rect 17388 26908 17444 26964
rect 16716 25452 16772 25508
rect 16940 25340 16996 25396
rect 16716 25228 16772 25284
rect 16156 24834 16212 24836
rect 16156 24782 16158 24834
rect 16158 24782 16210 24834
rect 16210 24782 16212 24834
rect 16156 24780 16212 24782
rect 16044 23772 16100 23828
rect 17052 25228 17108 25284
rect 17276 25452 17332 25508
rect 17276 25004 17332 25060
rect 16940 24722 16996 24724
rect 16940 24670 16942 24722
rect 16942 24670 16994 24722
rect 16994 24670 16996 24722
rect 16940 24668 16996 24670
rect 18284 35532 18340 35588
rect 17948 35084 18004 35140
rect 17948 34748 18004 34804
rect 17948 34130 18004 34132
rect 17948 34078 17950 34130
rect 17950 34078 18002 34130
rect 18002 34078 18004 34130
rect 17948 34076 18004 34078
rect 17836 30940 17892 30996
rect 17836 29820 17892 29876
rect 17724 28700 17780 28756
rect 18060 30156 18116 30212
rect 18508 35084 18564 35140
rect 18508 34636 18564 34692
rect 18508 33346 18564 33348
rect 18508 33294 18510 33346
rect 18510 33294 18562 33346
rect 18562 33294 18564 33346
rect 18508 33292 18564 33294
rect 18060 29596 18116 29652
rect 17948 28588 18004 28644
rect 17948 28364 18004 28420
rect 18956 38108 19012 38164
rect 19404 39506 19460 39508
rect 19404 39454 19406 39506
rect 19406 39454 19458 39506
rect 19458 39454 19460 39506
rect 19404 39452 19460 39454
rect 19516 38946 19572 38948
rect 19516 38894 19518 38946
rect 19518 38894 19570 38946
rect 19570 38894 19572 38946
rect 19516 38892 19572 38894
rect 19404 38162 19460 38164
rect 19404 38110 19406 38162
rect 19406 38110 19458 38162
rect 19458 38110 19460 38162
rect 19404 38108 19460 38110
rect 19292 37436 19348 37492
rect 19516 37490 19572 37492
rect 19516 37438 19518 37490
rect 19518 37438 19570 37490
rect 19570 37438 19572 37490
rect 19516 37436 19572 37438
rect 18956 35980 19012 36036
rect 19180 36764 19236 36820
rect 18732 34972 18788 35028
rect 18956 34972 19012 35028
rect 18732 34300 18788 34356
rect 19516 36764 19572 36820
rect 19180 35084 19236 35140
rect 19404 35810 19460 35812
rect 19404 35758 19406 35810
rect 19406 35758 19458 35810
rect 19458 35758 19460 35810
rect 19404 35756 19460 35758
rect 19292 34972 19348 35028
rect 19852 40124 19908 40180
rect 19836 39226 19892 39228
rect 19836 39174 19838 39226
rect 19838 39174 19890 39226
rect 19890 39174 19892 39226
rect 19836 39172 19892 39174
rect 19940 39226 19996 39228
rect 19940 39174 19942 39226
rect 19942 39174 19994 39226
rect 19994 39174 19996 39226
rect 19940 39172 19996 39174
rect 20044 39226 20100 39228
rect 20044 39174 20046 39226
rect 20046 39174 20098 39226
rect 20098 39174 20100 39226
rect 20044 39172 20100 39174
rect 20188 38892 20244 38948
rect 20300 39340 20356 39396
rect 20300 38780 20356 38836
rect 20636 40236 20692 40292
rect 19852 38220 19908 38276
rect 19836 37658 19892 37660
rect 19836 37606 19838 37658
rect 19838 37606 19890 37658
rect 19890 37606 19892 37658
rect 19836 37604 19892 37606
rect 19940 37658 19996 37660
rect 19940 37606 19942 37658
rect 19942 37606 19994 37658
rect 19994 37606 19996 37658
rect 19940 37604 19996 37606
rect 20044 37658 20100 37660
rect 20044 37606 20046 37658
rect 20046 37606 20098 37658
rect 20098 37606 20100 37658
rect 20044 37604 20100 37606
rect 20188 37436 20244 37492
rect 20300 37212 20356 37268
rect 20412 37884 20468 37940
rect 21644 41804 21700 41860
rect 20972 40236 21028 40292
rect 22316 41020 22372 41076
rect 24556 45778 24612 45780
rect 24556 45726 24558 45778
rect 24558 45726 24610 45778
rect 24610 45726 24612 45778
rect 24556 45724 24612 45726
rect 25340 45724 25396 45780
rect 23884 45164 23940 45220
rect 24444 45106 24500 45108
rect 24444 45054 24446 45106
rect 24446 45054 24498 45106
rect 24498 45054 24500 45106
rect 24444 45052 24500 45054
rect 23212 42700 23268 42756
rect 23100 41858 23156 41860
rect 23100 41806 23102 41858
rect 23102 41806 23154 41858
rect 23154 41806 23156 41858
rect 23100 41804 23156 41806
rect 23548 41692 23604 41748
rect 22876 40572 22932 40628
rect 21756 40236 21812 40292
rect 20860 37324 20916 37380
rect 21084 37266 21140 37268
rect 21084 37214 21086 37266
rect 21086 37214 21138 37266
rect 21138 37214 21140 37266
rect 21084 37212 21140 37214
rect 20748 36764 20804 36820
rect 19836 36090 19892 36092
rect 19836 36038 19838 36090
rect 19838 36038 19890 36090
rect 19890 36038 19892 36090
rect 19836 36036 19892 36038
rect 19940 36090 19996 36092
rect 19940 36038 19942 36090
rect 19942 36038 19994 36090
rect 19994 36038 19996 36090
rect 19940 36036 19996 36038
rect 20044 36090 20100 36092
rect 20044 36038 20046 36090
rect 20046 36038 20098 36090
rect 20098 36038 20100 36090
rect 20044 36036 20100 36038
rect 19964 35922 20020 35924
rect 19964 35870 19966 35922
rect 19966 35870 20018 35922
rect 20018 35870 20020 35922
rect 19964 35868 20020 35870
rect 19740 35084 19796 35140
rect 19628 34914 19684 34916
rect 19628 34862 19630 34914
rect 19630 34862 19682 34914
rect 19682 34862 19684 34914
rect 19628 34860 19684 34862
rect 18844 34748 18900 34804
rect 18956 34690 19012 34692
rect 18956 34638 18958 34690
rect 18958 34638 19010 34690
rect 19010 34638 19012 34690
rect 18956 34636 19012 34638
rect 18956 34242 19012 34244
rect 18956 34190 18958 34242
rect 18958 34190 19010 34242
rect 19010 34190 19012 34242
rect 18956 34188 19012 34190
rect 19292 34636 19348 34692
rect 19180 34130 19236 34132
rect 19180 34078 19182 34130
rect 19182 34078 19234 34130
rect 19234 34078 19236 34130
rect 19180 34076 19236 34078
rect 20076 34914 20132 34916
rect 20076 34862 20078 34914
rect 20078 34862 20130 34914
rect 20130 34862 20132 34914
rect 20076 34860 20132 34862
rect 19852 34748 19908 34804
rect 20188 34748 20244 34804
rect 19740 34636 19796 34692
rect 19836 34522 19892 34524
rect 19836 34470 19838 34522
rect 19838 34470 19890 34522
rect 19890 34470 19892 34522
rect 19836 34468 19892 34470
rect 19940 34522 19996 34524
rect 19940 34470 19942 34522
rect 19942 34470 19994 34522
rect 19994 34470 19996 34522
rect 19940 34468 19996 34470
rect 20044 34522 20100 34524
rect 20044 34470 20046 34522
rect 20046 34470 20098 34522
rect 20098 34470 20100 34522
rect 20044 34468 20100 34470
rect 19852 34300 19908 34356
rect 19516 33740 19572 33796
rect 19628 34188 19684 34244
rect 19292 33628 19348 33684
rect 18956 32786 19012 32788
rect 18956 32734 18958 32786
rect 18958 32734 19010 32786
rect 19010 32734 19012 32786
rect 18956 32732 19012 32734
rect 18844 32172 18900 32228
rect 18508 30268 18564 30324
rect 18620 31612 18676 31668
rect 18284 30044 18340 30100
rect 18396 29596 18452 29652
rect 18508 29932 18564 29988
rect 18172 28588 18228 28644
rect 17836 28082 17892 28084
rect 17836 28030 17838 28082
rect 17838 28030 17890 28082
rect 17890 28030 17892 28082
rect 17836 28028 17892 28030
rect 17724 27916 17780 27972
rect 18396 27858 18452 27860
rect 18396 27806 18398 27858
rect 18398 27806 18450 27858
rect 18450 27806 18452 27858
rect 18396 27804 18452 27806
rect 18060 27468 18116 27524
rect 17836 26962 17892 26964
rect 17836 26910 17838 26962
rect 17838 26910 17890 26962
rect 17890 26910 17892 26962
rect 17836 26908 17892 26910
rect 17500 25340 17556 25396
rect 17612 25116 17668 25172
rect 17500 24892 17556 24948
rect 17836 25506 17892 25508
rect 17836 25454 17838 25506
rect 17838 25454 17890 25506
rect 17890 25454 17892 25506
rect 17836 25452 17892 25454
rect 18284 26402 18340 26404
rect 18284 26350 18286 26402
rect 18286 26350 18338 26402
rect 18338 26350 18340 26402
rect 18284 26348 18340 26350
rect 20188 33404 20244 33460
rect 19836 32954 19892 32956
rect 19836 32902 19838 32954
rect 19838 32902 19890 32954
rect 19890 32902 19892 32954
rect 19836 32900 19892 32902
rect 19940 32954 19996 32956
rect 19940 32902 19942 32954
rect 19942 32902 19994 32954
rect 19994 32902 19996 32954
rect 19940 32900 19996 32902
rect 20044 32954 20100 32956
rect 20044 32902 20046 32954
rect 20046 32902 20098 32954
rect 20098 32902 20100 32954
rect 20044 32900 20100 32902
rect 19516 32620 19572 32676
rect 19292 31948 19348 32004
rect 20188 32450 20244 32452
rect 20188 32398 20190 32450
rect 20190 32398 20242 32450
rect 20242 32398 20244 32450
rect 20188 32396 20244 32398
rect 19852 31948 19908 32004
rect 19516 31554 19572 31556
rect 19516 31502 19518 31554
rect 19518 31502 19570 31554
rect 19570 31502 19572 31554
rect 19516 31500 19572 31502
rect 20412 36540 20468 36596
rect 20860 35644 20916 35700
rect 20972 32450 21028 32452
rect 20972 32398 20974 32450
rect 20974 32398 21026 32450
rect 21026 32398 21028 32450
rect 20972 32396 21028 32398
rect 21532 38556 21588 38612
rect 23212 40012 23268 40068
rect 22652 39058 22708 39060
rect 22652 39006 22654 39058
rect 22654 39006 22706 39058
rect 22706 39006 22708 39058
rect 22652 39004 22708 39006
rect 22092 38780 22148 38836
rect 21980 38556 22036 38612
rect 23660 40012 23716 40068
rect 24108 39564 24164 39620
rect 21644 37938 21700 37940
rect 21644 37886 21646 37938
rect 21646 37886 21698 37938
rect 21698 37886 21700 37938
rect 21644 37884 21700 37886
rect 21644 37378 21700 37380
rect 21644 37326 21646 37378
rect 21646 37326 21698 37378
rect 21698 37326 21700 37378
rect 21644 37324 21700 37326
rect 21532 37100 21588 37156
rect 21308 34972 21364 35028
rect 21868 37212 21924 37268
rect 22764 37996 22820 38052
rect 22876 38332 22932 38388
rect 22540 37324 22596 37380
rect 21532 35756 21588 35812
rect 21532 35196 21588 35252
rect 21868 36258 21924 36260
rect 21868 36206 21870 36258
rect 21870 36206 21922 36258
rect 21922 36206 21924 36258
rect 21868 36204 21924 36206
rect 21756 35196 21812 35252
rect 21868 34300 21924 34356
rect 22876 37772 22932 37828
rect 22652 36204 22708 36260
rect 22764 37436 22820 37492
rect 22540 35084 22596 35140
rect 22428 34860 22484 34916
rect 22540 34802 22596 34804
rect 22540 34750 22542 34802
rect 22542 34750 22594 34802
rect 22594 34750 22596 34802
rect 22540 34748 22596 34750
rect 22988 36764 23044 36820
rect 22988 35196 23044 35252
rect 22876 34860 22932 34916
rect 22764 34524 22820 34580
rect 23324 38556 23380 38612
rect 25340 45052 25396 45108
rect 24892 43372 24948 43428
rect 24556 41804 24612 41860
rect 24892 41692 24948 41748
rect 25116 41916 25172 41972
rect 26236 46060 26292 46116
rect 29372 46114 29428 46116
rect 29372 46062 29374 46114
rect 29374 46062 29426 46114
rect 29426 46062 29428 46114
rect 29372 46060 29428 46062
rect 30268 46060 30324 46116
rect 25564 45276 25620 45332
rect 25676 45164 25732 45220
rect 25900 42476 25956 42532
rect 26124 43708 26180 43764
rect 27356 45052 27412 45108
rect 26572 44716 26628 44772
rect 26908 44492 26964 44548
rect 28588 44716 28644 44772
rect 27692 44546 27748 44548
rect 27692 44494 27694 44546
rect 27694 44494 27746 44546
rect 27746 44494 27748 44546
rect 27692 44492 27748 44494
rect 28700 44268 28756 44324
rect 30380 45106 30436 45108
rect 30380 45054 30382 45106
rect 30382 45054 30434 45106
rect 30434 45054 30436 45106
rect 30380 45052 30436 45054
rect 29932 44322 29988 44324
rect 29932 44270 29934 44322
rect 29934 44270 29986 44322
rect 29986 44270 29988 44322
rect 29932 44268 29988 44270
rect 28364 44044 28420 44100
rect 26572 43708 26628 43764
rect 29372 44098 29428 44100
rect 29372 44046 29374 44098
rect 29374 44046 29426 44098
rect 29426 44046 29428 44098
rect 29372 44044 29428 44046
rect 29148 43762 29204 43764
rect 29148 43710 29150 43762
rect 29150 43710 29202 43762
rect 29202 43710 29204 43762
rect 29148 43708 29204 43710
rect 29820 43708 29876 43764
rect 30380 44322 30436 44324
rect 30380 44270 30382 44322
rect 30382 44270 30434 44322
rect 30434 44270 30436 44322
rect 30380 44268 30436 44270
rect 30268 44044 30324 44100
rect 28476 42700 28532 42756
rect 27356 42642 27412 42644
rect 27356 42590 27358 42642
rect 27358 42590 27410 42642
rect 27410 42590 27412 42642
rect 27356 42588 27412 42590
rect 29260 42642 29316 42644
rect 29260 42590 29262 42642
rect 29262 42590 29314 42642
rect 29314 42590 29316 42642
rect 29260 42588 29316 42590
rect 26572 42530 26628 42532
rect 26572 42478 26574 42530
rect 26574 42478 26626 42530
rect 26626 42478 26628 42530
rect 26572 42476 26628 42478
rect 24668 39506 24724 39508
rect 24668 39454 24670 39506
rect 24670 39454 24722 39506
rect 24722 39454 24724 39506
rect 24668 39452 24724 39454
rect 24220 37772 24276 37828
rect 23772 37548 23828 37604
rect 23436 37436 23492 37492
rect 23548 37378 23604 37380
rect 23548 37326 23550 37378
rect 23550 37326 23602 37378
rect 23602 37326 23604 37378
rect 23548 37324 23604 37326
rect 24668 37436 24724 37492
rect 23324 37212 23380 37268
rect 23436 35868 23492 35924
rect 23884 37100 23940 37156
rect 23324 35644 23380 35700
rect 23772 35308 23828 35364
rect 23212 34860 23268 34916
rect 21196 32172 21252 32228
rect 20300 31778 20356 31780
rect 20300 31726 20302 31778
rect 20302 31726 20354 31778
rect 20354 31726 20356 31778
rect 20300 31724 20356 31726
rect 19836 31386 19892 31388
rect 19836 31334 19838 31386
rect 19838 31334 19890 31386
rect 19890 31334 19892 31386
rect 19836 31332 19892 31334
rect 19940 31386 19996 31388
rect 19940 31334 19942 31386
rect 19942 31334 19994 31386
rect 19994 31334 19996 31386
rect 19940 31332 19996 31334
rect 20044 31386 20100 31388
rect 20044 31334 20046 31386
rect 20046 31334 20098 31386
rect 20098 31334 20100 31386
rect 20044 31332 20100 31334
rect 18956 31052 19012 31108
rect 19516 30882 19572 30884
rect 19516 30830 19518 30882
rect 19518 30830 19570 30882
rect 19570 30830 19572 30882
rect 19516 30828 19572 30830
rect 18956 30268 19012 30324
rect 19180 30268 19236 30324
rect 19180 29932 19236 29988
rect 18956 29314 19012 29316
rect 18956 29262 18958 29314
rect 18958 29262 19010 29314
rect 19010 29262 19012 29314
rect 18956 29260 19012 29262
rect 18956 28642 19012 28644
rect 18956 28590 18958 28642
rect 18958 28590 19010 28642
rect 19010 28590 19012 28642
rect 18956 28588 19012 28590
rect 19180 28028 19236 28084
rect 18508 26124 18564 26180
rect 18396 26066 18452 26068
rect 18396 26014 18398 26066
rect 18398 26014 18450 26066
rect 18450 26014 18452 26066
rect 18396 26012 18452 26014
rect 18060 25564 18116 25620
rect 18172 25676 18228 25732
rect 18396 25452 18452 25508
rect 17836 25228 17892 25284
rect 16940 23996 16996 24052
rect 16156 23212 16212 23268
rect 16044 22876 16100 22932
rect 17276 23938 17332 23940
rect 17276 23886 17278 23938
rect 17278 23886 17330 23938
rect 17330 23886 17332 23938
rect 17276 23884 17332 23886
rect 17388 23714 17444 23716
rect 17388 23662 17390 23714
rect 17390 23662 17442 23714
rect 17442 23662 17444 23714
rect 17388 23660 17444 23662
rect 17836 23996 17892 24052
rect 17836 23324 17892 23380
rect 18284 25004 18340 25060
rect 18060 24668 18116 24724
rect 18284 23826 18340 23828
rect 18284 23774 18286 23826
rect 18286 23774 18338 23826
rect 18338 23774 18340 23826
rect 18284 23772 18340 23774
rect 16492 21474 16548 21476
rect 16492 21422 16494 21474
rect 16494 21422 16546 21474
rect 16546 21422 16548 21474
rect 16492 21420 16548 21422
rect 17836 22652 17892 22708
rect 15820 20636 15876 20692
rect 15708 20242 15764 20244
rect 15708 20190 15710 20242
rect 15710 20190 15762 20242
rect 15762 20190 15764 20242
rect 15708 20188 15764 20190
rect 16604 20636 16660 20692
rect 16380 20578 16436 20580
rect 16380 20526 16382 20578
rect 16382 20526 16434 20578
rect 16434 20526 16436 20578
rect 16380 20524 16436 20526
rect 16044 20018 16100 20020
rect 16044 19966 16046 20018
rect 16046 19966 16098 20018
rect 16098 19966 16100 20018
rect 16044 19964 16100 19966
rect 16044 18956 16100 19012
rect 15932 18620 15988 18676
rect 15820 17388 15876 17444
rect 15148 16828 15204 16884
rect 15372 16716 15428 16772
rect 15820 15202 15876 15204
rect 15820 15150 15822 15202
rect 15822 15150 15874 15202
rect 15874 15150 15876 15202
rect 15820 15148 15876 15150
rect 16044 16770 16100 16772
rect 16044 16718 16046 16770
rect 16046 16718 16098 16770
rect 16098 16718 16100 16770
rect 16044 16716 16100 16718
rect 15036 12796 15092 12852
rect 15372 12796 15428 12852
rect 14028 12066 14084 12068
rect 14028 12014 14030 12066
rect 14030 12014 14082 12066
rect 14082 12014 14084 12066
rect 14028 12012 14084 12014
rect 13692 11676 13748 11732
rect 13020 8370 13076 8372
rect 13020 8318 13022 8370
rect 13022 8318 13074 8370
rect 13074 8318 13076 8370
rect 13020 8316 13076 8318
rect 12908 8204 12964 8260
rect 12572 7532 12628 7588
rect 12348 6860 12404 6916
rect 12572 6972 12628 7028
rect 11900 6018 11956 6020
rect 11900 5966 11902 6018
rect 11902 5966 11954 6018
rect 11954 5966 11956 6018
rect 11900 5964 11956 5966
rect 11900 5682 11956 5684
rect 11900 5630 11902 5682
rect 11902 5630 11954 5682
rect 11954 5630 11956 5682
rect 11900 5628 11956 5630
rect 11788 5180 11844 5236
rect 11788 5010 11844 5012
rect 11788 4958 11790 5010
rect 11790 4958 11842 5010
rect 11842 4958 11844 5010
rect 11788 4956 11844 4958
rect 11564 4732 11620 4788
rect 10780 4396 10836 4452
rect 10668 4114 10724 4116
rect 10668 4062 10670 4114
rect 10670 4062 10722 4114
rect 10722 4062 10724 4114
rect 10668 4060 10724 4062
rect 10780 3836 10836 3892
rect 13468 8316 13524 8372
rect 13692 9548 13748 9604
rect 14364 9212 14420 9268
rect 14476 9100 14532 9156
rect 15148 12684 15204 12740
rect 15932 12178 15988 12180
rect 15932 12126 15934 12178
rect 15934 12126 15986 12178
rect 15986 12126 15988 12178
rect 15932 12124 15988 12126
rect 15148 11900 15204 11956
rect 15708 12012 15764 12068
rect 15484 10108 15540 10164
rect 14924 9324 14980 9380
rect 14812 9100 14868 9156
rect 13580 8204 13636 8260
rect 13132 7756 13188 7812
rect 12572 6578 12628 6580
rect 12572 6526 12574 6578
rect 12574 6526 12626 6578
rect 12626 6526 12628 6578
rect 12572 6524 12628 6526
rect 12684 6466 12740 6468
rect 12684 6414 12686 6466
rect 12686 6414 12738 6466
rect 12738 6414 12740 6466
rect 12684 6412 12740 6414
rect 12460 6076 12516 6132
rect 12124 3500 12180 3556
rect 12236 5740 12292 5796
rect 12684 5740 12740 5796
rect 12572 5068 12628 5124
rect 12684 4956 12740 5012
rect 12908 6690 12964 6692
rect 12908 6638 12910 6690
rect 12910 6638 12962 6690
rect 12962 6638 12964 6690
rect 12908 6636 12964 6638
rect 13020 6860 13076 6916
rect 12908 6130 12964 6132
rect 12908 6078 12910 6130
rect 12910 6078 12962 6130
rect 12962 6078 12964 6130
rect 12908 6076 12964 6078
rect 13132 6412 13188 6468
rect 13244 6076 13300 6132
rect 13132 6018 13188 6020
rect 13132 5966 13134 6018
rect 13134 5966 13186 6018
rect 13186 5966 13188 6018
rect 13132 5964 13188 5966
rect 12908 4732 12964 4788
rect 14028 8146 14084 8148
rect 14028 8094 14030 8146
rect 14030 8094 14082 8146
rect 14082 8094 14084 8146
rect 14028 8092 14084 8094
rect 14252 7644 14308 7700
rect 14588 7868 14644 7924
rect 13580 6748 13636 6804
rect 13692 6690 13748 6692
rect 13692 6638 13694 6690
rect 13694 6638 13746 6690
rect 13746 6638 13748 6690
rect 13692 6636 13748 6638
rect 13692 6412 13748 6468
rect 13468 5628 13524 5684
rect 13580 5292 13636 5348
rect 13916 5740 13972 5796
rect 13804 5292 13860 5348
rect 14476 5180 14532 5236
rect 13916 4956 13972 5012
rect 13468 3554 13524 3556
rect 13468 3502 13470 3554
rect 13470 3502 13522 3554
rect 13522 3502 13524 3554
rect 13468 3500 13524 3502
rect 14140 4898 14196 4900
rect 14140 4846 14142 4898
rect 14142 4846 14194 4898
rect 14194 4846 14196 4898
rect 14140 4844 14196 4846
rect 13692 4226 13748 4228
rect 13692 4174 13694 4226
rect 13694 4174 13746 4226
rect 13746 4174 13748 4226
rect 13692 4172 13748 4174
rect 14252 4172 14308 4228
rect 14140 3500 14196 3556
rect 14700 6466 14756 6468
rect 14700 6414 14702 6466
rect 14702 6414 14754 6466
rect 14754 6414 14756 6466
rect 14700 6412 14756 6414
rect 15932 9324 15988 9380
rect 15036 9266 15092 9268
rect 15036 9214 15038 9266
rect 15038 9214 15090 9266
rect 15090 9214 15092 9266
rect 15036 9212 15092 9214
rect 16380 20300 16436 20356
rect 16716 20524 16772 20580
rect 17276 20578 17332 20580
rect 17276 20526 17278 20578
rect 17278 20526 17330 20578
rect 17330 20526 17332 20578
rect 17276 20524 17332 20526
rect 16940 20300 16996 20356
rect 16828 19516 16884 19572
rect 17388 19404 17444 19460
rect 16268 18620 16324 18676
rect 16268 18226 16324 18228
rect 16268 18174 16270 18226
rect 16270 18174 16322 18226
rect 16322 18174 16324 18226
rect 16268 18172 16324 18174
rect 16380 17724 16436 17780
rect 16268 17388 16324 17444
rect 16716 19010 16772 19012
rect 16716 18958 16718 19010
rect 16718 18958 16770 19010
rect 16770 18958 16772 19010
rect 16716 18956 16772 18958
rect 18060 20524 18116 20580
rect 16940 18956 16996 19012
rect 17276 18732 17332 18788
rect 16828 17778 16884 17780
rect 16828 17726 16830 17778
rect 16830 17726 16882 17778
rect 16882 17726 16884 17778
rect 16828 17724 16884 17726
rect 16940 17500 16996 17556
rect 16828 16828 16884 16884
rect 16940 16716 16996 16772
rect 16492 15874 16548 15876
rect 16492 15822 16494 15874
rect 16494 15822 16546 15874
rect 16546 15822 16548 15874
rect 16492 15820 16548 15822
rect 16380 15426 16436 15428
rect 16380 15374 16382 15426
rect 16382 15374 16434 15426
rect 16434 15374 16436 15426
rect 16380 15372 16436 15374
rect 17500 17612 17556 17668
rect 17500 17442 17556 17444
rect 17500 17390 17502 17442
rect 17502 17390 17554 17442
rect 17554 17390 17556 17442
rect 17500 17388 17556 17390
rect 17836 17554 17892 17556
rect 17836 17502 17838 17554
rect 17838 17502 17890 17554
rect 17890 17502 17892 17554
rect 17836 17500 17892 17502
rect 17612 17164 17668 17220
rect 17948 17388 18004 17444
rect 17500 16716 17556 16772
rect 17276 16156 17332 16212
rect 17388 15932 17444 15988
rect 16492 14476 16548 14532
rect 16716 14306 16772 14308
rect 16716 14254 16718 14306
rect 16718 14254 16770 14306
rect 16770 14254 16772 14306
rect 16716 14252 16772 14254
rect 16604 13468 16660 13524
rect 16268 13020 16324 13076
rect 16716 12796 16772 12852
rect 16604 12066 16660 12068
rect 16604 12014 16606 12066
rect 16606 12014 16658 12066
rect 16658 12014 16660 12066
rect 16604 12012 16660 12014
rect 16492 11954 16548 11956
rect 16492 11902 16494 11954
rect 16494 11902 16546 11954
rect 16546 11902 16548 11954
rect 16492 11900 16548 11902
rect 17276 15596 17332 15652
rect 16940 15148 16996 15204
rect 17388 15314 17444 15316
rect 17388 15262 17390 15314
rect 17390 15262 17442 15314
rect 17442 15262 17444 15314
rect 17388 15260 17444 15262
rect 17724 15426 17780 15428
rect 17724 15374 17726 15426
rect 17726 15374 17778 15426
rect 17778 15374 17780 15426
rect 17724 15372 17780 15374
rect 17724 14588 17780 14644
rect 17500 14476 17556 14532
rect 18396 22876 18452 22932
rect 18284 20412 18340 20468
rect 18844 26124 18900 26180
rect 18732 25340 18788 25396
rect 19628 30268 19684 30324
rect 19740 30828 19796 30884
rect 19404 30156 19460 30212
rect 19964 30210 20020 30212
rect 19964 30158 19966 30210
rect 19966 30158 20018 30210
rect 20018 30158 20020 30210
rect 19964 30156 20020 30158
rect 19404 29986 19460 29988
rect 19404 29934 19406 29986
rect 19406 29934 19458 29986
rect 19458 29934 19460 29986
rect 19404 29932 19460 29934
rect 19404 29650 19460 29652
rect 19404 29598 19406 29650
rect 19406 29598 19458 29650
rect 19458 29598 19460 29650
rect 19404 29596 19460 29598
rect 19836 29818 19892 29820
rect 19836 29766 19838 29818
rect 19838 29766 19890 29818
rect 19890 29766 19892 29818
rect 19836 29764 19892 29766
rect 19940 29818 19996 29820
rect 19940 29766 19942 29818
rect 19942 29766 19994 29818
rect 19994 29766 19996 29818
rect 19940 29764 19996 29766
rect 20044 29818 20100 29820
rect 20044 29766 20046 29818
rect 20046 29766 20098 29818
rect 20098 29766 20100 29818
rect 20044 29764 20100 29766
rect 20300 30434 20356 30436
rect 20300 30382 20302 30434
rect 20302 30382 20354 30434
rect 20354 30382 20356 30434
rect 20300 30380 20356 30382
rect 20524 31164 20580 31220
rect 20524 30940 20580 30996
rect 21756 33516 21812 33572
rect 21420 31890 21476 31892
rect 21420 31838 21422 31890
rect 21422 31838 21474 31890
rect 21474 31838 21476 31890
rect 21420 31836 21476 31838
rect 21756 31836 21812 31892
rect 21308 31052 21364 31108
rect 20748 30492 20804 30548
rect 21308 30492 21364 30548
rect 21532 30828 21588 30884
rect 22540 34076 22596 34132
rect 22316 33516 22372 33572
rect 21980 32674 22036 32676
rect 21980 32622 21982 32674
rect 21982 32622 22034 32674
rect 22034 32622 22036 32674
rect 21980 32620 22036 32622
rect 22092 32562 22148 32564
rect 22092 32510 22094 32562
rect 22094 32510 22146 32562
rect 22146 32510 22148 32562
rect 22092 32508 22148 32510
rect 22316 32620 22372 32676
rect 22428 31836 22484 31892
rect 22204 30604 22260 30660
rect 20524 29932 20580 29988
rect 20636 30044 20692 30100
rect 20412 29596 20468 29652
rect 20188 29372 20244 29428
rect 20076 29314 20132 29316
rect 20076 29262 20078 29314
rect 20078 29262 20130 29314
rect 20130 29262 20132 29314
rect 20076 29260 20132 29262
rect 20636 29036 20692 29092
rect 21084 29260 21140 29316
rect 19740 28924 19796 28980
rect 20412 28924 20468 28980
rect 20188 28812 20244 28868
rect 19836 28250 19892 28252
rect 19836 28198 19838 28250
rect 19838 28198 19890 28250
rect 19890 28198 19892 28250
rect 19836 28196 19892 28198
rect 19940 28250 19996 28252
rect 19940 28198 19942 28250
rect 19942 28198 19994 28250
rect 19994 28198 19996 28250
rect 19940 28196 19996 28198
rect 20044 28250 20100 28252
rect 20044 28198 20046 28250
rect 20046 28198 20098 28250
rect 20098 28198 20100 28250
rect 20044 28196 20100 28198
rect 19836 26682 19892 26684
rect 19836 26630 19838 26682
rect 19838 26630 19890 26682
rect 19890 26630 19892 26682
rect 19836 26628 19892 26630
rect 19940 26682 19996 26684
rect 19940 26630 19942 26682
rect 19942 26630 19994 26682
rect 19994 26630 19996 26682
rect 19940 26628 19996 26630
rect 20044 26682 20100 26684
rect 20044 26630 20046 26682
rect 20046 26630 20098 26682
rect 20098 26630 20100 26682
rect 20044 26628 20100 26630
rect 20188 26124 20244 26180
rect 19292 25564 19348 25620
rect 19852 25788 19908 25844
rect 19852 25506 19908 25508
rect 19852 25454 19854 25506
rect 19854 25454 19906 25506
rect 19906 25454 19908 25506
rect 19852 25452 19908 25454
rect 20188 25340 20244 25396
rect 18844 25116 18900 25172
rect 20412 25788 20468 25844
rect 20748 27186 20804 27188
rect 20748 27134 20750 27186
rect 20750 27134 20802 27186
rect 20802 27134 20804 27186
rect 20748 27132 20804 27134
rect 20412 25394 20468 25396
rect 20412 25342 20414 25394
rect 20414 25342 20466 25394
rect 20466 25342 20468 25394
rect 20412 25340 20468 25342
rect 20300 25228 20356 25284
rect 19404 25116 19460 25172
rect 19836 25114 19892 25116
rect 19836 25062 19838 25114
rect 19838 25062 19890 25114
rect 19890 25062 19892 25114
rect 19836 25060 19892 25062
rect 19940 25114 19996 25116
rect 19940 25062 19942 25114
rect 19942 25062 19994 25114
rect 19994 25062 19996 25114
rect 19940 25060 19996 25062
rect 20044 25114 20100 25116
rect 20044 25062 20046 25114
rect 20046 25062 20098 25114
rect 20098 25062 20100 25114
rect 20044 25060 20100 25062
rect 19852 24556 19908 24612
rect 20748 24556 20804 24612
rect 19836 23546 19892 23548
rect 19836 23494 19838 23546
rect 19838 23494 19890 23546
rect 19890 23494 19892 23546
rect 19836 23492 19892 23494
rect 19940 23546 19996 23548
rect 19940 23494 19942 23546
rect 19942 23494 19994 23546
rect 19994 23494 19996 23546
rect 19940 23492 19996 23494
rect 20044 23546 20100 23548
rect 20044 23494 20046 23546
rect 20046 23494 20098 23546
rect 20098 23494 20100 23546
rect 20044 23492 20100 23494
rect 19068 22540 19124 22596
rect 21308 29372 21364 29428
rect 21196 28476 21252 28532
rect 21308 29036 21364 29092
rect 21756 30322 21812 30324
rect 21756 30270 21758 30322
rect 21758 30270 21810 30322
rect 21810 30270 21812 30322
rect 21756 30268 21812 30270
rect 21980 30156 22036 30212
rect 21644 30098 21700 30100
rect 21644 30046 21646 30098
rect 21646 30046 21698 30098
rect 21698 30046 21700 30098
rect 21644 30044 21700 30046
rect 21756 29426 21812 29428
rect 21756 29374 21758 29426
rect 21758 29374 21810 29426
rect 21810 29374 21812 29426
rect 21756 29372 21812 29374
rect 21308 27858 21364 27860
rect 21308 27806 21310 27858
rect 21310 27806 21362 27858
rect 21362 27806 21364 27858
rect 21308 27804 21364 27806
rect 21196 27244 21252 27300
rect 22988 34130 23044 34132
rect 22988 34078 22990 34130
rect 22990 34078 23042 34130
rect 23042 34078 23044 34130
rect 22988 34076 23044 34078
rect 23100 33628 23156 33684
rect 23100 33346 23156 33348
rect 23100 33294 23102 33346
rect 23102 33294 23154 33346
rect 23154 33294 23156 33346
rect 23100 33292 23156 33294
rect 22988 33122 23044 33124
rect 22988 33070 22990 33122
rect 22990 33070 23042 33122
rect 23042 33070 23044 33122
rect 22988 33068 23044 33070
rect 24332 37266 24388 37268
rect 24332 37214 24334 37266
rect 24334 37214 24386 37266
rect 24386 37214 24388 37266
rect 24332 37212 24388 37214
rect 24108 36482 24164 36484
rect 24108 36430 24110 36482
rect 24110 36430 24162 36482
rect 24162 36430 24164 36482
rect 24108 36428 24164 36430
rect 24332 35922 24388 35924
rect 24332 35870 24334 35922
rect 24334 35870 24386 35922
rect 24386 35870 24388 35922
rect 24332 35868 24388 35870
rect 23996 35308 24052 35364
rect 24108 34690 24164 34692
rect 24108 34638 24110 34690
rect 24110 34638 24162 34690
rect 24162 34638 24164 34690
rect 24108 34636 24164 34638
rect 24668 34636 24724 34692
rect 23772 33628 23828 33684
rect 22988 32284 23044 32340
rect 22764 31836 22820 31892
rect 22652 30828 22708 30884
rect 22540 30156 22596 30212
rect 23100 31836 23156 31892
rect 23436 32562 23492 32564
rect 23436 32510 23438 32562
rect 23438 32510 23490 32562
rect 23490 32510 23492 32562
rect 23436 32508 23492 32510
rect 23324 32396 23380 32452
rect 23660 32172 23716 32228
rect 23884 33346 23940 33348
rect 23884 33294 23886 33346
rect 23886 33294 23938 33346
rect 23938 33294 23940 33346
rect 23884 33292 23940 33294
rect 24220 34018 24276 34020
rect 24220 33966 24222 34018
rect 24222 33966 24274 34018
rect 24274 33966 24276 34018
rect 24220 33964 24276 33966
rect 24668 34076 24724 34132
rect 24332 33628 24388 33684
rect 24892 33628 24948 33684
rect 24220 33234 24276 33236
rect 24220 33182 24222 33234
rect 24222 33182 24274 33234
rect 24274 33182 24276 33234
rect 24220 33180 24276 33182
rect 23772 33068 23828 33124
rect 24444 33122 24500 33124
rect 24444 33070 24446 33122
rect 24446 33070 24498 33122
rect 24498 33070 24500 33122
rect 24444 33068 24500 33070
rect 23884 32674 23940 32676
rect 23884 32622 23886 32674
rect 23886 32622 23938 32674
rect 23938 32622 23940 32674
rect 23884 32620 23940 32622
rect 23996 31836 24052 31892
rect 24220 31890 24276 31892
rect 24220 31838 24222 31890
rect 24222 31838 24274 31890
rect 24274 31838 24276 31890
rect 24220 31836 24276 31838
rect 22876 30828 22932 30884
rect 22652 29986 22708 29988
rect 22652 29934 22654 29986
rect 22654 29934 22706 29986
rect 22706 29934 22708 29986
rect 22652 29932 22708 29934
rect 22092 29372 22148 29428
rect 22652 29148 22708 29204
rect 22764 28476 22820 28532
rect 22204 27970 22260 27972
rect 22204 27918 22206 27970
rect 22206 27918 22258 27970
rect 22258 27918 22260 27970
rect 22204 27916 22260 27918
rect 22988 28588 23044 28644
rect 22764 27132 22820 27188
rect 22092 27020 22148 27076
rect 21308 26796 21364 26852
rect 21196 26460 21252 26516
rect 22092 26178 22148 26180
rect 22092 26126 22094 26178
rect 22094 26126 22146 26178
rect 22146 26126 22148 26178
rect 22092 26124 22148 26126
rect 21420 25788 21476 25844
rect 22316 25618 22372 25620
rect 22316 25566 22318 25618
rect 22318 25566 22370 25618
rect 22370 25566 22372 25618
rect 22316 25564 22372 25566
rect 21420 25506 21476 25508
rect 21420 25454 21422 25506
rect 21422 25454 21474 25506
rect 21474 25454 21476 25506
rect 21420 25452 21476 25454
rect 22428 25228 22484 25284
rect 21868 24610 21924 24612
rect 21868 24558 21870 24610
rect 21870 24558 21922 24610
rect 21922 24558 21924 24610
rect 21868 24556 21924 24558
rect 22428 23436 22484 23492
rect 21084 22316 21140 22372
rect 21756 22258 21812 22260
rect 21756 22206 21758 22258
rect 21758 22206 21810 22258
rect 21810 22206 21812 22258
rect 21756 22204 21812 22206
rect 20188 22092 20244 22148
rect 19836 21978 19892 21980
rect 19836 21926 19838 21978
rect 19838 21926 19890 21978
rect 19890 21926 19892 21978
rect 19836 21924 19892 21926
rect 19940 21978 19996 21980
rect 19940 21926 19942 21978
rect 19942 21926 19994 21978
rect 19994 21926 19996 21978
rect 19940 21924 19996 21926
rect 20044 21978 20100 21980
rect 20044 21926 20046 21978
rect 20046 21926 20098 21978
rect 20098 21926 20100 21978
rect 20044 21924 20100 21926
rect 18956 20748 19012 20804
rect 19836 20410 19892 20412
rect 19836 20358 19838 20410
rect 19838 20358 19890 20410
rect 19890 20358 19892 20410
rect 19836 20356 19892 20358
rect 19940 20410 19996 20412
rect 19940 20358 19942 20410
rect 19942 20358 19994 20410
rect 19994 20358 19996 20410
rect 19940 20356 19996 20358
rect 20044 20410 20100 20412
rect 20044 20358 20046 20410
rect 20046 20358 20098 20410
rect 20098 20358 20100 20410
rect 20044 20356 20100 20358
rect 18844 19292 18900 19348
rect 18956 20076 19012 20132
rect 19740 20076 19796 20132
rect 19516 18620 19572 18676
rect 19836 18842 19892 18844
rect 19836 18790 19838 18842
rect 19838 18790 19890 18842
rect 19890 18790 19892 18842
rect 19836 18788 19892 18790
rect 19940 18842 19996 18844
rect 19940 18790 19942 18842
rect 19942 18790 19994 18842
rect 19994 18790 19996 18842
rect 19940 18788 19996 18790
rect 20044 18842 20100 18844
rect 20044 18790 20046 18842
rect 20046 18790 20098 18842
rect 20098 18790 20100 18842
rect 20044 18788 20100 18790
rect 20636 21810 20692 21812
rect 20636 21758 20638 21810
rect 20638 21758 20690 21810
rect 20690 21758 20692 21810
rect 20636 21756 20692 21758
rect 22540 22258 22596 22260
rect 22540 22206 22542 22258
rect 22542 22206 22594 22258
rect 22594 22206 22596 22258
rect 22540 22204 22596 22206
rect 20300 21532 20356 21588
rect 20748 19794 20804 19796
rect 20748 19742 20750 19794
rect 20750 19742 20802 19794
rect 20802 19742 20804 19794
rect 20748 19740 20804 19742
rect 20412 19180 20468 19236
rect 19740 17666 19796 17668
rect 19740 17614 19742 17666
rect 19742 17614 19794 17666
rect 19794 17614 19796 17666
rect 19740 17612 19796 17614
rect 18284 17442 18340 17444
rect 18284 17390 18286 17442
rect 18286 17390 18338 17442
rect 18338 17390 18340 17442
rect 18284 17388 18340 17390
rect 18284 16044 18340 16100
rect 19292 17164 19348 17220
rect 19836 17274 19892 17276
rect 19836 17222 19838 17274
rect 19838 17222 19890 17274
rect 19890 17222 19892 17274
rect 19836 17220 19892 17222
rect 19940 17274 19996 17276
rect 19940 17222 19942 17274
rect 19942 17222 19994 17274
rect 19994 17222 19996 17274
rect 19940 17220 19996 17222
rect 20044 17274 20100 17276
rect 20044 17222 20046 17274
rect 20046 17222 20098 17274
rect 20098 17222 20100 17274
rect 20044 17220 20100 17222
rect 19628 17052 19684 17108
rect 18396 15596 18452 15652
rect 18172 13020 18228 13076
rect 17724 12908 17780 12964
rect 16044 9212 16100 9268
rect 15708 9042 15764 9044
rect 15708 8990 15710 9042
rect 15710 8990 15762 9042
rect 15762 8990 15764 9042
rect 15708 8988 15764 8990
rect 16492 8988 16548 9044
rect 16268 8818 16324 8820
rect 16268 8766 16270 8818
rect 16270 8766 16322 8818
rect 16322 8766 16324 8818
rect 16268 8764 16324 8766
rect 15148 8540 15204 8596
rect 16940 9548 16996 9604
rect 16716 9212 16772 9268
rect 16492 8540 16548 8596
rect 16268 8204 16324 8260
rect 15596 8146 15652 8148
rect 15596 8094 15598 8146
rect 15598 8094 15650 8146
rect 15650 8094 15652 8146
rect 15596 8092 15652 8094
rect 14924 7644 14980 7700
rect 14700 6076 14756 6132
rect 14924 5740 14980 5796
rect 15036 5292 15092 5348
rect 15148 5234 15204 5236
rect 15148 5182 15150 5234
rect 15150 5182 15202 5234
rect 15202 5182 15204 5234
rect 15148 5180 15204 5182
rect 15596 7868 15652 7924
rect 15484 6076 15540 6132
rect 16604 8092 16660 8148
rect 16268 6524 16324 6580
rect 15484 4508 15540 4564
rect 15820 4226 15876 4228
rect 15820 4174 15822 4226
rect 15822 4174 15874 4226
rect 15874 4174 15876 4226
rect 15820 4172 15876 4174
rect 18172 12178 18228 12180
rect 18172 12126 18174 12178
rect 18174 12126 18226 12178
rect 18226 12126 18228 12178
rect 18172 12124 18228 12126
rect 17724 9996 17780 10052
rect 17612 9714 17668 9716
rect 17612 9662 17614 9714
rect 17614 9662 17666 9714
rect 17666 9662 17668 9714
rect 17612 9660 17668 9662
rect 17948 9548 18004 9604
rect 19964 15986 20020 15988
rect 19964 15934 19966 15986
rect 19966 15934 20018 15986
rect 20018 15934 20020 15986
rect 19964 15932 20020 15934
rect 19836 15706 19892 15708
rect 19836 15654 19838 15706
rect 19838 15654 19890 15706
rect 19890 15654 19892 15706
rect 19836 15652 19892 15654
rect 19940 15706 19996 15708
rect 19940 15654 19942 15706
rect 19942 15654 19994 15706
rect 19994 15654 19996 15706
rect 19940 15652 19996 15654
rect 20044 15706 20100 15708
rect 20044 15654 20046 15706
rect 20046 15654 20098 15706
rect 20098 15654 20100 15706
rect 20044 15652 20100 15654
rect 18620 15202 18676 15204
rect 18620 15150 18622 15202
rect 18622 15150 18674 15202
rect 18674 15150 18676 15202
rect 18620 15148 18676 15150
rect 19836 14138 19892 14140
rect 19836 14086 19838 14138
rect 19838 14086 19890 14138
rect 19890 14086 19892 14138
rect 19836 14084 19892 14086
rect 19940 14138 19996 14140
rect 19940 14086 19942 14138
rect 19942 14086 19994 14138
rect 19994 14086 19996 14138
rect 19940 14084 19996 14086
rect 20044 14138 20100 14140
rect 20044 14086 20046 14138
rect 20046 14086 20098 14138
rect 20098 14086 20100 14138
rect 20044 14084 20100 14086
rect 18732 13970 18788 13972
rect 18732 13918 18734 13970
rect 18734 13918 18786 13970
rect 18786 13918 18788 13970
rect 18732 13916 18788 13918
rect 20076 13804 20132 13860
rect 19180 13634 19236 13636
rect 19180 13582 19182 13634
rect 19182 13582 19234 13634
rect 19234 13582 19236 13634
rect 19180 13580 19236 13582
rect 19068 13468 19124 13524
rect 19404 13522 19460 13524
rect 19404 13470 19406 13522
rect 19406 13470 19458 13522
rect 19458 13470 19460 13522
rect 19404 13468 19460 13470
rect 20076 13580 20132 13636
rect 19628 13074 19684 13076
rect 19628 13022 19630 13074
rect 19630 13022 19682 13074
rect 19682 13022 19684 13074
rect 19628 13020 19684 13022
rect 19180 12738 19236 12740
rect 19180 12686 19182 12738
rect 19182 12686 19234 12738
rect 19234 12686 19236 12738
rect 19180 12684 19236 12686
rect 18508 12066 18564 12068
rect 18508 12014 18510 12066
rect 18510 12014 18562 12066
rect 18562 12014 18564 12066
rect 18508 12012 18564 12014
rect 18732 12348 18788 12404
rect 17724 9212 17780 9268
rect 18396 9154 18452 9156
rect 18396 9102 18398 9154
rect 18398 9102 18450 9154
rect 18450 9102 18452 9154
rect 18396 9100 18452 9102
rect 17948 8764 18004 8820
rect 17836 8316 17892 8372
rect 17388 8092 17444 8148
rect 18956 11900 19012 11956
rect 19516 12066 19572 12068
rect 19516 12014 19518 12066
rect 19518 12014 19570 12066
rect 19570 12014 19572 12066
rect 19516 12012 19572 12014
rect 19516 11340 19572 11396
rect 20188 12684 20244 12740
rect 19836 12570 19892 12572
rect 19836 12518 19838 12570
rect 19838 12518 19890 12570
rect 19890 12518 19892 12570
rect 19836 12516 19892 12518
rect 19940 12570 19996 12572
rect 19940 12518 19942 12570
rect 19942 12518 19994 12570
rect 19994 12518 19996 12570
rect 19940 12516 19996 12518
rect 20044 12570 20100 12572
rect 20044 12518 20046 12570
rect 20046 12518 20098 12570
rect 20098 12518 20100 12570
rect 20044 12516 20100 12518
rect 20076 12402 20132 12404
rect 20076 12350 20078 12402
rect 20078 12350 20130 12402
rect 20130 12350 20132 12402
rect 20076 12348 20132 12350
rect 20188 11788 20244 11844
rect 20748 18620 20804 18676
rect 20748 16380 20804 16436
rect 20748 16210 20804 16212
rect 20748 16158 20750 16210
rect 20750 16158 20802 16210
rect 20802 16158 20804 16210
rect 20748 16156 20804 16158
rect 20412 15596 20468 15652
rect 20412 15260 20468 15316
rect 21644 21308 21700 21364
rect 20972 20130 21028 20132
rect 20972 20078 20974 20130
rect 20974 20078 21026 20130
rect 21026 20078 21028 20130
rect 20972 20076 21028 20078
rect 21308 19234 21364 19236
rect 21308 19182 21310 19234
rect 21310 19182 21362 19234
rect 21362 19182 21364 19234
rect 21308 19180 21364 19182
rect 21084 18450 21140 18452
rect 21084 18398 21086 18450
rect 21086 18398 21138 18450
rect 21138 18398 21140 18450
rect 21084 18396 21140 18398
rect 21980 20802 22036 20804
rect 21980 20750 21982 20802
rect 21982 20750 22034 20802
rect 22034 20750 22036 20802
rect 21980 20748 22036 20750
rect 21980 18956 22036 19012
rect 21532 18284 21588 18340
rect 21420 17948 21476 18004
rect 22764 25900 22820 25956
rect 23100 27916 23156 27972
rect 22988 27074 23044 27076
rect 22988 27022 22990 27074
rect 22990 27022 23042 27074
rect 23042 27022 23044 27074
rect 22988 27020 23044 27022
rect 22876 25788 22932 25844
rect 23772 30604 23828 30660
rect 23996 31500 24052 31556
rect 23996 30380 24052 30436
rect 24108 30492 24164 30548
rect 24556 32172 24612 32228
rect 24892 31836 24948 31892
rect 24556 31500 24612 31556
rect 25004 30940 25060 30996
rect 24780 30828 24836 30884
rect 24444 30268 24500 30324
rect 24556 30210 24612 30212
rect 24556 30158 24558 30210
rect 24558 30158 24610 30210
rect 24610 30158 24612 30210
rect 24556 30156 24612 30158
rect 24108 29260 24164 29316
rect 23436 28642 23492 28644
rect 23436 28590 23438 28642
rect 23438 28590 23490 28642
rect 23490 28590 23492 28642
rect 23436 28588 23492 28590
rect 23660 28588 23716 28644
rect 23436 27858 23492 27860
rect 23436 27806 23438 27858
rect 23438 27806 23490 27858
rect 23490 27806 23492 27858
rect 23436 27804 23492 27806
rect 23212 25900 23268 25956
rect 23548 26908 23604 26964
rect 23212 25228 23268 25284
rect 22876 23266 22932 23268
rect 22876 23214 22878 23266
rect 22878 23214 22930 23266
rect 22930 23214 22932 23266
rect 22876 23212 22932 23214
rect 22876 22204 22932 22260
rect 22428 21308 22484 21364
rect 22988 21756 23044 21812
rect 23436 23548 23492 23604
rect 23884 28924 23940 28980
rect 23996 28530 24052 28532
rect 23996 28478 23998 28530
rect 23998 28478 24050 28530
rect 24050 28478 24052 28530
rect 23996 28476 24052 28478
rect 23996 27244 24052 27300
rect 24444 27020 24500 27076
rect 24556 26962 24612 26964
rect 24556 26910 24558 26962
rect 24558 26910 24610 26962
rect 24610 26910 24612 26962
rect 24556 26908 24612 26910
rect 23772 26236 23828 26292
rect 23772 25676 23828 25732
rect 24444 26348 24500 26404
rect 24556 25564 24612 25620
rect 25340 41858 25396 41860
rect 25340 41806 25342 41858
rect 25342 41806 25394 41858
rect 25394 41806 25396 41858
rect 25340 41804 25396 41806
rect 25228 39452 25284 39508
rect 26348 41692 26404 41748
rect 26460 40572 26516 40628
rect 31724 44492 31780 44548
rect 31612 44380 31668 44436
rect 31948 43708 32004 43764
rect 30940 43596 30996 43652
rect 30268 42700 30324 42756
rect 26012 40124 26068 40180
rect 26124 39564 26180 39620
rect 26124 39340 26180 39396
rect 26796 39340 26852 39396
rect 29148 40402 29204 40404
rect 29148 40350 29150 40402
rect 29150 40350 29202 40402
rect 29202 40350 29204 40402
rect 29148 40348 29204 40350
rect 27244 39394 27300 39396
rect 27244 39342 27246 39394
rect 27246 39342 27298 39394
rect 27298 39342 27300 39394
rect 27244 39340 27300 39342
rect 28588 40178 28644 40180
rect 28588 40126 28590 40178
rect 28590 40126 28642 40178
rect 28642 40126 28644 40178
rect 28588 40124 28644 40126
rect 29260 39564 29316 39620
rect 28476 39340 28532 39396
rect 29260 39394 29316 39396
rect 29260 39342 29262 39394
rect 29262 39342 29314 39394
rect 29314 39342 29316 39394
rect 29260 39340 29316 39342
rect 29932 40402 29988 40404
rect 29932 40350 29934 40402
rect 29934 40350 29986 40402
rect 29986 40350 29988 40402
rect 29932 40348 29988 40350
rect 27020 39228 27076 39284
rect 29036 39228 29092 39284
rect 26012 37996 26068 38052
rect 25340 37324 25396 37380
rect 27692 38668 27748 38724
rect 29820 39228 29876 39284
rect 29484 38722 29540 38724
rect 29484 38670 29486 38722
rect 29486 38670 29538 38722
rect 29538 38670 29540 38722
rect 29484 38668 29540 38670
rect 28028 36594 28084 36596
rect 28028 36542 28030 36594
rect 28030 36542 28082 36594
rect 28082 36542 28084 36594
rect 28028 36540 28084 36542
rect 26124 36204 26180 36260
rect 25900 35532 25956 35588
rect 27244 36258 27300 36260
rect 27244 36206 27246 36258
rect 27246 36206 27298 36258
rect 27298 36206 27300 36258
rect 27244 36204 27300 36206
rect 26124 35196 26180 35252
rect 30380 39564 30436 39620
rect 30044 38892 30100 38948
rect 31836 42700 31892 42756
rect 31612 42476 31668 42532
rect 31276 41244 31332 41300
rect 30492 39004 30548 39060
rect 30380 38668 30436 38724
rect 29484 36764 29540 36820
rect 29484 36540 29540 36596
rect 29820 36594 29876 36596
rect 29820 36542 29822 36594
rect 29822 36542 29874 36594
rect 29874 36542 29876 36594
rect 29820 36540 29876 36542
rect 29260 36482 29316 36484
rect 29260 36430 29262 36482
rect 29262 36430 29314 36482
rect 29314 36430 29316 36482
rect 29260 36428 29316 36430
rect 26460 34802 26516 34804
rect 26460 34750 26462 34802
rect 26462 34750 26514 34802
rect 26514 34750 26516 34802
rect 26460 34748 26516 34750
rect 25340 34300 25396 34356
rect 25788 34076 25844 34132
rect 25452 33180 25508 33236
rect 26012 34018 26068 34020
rect 26012 33966 26014 34018
rect 26014 33966 26066 34018
rect 26066 33966 26068 34018
rect 26012 33964 26068 33966
rect 25340 33122 25396 33124
rect 25340 33070 25342 33122
rect 25342 33070 25394 33122
rect 25394 33070 25396 33122
rect 25340 33068 25396 33070
rect 25340 30994 25396 30996
rect 25340 30942 25342 30994
rect 25342 30942 25394 30994
rect 25394 30942 25396 30994
rect 25340 30940 25396 30942
rect 25340 30268 25396 30324
rect 26236 32396 26292 32452
rect 28028 34972 28084 35028
rect 29148 34972 29204 35028
rect 26572 31836 26628 31892
rect 25788 31778 25844 31780
rect 25788 31726 25790 31778
rect 25790 31726 25842 31778
rect 25842 31726 25844 31778
rect 25788 31724 25844 31726
rect 26012 30882 26068 30884
rect 26012 30830 26014 30882
rect 26014 30830 26066 30882
rect 26066 30830 26068 30882
rect 26012 30828 26068 30830
rect 28140 34748 28196 34804
rect 28812 34242 28868 34244
rect 28812 34190 28814 34242
rect 28814 34190 28866 34242
rect 28866 34190 28868 34242
rect 28812 34188 28868 34190
rect 28364 33852 28420 33908
rect 27916 31890 27972 31892
rect 27916 31838 27918 31890
rect 27918 31838 27970 31890
rect 27970 31838 27972 31890
rect 27916 31836 27972 31838
rect 26908 30492 26964 30548
rect 28140 30492 28196 30548
rect 25452 29820 25508 29876
rect 26236 29932 26292 29988
rect 25900 29484 25956 29540
rect 26236 28642 26292 28644
rect 26236 28590 26238 28642
rect 26238 28590 26290 28642
rect 26290 28590 26292 28642
rect 26236 28588 26292 28590
rect 25788 28476 25844 28532
rect 25788 27916 25844 27972
rect 26572 28588 26628 28644
rect 26908 29986 26964 29988
rect 26908 29934 26910 29986
rect 26910 29934 26962 29986
rect 26962 29934 26964 29986
rect 26908 29932 26964 29934
rect 27132 29986 27188 29988
rect 27132 29934 27134 29986
rect 27134 29934 27186 29986
rect 27186 29934 27188 29986
rect 27132 29932 27188 29934
rect 27020 29538 27076 29540
rect 27020 29486 27022 29538
rect 27022 29486 27074 29538
rect 27074 29486 27076 29538
rect 27020 29484 27076 29486
rect 27692 29538 27748 29540
rect 27692 29486 27694 29538
rect 27694 29486 27746 29538
rect 27746 29486 27748 29538
rect 27692 29484 27748 29486
rect 26908 28530 26964 28532
rect 26908 28478 26910 28530
rect 26910 28478 26962 28530
rect 26962 28478 26964 28530
rect 26908 28476 26964 28478
rect 27468 28530 27524 28532
rect 27468 28478 27470 28530
rect 27470 28478 27522 28530
rect 27522 28478 27524 28530
rect 27468 28476 27524 28478
rect 26124 25618 26180 25620
rect 26124 25566 26126 25618
rect 26126 25566 26178 25618
rect 26178 25566 26180 25618
rect 26124 25564 26180 25566
rect 24332 23548 24388 23604
rect 24220 23212 24276 23268
rect 23660 22930 23716 22932
rect 23660 22878 23662 22930
rect 23662 22878 23714 22930
rect 23714 22878 23716 22930
rect 23660 22876 23716 22878
rect 23436 22652 23492 22708
rect 23100 21586 23156 21588
rect 23100 21534 23102 21586
rect 23102 21534 23154 21586
rect 23154 21534 23156 21586
rect 23100 21532 23156 21534
rect 23212 21756 23268 21812
rect 22764 20748 22820 20804
rect 22988 20860 23044 20916
rect 23660 21308 23716 21364
rect 24332 23100 24388 23156
rect 24220 21308 24276 21364
rect 23996 20914 24052 20916
rect 23996 20862 23998 20914
rect 23998 20862 24050 20914
rect 24050 20862 24052 20914
rect 23996 20860 24052 20862
rect 23212 20802 23268 20804
rect 23212 20750 23214 20802
rect 23214 20750 23266 20802
rect 23266 20750 23268 20802
rect 23212 20748 23268 20750
rect 23100 20188 23156 20244
rect 22652 18508 22708 18564
rect 22092 17612 22148 17668
rect 21980 17500 22036 17556
rect 22092 17052 22148 17108
rect 22540 17276 22596 17332
rect 22316 16882 22372 16884
rect 22316 16830 22318 16882
rect 22318 16830 22370 16882
rect 22370 16830 22372 16882
rect 22316 16828 22372 16830
rect 21868 16716 21924 16772
rect 21756 16210 21812 16212
rect 21756 16158 21758 16210
rect 21758 16158 21810 16210
rect 21810 16158 21812 16210
rect 21756 16156 21812 16158
rect 21644 15932 21700 15988
rect 22204 16716 22260 16772
rect 22876 16658 22932 16660
rect 22876 16606 22878 16658
rect 22878 16606 22930 16658
rect 22930 16606 22932 16658
rect 22876 16604 22932 16606
rect 22204 16044 22260 16100
rect 22428 16380 22484 16436
rect 21084 15484 21140 15540
rect 19836 11002 19892 11004
rect 19836 10950 19838 11002
rect 19838 10950 19890 11002
rect 19890 10950 19892 11002
rect 19836 10948 19892 10950
rect 19940 11002 19996 11004
rect 19940 10950 19942 11002
rect 19942 10950 19994 11002
rect 19994 10950 19996 11002
rect 19940 10948 19996 10950
rect 20044 11002 20100 11004
rect 20044 10950 20046 11002
rect 20046 10950 20098 11002
rect 20098 10950 20100 11002
rect 20044 10948 20100 10950
rect 20636 14588 20692 14644
rect 20636 13916 20692 13972
rect 20636 13468 20692 13524
rect 20636 12572 20692 12628
rect 21196 14588 21252 14644
rect 24108 20188 24164 20244
rect 23436 18396 23492 18452
rect 23996 18620 24052 18676
rect 23884 18338 23940 18340
rect 23884 18286 23886 18338
rect 23886 18286 23938 18338
rect 23938 18286 23940 18338
rect 23884 18284 23940 18286
rect 23772 17106 23828 17108
rect 23772 17054 23774 17106
rect 23774 17054 23826 17106
rect 23826 17054 23828 17106
rect 23772 17052 23828 17054
rect 23324 16940 23380 16996
rect 23212 15986 23268 15988
rect 23212 15934 23214 15986
rect 23214 15934 23266 15986
rect 23266 15934 23268 15986
rect 23212 15932 23268 15934
rect 22764 15596 22820 15652
rect 21868 15484 21924 15540
rect 21308 14476 21364 14532
rect 20188 9884 20244 9940
rect 19628 9548 19684 9604
rect 18844 9266 18900 9268
rect 18844 9214 18846 9266
rect 18846 9214 18898 9266
rect 18898 9214 18900 9266
rect 18844 9212 18900 9214
rect 20188 9602 20244 9604
rect 20188 9550 20190 9602
rect 20190 9550 20242 9602
rect 20242 9550 20244 9602
rect 20188 9548 20244 9550
rect 19836 9434 19892 9436
rect 19836 9382 19838 9434
rect 19838 9382 19890 9434
rect 19890 9382 19892 9434
rect 19836 9380 19892 9382
rect 19940 9434 19996 9436
rect 19940 9382 19942 9434
rect 19942 9382 19994 9434
rect 19994 9382 19996 9434
rect 19940 9380 19996 9382
rect 20044 9434 20100 9436
rect 20044 9382 20046 9434
rect 20046 9382 20098 9434
rect 20098 9382 20100 9434
rect 20044 9380 20100 9382
rect 20188 9042 20244 9044
rect 20188 8990 20190 9042
rect 20190 8990 20242 9042
rect 20242 8990 20244 9042
rect 20188 8988 20244 8990
rect 18732 8092 18788 8148
rect 16828 7756 16884 7812
rect 17052 7644 17108 7700
rect 17500 7756 17556 7812
rect 18844 8034 18900 8036
rect 18844 7982 18846 8034
rect 18846 7982 18898 8034
rect 18898 7982 18900 8034
rect 18844 7980 18900 7982
rect 20748 11340 20804 11396
rect 21980 13580 22036 13636
rect 22540 14476 22596 14532
rect 21868 13020 21924 13076
rect 21980 12236 22036 12292
rect 22764 12572 22820 12628
rect 22764 12402 22820 12404
rect 22764 12350 22766 12402
rect 22766 12350 22818 12402
rect 22818 12350 22820 12402
rect 22764 12348 22820 12350
rect 21196 9660 21252 9716
rect 22428 10444 22484 10500
rect 23884 16828 23940 16884
rect 23660 16604 23716 16660
rect 23660 16098 23716 16100
rect 23660 16046 23662 16098
rect 23662 16046 23714 16098
rect 23714 16046 23716 16098
rect 23660 16044 23716 16046
rect 24220 18450 24276 18452
rect 24220 18398 24222 18450
rect 24222 18398 24274 18450
rect 24274 18398 24276 18450
rect 24220 18396 24276 18398
rect 24332 18338 24388 18340
rect 24332 18286 24334 18338
rect 24334 18286 24386 18338
rect 24386 18286 24388 18338
rect 24332 18284 24388 18286
rect 25228 23436 25284 23492
rect 25340 23100 25396 23156
rect 25452 23436 25508 23492
rect 25564 23212 25620 23268
rect 25676 23154 25732 23156
rect 25676 23102 25678 23154
rect 25678 23102 25730 23154
rect 25730 23102 25732 23154
rect 25676 23100 25732 23102
rect 26012 22540 26068 22596
rect 26684 27804 26740 27860
rect 26460 27186 26516 27188
rect 26460 27134 26462 27186
rect 26462 27134 26514 27186
rect 26514 27134 26516 27186
rect 26460 27132 26516 27134
rect 27356 27858 27412 27860
rect 27356 27806 27358 27858
rect 27358 27806 27410 27858
rect 27410 27806 27412 27858
rect 27356 27804 27412 27806
rect 27132 27132 27188 27188
rect 27804 26402 27860 26404
rect 27804 26350 27806 26402
rect 27806 26350 27858 26402
rect 27858 26350 27860 26402
rect 27804 26348 27860 26350
rect 27468 26290 27524 26292
rect 27468 26238 27470 26290
rect 27470 26238 27522 26290
rect 27522 26238 27524 26290
rect 27468 26236 27524 26238
rect 27020 26066 27076 26068
rect 27020 26014 27022 26066
rect 27022 26014 27074 26066
rect 27074 26014 27076 26066
rect 27020 26012 27076 26014
rect 26796 23996 26852 24052
rect 26572 23324 26628 23380
rect 27804 24050 27860 24052
rect 27804 23998 27806 24050
rect 27806 23998 27858 24050
rect 27858 23998 27860 24050
rect 27804 23996 27860 23998
rect 27580 23266 27636 23268
rect 27580 23214 27582 23266
rect 27582 23214 27634 23266
rect 27634 23214 27636 23266
rect 27580 23212 27636 23214
rect 28588 33292 28644 33348
rect 29260 33964 29316 34020
rect 28588 33122 28644 33124
rect 28588 33070 28590 33122
rect 28590 33070 28642 33122
rect 28642 33070 28644 33122
rect 28588 33068 28644 33070
rect 28588 31724 28644 31780
rect 28588 30156 28644 30212
rect 28588 29372 28644 29428
rect 28588 26348 28644 26404
rect 29932 34802 29988 34804
rect 29932 34750 29934 34802
rect 29934 34750 29986 34802
rect 29986 34750 29988 34802
rect 29932 34748 29988 34750
rect 29932 34188 29988 34244
rect 29372 33068 29428 33124
rect 29148 31778 29204 31780
rect 29148 31726 29150 31778
rect 29150 31726 29202 31778
rect 29202 31726 29204 31778
rect 29148 31724 29204 31726
rect 29596 31164 29652 31220
rect 29260 29932 29316 29988
rect 29596 29986 29652 29988
rect 29596 29934 29598 29986
rect 29598 29934 29650 29986
rect 29650 29934 29652 29986
rect 29596 29932 29652 29934
rect 29484 29372 29540 29428
rect 29596 29036 29652 29092
rect 30828 35644 30884 35700
rect 30268 34018 30324 34020
rect 30268 33966 30270 34018
rect 30270 33966 30322 34018
rect 30322 33966 30324 34018
rect 30268 33964 30324 33966
rect 31052 38946 31108 38948
rect 31052 38894 31054 38946
rect 31054 38894 31106 38946
rect 31106 38894 31108 38946
rect 31052 38892 31108 38894
rect 31388 38556 31444 38612
rect 31948 39676 32004 39732
rect 31836 39058 31892 39060
rect 31836 39006 31838 39058
rect 31838 39006 31890 39058
rect 31890 39006 31892 39058
rect 31836 39004 31892 39006
rect 31276 36764 31332 36820
rect 31612 36482 31668 36484
rect 31612 36430 31614 36482
rect 31614 36430 31666 36482
rect 31666 36430 31668 36482
rect 31612 36428 31668 36430
rect 31388 36204 31444 36260
rect 31612 35698 31668 35700
rect 31612 35646 31614 35698
rect 31614 35646 31666 35698
rect 31666 35646 31668 35698
rect 31612 35644 31668 35646
rect 31164 33292 31220 33348
rect 31052 31836 31108 31892
rect 30716 31218 30772 31220
rect 30716 31166 30718 31218
rect 30718 31166 30770 31218
rect 30770 31166 30772 31218
rect 30716 31164 30772 31166
rect 30044 29036 30100 29092
rect 29708 28812 29764 28868
rect 31388 34860 31444 34916
rect 32172 43596 32228 43652
rect 32956 46956 33012 47012
rect 33180 46114 33236 46116
rect 33180 46062 33182 46114
rect 33182 46062 33234 46114
rect 33234 46062 33236 46114
rect 33180 46060 33236 46062
rect 33068 44380 33124 44436
rect 33180 44156 33236 44212
rect 36988 46956 37044 47012
rect 35196 46282 35252 46284
rect 35196 46230 35198 46282
rect 35198 46230 35250 46282
rect 35250 46230 35252 46282
rect 35196 46228 35252 46230
rect 35300 46282 35356 46284
rect 35300 46230 35302 46282
rect 35302 46230 35354 46282
rect 35354 46230 35356 46282
rect 35300 46228 35356 46230
rect 35404 46282 35460 46284
rect 35404 46230 35406 46282
rect 35406 46230 35458 46282
rect 35458 46230 35460 46282
rect 35404 46228 35460 46230
rect 35196 45276 35252 45332
rect 33964 45106 34020 45108
rect 33964 45054 33966 45106
rect 33966 45054 34018 45106
rect 34018 45054 34020 45106
rect 33964 45052 34020 45054
rect 35420 44828 35476 44884
rect 35196 44714 35252 44716
rect 35196 44662 35198 44714
rect 35198 44662 35250 44714
rect 35250 44662 35252 44714
rect 35196 44660 35252 44662
rect 35300 44714 35356 44716
rect 35300 44662 35302 44714
rect 35302 44662 35354 44714
rect 35354 44662 35356 44714
rect 35300 44660 35356 44662
rect 35404 44714 35460 44716
rect 35404 44662 35406 44714
rect 35406 44662 35458 44714
rect 35458 44662 35460 44714
rect 35404 44660 35460 44662
rect 33292 44380 33348 44436
rect 32284 43372 32340 43428
rect 32508 42924 32564 42980
rect 32284 41916 32340 41972
rect 32284 41298 32340 41300
rect 32284 41246 32286 41298
rect 32286 41246 32338 41298
rect 32338 41246 32340 41298
rect 32284 41244 32340 41246
rect 32732 39676 32788 39732
rect 32284 38668 32340 38724
rect 32172 38556 32228 38612
rect 32172 37436 32228 37492
rect 32620 35868 32676 35924
rect 32060 35644 32116 35700
rect 32060 34748 32116 34804
rect 32060 33852 32116 33908
rect 33628 41020 33684 41076
rect 33516 40796 33572 40852
rect 33404 38834 33460 38836
rect 33404 38782 33406 38834
rect 33406 38782 33458 38834
rect 33458 38782 33460 38834
rect 33404 38780 33460 38782
rect 33292 38556 33348 38612
rect 34524 44546 34580 44548
rect 34524 44494 34526 44546
rect 34526 44494 34578 44546
rect 34578 44494 34580 44546
rect 34524 44492 34580 44494
rect 33964 43596 34020 43652
rect 34412 43708 34468 43764
rect 34076 43426 34132 43428
rect 34076 43374 34078 43426
rect 34078 43374 34130 43426
rect 34130 43374 34132 43426
rect 34076 43372 34132 43374
rect 34188 42530 34244 42532
rect 34188 42478 34190 42530
rect 34190 42478 34242 42530
rect 34242 42478 34244 42530
rect 34188 42476 34244 42478
rect 34300 41074 34356 41076
rect 34300 41022 34302 41074
rect 34302 41022 34354 41074
rect 34354 41022 34356 41074
rect 34300 41020 34356 41022
rect 35196 43146 35252 43148
rect 35196 43094 35198 43146
rect 35198 43094 35250 43146
rect 35250 43094 35252 43146
rect 35196 43092 35252 43094
rect 35300 43146 35356 43148
rect 35300 43094 35302 43146
rect 35302 43094 35354 43146
rect 35354 43094 35356 43146
rect 35300 43092 35356 43094
rect 35404 43146 35460 43148
rect 35404 43094 35406 43146
rect 35406 43094 35458 43146
rect 35458 43094 35460 43146
rect 35404 43092 35460 43094
rect 34524 42978 34580 42980
rect 34524 42926 34526 42978
rect 34526 42926 34578 42978
rect 34578 42926 34580 42978
rect 34524 42924 34580 42926
rect 35084 42700 35140 42756
rect 34636 41804 34692 41860
rect 34748 40796 34804 40852
rect 33964 40236 34020 40292
rect 33964 40012 34020 40068
rect 34076 38834 34132 38836
rect 34076 38782 34078 38834
rect 34078 38782 34130 38834
rect 34130 38782 34132 38834
rect 34076 38780 34132 38782
rect 34972 40572 35028 40628
rect 34860 40124 34916 40180
rect 36316 45052 36372 45108
rect 35980 44156 36036 44212
rect 35868 41916 35924 41972
rect 35980 41858 36036 41860
rect 35980 41806 35982 41858
rect 35982 41806 36034 41858
rect 36034 41806 36036 41858
rect 35980 41804 36036 41806
rect 35196 41578 35252 41580
rect 35196 41526 35198 41578
rect 35198 41526 35250 41578
rect 35250 41526 35252 41578
rect 35196 41524 35252 41526
rect 35300 41578 35356 41580
rect 35300 41526 35302 41578
rect 35302 41526 35354 41578
rect 35354 41526 35356 41578
rect 35300 41524 35356 41526
rect 35404 41578 35460 41580
rect 35404 41526 35406 41578
rect 35406 41526 35458 41578
rect 35458 41526 35460 41578
rect 35404 41524 35460 41526
rect 37324 45836 37380 45892
rect 37100 45106 37156 45108
rect 37100 45054 37102 45106
rect 37102 45054 37154 45106
rect 37154 45054 37156 45106
rect 37100 45052 37156 45054
rect 37100 44434 37156 44436
rect 37100 44382 37102 44434
rect 37102 44382 37154 44434
rect 37154 44382 37156 44434
rect 37100 44380 37156 44382
rect 36764 43484 36820 43540
rect 36988 43596 37044 43652
rect 36428 42924 36484 42980
rect 37212 42978 37268 42980
rect 37212 42926 37214 42978
rect 37214 42926 37266 42978
rect 37266 42926 37268 42978
rect 37212 42924 37268 42926
rect 36204 41356 36260 41412
rect 36204 41186 36260 41188
rect 36204 41134 36206 41186
rect 36206 41134 36258 41186
rect 36258 41134 36260 41186
rect 36204 41132 36260 41134
rect 35196 40796 35252 40852
rect 35196 40236 35252 40292
rect 35196 40010 35252 40012
rect 35196 39958 35198 40010
rect 35198 39958 35250 40010
rect 35250 39958 35252 40010
rect 35196 39956 35252 39958
rect 35300 40010 35356 40012
rect 35300 39958 35302 40010
rect 35302 39958 35354 40010
rect 35354 39958 35356 40010
rect 35300 39956 35356 39958
rect 35404 40010 35460 40012
rect 35404 39958 35406 40010
rect 35406 39958 35458 40010
rect 35458 39958 35460 40010
rect 35404 39956 35460 39958
rect 36428 40962 36484 40964
rect 36428 40910 36430 40962
rect 36430 40910 36482 40962
rect 36482 40910 36484 40962
rect 36428 40908 36484 40910
rect 36316 40626 36372 40628
rect 36316 40574 36318 40626
rect 36318 40574 36370 40626
rect 36370 40574 36372 40626
rect 36316 40572 36372 40574
rect 35644 40514 35700 40516
rect 35644 40462 35646 40514
rect 35646 40462 35698 40514
rect 35698 40462 35700 40514
rect 35644 40460 35700 40462
rect 37212 41410 37268 41412
rect 37212 41358 37214 41410
rect 37214 41358 37266 41410
rect 37266 41358 37268 41410
rect 37212 41356 37268 41358
rect 35868 39676 35924 39732
rect 34524 39004 34580 39060
rect 34412 38556 34468 38612
rect 33292 35922 33348 35924
rect 33292 35870 33294 35922
rect 33294 35870 33346 35922
rect 33346 35870 33348 35922
rect 33292 35868 33348 35870
rect 33404 34802 33460 34804
rect 33404 34750 33406 34802
rect 33406 34750 33458 34802
rect 33458 34750 33460 34802
rect 33404 34748 33460 34750
rect 32956 33404 33012 33460
rect 32284 32674 32340 32676
rect 32284 32622 32286 32674
rect 32286 32622 32338 32674
rect 32338 32622 32340 32674
rect 32284 32620 32340 32622
rect 31388 31106 31444 31108
rect 31388 31054 31390 31106
rect 31390 31054 31442 31106
rect 31442 31054 31444 31106
rect 31388 31052 31444 31054
rect 32060 31890 32116 31892
rect 32060 31838 32062 31890
rect 32062 31838 32114 31890
rect 32114 31838 32116 31890
rect 32060 31836 32116 31838
rect 32396 31778 32452 31780
rect 32396 31726 32398 31778
rect 32398 31726 32450 31778
rect 32450 31726 32452 31778
rect 32396 31724 32452 31726
rect 31276 29484 31332 29540
rect 30716 28866 30772 28868
rect 30716 28814 30718 28866
rect 30718 28814 30770 28866
rect 30770 28814 30772 28866
rect 30716 28812 30772 28814
rect 30268 28754 30324 28756
rect 30268 28702 30270 28754
rect 30270 28702 30322 28754
rect 30322 28702 30324 28754
rect 30268 28700 30324 28702
rect 31836 30044 31892 30100
rect 33516 34018 33572 34020
rect 33516 33966 33518 34018
rect 33518 33966 33570 34018
rect 33570 33966 33572 34018
rect 33516 33964 33572 33966
rect 34860 36204 34916 36260
rect 35196 38556 35252 38612
rect 35196 38442 35252 38444
rect 35196 38390 35198 38442
rect 35198 38390 35250 38442
rect 35250 38390 35252 38442
rect 35196 38388 35252 38390
rect 35300 38442 35356 38444
rect 35300 38390 35302 38442
rect 35302 38390 35354 38442
rect 35354 38390 35356 38442
rect 35300 38388 35356 38390
rect 35404 38442 35460 38444
rect 35404 38390 35406 38442
rect 35406 38390 35458 38442
rect 35458 38390 35460 38442
rect 35404 38388 35460 38390
rect 35420 37490 35476 37492
rect 35420 37438 35422 37490
rect 35422 37438 35474 37490
rect 35474 37438 35476 37490
rect 35420 37436 35476 37438
rect 35196 36874 35252 36876
rect 35196 36822 35198 36874
rect 35198 36822 35250 36874
rect 35250 36822 35252 36874
rect 35196 36820 35252 36822
rect 35300 36874 35356 36876
rect 35300 36822 35302 36874
rect 35302 36822 35354 36874
rect 35354 36822 35356 36874
rect 35300 36820 35356 36822
rect 35404 36874 35460 36876
rect 35404 36822 35406 36874
rect 35406 36822 35458 36874
rect 35458 36822 35460 36874
rect 35404 36820 35460 36822
rect 35308 36428 35364 36484
rect 35196 35306 35252 35308
rect 35196 35254 35198 35306
rect 35198 35254 35250 35306
rect 35250 35254 35252 35306
rect 35196 35252 35252 35254
rect 35300 35306 35356 35308
rect 35300 35254 35302 35306
rect 35302 35254 35354 35306
rect 35354 35254 35356 35306
rect 35300 35252 35356 35254
rect 35404 35306 35460 35308
rect 35404 35254 35406 35306
rect 35406 35254 35458 35306
rect 35458 35254 35460 35306
rect 35404 35252 35460 35254
rect 33852 33852 33908 33908
rect 33404 33458 33460 33460
rect 33404 33406 33406 33458
rect 33406 33406 33458 33458
rect 33458 33406 33460 33458
rect 33404 33404 33460 33406
rect 35532 34748 35588 34804
rect 34860 34690 34916 34692
rect 34860 34638 34862 34690
rect 34862 34638 34914 34690
rect 34914 34638 34916 34690
rect 34860 34636 34916 34638
rect 35532 33852 35588 33908
rect 35196 33738 35252 33740
rect 35196 33686 35198 33738
rect 35198 33686 35250 33738
rect 35250 33686 35252 33738
rect 35196 33684 35252 33686
rect 35300 33738 35356 33740
rect 35300 33686 35302 33738
rect 35302 33686 35354 33738
rect 35354 33686 35356 33738
rect 35300 33684 35356 33686
rect 35404 33738 35460 33740
rect 35404 33686 35406 33738
rect 35406 33686 35458 33738
rect 35458 33686 35460 33738
rect 35404 33684 35460 33686
rect 33964 33292 34020 33348
rect 35196 33346 35252 33348
rect 35196 33294 35198 33346
rect 35198 33294 35250 33346
rect 35250 33294 35252 33346
rect 35196 33292 35252 33294
rect 33964 32620 34020 32676
rect 35532 33180 35588 33236
rect 35196 32170 35252 32172
rect 35196 32118 35198 32170
rect 35198 32118 35250 32170
rect 35250 32118 35252 32170
rect 35196 32116 35252 32118
rect 35300 32170 35356 32172
rect 35300 32118 35302 32170
rect 35302 32118 35354 32170
rect 35354 32118 35356 32170
rect 35300 32116 35356 32118
rect 35404 32170 35460 32172
rect 35404 32118 35406 32170
rect 35406 32118 35458 32170
rect 35458 32118 35460 32170
rect 35404 32116 35460 32118
rect 32732 28924 32788 28980
rect 31836 28700 31892 28756
rect 34636 31612 34692 31668
rect 35308 31612 35364 31668
rect 34860 31106 34916 31108
rect 34860 31054 34862 31106
rect 34862 31054 34914 31106
rect 34914 31054 34916 31106
rect 34860 31052 34916 31054
rect 37660 45164 37716 45220
rect 37884 45612 37940 45668
rect 37772 45052 37828 45108
rect 39788 45890 39844 45892
rect 39788 45838 39790 45890
rect 39790 45838 39842 45890
rect 39842 45838 39844 45890
rect 39788 45836 39844 45838
rect 38892 45666 38948 45668
rect 38892 45614 38894 45666
rect 38894 45614 38946 45666
rect 38946 45614 38948 45666
rect 38892 45612 38948 45614
rect 38332 45052 38388 45108
rect 39004 44828 39060 44884
rect 38556 43596 38612 43652
rect 38668 43820 38724 43876
rect 37548 41916 37604 41972
rect 39228 44492 39284 44548
rect 40012 43932 40068 43988
rect 39564 43708 39620 43764
rect 39340 43538 39396 43540
rect 39340 43486 39342 43538
rect 39342 43486 39394 43538
rect 39394 43486 39396 43538
rect 39340 43484 39396 43486
rect 39228 41916 39284 41972
rect 39228 41692 39284 41748
rect 39676 41970 39732 41972
rect 39676 41918 39678 41970
rect 39678 41918 39730 41970
rect 39730 41918 39732 41970
rect 39676 41916 39732 41918
rect 37436 40908 37492 40964
rect 38220 41074 38276 41076
rect 38220 41022 38222 41074
rect 38222 41022 38274 41074
rect 38274 41022 38276 41074
rect 38220 41020 38276 41022
rect 37772 40460 37828 40516
rect 37324 40124 37380 40180
rect 37772 40124 37828 40180
rect 36428 39730 36484 39732
rect 36428 39678 36430 39730
rect 36430 39678 36482 39730
rect 36482 39678 36484 39730
rect 36428 39676 36484 39678
rect 37100 39730 37156 39732
rect 37100 39678 37102 39730
rect 37102 39678 37154 39730
rect 37154 39678 37156 39730
rect 37100 39676 37156 39678
rect 38892 41186 38948 41188
rect 38892 41134 38894 41186
rect 38894 41134 38946 41186
rect 38946 41134 38948 41186
rect 38892 41132 38948 41134
rect 40796 45276 40852 45332
rect 42028 45164 42084 45220
rect 40684 44434 40740 44436
rect 40684 44382 40686 44434
rect 40686 44382 40738 44434
rect 40738 44382 40740 44434
rect 40684 44380 40740 44382
rect 39900 41804 39956 41860
rect 40124 41858 40180 41860
rect 40124 41806 40126 41858
rect 40126 41806 40178 41858
rect 40178 41806 40180 41858
rect 40124 41804 40180 41806
rect 39228 41020 39284 41076
rect 39340 40572 39396 40628
rect 38780 40348 38836 40404
rect 38668 39842 38724 39844
rect 38668 39790 38670 39842
rect 38670 39790 38722 39842
rect 38722 39790 38724 39842
rect 38668 39788 38724 39790
rect 38108 38892 38164 38948
rect 36204 37884 36260 37940
rect 37548 38668 37604 38724
rect 38668 38722 38724 38724
rect 38668 38670 38670 38722
rect 38670 38670 38722 38722
rect 38722 38670 38724 38722
rect 38668 38668 38724 38670
rect 37772 38556 37828 38612
rect 37212 37938 37268 37940
rect 37212 37886 37214 37938
rect 37214 37886 37266 37938
rect 37266 37886 37268 37938
rect 37212 37884 37268 37886
rect 36316 36482 36372 36484
rect 36316 36430 36318 36482
rect 36318 36430 36370 36482
rect 36370 36430 36372 36482
rect 36316 36428 36372 36430
rect 35756 36258 35812 36260
rect 35756 36206 35758 36258
rect 35758 36206 35810 36258
rect 35810 36206 35812 36258
rect 35756 36204 35812 36206
rect 36092 34636 36148 34692
rect 35756 33964 35812 34020
rect 35980 33234 36036 33236
rect 35980 33182 35982 33234
rect 35982 33182 36034 33234
rect 36034 33182 36036 33234
rect 35980 33180 36036 33182
rect 35756 32620 35812 32676
rect 35196 30602 35252 30604
rect 35196 30550 35198 30602
rect 35198 30550 35250 30602
rect 35250 30550 35252 30602
rect 35196 30548 35252 30550
rect 35300 30602 35356 30604
rect 35300 30550 35302 30602
rect 35302 30550 35354 30602
rect 35354 30550 35356 30602
rect 35300 30548 35356 30550
rect 35404 30602 35460 30604
rect 35404 30550 35406 30602
rect 35406 30550 35458 30602
rect 35458 30550 35460 30602
rect 35404 30548 35460 30550
rect 33180 29932 33236 29988
rect 33068 29148 33124 29204
rect 34524 29986 34580 29988
rect 34524 29934 34526 29986
rect 34526 29934 34578 29986
rect 34578 29934 34580 29986
rect 34524 29932 34580 29934
rect 34076 29708 34132 29764
rect 33404 29260 33460 29316
rect 32844 28476 32900 28532
rect 35196 29314 35252 29316
rect 35196 29262 35198 29314
rect 35198 29262 35250 29314
rect 35250 29262 35252 29314
rect 35196 29260 35252 29262
rect 35644 29708 35700 29764
rect 35980 29426 36036 29428
rect 35980 29374 35982 29426
rect 35982 29374 36034 29426
rect 36034 29374 36036 29426
rect 35980 29372 36036 29374
rect 35420 29260 35476 29316
rect 34860 29148 34916 29204
rect 35196 29034 35252 29036
rect 35196 28982 35198 29034
rect 35198 28982 35250 29034
rect 35250 28982 35252 29034
rect 35196 28980 35252 28982
rect 35300 29034 35356 29036
rect 35300 28982 35302 29034
rect 35302 28982 35354 29034
rect 35354 28982 35356 29034
rect 35300 28980 35356 28982
rect 35404 29034 35460 29036
rect 35404 28982 35406 29034
rect 35406 28982 35458 29034
rect 35458 28982 35460 29034
rect 35404 28980 35460 28982
rect 32396 27244 32452 27300
rect 31612 27020 31668 27076
rect 29484 26348 29540 26404
rect 28588 23938 28644 23940
rect 28588 23886 28590 23938
rect 28590 23886 28642 23938
rect 28642 23886 28644 23938
rect 28588 23884 28644 23886
rect 29372 25506 29428 25508
rect 29372 25454 29374 25506
rect 29374 25454 29426 25506
rect 29426 25454 29428 25506
rect 29372 25452 29428 25454
rect 29260 24668 29316 24724
rect 28700 23548 28756 23604
rect 29372 23884 29428 23940
rect 35196 27466 35252 27468
rect 35196 27414 35198 27466
rect 35198 27414 35250 27466
rect 35250 27414 35252 27466
rect 35196 27412 35252 27414
rect 35300 27466 35356 27468
rect 35300 27414 35302 27466
rect 35302 27414 35354 27466
rect 35354 27414 35356 27466
rect 35300 27412 35356 27414
rect 35404 27466 35460 27468
rect 35404 27414 35406 27466
rect 35406 27414 35458 27466
rect 35458 27414 35460 27466
rect 35404 27412 35460 27414
rect 35868 27020 35924 27076
rect 30380 25564 30436 25620
rect 30044 24892 30100 24948
rect 29036 23436 29092 23492
rect 29372 23378 29428 23380
rect 29372 23326 29374 23378
rect 29374 23326 29426 23378
rect 29426 23326 29428 23378
rect 29372 23324 29428 23326
rect 29484 23266 29540 23268
rect 29484 23214 29486 23266
rect 29486 23214 29538 23266
rect 29538 23214 29540 23266
rect 29484 23212 29540 23214
rect 28364 22764 28420 22820
rect 26348 22652 26404 22708
rect 23436 15932 23492 15988
rect 24332 15986 24388 15988
rect 24332 15934 24334 15986
rect 24334 15934 24386 15986
rect 24386 15934 24388 15986
rect 24332 15932 24388 15934
rect 24108 15874 24164 15876
rect 24108 15822 24110 15874
rect 24110 15822 24162 15874
rect 24162 15822 24164 15874
rect 24108 15820 24164 15822
rect 24444 15708 24500 15764
rect 23996 15260 24052 15316
rect 23548 15148 23604 15204
rect 24220 15314 24276 15316
rect 24220 15262 24222 15314
rect 24222 15262 24274 15314
rect 24274 15262 24276 15314
rect 24220 15260 24276 15262
rect 24108 15148 24164 15204
rect 23660 14642 23716 14644
rect 23660 14590 23662 14642
rect 23662 14590 23714 14642
rect 23714 14590 23716 14642
rect 23660 14588 23716 14590
rect 25564 19346 25620 19348
rect 25564 19294 25566 19346
rect 25566 19294 25618 19346
rect 25618 19294 25620 19346
rect 25564 19292 25620 19294
rect 25452 18674 25508 18676
rect 25452 18622 25454 18674
rect 25454 18622 25506 18674
rect 25506 18622 25508 18674
rect 25452 18620 25508 18622
rect 25788 18508 25844 18564
rect 25228 17612 25284 17668
rect 25676 18450 25732 18452
rect 25676 18398 25678 18450
rect 25678 18398 25730 18450
rect 25730 18398 25732 18450
rect 25676 18396 25732 18398
rect 25564 18338 25620 18340
rect 25564 18286 25566 18338
rect 25566 18286 25618 18338
rect 25618 18286 25620 18338
rect 25564 18284 25620 18286
rect 25900 19292 25956 19348
rect 30268 23436 30324 23492
rect 32172 25618 32228 25620
rect 32172 25566 32174 25618
rect 32174 25566 32226 25618
rect 32226 25566 32228 25618
rect 32172 25564 32228 25566
rect 36204 28530 36260 28532
rect 36204 28478 36206 28530
rect 36206 28478 36258 28530
rect 36258 28478 36260 28530
rect 36204 28476 36260 28478
rect 33068 25452 33124 25508
rect 36316 26178 36372 26180
rect 36316 26126 36318 26178
rect 36318 26126 36370 26178
rect 36370 26126 36372 26178
rect 36316 26124 36372 26126
rect 35196 25898 35252 25900
rect 35196 25846 35198 25898
rect 35198 25846 35250 25898
rect 35250 25846 35252 25898
rect 35196 25844 35252 25846
rect 35300 25898 35356 25900
rect 35300 25846 35302 25898
rect 35302 25846 35354 25898
rect 35354 25846 35356 25898
rect 35300 25844 35356 25846
rect 35404 25898 35460 25900
rect 35404 25846 35406 25898
rect 35406 25846 35458 25898
rect 35458 25846 35460 25898
rect 35404 25844 35460 25846
rect 30940 24946 30996 24948
rect 30940 24894 30942 24946
rect 30942 24894 30994 24946
rect 30994 24894 30996 24946
rect 30940 24892 30996 24894
rect 30828 24722 30884 24724
rect 30828 24670 30830 24722
rect 30830 24670 30882 24722
rect 30882 24670 30884 24722
rect 30828 24668 30884 24670
rect 30828 23938 30884 23940
rect 30828 23886 30830 23938
rect 30830 23886 30882 23938
rect 30882 23886 30884 23938
rect 30828 23884 30884 23886
rect 29708 23154 29764 23156
rect 29708 23102 29710 23154
rect 29710 23102 29762 23154
rect 29762 23102 29764 23154
rect 29708 23100 29764 23102
rect 29596 22428 29652 22484
rect 26796 21586 26852 21588
rect 26796 21534 26798 21586
rect 26798 21534 26850 21586
rect 26850 21534 26852 21586
rect 26796 21532 26852 21534
rect 27692 21586 27748 21588
rect 27692 21534 27694 21586
rect 27694 21534 27746 21586
rect 27746 21534 27748 21586
rect 27692 21532 27748 21534
rect 26572 20690 26628 20692
rect 26572 20638 26574 20690
rect 26574 20638 26626 20690
rect 26626 20638 26628 20690
rect 26572 20636 26628 20638
rect 27580 20524 27636 20580
rect 25900 18620 25956 18676
rect 27020 19740 27076 19796
rect 25228 17106 25284 17108
rect 25228 17054 25230 17106
rect 25230 17054 25282 17106
rect 25282 17054 25284 17106
rect 25228 17052 25284 17054
rect 24780 16380 24836 16436
rect 24668 16098 24724 16100
rect 24668 16046 24670 16098
rect 24670 16046 24722 16098
rect 24722 16046 24724 16098
rect 24668 16044 24724 16046
rect 24556 14476 24612 14532
rect 25340 15426 25396 15428
rect 25340 15374 25342 15426
rect 25342 15374 25394 15426
rect 25394 15374 25396 15426
rect 25340 15372 25396 15374
rect 26572 18620 26628 18676
rect 26460 18396 26516 18452
rect 27020 18284 27076 18340
rect 27244 18396 27300 18452
rect 29148 21868 29204 21924
rect 29260 21756 29316 21812
rect 29708 21868 29764 21924
rect 28028 19964 28084 20020
rect 28252 21308 28308 21364
rect 27916 19404 27972 19460
rect 28364 20524 28420 20580
rect 28588 19010 28644 19012
rect 28588 18958 28590 19010
rect 28590 18958 28642 19010
rect 28642 18958 28644 19010
rect 28588 18956 28644 18958
rect 28924 20018 28980 20020
rect 28924 19966 28926 20018
rect 28926 19966 28978 20018
rect 28978 19966 28980 20018
rect 28924 19964 28980 19966
rect 28812 19794 28868 19796
rect 28812 19742 28814 19794
rect 28814 19742 28866 19794
rect 28866 19742 28868 19794
rect 28812 19740 28868 19742
rect 28700 18732 28756 18788
rect 28364 18562 28420 18564
rect 28364 18510 28366 18562
rect 28366 18510 28418 18562
rect 28418 18510 28420 18562
rect 28364 18508 28420 18510
rect 29260 19740 29316 19796
rect 29260 19122 29316 19124
rect 29260 19070 29262 19122
rect 29262 19070 29314 19122
rect 29314 19070 29316 19122
rect 29260 19068 29316 19070
rect 30156 21586 30212 21588
rect 30156 21534 30158 21586
rect 30158 21534 30210 21586
rect 30210 21534 30212 21586
rect 30156 21532 30212 21534
rect 30716 22316 30772 22372
rect 30940 23378 30996 23380
rect 30940 23326 30942 23378
rect 30942 23326 30994 23378
rect 30994 23326 30996 23378
rect 30940 23324 30996 23326
rect 31052 23266 31108 23268
rect 31052 23214 31054 23266
rect 31054 23214 31106 23266
rect 31106 23214 31108 23266
rect 31052 23212 31108 23214
rect 32732 23548 32788 23604
rect 32060 23436 32116 23492
rect 31500 23212 31556 23268
rect 31948 23266 32004 23268
rect 31948 23214 31950 23266
rect 31950 23214 32002 23266
rect 32002 23214 32004 23266
rect 31948 23212 32004 23214
rect 32060 22316 32116 22372
rect 32508 22540 32564 22596
rect 32284 22316 32340 22372
rect 31388 21868 31444 21924
rect 30828 21756 30884 21812
rect 30492 21586 30548 21588
rect 30492 21534 30494 21586
rect 30494 21534 30546 21586
rect 30546 21534 30548 21586
rect 30492 21532 30548 21534
rect 30828 21586 30884 21588
rect 30828 21534 30830 21586
rect 30830 21534 30882 21586
rect 30882 21534 30884 21586
rect 30828 21532 30884 21534
rect 30940 20748 30996 20804
rect 31052 20578 31108 20580
rect 31052 20526 31054 20578
rect 31054 20526 31106 20578
rect 31106 20526 31108 20578
rect 31052 20524 31108 20526
rect 30380 20188 30436 20244
rect 30156 20130 30212 20132
rect 30156 20078 30158 20130
rect 30158 20078 30210 20130
rect 30210 20078 30212 20130
rect 30156 20076 30212 20078
rect 29708 18956 29764 19012
rect 29820 19068 29876 19124
rect 29036 18620 29092 18676
rect 29484 18844 29540 18900
rect 26236 16716 26292 16772
rect 27916 16380 27972 16436
rect 25676 15708 25732 15764
rect 27916 15820 27972 15876
rect 26012 15372 26068 15428
rect 26684 15372 26740 15428
rect 26124 15314 26180 15316
rect 26124 15262 26126 15314
rect 26126 15262 26178 15314
rect 26178 15262 26180 15314
rect 26124 15260 26180 15262
rect 25564 14700 25620 14756
rect 26012 15148 26068 15204
rect 24556 14306 24612 14308
rect 24556 14254 24558 14306
rect 24558 14254 24610 14306
rect 24610 14254 24612 14306
rect 24556 14252 24612 14254
rect 24444 13858 24500 13860
rect 24444 13806 24446 13858
rect 24446 13806 24498 13858
rect 24498 13806 24500 13858
rect 24444 13804 24500 13806
rect 23100 13244 23156 13300
rect 23324 13580 23380 13636
rect 23772 13746 23828 13748
rect 23772 13694 23774 13746
rect 23774 13694 23826 13746
rect 23826 13694 23828 13746
rect 23772 13692 23828 13694
rect 23660 13634 23716 13636
rect 23660 13582 23662 13634
rect 23662 13582 23714 13634
rect 23714 13582 23716 13634
rect 23660 13580 23716 13582
rect 23996 13580 24052 13636
rect 23548 13020 23604 13076
rect 23996 13244 24052 13300
rect 24332 13074 24388 13076
rect 24332 13022 24334 13074
rect 24334 13022 24386 13074
rect 24386 13022 24388 13074
rect 24332 13020 24388 13022
rect 24220 12348 24276 12404
rect 23436 12290 23492 12292
rect 23436 12238 23438 12290
rect 23438 12238 23490 12290
rect 23490 12238 23492 12290
rect 23436 12236 23492 12238
rect 22988 10444 23044 10500
rect 23212 10220 23268 10276
rect 24780 14140 24836 14196
rect 25004 13804 25060 13860
rect 25340 14476 25396 14532
rect 27692 15426 27748 15428
rect 27692 15374 27694 15426
rect 27694 15374 27746 15426
rect 27746 15374 27748 15426
rect 27692 15372 27748 15374
rect 27580 15314 27636 15316
rect 27580 15262 27582 15314
rect 27582 15262 27634 15314
rect 27634 15262 27636 15314
rect 27580 15260 27636 15262
rect 26236 14642 26292 14644
rect 26236 14590 26238 14642
rect 26238 14590 26290 14642
rect 26290 14590 26292 14642
rect 26236 14588 26292 14590
rect 25116 13580 25172 13636
rect 27244 14418 27300 14420
rect 27244 14366 27246 14418
rect 27246 14366 27298 14418
rect 27298 14366 27300 14418
rect 27244 14364 27300 14366
rect 26124 14140 26180 14196
rect 27356 14306 27412 14308
rect 27356 14254 27358 14306
rect 27358 14254 27410 14306
rect 27410 14254 27412 14306
rect 27356 14252 27412 14254
rect 27244 14140 27300 14196
rect 27468 14140 27524 14196
rect 28924 16994 28980 16996
rect 28924 16942 28926 16994
rect 28926 16942 28978 16994
rect 28978 16942 28980 16994
rect 28924 16940 28980 16942
rect 28700 16156 28756 16212
rect 28588 15986 28644 15988
rect 28588 15934 28590 15986
rect 28590 15934 28642 15986
rect 28642 15934 28644 15986
rect 28588 15932 28644 15934
rect 28476 14588 28532 14644
rect 29596 18620 29652 18676
rect 30156 19346 30212 19348
rect 30156 19294 30158 19346
rect 30158 19294 30210 19346
rect 30210 19294 30212 19346
rect 30156 19292 30212 19294
rect 30268 19234 30324 19236
rect 30268 19182 30270 19234
rect 30270 19182 30322 19234
rect 30322 19182 30324 19234
rect 30268 19180 30324 19182
rect 30604 18956 30660 19012
rect 30940 19010 30996 19012
rect 30940 18958 30942 19010
rect 30942 18958 30994 19010
rect 30994 18958 30996 19010
rect 30940 18956 30996 18958
rect 32060 21532 32116 21588
rect 31276 20860 31332 20916
rect 32172 20914 32228 20916
rect 32172 20862 32174 20914
rect 32174 20862 32226 20914
rect 32226 20862 32228 20914
rect 32172 20860 32228 20862
rect 31500 20802 31556 20804
rect 31500 20750 31502 20802
rect 31502 20750 31554 20802
rect 31554 20750 31556 20802
rect 31500 20748 31556 20750
rect 31948 20636 32004 20692
rect 32396 20188 32452 20244
rect 32284 20076 32340 20132
rect 31276 19292 31332 19348
rect 31164 18844 31220 18900
rect 31276 18956 31332 19012
rect 30940 18732 30996 18788
rect 30380 18674 30436 18676
rect 30380 18622 30382 18674
rect 30382 18622 30434 18674
rect 30434 18622 30436 18674
rect 30380 18620 30436 18622
rect 29932 18562 29988 18564
rect 29932 18510 29934 18562
rect 29934 18510 29986 18562
rect 29986 18510 29988 18562
rect 29932 18508 29988 18510
rect 29820 18396 29876 18452
rect 30156 18562 30212 18564
rect 30156 18510 30158 18562
rect 30158 18510 30210 18562
rect 30210 18510 30212 18562
rect 30156 18508 30212 18510
rect 30156 17724 30212 17780
rect 31276 18732 31332 18788
rect 31164 18562 31220 18564
rect 31164 18510 31166 18562
rect 31166 18510 31218 18562
rect 31218 18510 31220 18562
rect 31164 18508 31220 18510
rect 30940 17948 30996 18004
rect 31276 17836 31332 17892
rect 30828 17778 30884 17780
rect 30828 17726 30830 17778
rect 30830 17726 30882 17778
rect 30882 17726 30884 17778
rect 30828 17724 30884 17726
rect 31836 19404 31892 19460
rect 32284 19068 32340 19124
rect 32060 19010 32116 19012
rect 32060 18958 32062 19010
rect 32062 18958 32114 19010
rect 32114 18958 32116 19010
rect 32060 18956 32116 18958
rect 31612 18732 31668 18788
rect 31500 17612 31556 17668
rect 31836 18732 31892 18788
rect 32508 18620 32564 18676
rect 31724 18284 31780 18340
rect 31836 17948 31892 18004
rect 31836 17666 31892 17668
rect 31836 17614 31838 17666
rect 31838 17614 31890 17666
rect 31890 17614 31892 17666
rect 31836 17612 31892 17614
rect 29260 16994 29316 16996
rect 29260 16942 29262 16994
rect 29262 16942 29314 16994
rect 29314 16942 29316 16994
rect 29260 16940 29316 16942
rect 29484 16882 29540 16884
rect 29484 16830 29486 16882
rect 29486 16830 29538 16882
rect 29538 16830 29540 16882
rect 29484 16828 29540 16830
rect 28700 14476 28756 14532
rect 26348 13356 26404 13412
rect 26236 12908 26292 12964
rect 26124 12124 26180 12180
rect 25116 11004 25172 11060
rect 25340 12012 25396 12068
rect 24892 10668 24948 10724
rect 24668 10498 24724 10500
rect 24668 10446 24670 10498
rect 24670 10446 24722 10498
rect 24722 10446 24724 10498
rect 24668 10444 24724 10446
rect 25228 10444 25284 10500
rect 24444 10220 24500 10276
rect 26796 12348 26852 12404
rect 28028 14364 28084 14420
rect 28028 13580 28084 13636
rect 28476 13634 28532 13636
rect 28476 13582 28478 13634
rect 28478 13582 28530 13634
rect 28530 13582 28532 13634
rect 28476 13580 28532 13582
rect 28924 13634 28980 13636
rect 28924 13582 28926 13634
rect 28926 13582 28978 13634
rect 28978 13582 28980 13634
rect 28924 13580 28980 13582
rect 27244 13356 27300 13412
rect 26908 13020 26964 13076
rect 27468 12962 27524 12964
rect 27468 12910 27470 12962
rect 27470 12910 27522 12962
rect 27522 12910 27524 12962
rect 27468 12908 27524 12910
rect 28700 13074 28756 13076
rect 28700 13022 28702 13074
rect 28702 13022 28754 13074
rect 28754 13022 28756 13074
rect 28700 13020 28756 13022
rect 28252 12908 28308 12964
rect 27244 12348 27300 12404
rect 27244 12012 27300 12068
rect 26012 10722 26068 10724
rect 26012 10670 26014 10722
rect 26014 10670 26066 10722
rect 26066 10670 26068 10722
rect 26012 10668 26068 10670
rect 27468 10220 27524 10276
rect 25676 9938 25732 9940
rect 25676 9886 25678 9938
rect 25678 9886 25730 9938
rect 25730 9886 25732 9938
rect 25676 9884 25732 9886
rect 21420 9548 21476 9604
rect 22092 9602 22148 9604
rect 22092 9550 22094 9602
rect 22094 9550 22146 9602
rect 22146 9550 22148 9602
rect 22092 9548 22148 9550
rect 26236 9660 26292 9716
rect 21196 8988 21252 9044
rect 18396 7644 18452 7700
rect 17948 7308 18004 7364
rect 16604 5740 16660 5796
rect 16940 5628 16996 5684
rect 17724 6412 17780 6468
rect 19068 7586 19124 7588
rect 19068 7534 19070 7586
rect 19070 7534 19122 7586
rect 19122 7534 19124 7586
rect 19068 7532 19124 7534
rect 17052 5180 17108 5236
rect 18956 7362 19012 7364
rect 18956 7310 18958 7362
rect 18958 7310 19010 7362
rect 19010 7310 19012 7362
rect 18956 7308 19012 7310
rect 16716 4172 16772 4228
rect 17500 6018 17556 6020
rect 17500 5966 17502 6018
rect 17502 5966 17554 6018
rect 17554 5966 17556 6018
rect 17500 5964 17556 5966
rect 17724 5292 17780 5348
rect 17500 3612 17556 3668
rect 17836 5068 17892 5124
rect 18060 5068 18116 5124
rect 17948 4562 18004 4564
rect 17948 4510 17950 4562
rect 17950 4510 18002 4562
rect 18002 4510 18004 4562
rect 17948 4508 18004 4510
rect 18396 5682 18452 5684
rect 18396 5630 18398 5682
rect 18398 5630 18450 5682
rect 18450 5630 18452 5682
rect 18396 5628 18452 5630
rect 19836 7866 19892 7868
rect 19404 7756 19460 7812
rect 19836 7814 19838 7866
rect 19838 7814 19890 7866
rect 19890 7814 19892 7866
rect 19836 7812 19892 7814
rect 19940 7866 19996 7868
rect 19940 7814 19942 7866
rect 19942 7814 19994 7866
rect 19994 7814 19996 7866
rect 19940 7812 19996 7814
rect 20044 7866 20100 7868
rect 20044 7814 20046 7866
rect 20046 7814 20098 7866
rect 20098 7814 20100 7866
rect 20044 7812 20100 7814
rect 19740 7586 19796 7588
rect 19740 7534 19742 7586
rect 19742 7534 19794 7586
rect 19794 7534 19796 7586
rect 19740 7532 19796 7534
rect 19836 6298 19892 6300
rect 19836 6246 19838 6298
rect 19838 6246 19890 6298
rect 19890 6246 19892 6298
rect 19836 6244 19892 6246
rect 19940 6298 19996 6300
rect 19940 6246 19942 6298
rect 19942 6246 19994 6298
rect 19994 6246 19996 6298
rect 19940 6244 19996 6246
rect 20044 6298 20100 6300
rect 20044 6246 20046 6298
rect 20046 6246 20098 6298
rect 20098 6246 20100 6298
rect 20044 6244 20100 6246
rect 19068 5292 19124 5348
rect 18508 5068 18564 5124
rect 18732 5180 18788 5236
rect 18844 5068 18900 5124
rect 18620 3666 18676 3668
rect 18620 3614 18622 3666
rect 18622 3614 18674 3666
rect 18674 3614 18676 3666
rect 18620 3612 18676 3614
rect 19852 5906 19908 5908
rect 19852 5854 19854 5906
rect 19854 5854 19906 5906
rect 19906 5854 19908 5906
rect 19852 5852 19908 5854
rect 19516 5628 19572 5684
rect 19740 5010 19796 5012
rect 19740 4958 19742 5010
rect 19742 4958 19794 5010
rect 19794 4958 19796 5010
rect 19740 4956 19796 4958
rect 19836 4730 19892 4732
rect 19836 4678 19838 4730
rect 19838 4678 19890 4730
rect 19890 4678 19892 4730
rect 19836 4676 19892 4678
rect 19940 4730 19996 4732
rect 19940 4678 19942 4730
rect 19942 4678 19994 4730
rect 19994 4678 19996 4730
rect 19940 4676 19996 4678
rect 20044 4730 20100 4732
rect 20044 4678 20046 4730
rect 20046 4678 20098 4730
rect 20098 4678 20100 4730
rect 20044 4676 20100 4678
rect 20188 4508 20244 4564
rect 20524 5906 20580 5908
rect 20524 5854 20526 5906
rect 20526 5854 20578 5906
rect 20578 5854 20580 5906
rect 20524 5852 20580 5854
rect 20748 5740 20804 5796
rect 20748 5234 20804 5236
rect 20748 5182 20750 5234
rect 20750 5182 20802 5234
rect 20802 5182 20804 5234
rect 20748 5180 20804 5182
rect 21644 8988 21700 9044
rect 21532 8428 21588 8484
rect 21420 7586 21476 7588
rect 21420 7534 21422 7586
rect 21422 7534 21474 7586
rect 21474 7534 21476 7586
rect 21420 7532 21476 7534
rect 22092 8428 22148 8484
rect 21980 8258 22036 8260
rect 21980 8206 21982 8258
rect 21982 8206 22034 8258
rect 22034 8206 22036 8258
rect 21980 8204 22036 8206
rect 22428 8428 22484 8484
rect 28252 12460 28308 12516
rect 28252 12124 28308 12180
rect 28140 11506 28196 11508
rect 28140 11454 28142 11506
rect 28142 11454 28194 11506
rect 28194 11454 28196 11506
rect 28140 11452 28196 11454
rect 28028 10556 28084 10612
rect 27692 9996 27748 10052
rect 27804 10444 27860 10500
rect 27580 9548 27636 9604
rect 31500 17164 31556 17220
rect 31724 16940 31780 16996
rect 31836 17052 31892 17108
rect 30268 15986 30324 15988
rect 30268 15934 30270 15986
rect 30270 15934 30322 15986
rect 30322 15934 30324 15986
rect 30268 15932 30324 15934
rect 29260 13858 29316 13860
rect 29260 13806 29262 13858
rect 29262 13806 29314 13858
rect 29314 13806 29316 13858
rect 29260 13804 29316 13806
rect 29484 14530 29540 14532
rect 29484 14478 29486 14530
rect 29486 14478 29538 14530
rect 29538 14478 29540 14530
rect 29484 14476 29540 14478
rect 31164 15874 31220 15876
rect 31164 15822 31166 15874
rect 31166 15822 31218 15874
rect 31218 15822 31220 15874
rect 31164 15820 31220 15822
rect 32060 17388 32116 17444
rect 32060 17164 32116 17220
rect 32284 17666 32340 17668
rect 32284 17614 32286 17666
rect 32286 17614 32338 17666
rect 32338 17614 32340 17666
rect 32284 17612 32340 17614
rect 35196 24330 35252 24332
rect 35196 24278 35198 24330
rect 35198 24278 35250 24330
rect 35250 24278 35252 24330
rect 35196 24276 35252 24278
rect 35300 24330 35356 24332
rect 35300 24278 35302 24330
rect 35302 24278 35354 24330
rect 35354 24278 35356 24330
rect 35300 24276 35356 24278
rect 35404 24330 35460 24332
rect 35404 24278 35406 24330
rect 35406 24278 35458 24330
rect 35458 24278 35460 24330
rect 35404 24276 35460 24278
rect 36316 23996 36372 24052
rect 35532 23660 35588 23716
rect 33740 23212 33796 23268
rect 33180 19404 33236 19460
rect 33292 20188 33348 20244
rect 33180 19234 33236 19236
rect 33180 19182 33182 19234
rect 33182 19182 33234 19234
rect 33234 19182 33236 19234
rect 33180 19180 33236 19182
rect 35532 23154 35588 23156
rect 35532 23102 35534 23154
rect 35534 23102 35586 23154
rect 35586 23102 35588 23154
rect 35532 23100 35588 23102
rect 35196 22762 35252 22764
rect 35196 22710 35198 22762
rect 35198 22710 35250 22762
rect 35250 22710 35252 22762
rect 35196 22708 35252 22710
rect 35300 22762 35356 22764
rect 35300 22710 35302 22762
rect 35302 22710 35354 22762
rect 35354 22710 35356 22762
rect 35300 22708 35356 22710
rect 35404 22762 35460 22764
rect 35404 22710 35406 22762
rect 35406 22710 35458 22762
rect 35458 22710 35460 22762
rect 35404 22708 35460 22710
rect 34412 20412 34468 20468
rect 34636 21308 34692 21364
rect 35980 23884 36036 23940
rect 35868 23548 35924 23604
rect 35196 21308 35252 21364
rect 35196 21194 35252 21196
rect 35196 21142 35198 21194
rect 35198 21142 35250 21194
rect 35250 21142 35252 21194
rect 35196 21140 35252 21142
rect 35300 21194 35356 21196
rect 35300 21142 35302 21194
rect 35302 21142 35354 21194
rect 35354 21142 35356 21194
rect 35300 21140 35356 21142
rect 35404 21194 35460 21196
rect 35404 21142 35406 21194
rect 35406 21142 35458 21194
rect 35458 21142 35460 21194
rect 35404 21140 35460 21142
rect 34636 20748 34692 20804
rect 34300 20188 34356 20244
rect 33964 19346 34020 19348
rect 33964 19294 33966 19346
rect 33966 19294 34018 19346
rect 34018 19294 34020 19346
rect 33964 19292 34020 19294
rect 33068 18732 33124 18788
rect 35756 20860 35812 20916
rect 37100 36876 37156 36932
rect 39004 39676 39060 39732
rect 39676 40684 39732 40740
rect 39788 41074 39844 41076
rect 39788 41022 39790 41074
rect 39790 41022 39842 41074
rect 39842 41022 39844 41074
rect 39788 41020 39844 41022
rect 39788 40348 39844 40404
rect 39900 39506 39956 39508
rect 39900 39454 39902 39506
rect 39902 39454 39954 39506
rect 39954 39454 39956 39506
rect 39900 39452 39956 39454
rect 39564 39004 39620 39060
rect 40908 43650 40964 43652
rect 40908 43598 40910 43650
rect 40910 43598 40962 43650
rect 40962 43598 40964 43650
rect 40908 43596 40964 43598
rect 42028 43932 42084 43988
rect 41244 43538 41300 43540
rect 41244 43486 41246 43538
rect 41246 43486 41298 43538
rect 41298 43486 41300 43538
rect 41244 43484 41300 43486
rect 41020 41858 41076 41860
rect 41020 41806 41022 41858
rect 41022 41806 41074 41858
rect 41074 41806 41076 41858
rect 41020 41804 41076 41806
rect 40124 39676 40180 39732
rect 40236 40348 40292 40404
rect 40012 39004 40068 39060
rect 40348 39004 40404 39060
rect 39900 38834 39956 38836
rect 39900 38782 39902 38834
rect 39902 38782 39954 38834
rect 39954 38782 39956 38834
rect 39900 38780 39956 38782
rect 39900 37490 39956 37492
rect 39900 37438 39902 37490
rect 39902 37438 39954 37490
rect 39954 37438 39956 37490
rect 39900 37436 39956 37438
rect 39452 36876 39508 36932
rect 38220 36540 38276 36596
rect 39004 36428 39060 36484
rect 37100 33852 37156 33908
rect 37436 33628 37492 33684
rect 37772 34636 37828 34692
rect 37772 33404 37828 33460
rect 37212 33122 37268 33124
rect 37212 33070 37214 33122
rect 37214 33070 37266 33122
rect 37266 33070 37268 33122
rect 37212 33068 37268 33070
rect 38780 33180 38836 33236
rect 38108 33068 38164 33124
rect 37212 30156 37268 30212
rect 37212 29484 37268 29540
rect 37324 29372 37380 29428
rect 36540 28476 36596 28532
rect 37996 30828 38052 30884
rect 39900 36594 39956 36596
rect 39900 36542 39902 36594
rect 39902 36542 39954 36594
rect 39954 36542 39956 36594
rect 39900 36540 39956 36542
rect 41020 40962 41076 40964
rect 41020 40910 41022 40962
rect 41022 40910 41074 40962
rect 41074 40910 41076 40962
rect 41020 40908 41076 40910
rect 41804 40572 41860 40628
rect 41692 40514 41748 40516
rect 41692 40462 41694 40514
rect 41694 40462 41746 40514
rect 41746 40462 41748 40514
rect 41692 40460 41748 40462
rect 40908 39452 40964 39508
rect 42364 41074 42420 41076
rect 42364 41022 42366 41074
rect 42366 41022 42418 41074
rect 42418 41022 42420 41074
rect 42364 41020 42420 41022
rect 42028 40796 42084 40852
rect 42700 40796 42756 40852
rect 41804 40124 41860 40180
rect 41356 40012 41412 40068
rect 42028 40012 42084 40068
rect 43260 44380 43316 44436
rect 42924 43484 42980 43540
rect 42812 39788 42868 39844
rect 42924 42588 42980 42644
rect 43820 42642 43876 42644
rect 43820 42590 43822 42642
rect 43822 42590 43874 42642
rect 43874 42590 43876 42642
rect 43820 42588 43876 42590
rect 43596 41916 43652 41972
rect 41692 39058 41748 39060
rect 41692 39006 41694 39058
rect 41694 39006 41746 39058
rect 41746 39006 41748 39058
rect 41692 39004 41748 39006
rect 40684 38668 40740 38724
rect 43708 40908 43764 40964
rect 43932 41804 43988 41860
rect 45276 46396 45332 46452
rect 45052 45724 45108 45780
rect 44380 45276 44436 45332
rect 44604 45052 44660 45108
rect 44716 44994 44772 44996
rect 44716 44942 44718 44994
rect 44718 44942 44770 44994
rect 44770 44942 44772 44994
rect 44716 44940 44772 44942
rect 45052 44940 45108 44996
rect 44940 44546 44996 44548
rect 44940 44494 44942 44546
rect 44942 44494 44994 44546
rect 44994 44494 44996 44546
rect 44940 44492 44996 44494
rect 44716 43820 44772 43876
rect 46060 45330 46116 45332
rect 46060 45278 46062 45330
rect 46062 45278 46114 45330
rect 46114 45278 46116 45330
rect 46060 45276 46116 45278
rect 46844 45052 46900 45108
rect 45836 44380 45892 44436
rect 45276 43932 45332 43988
rect 45052 42140 45108 42196
rect 44492 41804 44548 41860
rect 44268 41692 44324 41748
rect 44156 41132 44212 41188
rect 44156 40460 44212 40516
rect 43484 40178 43540 40180
rect 43484 40126 43486 40178
rect 43486 40126 43538 40178
rect 43538 40126 43540 40178
rect 43484 40124 43540 40126
rect 43372 39842 43428 39844
rect 43372 39790 43374 39842
rect 43374 39790 43426 39842
rect 43426 39790 43428 39842
rect 43372 39788 43428 39790
rect 44940 40348 44996 40404
rect 45276 39676 45332 39732
rect 47740 44380 47796 44436
rect 45724 41132 45780 41188
rect 46844 42140 46900 42196
rect 45836 41804 45892 41860
rect 45612 40012 45668 40068
rect 45500 39788 45556 39844
rect 41692 37884 41748 37940
rect 41468 37772 41524 37828
rect 41020 37490 41076 37492
rect 41020 37438 41022 37490
rect 41022 37438 41074 37490
rect 41074 37438 41076 37490
rect 41020 37436 41076 37438
rect 42140 37436 42196 37492
rect 42028 37154 42084 37156
rect 42028 37102 42030 37154
rect 42030 37102 42082 37154
rect 42082 37102 42084 37154
rect 42028 37100 42084 37102
rect 42476 36482 42532 36484
rect 42476 36430 42478 36482
rect 42478 36430 42530 36482
rect 42530 36430 42532 36482
rect 42476 36428 42532 36430
rect 40124 35922 40180 35924
rect 40124 35870 40126 35922
rect 40126 35870 40178 35922
rect 40178 35870 40180 35922
rect 40124 35868 40180 35870
rect 40236 35756 40292 35812
rect 39788 35308 39844 35364
rect 41692 35922 41748 35924
rect 41692 35870 41694 35922
rect 41694 35870 41746 35922
rect 41746 35870 41748 35922
rect 41692 35868 41748 35870
rect 41356 34972 41412 35028
rect 41132 34914 41188 34916
rect 41132 34862 41134 34914
rect 41134 34862 41186 34914
rect 41186 34862 41188 34914
rect 41132 34860 41188 34862
rect 40908 34690 40964 34692
rect 40908 34638 40910 34690
rect 40910 34638 40962 34690
rect 40962 34638 40964 34690
rect 40908 34636 40964 34638
rect 43148 38108 43204 38164
rect 43036 37826 43092 37828
rect 43036 37774 43038 37826
rect 43038 37774 43090 37826
rect 43090 37774 43092 37826
rect 43036 37772 43092 37774
rect 43372 38050 43428 38052
rect 43372 37998 43374 38050
rect 43374 37998 43426 38050
rect 43426 37998 43428 38050
rect 43372 37996 43428 37998
rect 42252 34972 42308 35028
rect 43148 36482 43204 36484
rect 43148 36430 43150 36482
rect 43150 36430 43202 36482
rect 43202 36430 43204 36482
rect 43148 36428 43204 36430
rect 42252 34748 42308 34804
rect 41356 34524 41412 34580
rect 39340 33628 39396 33684
rect 39340 32060 39396 32116
rect 38668 31836 38724 31892
rect 40908 33628 40964 33684
rect 40460 33122 40516 33124
rect 40460 33070 40462 33122
rect 40462 33070 40514 33122
rect 40514 33070 40516 33122
rect 40460 33068 40516 33070
rect 41580 32674 41636 32676
rect 41580 32622 41582 32674
rect 41582 32622 41634 32674
rect 41634 32622 41636 32674
rect 41580 32620 41636 32622
rect 40124 32508 40180 32564
rect 39676 31948 39732 32004
rect 39788 31836 39844 31892
rect 38444 31164 38500 31220
rect 38220 30156 38276 30212
rect 38780 30882 38836 30884
rect 38780 30830 38782 30882
rect 38782 30830 38834 30882
rect 38834 30830 38836 30882
rect 38780 30828 38836 30830
rect 41020 32060 41076 32116
rect 38332 28924 38388 28980
rect 37772 27074 37828 27076
rect 37772 27022 37774 27074
rect 37774 27022 37826 27074
rect 37826 27022 37828 27074
rect 37772 27020 37828 27022
rect 39116 28924 39172 28980
rect 39340 29260 39396 29316
rect 39900 28924 39956 28980
rect 40684 30156 40740 30212
rect 42364 34690 42420 34692
rect 42364 34638 42366 34690
rect 42366 34638 42418 34690
rect 42418 34638 42420 34690
rect 42364 34636 42420 34638
rect 41916 32338 41972 32340
rect 41916 32286 41918 32338
rect 41918 32286 41970 32338
rect 41970 32286 41972 32338
rect 41916 32284 41972 32286
rect 42812 34914 42868 34916
rect 42812 34862 42814 34914
rect 42814 34862 42866 34914
rect 42866 34862 42868 34914
rect 42812 34860 42868 34862
rect 41132 31218 41188 31220
rect 41132 31166 41134 31218
rect 41134 31166 41186 31218
rect 41186 31166 41188 31218
rect 41132 31164 41188 31166
rect 41692 31724 41748 31780
rect 42588 31612 42644 31668
rect 43260 35196 43316 35252
rect 44156 38108 44212 38164
rect 44940 38162 44996 38164
rect 44940 38110 44942 38162
rect 44942 38110 44994 38162
rect 44994 38110 44996 38162
rect 44940 38108 44996 38110
rect 47404 42700 47460 42756
rect 46956 40348 47012 40404
rect 46060 39730 46116 39732
rect 46060 39678 46062 39730
rect 46062 39678 46114 39730
rect 46114 39678 46116 39730
rect 46060 39676 46116 39678
rect 47740 41858 47796 41860
rect 47740 41806 47742 41858
rect 47742 41806 47794 41858
rect 47794 41806 47796 41858
rect 47740 41804 47796 41806
rect 47964 41692 48020 41748
rect 47852 39676 47908 39732
rect 47516 39004 47572 39060
rect 45836 38780 45892 38836
rect 47964 39004 48020 39060
rect 44940 37266 44996 37268
rect 44940 37214 44942 37266
rect 44942 37214 44994 37266
rect 44994 37214 44996 37266
rect 44940 37212 44996 37214
rect 43932 37100 43988 37156
rect 44156 36370 44212 36372
rect 44156 36318 44158 36370
rect 44158 36318 44210 36370
rect 44210 36318 44212 36370
rect 44156 36316 44212 36318
rect 44604 35698 44660 35700
rect 44604 35646 44606 35698
rect 44606 35646 44658 35698
rect 44658 35646 44660 35698
rect 44604 35644 44660 35646
rect 45052 36316 45108 36372
rect 45612 35868 45668 35924
rect 46060 37938 46116 37940
rect 46060 37886 46062 37938
rect 46062 37886 46114 37938
rect 46114 37886 46116 37938
rect 46060 37884 46116 37886
rect 43484 35084 43540 35140
rect 44268 35196 44324 35252
rect 43148 34188 43204 34244
rect 43484 33234 43540 33236
rect 43484 33182 43486 33234
rect 43486 33182 43538 33234
rect 43538 33182 43540 33234
rect 43484 33180 43540 33182
rect 43820 34524 43876 34580
rect 43820 34018 43876 34020
rect 43820 33966 43822 34018
rect 43822 33966 43874 34018
rect 43874 33966 43876 34018
rect 43820 33964 43876 33966
rect 43708 32620 43764 32676
rect 43148 31778 43204 31780
rect 43148 31726 43150 31778
rect 43150 31726 43202 31778
rect 43202 31726 43204 31778
rect 43148 31724 43204 31726
rect 43820 31778 43876 31780
rect 43820 31726 43822 31778
rect 43822 31726 43874 31778
rect 43874 31726 43876 31778
rect 43820 31724 43876 31726
rect 41020 29426 41076 29428
rect 41020 29374 41022 29426
rect 41022 29374 41074 29426
rect 41074 29374 41076 29426
rect 41020 29372 41076 29374
rect 41468 28866 41524 28868
rect 41468 28814 41470 28866
rect 41470 28814 41522 28866
rect 41522 28814 41524 28866
rect 41468 28812 41524 28814
rect 39676 27692 39732 27748
rect 38220 26460 38276 26516
rect 38332 26908 38388 26964
rect 37548 26124 37604 26180
rect 37324 25900 37380 25956
rect 37100 23996 37156 24052
rect 36428 23772 36484 23828
rect 35980 20972 36036 21028
rect 36092 22988 36148 23044
rect 35308 20412 35364 20468
rect 39676 26962 39732 26964
rect 39676 26910 39678 26962
rect 39678 26910 39730 26962
rect 39730 26910 39732 26962
rect 39676 26908 39732 26910
rect 40348 27746 40404 27748
rect 40348 27694 40350 27746
rect 40350 27694 40402 27746
rect 40402 27694 40404 27746
rect 40348 27692 40404 27694
rect 39676 26514 39732 26516
rect 39676 26462 39678 26514
rect 39678 26462 39730 26514
rect 39730 26462 39732 26514
rect 39676 26460 39732 26462
rect 39228 26290 39284 26292
rect 39228 26238 39230 26290
rect 39230 26238 39282 26290
rect 39282 26238 39284 26290
rect 39228 26236 39284 26238
rect 37548 25394 37604 25396
rect 37548 25342 37550 25394
rect 37550 25342 37602 25394
rect 37602 25342 37604 25394
rect 37548 25340 37604 25342
rect 38332 25676 38388 25732
rect 39116 25676 39172 25732
rect 38780 25564 38836 25620
rect 38780 25340 38836 25396
rect 38668 24444 38724 24500
rect 37996 24332 38052 24388
rect 40684 28588 40740 28644
rect 41916 28642 41972 28644
rect 41916 28590 41918 28642
rect 41918 28590 41970 28642
rect 41970 28590 41972 28642
rect 41916 28588 41972 28590
rect 41580 28476 41636 28532
rect 42812 30882 42868 30884
rect 42812 30830 42814 30882
rect 42814 30830 42866 30882
rect 42866 30830 42868 30882
rect 42812 30828 42868 30830
rect 42700 30156 42756 30212
rect 43820 30828 43876 30884
rect 42700 29372 42756 29428
rect 42252 28530 42308 28532
rect 42252 28478 42254 28530
rect 42254 28478 42306 28530
rect 42306 28478 42308 28530
rect 42252 28476 42308 28478
rect 42364 28924 42420 28980
rect 39788 25676 39844 25732
rect 40124 26124 40180 26180
rect 39564 25506 39620 25508
rect 39564 25454 39566 25506
rect 39566 25454 39618 25506
rect 39618 25454 39620 25506
rect 39564 25452 39620 25454
rect 39340 25228 39396 25284
rect 40348 25676 40404 25732
rect 40572 25618 40628 25620
rect 40572 25566 40574 25618
rect 40574 25566 40626 25618
rect 40626 25566 40628 25618
rect 40572 25564 40628 25566
rect 40460 25452 40516 25508
rect 39788 25228 39844 25284
rect 40012 24556 40068 24612
rect 37436 23660 37492 23716
rect 37436 23324 37492 23380
rect 38892 23548 38948 23604
rect 37548 22146 37604 22148
rect 37548 22094 37550 22146
rect 37550 22094 37602 22146
rect 37602 22094 37604 22146
rect 37548 22092 37604 22094
rect 36428 20914 36484 20916
rect 36428 20862 36430 20914
rect 36430 20862 36482 20914
rect 36482 20862 36484 20914
rect 36428 20860 36484 20862
rect 37548 21698 37604 21700
rect 37548 21646 37550 21698
rect 37550 21646 37602 21698
rect 37602 21646 37604 21698
rect 37548 21644 37604 21646
rect 36092 19740 36148 19796
rect 35196 19626 35252 19628
rect 35196 19574 35198 19626
rect 35198 19574 35250 19626
rect 35250 19574 35252 19626
rect 35196 19572 35252 19574
rect 35300 19626 35356 19628
rect 35300 19574 35302 19626
rect 35302 19574 35354 19626
rect 35354 19574 35356 19626
rect 35300 19572 35356 19574
rect 35404 19626 35460 19628
rect 35404 19574 35406 19626
rect 35406 19574 35458 19626
rect 35458 19574 35460 19626
rect 35404 19572 35460 19574
rect 35308 19404 35364 19460
rect 33516 18956 33572 19012
rect 32844 18620 32900 18676
rect 32620 17612 32676 17668
rect 32956 18508 33012 18564
rect 32956 17554 33012 17556
rect 32956 17502 32958 17554
rect 32958 17502 33010 17554
rect 33010 17502 33012 17554
rect 32956 17500 33012 17502
rect 33068 18284 33124 18340
rect 31612 15986 31668 15988
rect 31612 15934 31614 15986
rect 31614 15934 31666 15986
rect 31666 15934 31668 15986
rect 31612 15932 31668 15934
rect 32844 16940 32900 16996
rect 33068 17052 33124 17108
rect 33516 16882 33572 16884
rect 33516 16830 33518 16882
rect 33518 16830 33570 16882
rect 33570 16830 33572 16882
rect 33516 16828 33572 16830
rect 33068 16604 33124 16660
rect 33068 15932 33124 15988
rect 29820 14476 29876 14532
rect 29932 14700 29988 14756
rect 29596 14140 29652 14196
rect 29372 13692 29428 13748
rect 29484 13804 29540 13860
rect 29596 12850 29652 12852
rect 29596 12798 29598 12850
rect 29598 12798 29650 12850
rect 29650 12798 29652 12850
rect 29596 12796 29652 12798
rect 29820 12796 29876 12852
rect 29036 11452 29092 11508
rect 28476 11394 28532 11396
rect 28476 11342 28478 11394
rect 28478 11342 28530 11394
rect 28530 11342 28532 11394
rect 28476 11340 28532 11342
rect 29260 12460 29316 12516
rect 29372 12402 29428 12404
rect 29372 12350 29374 12402
rect 29374 12350 29426 12402
rect 29426 12350 29428 12402
rect 29372 12348 29428 12350
rect 30156 14530 30212 14532
rect 30156 14478 30158 14530
rect 30158 14478 30210 14530
rect 30210 14478 30212 14530
rect 30156 14476 30212 14478
rect 30380 14028 30436 14084
rect 30380 13020 30436 13076
rect 30268 12850 30324 12852
rect 30268 12798 30270 12850
rect 30270 12798 30322 12850
rect 30322 12798 30324 12850
rect 30268 12796 30324 12798
rect 30044 12124 30100 12180
rect 29372 11394 29428 11396
rect 29372 11342 29374 11394
rect 29374 11342 29426 11394
rect 29426 11342 29428 11394
rect 29372 11340 29428 11342
rect 29708 11282 29764 11284
rect 29708 11230 29710 11282
rect 29710 11230 29762 11282
rect 29762 11230 29764 11282
rect 29708 11228 29764 11230
rect 30268 12236 30324 12292
rect 29372 10780 29428 10836
rect 28028 10332 28084 10388
rect 28700 10610 28756 10612
rect 28700 10558 28702 10610
rect 28702 10558 28754 10610
rect 28754 10558 28756 10610
rect 28700 10556 28756 10558
rect 29484 10556 29540 10612
rect 28588 10498 28644 10500
rect 28588 10446 28590 10498
rect 28590 10446 28642 10498
rect 28642 10446 28644 10498
rect 28588 10444 28644 10446
rect 28588 9826 28644 9828
rect 28588 9774 28590 9826
rect 28590 9774 28642 9826
rect 28642 9774 28644 9826
rect 28588 9772 28644 9774
rect 28252 8652 28308 8708
rect 27468 8540 27524 8596
rect 21980 6690 22036 6692
rect 21980 6638 21982 6690
rect 21982 6638 22034 6690
rect 22034 6638 22036 6690
rect 21980 6636 22036 6638
rect 21308 6300 21364 6356
rect 21420 5964 21476 6020
rect 20972 5180 21028 5236
rect 21532 5740 21588 5796
rect 21532 5346 21588 5348
rect 21532 5294 21534 5346
rect 21534 5294 21586 5346
rect 21586 5294 21588 5346
rect 21532 5292 21588 5294
rect 20412 5068 20468 5124
rect 21980 5852 22036 5908
rect 22204 6300 22260 6356
rect 25452 7532 25508 7588
rect 23436 7308 23492 7364
rect 23100 6636 23156 6692
rect 22988 6412 23044 6468
rect 22764 6188 22820 6244
rect 22764 5906 22820 5908
rect 22764 5854 22766 5906
rect 22766 5854 22818 5906
rect 22818 5854 22820 5906
rect 22764 5852 22820 5854
rect 22316 5516 22372 5572
rect 22764 5180 22820 5236
rect 22428 5068 22484 5124
rect 22204 4620 22260 4676
rect 22092 4562 22148 4564
rect 22092 4510 22094 4562
rect 22094 4510 22146 4562
rect 22146 4510 22148 4562
rect 22092 4508 22148 4510
rect 22316 4844 22372 4900
rect 20300 3500 20356 3556
rect 20860 3612 20916 3668
rect 19836 3162 19892 3164
rect 19836 3110 19838 3162
rect 19838 3110 19890 3162
rect 19890 3110 19892 3162
rect 19836 3108 19892 3110
rect 19940 3162 19996 3164
rect 19940 3110 19942 3162
rect 19942 3110 19994 3162
rect 19994 3110 19996 3162
rect 19940 3108 19996 3110
rect 20044 3162 20100 3164
rect 20044 3110 20046 3162
rect 20046 3110 20098 3162
rect 20098 3110 20100 3162
rect 20044 3108 20100 3110
rect 22092 3666 22148 3668
rect 22092 3614 22094 3666
rect 22094 3614 22146 3666
rect 22146 3614 22148 3666
rect 22092 3612 22148 3614
rect 21084 3554 21140 3556
rect 21084 3502 21086 3554
rect 21086 3502 21138 3554
rect 21138 3502 21140 3554
rect 21084 3500 21140 3502
rect 22876 4956 22932 5012
rect 22764 4396 22820 4452
rect 23100 6018 23156 6020
rect 23100 5966 23102 6018
rect 23102 5966 23154 6018
rect 23154 5966 23156 6018
rect 23100 5964 23156 5966
rect 23324 5964 23380 6020
rect 23324 5628 23380 5684
rect 24444 7362 24500 7364
rect 24444 7310 24446 7362
rect 24446 7310 24498 7362
rect 24498 7310 24500 7362
rect 24444 7308 24500 7310
rect 23660 6524 23716 6580
rect 24332 6578 24388 6580
rect 24332 6526 24334 6578
rect 24334 6526 24386 6578
rect 24386 6526 24388 6578
rect 24332 6524 24388 6526
rect 23996 6412 24052 6468
rect 23100 5516 23156 5572
rect 23436 5068 23492 5124
rect 23548 5740 23604 5796
rect 23772 5292 23828 5348
rect 23996 4732 24052 4788
rect 24444 5794 24500 5796
rect 24444 5742 24446 5794
rect 24446 5742 24498 5794
rect 24498 5742 24500 5794
rect 24444 5740 24500 5742
rect 27916 8316 27972 8372
rect 27132 8146 27188 8148
rect 27132 8094 27134 8146
rect 27134 8094 27186 8146
rect 27186 8094 27188 8146
rect 27132 8092 27188 8094
rect 27580 8146 27636 8148
rect 27580 8094 27582 8146
rect 27582 8094 27634 8146
rect 27634 8094 27636 8146
rect 27580 8092 27636 8094
rect 26012 7980 26068 8036
rect 26012 7698 26068 7700
rect 26012 7646 26014 7698
rect 26014 7646 26066 7698
rect 26066 7646 26068 7698
rect 26012 7644 26068 7646
rect 27468 7868 27524 7924
rect 27132 7586 27188 7588
rect 27132 7534 27134 7586
rect 27134 7534 27186 7586
rect 27186 7534 27188 7586
rect 27132 7532 27188 7534
rect 26348 6412 26404 6468
rect 25676 6188 25732 6244
rect 24780 5740 24836 5796
rect 24220 5628 24276 5684
rect 25228 5682 25284 5684
rect 25228 5630 25230 5682
rect 25230 5630 25282 5682
rect 25282 5630 25284 5682
rect 25228 5628 25284 5630
rect 25452 5516 25508 5572
rect 24780 5292 24836 5348
rect 24668 5068 24724 5124
rect 24556 4732 24612 4788
rect 23884 4396 23940 4452
rect 24556 4172 24612 4228
rect 24892 5180 24948 5236
rect 25228 4172 25284 4228
rect 26572 6188 26628 6244
rect 26684 6412 26740 6468
rect 26236 5906 26292 5908
rect 26236 5854 26238 5906
rect 26238 5854 26290 5906
rect 26290 5854 26292 5906
rect 26236 5852 26292 5854
rect 25676 5516 25732 5572
rect 25676 4956 25732 5012
rect 25788 4844 25844 4900
rect 25788 4620 25844 4676
rect 26236 5628 26292 5684
rect 29148 9772 29204 9828
rect 30268 10556 30324 10612
rect 30380 12348 30436 12404
rect 29932 10332 29988 10388
rect 30156 10498 30212 10500
rect 30156 10446 30158 10498
rect 30158 10446 30210 10498
rect 30210 10446 30212 10498
rect 30156 10444 30212 10446
rect 29596 10220 29652 10276
rect 30156 10220 30212 10276
rect 30156 9996 30212 10052
rect 29260 9602 29316 9604
rect 29260 9550 29262 9602
rect 29262 9550 29314 9602
rect 29314 9550 29316 9602
rect 29260 9548 29316 9550
rect 28700 8652 28756 8708
rect 29932 8930 29988 8932
rect 29932 8878 29934 8930
rect 29934 8878 29986 8930
rect 29986 8878 29988 8930
rect 29932 8876 29988 8878
rect 29932 8428 29988 8484
rect 28700 8370 28756 8372
rect 28700 8318 28702 8370
rect 28702 8318 28754 8370
rect 28754 8318 28756 8370
rect 28700 8316 28756 8318
rect 30156 9714 30212 9716
rect 30156 9662 30158 9714
rect 30158 9662 30210 9714
rect 30210 9662 30212 9714
rect 30156 9660 30212 9662
rect 30044 8204 30100 8260
rect 29372 8092 29428 8148
rect 28924 7474 28980 7476
rect 28924 7422 28926 7474
rect 28926 7422 28978 7474
rect 28978 7422 28980 7474
rect 28924 7420 28980 7422
rect 27916 6860 27972 6916
rect 29596 7868 29652 7924
rect 29484 6300 29540 6356
rect 28700 5964 28756 6020
rect 29820 7980 29876 8036
rect 29820 7420 29876 7476
rect 29708 6690 29764 6692
rect 29708 6638 29710 6690
rect 29710 6638 29762 6690
rect 29762 6638 29764 6690
rect 29708 6636 29764 6638
rect 30044 7868 30100 7924
rect 30940 14700 30996 14756
rect 30716 14306 30772 14308
rect 30716 14254 30718 14306
rect 30718 14254 30770 14306
rect 30770 14254 30772 14306
rect 30716 14252 30772 14254
rect 30716 14028 30772 14084
rect 31276 14418 31332 14420
rect 31276 14366 31278 14418
rect 31278 14366 31330 14418
rect 31330 14366 31332 14418
rect 31276 14364 31332 14366
rect 31276 13858 31332 13860
rect 31276 13806 31278 13858
rect 31278 13806 31330 13858
rect 31330 13806 31332 13858
rect 31276 13804 31332 13806
rect 31164 13692 31220 13748
rect 31500 13468 31556 13524
rect 31164 13356 31220 13412
rect 30940 12178 30996 12180
rect 30940 12126 30942 12178
rect 30942 12126 30994 12178
rect 30994 12126 30996 12178
rect 30940 12124 30996 12126
rect 31052 11564 31108 11620
rect 31164 11900 31220 11956
rect 30604 11228 30660 11284
rect 30828 11340 30884 11396
rect 30604 11004 30660 11060
rect 30828 11170 30884 11172
rect 30828 11118 30830 11170
rect 30830 11118 30882 11170
rect 30882 11118 30884 11170
rect 30828 11116 30884 11118
rect 31164 10780 31220 10836
rect 31164 10610 31220 10612
rect 31164 10558 31166 10610
rect 31166 10558 31218 10610
rect 31218 10558 31220 10610
rect 31164 10556 31220 10558
rect 33292 14364 33348 14420
rect 33180 14140 33236 14196
rect 31724 14028 31780 14084
rect 32284 13580 32340 13636
rect 31724 12348 31780 12404
rect 31836 12290 31892 12292
rect 31836 12238 31838 12290
rect 31838 12238 31890 12290
rect 31890 12238 31892 12290
rect 31836 12236 31892 12238
rect 31948 11954 32004 11956
rect 31948 11902 31950 11954
rect 31950 11902 32002 11954
rect 32002 11902 32004 11954
rect 31948 11900 32004 11902
rect 32172 11900 32228 11956
rect 31836 11394 31892 11396
rect 31836 11342 31838 11394
rect 31838 11342 31890 11394
rect 31890 11342 31892 11394
rect 31836 11340 31892 11342
rect 31724 10834 31780 10836
rect 31724 10782 31726 10834
rect 31726 10782 31778 10834
rect 31778 10782 31780 10834
rect 31724 10780 31780 10782
rect 31388 10556 31444 10612
rect 32060 10556 32116 10612
rect 31052 10332 31108 10388
rect 31724 10332 31780 10388
rect 30828 9996 30884 10052
rect 30716 9826 30772 9828
rect 30716 9774 30718 9826
rect 30718 9774 30770 9826
rect 30770 9774 30772 9826
rect 30716 9772 30772 9774
rect 30716 8034 30772 8036
rect 30716 7982 30718 8034
rect 30718 7982 30770 8034
rect 30770 7982 30772 8034
rect 30716 7980 30772 7982
rect 31276 8428 31332 8484
rect 31612 8258 31668 8260
rect 31612 8206 31614 8258
rect 31614 8206 31666 8258
rect 31666 8206 31668 8258
rect 31612 8204 31668 8206
rect 31052 7868 31108 7924
rect 32284 8764 32340 8820
rect 32396 12012 32452 12068
rect 32508 11564 32564 11620
rect 32508 8764 32564 8820
rect 32508 8428 32564 8484
rect 31388 7532 31444 7588
rect 30380 6972 30436 7028
rect 30716 6300 30772 6356
rect 29708 6076 29764 6132
rect 26796 5906 26852 5908
rect 26796 5854 26798 5906
rect 26798 5854 26850 5906
rect 26850 5854 26852 5906
rect 26796 5852 26852 5854
rect 26684 5516 26740 5572
rect 26908 5740 26964 5796
rect 26796 5234 26852 5236
rect 26796 5182 26798 5234
rect 26798 5182 26850 5234
rect 26850 5182 26852 5234
rect 26796 5180 26852 5182
rect 26684 5122 26740 5124
rect 26684 5070 26686 5122
rect 26686 5070 26738 5122
rect 26738 5070 26740 5122
rect 26684 5068 26740 5070
rect 27580 5906 27636 5908
rect 27580 5854 27582 5906
rect 27582 5854 27634 5906
rect 27634 5854 27636 5906
rect 27580 5852 27636 5854
rect 28028 5852 28084 5908
rect 27020 5516 27076 5572
rect 27804 5068 27860 5124
rect 28588 5906 28644 5908
rect 28588 5854 28590 5906
rect 28590 5854 28642 5906
rect 28642 5854 28644 5906
rect 28588 5852 28644 5854
rect 29372 5740 29428 5796
rect 29260 5628 29316 5684
rect 29148 5404 29204 5460
rect 28140 5292 28196 5348
rect 29484 5122 29540 5124
rect 29484 5070 29486 5122
rect 29486 5070 29538 5122
rect 29538 5070 29540 5122
rect 29484 5068 29540 5070
rect 29820 5404 29876 5460
rect 31164 6018 31220 6020
rect 31164 5966 31166 6018
rect 31166 5966 31218 6018
rect 31218 5966 31220 6018
rect 31164 5964 31220 5966
rect 31388 5964 31444 6020
rect 30380 5682 30436 5684
rect 30380 5630 30382 5682
rect 30382 5630 30434 5682
rect 30434 5630 30436 5682
rect 30380 5628 30436 5630
rect 31724 6524 31780 6580
rect 31724 5740 31780 5796
rect 31612 5068 31668 5124
rect 30380 4956 30436 5012
rect 30268 4508 30324 4564
rect 29596 3724 29652 3780
rect 25900 3500 25956 3556
rect 26236 3612 26292 3668
rect 29372 3666 29428 3668
rect 29372 3614 29374 3666
rect 29374 3614 29426 3666
rect 29426 3614 29428 3666
rect 29372 3612 29428 3614
rect 28588 3554 28644 3556
rect 28588 3502 28590 3554
rect 28590 3502 28642 3554
rect 28642 3502 28644 3554
rect 28588 3500 28644 3502
rect 30940 3724 30996 3780
rect 30268 3500 30324 3556
rect 31836 5516 31892 5572
rect 31276 4898 31332 4900
rect 31276 4846 31278 4898
rect 31278 4846 31330 4898
rect 31330 4846 31332 4898
rect 31276 4844 31332 4846
rect 32620 8034 32676 8036
rect 32620 7982 32622 8034
rect 32622 7982 32674 8034
rect 32674 7982 32676 8034
rect 32620 7980 32676 7982
rect 33404 13746 33460 13748
rect 33404 13694 33406 13746
rect 33406 13694 33458 13746
rect 33458 13694 33460 13746
rect 33404 13692 33460 13694
rect 33292 12460 33348 12516
rect 33292 12066 33348 12068
rect 33292 12014 33294 12066
rect 33294 12014 33346 12066
rect 33346 12014 33348 12066
rect 33292 12012 33348 12014
rect 33180 10610 33236 10612
rect 33180 10558 33182 10610
rect 33182 10558 33234 10610
rect 33234 10558 33236 10610
rect 33180 10556 33236 10558
rect 34188 19068 34244 19124
rect 33964 16940 34020 16996
rect 33852 16716 33908 16772
rect 33852 16268 33908 16324
rect 33852 15484 33908 15540
rect 34860 19122 34916 19124
rect 34860 19070 34862 19122
rect 34862 19070 34914 19122
rect 34914 19070 34916 19122
rect 34860 19068 34916 19070
rect 34300 18732 34356 18788
rect 35420 19122 35476 19124
rect 35420 19070 35422 19122
rect 35422 19070 35474 19122
rect 35474 19070 35476 19122
rect 35420 19068 35476 19070
rect 36764 19068 36820 19124
rect 36428 18732 36484 18788
rect 35308 18508 35364 18564
rect 36204 18508 36260 18564
rect 35196 18058 35252 18060
rect 34412 17948 34468 18004
rect 35196 18006 35198 18058
rect 35198 18006 35250 18058
rect 35250 18006 35252 18058
rect 35196 18004 35252 18006
rect 35300 18058 35356 18060
rect 35300 18006 35302 18058
rect 35302 18006 35354 18058
rect 35354 18006 35356 18058
rect 35300 18004 35356 18006
rect 35404 18058 35460 18060
rect 35404 18006 35406 18058
rect 35406 18006 35458 18058
rect 35458 18006 35460 18058
rect 35404 18004 35460 18006
rect 36204 18060 36260 18116
rect 34972 17442 35028 17444
rect 34972 17390 34974 17442
rect 34974 17390 35026 17442
rect 35026 17390 35028 17442
rect 34972 17388 35028 17390
rect 34636 17052 34692 17108
rect 34188 16716 34244 16772
rect 34300 16098 34356 16100
rect 34300 16046 34302 16098
rect 34302 16046 34354 16098
rect 34354 16046 34356 16098
rect 34300 16044 34356 16046
rect 34972 16994 35028 16996
rect 34972 16942 34974 16994
rect 34974 16942 35026 16994
rect 35026 16942 35028 16994
rect 34972 16940 35028 16942
rect 34860 16828 34916 16884
rect 34860 16044 34916 16100
rect 36428 18284 36484 18340
rect 35644 17554 35700 17556
rect 35644 17502 35646 17554
rect 35646 17502 35698 17554
rect 35698 17502 35700 17554
rect 35644 17500 35700 17502
rect 35532 17388 35588 17444
rect 35420 17106 35476 17108
rect 35420 17054 35422 17106
rect 35422 17054 35474 17106
rect 35474 17054 35476 17106
rect 35420 17052 35476 17054
rect 35196 16490 35252 16492
rect 35196 16438 35198 16490
rect 35198 16438 35250 16490
rect 35250 16438 35252 16490
rect 35196 16436 35252 16438
rect 35300 16490 35356 16492
rect 35300 16438 35302 16490
rect 35302 16438 35354 16490
rect 35354 16438 35356 16490
rect 35300 16436 35356 16438
rect 35404 16490 35460 16492
rect 35404 16438 35406 16490
rect 35406 16438 35458 16490
rect 35458 16438 35460 16490
rect 35404 16436 35460 16438
rect 35196 16098 35252 16100
rect 35196 16046 35198 16098
rect 35198 16046 35250 16098
rect 35250 16046 35252 16098
rect 35196 16044 35252 16046
rect 34188 15820 34244 15876
rect 34412 15596 34468 15652
rect 34300 14700 34356 14756
rect 34524 15538 34580 15540
rect 34524 15486 34526 15538
rect 34526 15486 34578 15538
rect 34578 15486 34580 15538
rect 34524 15484 34580 15486
rect 36540 17164 36596 17220
rect 36652 18396 36708 18452
rect 36540 16994 36596 16996
rect 36540 16942 36542 16994
rect 36542 16942 36594 16994
rect 36594 16942 36596 16994
rect 36540 16940 36596 16942
rect 34972 15596 35028 15652
rect 35756 15596 35812 15652
rect 35868 15820 35924 15876
rect 36092 15260 36148 15316
rect 35196 14922 35252 14924
rect 35196 14870 35198 14922
rect 35198 14870 35250 14922
rect 35250 14870 35252 14922
rect 35196 14868 35252 14870
rect 35300 14922 35356 14924
rect 35300 14870 35302 14922
rect 35302 14870 35354 14922
rect 35354 14870 35356 14922
rect 35300 14868 35356 14870
rect 35404 14922 35460 14924
rect 35404 14870 35406 14922
rect 35406 14870 35458 14922
rect 35458 14870 35460 14922
rect 35404 14868 35460 14870
rect 35644 14812 35700 14868
rect 34636 14252 34692 14308
rect 33964 13746 34020 13748
rect 33964 13694 33966 13746
rect 33966 13694 34018 13746
rect 34018 13694 34020 13746
rect 33964 13692 34020 13694
rect 34300 13692 34356 13748
rect 33740 12066 33796 12068
rect 33740 12014 33742 12066
rect 33742 12014 33794 12066
rect 33794 12014 33796 12066
rect 33740 12012 33796 12014
rect 35644 13916 35700 13972
rect 35756 14700 35812 14756
rect 34636 13468 34692 13524
rect 34412 12796 34468 12852
rect 33852 11116 33908 11172
rect 33292 9324 33348 9380
rect 34076 10556 34132 10612
rect 33740 9996 33796 10052
rect 35196 13354 35252 13356
rect 35196 13302 35198 13354
rect 35198 13302 35250 13354
rect 35250 13302 35252 13354
rect 35196 13300 35252 13302
rect 35300 13354 35356 13356
rect 35300 13302 35302 13354
rect 35302 13302 35354 13354
rect 35354 13302 35356 13354
rect 35300 13300 35356 13302
rect 35404 13354 35460 13356
rect 35404 13302 35406 13354
rect 35406 13302 35458 13354
rect 35458 13302 35460 13354
rect 35404 13300 35460 13302
rect 35420 13186 35476 13188
rect 35420 13134 35422 13186
rect 35422 13134 35474 13186
rect 35474 13134 35476 13186
rect 35420 13132 35476 13134
rect 35868 13522 35924 13524
rect 35868 13470 35870 13522
rect 35870 13470 35922 13522
rect 35922 13470 35924 13522
rect 35868 13468 35924 13470
rect 35980 13356 36036 13412
rect 34972 12796 35028 12852
rect 36092 13916 36148 13972
rect 34748 12124 34804 12180
rect 35532 12178 35588 12180
rect 35532 12126 35534 12178
rect 35534 12126 35586 12178
rect 35586 12126 35588 12178
rect 35532 12124 35588 12126
rect 35084 12066 35140 12068
rect 35084 12014 35086 12066
rect 35086 12014 35138 12066
rect 35138 12014 35140 12066
rect 35084 12012 35140 12014
rect 35196 11786 35252 11788
rect 35196 11734 35198 11786
rect 35198 11734 35250 11786
rect 35250 11734 35252 11786
rect 35196 11732 35252 11734
rect 35300 11786 35356 11788
rect 35300 11734 35302 11786
rect 35302 11734 35354 11786
rect 35354 11734 35356 11786
rect 35300 11732 35356 11734
rect 35404 11786 35460 11788
rect 35404 11734 35406 11786
rect 35406 11734 35458 11786
rect 35458 11734 35460 11786
rect 35404 11732 35460 11734
rect 35084 11506 35140 11508
rect 35084 11454 35086 11506
rect 35086 11454 35138 11506
rect 35138 11454 35140 11506
rect 35084 11452 35140 11454
rect 35532 11116 35588 11172
rect 35644 11900 35700 11956
rect 35196 10218 35252 10220
rect 35196 10166 35198 10218
rect 35198 10166 35250 10218
rect 35250 10166 35252 10218
rect 35196 10164 35252 10166
rect 35300 10218 35356 10220
rect 35300 10166 35302 10218
rect 35302 10166 35354 10218
rect 35354 10166 35356 10218
rect 35300 10164 35356 10166
rect 35404 10218 35460 10220
rect 35404 10166 35406 10218
rect 35406 10166 35458 10218
rect 35458 10166 35460 10218
rect 35404 10164 35460 10166
rect 36540 14812 36596 14868
rect 36316 14476 36372 14532
rect 36428 13692 36484 13748
rect 36204 11676 36260 11732
rect 36316 12012 36372 12068
rect 36204 11506 36260 11508
rect 36204 11454 36206 11506
rect 36206 11454 36258 11506
rect 36258 11454 36260 11506
rect 36204 11452 36260 11454
rect 35980 11116 36036 11172
rect 35868 10220 35924 10276
rect 34300 9266 34356 9268
rect 34300 9214 34302 9266
rect 34302 9214 34354 9266
rect 34354 9214 34356 9266
rect 34300 9212 34356 9214
rect 33964 8370 34020 8372
rect 33964 8318 33966 8370
rect 33966 8318 34018 8370
rect 34018 8318 34020 8370
rect 33964 8316 34020 8318
rect 36092 9996 36148 10052
rect 34636 9660 34692 9716
rect 36876 21420 36932 21476
rect 38444 23436 38500 23492
rect 37884 23324 37940 23380
rect 37996 23042 38052 23044
rect 37996 22990 37998 23042
rect 37998 22990 38050 23042
rect 38050 22990 38052 23042
rect 37996 22988 38052 22990
rect 37884 22316 37940 22372
rect 38108 22146 38164 22148
rect 38108 22094 38110 22146
rect 38110 22094 38162 22146
rect 38162 22094 38164 22146
rect 38108 22092 38164 22094
rect 38444 22146 38500 22148
rect 38444 22094 38446 22146
rect 38446 22094 38498 22146
rect 38498 22094 38500 22146
rect 38444 22092 38500 22094
rect 39676 22876 39732 22932
rect 40348 24444 40404 24500
rect 40012 23826 40068 23828
rect 40012 23774 40014 23826
rect 40014 23774 40066 23826
rect 40066 23774 40068 23826
rect 40012 23772 40068 23774
rect 39900 22988 39956 23044
rect 40012 23324 40068 23380
rect 38892 21980 38948 22036
rect 39004 21698 39060 21700
rect 39004 21646 39006 21698
rect 39006 21646 39058 21698
rect 39058 21646 39060 21698
rect 39004 21644 39060 21646
rect 37660 21420 37716 21476
rect 37212 20972 37268 21028
rect 38332 21308 38388 21364
rect 37660 20914 37716 20916
rect 37660 20862 37662 20914
rect 37662 20862 37714 20914
rect 37714 20862 37716 20914
rect 37660 20860 37716 20862
rect 38444 20972 38500 21028
rect 37212 18508 37268 18564
rect 37660 18844 37716 18900
rect 37100 18450 37156 18452
rect 37100 18398 37102 18450
rect 37102 18398 37154 18450
rect 37154 18398 37156 18450
rect 37100 18396 37156 18398
rect 37324 18060 37380 18116
rect 37212 16268 37268 16324
rect 37212 16098 37268 16100
rect 37212 16046 37214 16098
rect 37214 16046 37266 16098
rect 37266 16046 37268 16098
rect 37212 16044 37268 16046
rect 37324 15484 37380 15540
rect 37548 17164 37604 17220
rect 37548 16492 37604 16548
rect 39564 22204 39620 22260
rect 39788 22258 39844 22260
rect 39788 22206 39790 22258
rect 39790 22206 39842 22258
rect 39842 22206 39844 22258
rect 39788 22204 39844 22206
rect 40012 22316 40068 22372
rect 40124 23212 40180 23268
rect 38444 18172 38500 18228
rect 38668 20412 38724 20468
rect 39004 20076 39060 20132
rect 39228 19852 39284 19908
rect 40012 21868 40068 21924
rect 40012 20748 40068 20804
rect 39900 19740 39956 19796
rect 40012 19964 40068 20020
rect 39900 19346 39956 19348
rect 39900 19294 39902 19346
rect 39902 19294 39954 19346
rect 39954 19294 39956 19346
rect 39900 19292 39956 19294
rect 37884 17164 37940 17220
rect 39228 17500 39284 17556
rect 38220 16940 38276 16996
rect 38444 17388 38500 17444
rect 38108 16268 38164 16324
rect 37996 15596 38052 15652
rect 37772 15538 37828 15540
rect 37772 15486 37774 15538
rect 37774 15486 37826 15538
rect 37826 15486 37828 15538
rect 37772 15484 37828 15486
rect 38220 15874 38276 15876
rect 38220 15822 38222 15874
rect 38222 15822 38274 15874
rect 38274 15822 38276 15874
rect 38220 15820 38276 15822
rect 38668 17276 38724 17332
rect 39004 16994 39060 16996
rect 39004 16942 39006 16994
rect 39006 16942 39058 16994
rect 39058 16942 39060 16994
rect 39004 16940 39060 16942
rect 40572 25340 40628 25396
rect 40908 26178 40964 26180
rect 40908 26126 40910 26178
rect 40910 26126 40962 26178
rect 40962 26126 40964 26178
rect 40908 26124 40964 26126
rect 40796 25228 40852 25284
rect 43484 29932 43540 29988
rect 43484 28924 43540 28980
rect 43372 28588 43428 28644
rect 43260 28252 43316 28308
rect 43372 26796 43428 26852
rect 41916 26178 41972 26180
rect 41916 26126 41918 26178
rect 41918 26126 41970 26178
rect 41970 26126 41972 26178
rect 41916 26124 41972 26126
rect 43260 26124 43316 26180
rect 41244 25452 41300 25508
rect 41692 25452 41748 25508
rect 40684 24444 40740 24500
rect 41132 24668 41188 24724
rect 41020 24610 41076 24612
rect 41020 24558 41022 24610
rect 41022 24558 41074 24610
rect 41074 24558 41076 24610
rect 41020 24556 41076 24558
rect 40796 23324 40852 23380
rect 42364 25506 42420 25508
rect 42364 25454 42366 25506
rect 42366 25454 42418 25506
rect 42418 25454 42420 25506
rect 42364 25452 42420 25454
rect 43036 25340 43092 25396
rect 43148 25228 43204 25284
rect 41804 24780 41860 24836
rect 42700 24780 42756 24836
rect 42476 24722 42532 24724
rect 42476 24670 42478 24722
rect 42478 24670 42530 24722
rect 42530 24670 42532 24722
rect 42476 24668 42532 24670
rect 42140 24498 42196 24500
rect 42140 24446 42142 24498
rect 42142 24446 42194 24498
rect 42194 24446 42196 24498
rect 42140 24444 42196 24446
rect 40908 22930 40964 22932
rect 40908 22878 40910 22930
rect 40910 22878 40962 22930
rect 40962 22878 40964 22930
rect 40908 22876 40964 22878
rect 41244 22930 41300 22932
rect 41244 22878 41246 22930
rect 41246 22878 41298 22930
rect 41298 22878 41300 22930
rect 41244 22876 41300 22878
rect 40572 22370 40628 22372
rect 40572 22318 40574 22370
rect 40574 22318 40626 22370
rect 40626 22318 40628 22370
rect 40572 22316 40628 22318
rect 40796 22258 40852 22260
rect 40796 22206 40798 22258
rect 40798 22206 40850 22258
rect 40850 22206 40852 22258
rect 40796 22204 40852 22206
rect 41916 23772 41972 23828
rect 41804 23436 41860 23492
rect 42364 23436 42420 23492
rect 42028 23100 42084 23156
rect 43820 28866 43876 28868
rect 43820 28814 43822 28866
rect 43822 28814 43874 28866
rect 43874 28814 43876 28866
rect 43820 28812 43876 28814
rect 44156 34242 44212 34244
rect 44156 34190 44158 34242
rect 44158 34190 44210 34242
rect 44210 34190 44212 34242
rect 44156 34188 44212 34190
rect 48300 43708 48356 43764
rect 48188 43036 48244 43092
rect 48188 42754 48244 42756
rect 48188 42702 48190 42754
rect 48190 42702 48242 42754
rect 48242 42702 48244 42754
rect 48188 42700 48244 42702
rect 48188 42364 48244 42420
rect 48188 37996 48244 38052
rect 47068 35644 47124 35700
rect 45836 35196 45892 35252
rect 45052 34972 45108 35028
rect 44940 34802 44996 34804
rect 44940 34750 44942 34802
rect 44942 34750 44994 34802
rect 44994 34750 44996 34802
rect 44940 34748 44996 34750
rect 44604 34636 44660 34692
rect 44268 33964 44324 34020
rect 45164 34636 45220 34692
rect 45276 33404 45332 33460
rect 45612 32562 45668 32564
rect 45612 32510 45614 32562
rect 45614 32510 45666 32562
rect 45666 32510 45668 32562
rect 45612 32508 45668 32510
rect 46060 33458 46116 33460
rect 46060 33406 46062 33458
rect 46062 33406 46114 33458
rect 46114 33406 46116 33458
rect 46060 33404 46116 33406
rect 45276 30940 45332 30996
rect 45388 30210 45444 30212
rect 45388 30158 45390 30210
rect 45390 30158 45442 30210
rect 45442 30158 45444 30210
rect 45388 30156 45444 30158
rect 44044 29932 44100 29988
rect 44940 29986 44996 29988
rect 44940 29934 44942 29986
rect 44942 29934 44994 29986
rect 44994 29934 44996 29986
rect 44940 29932 44996 29934
rect 45836 31724 45892 31780
rect 46284 30268 46340 30324
rect 46060 29708 46116 29764
rect 43932 27916 43988 27972
rect 43372 25564 43428 25620
rect 43484 25228 43540 25284
rect 44044 25564 44100 25620
rect 43708 25004 43764 25060
rect 43820 24780 43876 24836
rect 43036 24332 43092 24388
rect 42588 23772 42644 23828
rect 43148 23772 43204 23828
rect 43596 23826 43652 23828
rect 43596 23774 43598 23826
rect 43598 23774 43650 23826
rect 43650 23774 43652 23826
rect 43596 23772 43652 23774
rect 44044 24220 44100 24276
rect 42812 23100 42868 23156
rect 42924 23212 42980 23268
rect 44044 23436 44100 23492
rect 43484 23100 43540 23156
rect 43148 22876 43204 22932
rect 42252 22258 42308 22260
rect 42252 22206 42254 22258
rect 42254 22206 42306 22258
rect 42306 22206 42308 22258
rect 42252 22204 42308 22206
rect 42140 21810 42196 21812
rect 42140 21758 42142 21810
rect 42142 21758 42194 21810
rect 42194 21758 42196 21810
rect 42140 21756 42196 21758
rect 43484 21980 43540 22036
rect 42812 21756 42868 21812
rect 43260 21756 43316 21812
rect 41916 21196 41972 21252
rect 41244 20130 41300 20132
rect 41244 20078 41246 20130
rect 41246 20078 41298 20130
rect 41298 20078 41300 20130
rect 41244 20076 41300 20078
rect 39900 18450 39956 18452
rect 39900 18398 39902 18450
rect 39902 18398 39954 18450
rect 39954 18398 39956 18450
rect 39900 18396 39956 18398
rect 40460 18674 40516 18676
rect 40460 18622 40462 18674
rect 40462 18622 40514 18674
rect 40514 18622 40516 18674
rect 40460 18620 40516 18622
rect 39452 16940 39508 16996
rect 39116 16828 39172 16884
rect 38668 16322 38724 16324
rect 38668 16270 38670 16322
rect 38670 16270 38722 16322
rect 38722 16270 38724 16322
rect 38668 16268 38724 16270
rect 38444 15820 38500 15876
rect 38332 15484 38388 15540
rect 36876 15314 36932 15316
rect 36876 15262 36878 15314
rect 36878 15262 36930 15314
rect 36930 15262 36932 15314
rect 36876 15260 36932 15262
rect 37548 14476 37604 14532
rect 37884 14364 37940 14420
rect 38444 14306 38500 14308
rect 38444 14254 38446 14306
rect 38446 14254 38498 14306
rect 38498 14254 38500 14306
rect 38444 14252 38500 14254
rect 39116 14924 39172 14980
rect 39004 14530 39060 14532
rect 39004 14478 39006 14530
rect 39006 14478 39058 14530
rect 39058 14478 39060 14530
rect 39004 14476 39060 14478
rect 37884 13970 37940 13972
rect 37884 13918 37886 13970
rect 37886 13918 37938 13970
rect 37938 13918 37940 13970
rect 37884 13916 37940 13918
rect 36876 13746 36932 13748
rect 36876 13694 36878 13746
rect 36878 13694 36930 13746
rect 36930 13694 36932 13746
rect 36876 13692 36932 13694
rect 38556 13746 38612 13748
rect 38556 13694 38558 13746
rect 38558 13694 38610 13746
rect 38610 13694 38612 13746
rect 38556 13692 38612 13694
rect 37212 13356 37268 13412
rect 37660 13356 37716 13412
rect 36764 13020 36820 13076
rect 39564 16380 39620 16436
rect 39900 16994 39956 16996
rect 39900 16942 39902 16994
rect 39902 16942 39954 16994
rect 39954 16942 39956 16994
rect 39900 16940 39956 16942
rect 39900 16604 39956 16660
rect 40348 18450 40404 18452
rect 40348 18398 40350 18450
rect 40350 18398 40402 18450
rect 40402 18398 40404 18450
rect 40348 18396 40404 18398
rect 40572 18060 40628 18116
rect 40236 17836 40292 17892
rect 40348 17666 40404 17668
rect 40348 17614 40350 17666
rect 40350 17614 40402 17666
rect 40402 17614 40404 17666
rect 40348 17612 40404 17614
rect 40460 17276 40516 17332
rect 40572 17500 40628 17556
rect 40236 17164 40292 17220
rect 40124 16156 40180 16212
rect 40348 16268 40404 16324
rect 41020 19852 41076 19908
rect 42028 20860 42084 20916
rect 42140 20636 42196 20692
rect 42476 20018 42532 20020
rect 42476 19966 42478 20018
rect 42478 19966 42530 20018
rect 42530 19966 42532 20018
rect 42476 19964 42532 19966
rect 41244 19628 41300 19684
rect 43596 21756 43652 21812
rect 44828 28418 44884 28420
rect 44828 28366 44830 28418
rect 44830 28366 44882 28418
rect 44882 28366 44884 28418
rect 44828 28364 44884 28366
rect 45164 28028 45220 28084
rect 45612 28812 45668 28868
rect 45500 28252 45556 28308
rect 47852 35644 47908 35700
rect 47964 34300 48020 34356
rect 47404 33628 47460 33684
rect 47180 31948 47236 32004
rect 47068 29596 47124 29652
rect 45612 27244 45668 27300
rect 46620 27970 46676 27972
rect 46620 27918 46622 27970
rect 46622 27918 46674 27970
rect 46674 27918 46676 27970
rect 46620 27916 46676 27918
rect 45276 27132 45332 27188
rect 46060 27186 46116 27188
rect 46060 27134 46062 27186
rect 46062 27134 46114 27186
rect 46114 27134 46116 27186
rect 46060 27132 46116 27134
rect 44268 26850 44324 26852
rect 44268 26798 44270 26850
rect 44270 26798 44322 26850
rect 44322 26798 44324 26850
rect 44268 26796 44324 26798
rect 44716 26290 44772 26292
rect 44716 26238 44718 26290
rect 44718 26238 44770 26290
rect 44770 26238 44772 26290
rect 44716 26236 44772 26238
rect 47404 29932 47460 29988
rect 48188 32284 48244 32340
rect 47740 28924 47796 28980
rect 47628 28082 47684 28084
rect 47628 28030 47630 28082
rect 47630 28030 47682 28082
rect 47682 28030 47684 28082
rect 47628 28028 47684 28030
rect 47964 28252 48020 28308
rect 47852 28028 47908 28084
rect 45388 26236 45444 26292
rect 45612 25900 45668 25956
rect 44604 25340 44660 25396
rect 45276 25004 45332 25060
rect 45164 24892 45220 24948
rect 44940 24834 44996 24836
rect 44940 24782 44942 24834
rect 44942 24782 44994 24834
rect 44994 24782 44996 24834
rect 44940 24780 44996 24782
rect 44940 23996 44996 24052
rect 44380 23324 44436 23380
rect 44380 22482 44436 22484
rect 44380 22430 44382 22482
rect 44382 22430 44434 22482
rect 44434 22430 44436 22482
rect 44380 22428 44436 22430
rect 46060 25394 46116 25396
rect 46060 25342 46062 25394
rect 46062 25342 46114 25394
rect 46114 25342 46116 25394
rect 46060 25340 46116 25342
rect 45724 24780 45780 24836
rect 45612 23938 45668 23940
rect 45612 23886 45614 23938
rect 45614 23886 45666 23938
rect 45666 23886 45668 23938
rect 45612 23884 45668 23886
rect 45388 23212 45444 23268
rect 47964 25564 48020 25620
rect 47404 25004 47460 25060
rect 46508 23378 46564 23380
rect 46508 23326 46510 23378
rect 46510 23326 46562 23378
rect 46562 23326 46564 23378
rect 46508 23324 46564 23326
rect 46844 23212 46900 23268
rect 47404 23660 47460 23716
rect 46956 22876 47012 22932
rect 46284 22428 46340 22484
rect 47068 22428 47124 22484
rect 47180 23212 47236 23268
rect 44156 21532 44212 21588
rect 43260 21196 43316 21252
rect 43148 20860 43204 20916
rect 42700 19628 42756 19684
rect 41020 19180 41076 19236
rect 41692 19234 41748 19236
rect 41692 19182 41694 19234
rect 41694 19182 41746 19234
rect 41746 19182 41748 19234
rect 41692 19180 41748 19182
rect 41356 18620 41412 18676
rect 40908 17388 40964 17444
rect 41132 17164 41188 17220
rect 40796 16940 40852 16996
rect 40908 16882 40964 16884
rect 40908 16830 40910 16882
rect 40910 16830 40962 16882
rect 40962 16830 40964 16882
rect 40908 16828 40964 16830
rect 41356 17106 41412 17108
rect 41356 17054 41358 17106
rect 41358 17054 41410 17106
rect 41410 17054 41412 17106
rect 41356 17052 41412 17054
rect 42924 20690 42980 20692
rect 42924 20638 42926 20690
rect 42926 20638 42978 20690
rect 42978 20638 42980 20690
rect 42924 20636 42980 20638
rect 43708 20130 43764 20132
rect 43708 20078 43710 20130
rect 43710 20078 43762 20130
rect 43762 20078 43764 20130
rect 43708 20076 43764 20078
rect 43372 19740 43428 19796
rect 45276 22204 45332 22260
rect 45052 21308 45108 21364
rect 46060 22258 46116 22260
rect 46060 22206 46062 22258
rect 46062 22206 46114 22258
rect 46114 22206 46116 22258
rect 46060 22204 46116 22206
rect 45612 22092 45668 22148
rect 45388 21980 45444 22036
rect 45388 21756 45444 21812
rect 44156 20188 44212 20244
rect 45052 20188 45108 20244
rect 42588 19180 42644 19236
rect 42476 18620 42532 18676
rect 43484 18620 43540 18676
rect 43708 19628 43764 19684
rect 42252 18508 42308 18564
rect 43260 18450 43316 18452
rect 43260 18398 43262 18450
rect 43262 18398 43314 18450
rect 43314 18398 43316 18450
rect 43260 18396 43316 18398
rect 42028 17724 42084 17780
rect 41132 16882 41188 16884
rect 41132 16830 41134 16882
rect 41134 16830 41186 16882
rect 41186 16830 41188 16882
rect 41132 16828 41188 16830
rect 42140 18172 42196 18228
rect 42700 18226 42756 18228
rect 42700 18174 42702 18226
rect 42702 18174 42754 18226
rect 42754 18174 42756 18226
rect 42700 18172 42756 18174
rect 42700 17778 42756 17780
rect 42700 17726 42702 17778
rect 42702 17726 42754 17778
rect 42754 17726 42756 17778
rect 42700 17724 42756 17726
rect 42364 17554 42420 17556
rect 42364 17502 42366 17554
rect 42366 17502 42418 17554
rect 42418 17502 42420 17554
rect 42364 17500 42420 17502
rect 42700 17500 42756 17556
rect 41916 16828 41972 16884
rect 40796 16716 40852 16772
rect 40684 16604 40740 16660
rect 41020 16268 41076 16324
rect 42812 17164 42868 17220
rect 43484 18172 43540 18228
rect 43708 17836 43764 17892
rect 43708 17612 43764 17668
rect 43260 17052 43316 17108
rect 44268 19010 44324 19012
rect 44268 18958 44270 19010
rect 44270 18958 44322 19010
rect 44322 18958 44324 19010
rect 44268 18956 44324 18958
rect 46060 21980 46116 22036
rect 47964 23548 48020 23604
rect 48188 23212 48244 23268
rect 48300 23660 48356 23716
rect 47964 22204 48020 22260
rect 47516 21532 47572 21588
rect 46956 21362 47012 21364
rect 46956 21310 46958 21362
rect 46958 21310 47010 21362
rect 47010 21310 47012 21362
rect 46956 21308 47012 21310
rect 48300 21532 48356 21588
rect 47516 20860 47572 20916
rect 46620 20748 46676 20804
rect 44380 17948 44436 18004
rect 44716 18396 44772 18452
rect 44044 17724 44100 17780
rect 44044 17164 44100 17220
rect 43708 17106 43764 17108
rect 43708 17054 43710 17106
rect 43710 17054 43762 17106
rect 43762 17054 43764 17106
rect 43708 17052 43764 17054
rect 42700 16940 42756 16996
rect 40012 15986 40068 15988
rect 40012 15934 40014 15986
rect 40014 15934 40066 15986
rect 40066 15934 40068 15986
rect 40012 15932 40068 15934
rect 39788 15820 39844 15876
rect 40236 15874 40292 15876
rect 40236 15822 40238 15874
rect 40238 15822 40290 15874
rect 40290 15822 40292 15874
rect 40236 15820 40292 15822
rect 40012 15538 40068 15540
rect 40012 15486 40014 15538
rect 40014 15486 40066 15538
rect 40066 15486 40068 15538
rect 40012 15484 40068 15486
rect 39676 15260 39732 15316
rect 39340 14476 39396 14532
rect 39564 14588 39620 14644
rect 37772 12684 37828 12740
rect 37100 12290 37156 12292
rect 37100 12238 37102 12290
rect 37102 12238 37154 12290
rect 37154 12238 37156 12290
rect 37100 12236 37156 12238
rect 36540 11676 36596 11732
rect 34524 8876 34580 8932
rect 34524 8204 34580 8260
rect 32732 7868 32788 7924
rect 33404 7420 33460 7476
rect 32284 6860 32340 6916
rect 32172 6802 32228 6804
rect 32172 6750 32174 6802
rect 32174 6750 32226 6802
rect 32226 6750 32228 6802
rect 32172 6748 32228 6750
rect 33068 6860 33124 6916
rect 32956 6802 33012 6804
rect 32956 6750 32958 6802
rect 32958 6750 33010 6802
rect 33010 6750 33012 6802
rect 32956 6748 33012 6750
rect 32060 6300 32116 6356
rect 32060 6018 32116 6020
rect 32060 5966 32062 6018
rect 32062 5966 32114 6018
rect 32114 5966 32116 6018
rect 32060 5964 32116 5966
rect 31836 4844 31892 4900
rect 31500 4732 31556 4788
rect 30940 3388 30996 3444
rect 31724 4732 31780 4788
rect 32620 5628 32676 5684
rect 33180 6130 33236 6132
rect 33180 6078 33182 6130
rect 33182 6078 33234 6130
rect 33234 6078 33236 6130
rect 33180 6076 33236 6078
rect 34636 6690 34692 6692
rect 34636 6638 34638 6690
rect 34638 6638 34690 6690
rect 34690 6638 34692 6690
rect 34636 6636 34692 6638
rect 33740 6524 33796 6580
rect 35196 9324 35252 9380
rect 35196 8764 35252 8820
rect 35196 8650 35252 8652
rect 35196 8598 35198 8650
rect 35198 8598 35250 8650
rect 35250 8598 35252 8650
rect 35196 8596 35252 8598
rect 35300 8650 35356 8652
rect 35300 8598 35302 8650
rect 35302 8598 35354 8650
rect 35354 8598 35356 8650
rect 35300 8596 35356 8598
rect 35404 8650 35460 8652
rect 35404 8598 35406 8650
rect 35406 8598 35458 8650
rect 35458 8598 35460 8650
rect 35404 8596 35460 8598
rect 35644 8652 35700 8708
rect 34860 6412 34916 6468
rect 33852 5852 33908 5908
rect 33852 5292 33908 5348
rect 33068 4956 33124 5012
rect 32396 4396 32452 4452
rect 32284 3554 32340 3556
rect 32284 3502 32286 3554
rect 32286 3502 32338 3554
rect 32338 3502 32340 3554
rect 32284 3500 32340 3502
rect 32956 3612 33012 3668
rect 34524 5906 34580 5908
rect 34524 5854 34526 5906
rect 34526 5854 34578 5906
rect 34578 5854 34580 5906
rect 34524 5852 34580 5854
rect 34860 5682 34916 5684
rect 34860 5630 34862 5682
rect 34862 5630 34914 5682
rect 34914 5630 34916 5682
rect 34860 5628 34916 5630
rect 34188 4620 34244 4676
rect 34076 4562 34132 4564
rect 34076 4510 34078 4562
rect 34078 4510 34130 4562
rect 34130 4510 34132 4562
rect 34076 4508 34132 4510
rect 34636 4956 34692 5012
rect 33964 4450 34020 4452
rect 33964 4398 33966 4450
rect 33966 4398 34018 4450
rect 34018 4398 34020 4450
rect 33964 4396 34020 4398
rect 34972 4732 35028 4788
rect 33852 3666 33908 3668
rect 33852 3614 33854 3666
rect 33854 3614 33906 3666
rect 33906 3614 33908 3666
rect 33852 3612 33908 3614
rect 33628 3500 33684 3556
rect 35420 7474 35476 7476
rect 35420 7422 35422 7474
rect 35422 7422 35474 7474
rect 35474 7422 35476 7474
rect 35420 7420 35476 7422
rect 35196 7082 35252 7084
rect 35196 7030 35198 7082
rect 35198 7030 35250 7082
rect 35250 7030 35252 7082
rect 35196 7028 35252 7030
rect 35300 7082 35356 7084
rect 35300 7030 35302 7082
rect 35302 7030 35354 7082
rect 35354 7030 35356 7082
rect 35300 7028 35356 7030
rect 35404 7082 35460 7084
rect 35404 7030 35406 7082
rect 35406 7030 35458 7082
rect 35458 7030 35460 7082
rect 35404 7028 35460 7030
rect 35308 6914 35364 6916
rect 35308 6862 35310 6914
rect 35310 6862 35362 6914
rect 35362 6862 35364 6914
rect 35308 6860 35364 6862
rect 36988 11564 37044 11620
rect 37324 12178 37380 12180
rect 37324 12126 37326 12178
rect 37326 12126 37378 12178
rect 37378 12126 37380 12178
rect 37324 12124 37380 12126
rect 37996 12572 38052 12628
rect 37772 12012 37828 12068
rect 37436 11788 37492 11844
rect 36988 11228 37044 11284
rect 37100 10722 37156 10724
rect 37100 10670 37102 10722
rect 37102 10670 37154 10722
rect 37154 10670 37156 10722
rect 37100 10668 37156 10670
rect 36652 10444 36708 10500
rect 37548 11282 37604 11284
rect 37548 11230 37550 11282
rect 37550 11230 37602 11282
rect 37602 11230 37604 11282
rect 37548 11228 37604 11230
rect 37996 11788 38052 11844
rect 38220 11340 38276 11396
rect 38780 12236 38836 12292
rect 38332 11900 38388 11956
rect 38892 12012 38948 12068
rect 39004 13692 39060 13748
rect 39452 13020 39508 13076
rect 39340 12178 39396 12180
rect 39340 12126 39342 12178
rect 39342 12126 39394 12178
rect 39394 12126 39396 12178
rect 39340 12124 39396 12126
rect 40348 15426 40404 15428
rect 40348 15374 40350 15426
rect 40350 15374 40402 15426
rect 40402 15374 40404 15426
rect 40348 15372 40404 15374
rect 41916 16658 41972 16660
rect 41916 16606 41918 16658
rect 41918 16606 41970 16658
rect 41970 16606 41972 16658
rect 41916 16604 41972 16606
rect 40796 15484 40852 15540
rect 40908 15708 40964 15764
rect 40012 14924 40068 14980
rect 40124 14700 40180 14756
rect 40012 14530 40068 14532
rect 40012 14478 40014 14530
rect 40014 14478 40066 14530
rect 40066 14478 40068 14530
rect 40012 14476 40068 14478
rect 39676 14252 39732 14308
rect 39788 14028 39844 14084
rect 40012 13916 40068 13972
rect 39676 13580 39732 13636
rect 40572 14642 40628 14644
rect 40572 14590 40574 14642
rect 40574 14590 40626 14642
rect 40626 14590 40628 14642
rect 40572 14588 40628 14590
rect 41580 16380 41636 16436
rect 41244 15932 41300 15988
rect 41468 15986 41524 15988
rect 41468 15934 41470 15986
rect 41470 15934 41522 15986
rect 41522 15934 41524 15986
rect 41468 15932 41524 15934
rect 42028 16156 42084 16212
rect 42924 16492 42980 16548
rect 41020 15148 41076 15204
rect 42252 15874 42308 15876
rect 42252 15822 42254 15874
rect 42254 15822 42306 15874
rect 42306 15822 42308 15874
rect 42252 15820 42308 15822
rect 42140 15484 42196 15540
rect 41580 15314 41636 15316
rect 41580 15262 41582 15314
rect 41582 15262 41634 15314
rect 41634 15262 41636 15314
rect 41580 15260 41636 15262
rect 42364 15202 42420 15204
rect 42364 15150 42366 15202
rect 42366 15150 42418 15202
rect 42418 15150 42420 15202
rect 42364 15148 42420 15150
rect 41132 14476 41188 14532
rect 41468 14530 41524 14532
rect 41468 14478 41470 14530
rect 41470 14478 41522 14530
rect 41522 14478 41524 14530
rect 41468 14476 41524 14478
rect 40460 14306 40516 14308
rect 40460 14254 40462 14306
rect 40462 14254 40514 14306
rect 40514 14254 40516 14306
rect 40460 14252 40516 14254
rect 40796 14252 40852 14308
rect 40460 13692 40516 13748
rect 40684 14140 40740 14196
rect 41244 14140 41300 14196
rect 41020 14028 41076 14084
rect 40908 13356 40964 13412
rect 40012 12796 40068 12852
rect 40236 11676 40292 11732
rect 41132 13020 41188 13076
rect 40908 11564 40964 11620
rect 38444 11452 38500 11508
rect 39788 11452 39844 11508
rect 37996 10668 38052 10724
rect 38108 9996 38164 10052
rect 36876 9660 36932 9716
rect 37324 9154 37380 9156
rect 37324 9102 37326 9154
rect 37326 9102 37378 9154
rect 37378 9102 37380 9154
rect 37324 9100 37380 9102
rect 35980 8316 36036 8372
rect 35868 8092 35924 8148
rect 36540 8316 36596 8372
rect 35980 7644 36036 7700
rect 37324 8146 37380 8148
rect 37324 8094 37326 8146
rect 37326 8094 37378 8146
rect 37378 8094 37380 8146
rect 37324 8092 37380 8094
rect 35756 6748 35812 6804
rect 35196 6188 35252 6244
rect 35756 6076 35812 6132
rect 35308 5906 35364 5908
rect 35308 5854 35310 5906
rect 35310 5854 35362 5906
rect 35362 5854 35364 5906
rect 35308 5852 35364 5854
rect 37212 7698 37268 7700
rect 37212 7646 37214 7698
rect 37214 7646 37266 7698
rect 37266 7646 37268 7698
rect 37212 7644 37268 7646
rect 36428 6860 36484 6916
rect 37660 6748 37716 6804
rect 36652 6636 36708 6692
rect 35196 5514 35252 5516
rect 35196 5462 35198 5514
rect 35198 5462 35250 5514
rect 35250 5462 35252 5514
rect 35196 5460 35252 5462
rect 35300 5514 35356 5516
rect 35300 5462 35302 5514
rect 35302 5462 35354 5514
rect 35354 5462 35356 5514
rect 35300 5460 35356 5462
rect 35404 5514 35460 5516
rect 35404 5462 35406 5514
rect 35406 5462 35458 5514
rect 35458 5462 35460 5514
rect 35404 5460 35460 5462
rect 35644 5292 35700 5348
rect 35308 5010 35364 5012
rect 35308 4958 35310 5010
rect 35310 4958 35362 5010
rect 35362 4958 35364 5010
rect 35308 4956 35364 4958
rect 35196 4620 35252 4676
rect 36092 5516 36148 5572
rect 35868 5068 35924 5124
rect 36652 6412 36708 6468
rect 36764 6076 36820 6132
rect 37100 6524 37156 6580
rect 36652 5628 36708 5684
rect 36540 5292 36596 5348
rect 36092 4562 36148 4564
rect 36092 4510 36094 4562
rect 36094 4510 36146 4562
rect 36146 4510 36148 4562
rect 36092 4508 36148 4510
rect 37884 6748 37940 6804
rect 39228 11340 39284 11396
rect 39004 11282 39060 11284
rect 39004 11230 39006 11282
rect 39006 11230 39058 11282
rect 39058 11230 39060 11282
rect 39004 11228 39060 11230
rect 39676 11394 39732 11396
rect 39676 11342 39678 11394
rect 39678 11342 39730 11394
rect 39730 11342 39732 11394
rect 39676 11340 39732 11342
rect 40236 11452 40292 11508
rect 40684 11506 40740 11508
rect 40684 11454 40686 11506
rect 40686 11454 40738 11506
rect 40738 11454 40740 11506
rect 40684 11452 40740 11454
rect 41804 14588 41860 14644
rect 41692 14530 41748 14532
rect 41692 14478 41694 14530
rect 41694 14478 41746 14530
rect 41746 14478 41748 14530
rect 41692 14476 41748 14478
rect 41468 13804 41524 13860
rect 41580 13746 41636 13748
rect 41580 13694 41582 13746
rect 41582 13694 41634 13746
rect 41634 13694 41636 13746
rect 41580 13692 41636 13694
rect 41468 12908 41524 12964
rect 41692 13020 41748 13076
rect 42140 14364 42196 14420
rect 42028 14306 42084 14308
rect 42028 14254 42030 14306
rect 42030 14254 42082 14306
rect 42082 14254 42084 14306
rect 42028 14252 42084 14254
rect 42364 14140 42420 14196
rect 42252 13858 42308 13860
rect 42252 13806 42254 13858
rect 42254 13806 42306 13858
rect 42306 13806 42308 13858
rect 42252 13804 42308 13806
rect 42588 15372 42644 15428
rect 42812 16380 42868 16436
rect 43484 16828 43540 16884
rect 43036 16210 43092 16212
rect 43036 16158 43038 16210
rect 43038 16158 43090 16210
rect 43090 16158 43092 16210
rect 43036 16156 43092 16158
rect 43036 15596 43092 15652
rect 42700 14252 42756 14308
rect 43820 16882 43876 16884
rect 43820 16830 43822 16882
rect 43822 16830 43874 16882
rect 43874 16830 43876 16882
rect 43820 16828 43876 16830
rect 43148 14812 43204 14868
rect 44604 17388 44660 17444
rect 44380 17276 44436 17332
rect 44268 16994 44324 16996
rect 44268 16942 44270 16994
rect 44270 16942 44322 16994
rect 44322 16942 44324 16994
rect 44268 16940 44324 16942
rect 44156 16828 44212 16884
rect 44492 17052 44548 17108
rect 43596 14700 43652 14756
rect 43820 15314 43876 15316
rect 43820 15262 43822 15314
rect 43822 15262 43874 15314
rect 43874 15262 43876 15314
rect 43820 15260 43876 15262
rect 43484 14642 43540 14644
rect 43484 14590 43486 14642
rect 43486 14590 43538 14642
rect 43538 14590 43540 14642
rect 43484 14588 43540 14590
rect 44156 15036 44212 15092
rect 43484 14418 43540 14420
rect 43484 14366 43486 14418
rect 43486 14366 43538 14418
rect 43538 14366 43540 14418
rect 43484 14364 43540 14366
rect 42812 13804 42868 13860
rect 42476 13580 42532 13636
rect 42140 13132 42196 13188
rect 41468 12738 41524 12740
rect 41468 12686 41470 12738
rect 41470 12686 41522 12738
rect 41522 12686 41524 12738
rect 41468 12684 41524 12686
rect 38892 9884 38948 9940
rect 38780 9266 38836 9268
rect 38780 9214 38782 9266
rect 38782 9214 38834 9266
rect 38834 9214 38836 9266
rect 38780 9212 38836 9214
rect 39900 10108 39956 10164
rect 39004 8876 39060 8932
rect 38444 8540 38500 8596
rect 38108 7980 38164 8036
rect 38108 7644 38164 7700
rect 38220 8092 38276 8148
rect 38780 7532 38836 7588
rect 37996 6636 38052 6692
rect 39004 7084 39060 7140
rect 37772 6524 37828 6580
rect 37324 6076 37380 6132
rect 37996 6466 38052 6468
rect 37996 6414 37998 6466
rect 37998 6414 38050 6466
rect 38050 6414 38052 6466
rect 37996 6412 38052 6414
rect 38556 6636 38612 6692
rect 40684 9884 40740 9940
rect 39900 8876 39956 8932
rect 39452 7980 39508 8036
rect 39340 6802 39396 6804
rect 39340 6750 39342 6802
rect 39342 6750 39394 6802
rect 39394 6750 39396 6802
rect 39340 6748 39396 6750
rect 39564 8764 39620 8820
rect 40348 8930 40404 8932
rect 40348 8878 40350 8930
rect 40350 8878 40402 8930
rect 40402 8878 40404 8930
rect 40348 8876 40404 8878
rect 40012 8652 40068 8708
rect 40460 8316 40516 8372
rect 39900 7586 39956 7588
rect 39900 7534 39902 7586
rect 39902 7534 39954 7586
rect 39954 7534 39956 7586
rect 39900 7532 39956 7534
rect 39900 6860 39956 6916
rect 39564 6748 39620 6804
rect 39452 6524 39508 6580
rect 38892 5964 38948 6020
rect 38556 5740 38612 5796
rect 38668 5628 38724 5684
rect 37436 5292 37492 5348
rect 37660 5346 37716 5348
rect 37660 5294 37662 5346
rect 37662 5294 37714 5346
rect 37714 5294 37716 5346
rect 37660 5292 37716 5294
rect 39340 5852 39396 5908
rect 35980 4450 36036 4452
rect 35980 4398 35982 4450
rect 35982 4398 36034 4450
rect 36034 4398 36036 4450
rect 35980 4396 36036 4398
rect 35196 3946 35252 3948
rect 35196 3894 35198 3946
rect 35198 3894 35250 3946
rect 35250 3894 35252 3946
rect 35196 3892 35252 3894
rect 35300 3946 35356 3948
rect 35300 3894 35302 3946
rect 35302 3894 35354 3946
rect 35354 3894 35356 3946
rect 35300 3892 35356 3894
rect 35404 3946 35460 3948
rect 35404 3894 35406 3946
rect 35406 3894 35458 3946
rect 35458 3894 35460 3946
rect 35404 3892 35460 3894
rect 35084 3500 35140 3556
rect 36204 3554 36260 3556
rect 36204 3502 36206 3554
rect 36206 3502 36258 3554
rect 36258 3502 36260 3554
rect 36204 3500 36260 3502
rect 38108 5122 38164 5124
rect 38108 5070 38110 5122
rect 38110 5070 38162 5122
rect 38162 5070 38164 5122
rect 38108 5068 38164 5070
rect 38780 5010 38836 5012
rect 38780 4958 38782 5010
rect 38782 4958 38834 5010
rect 38834 4958 38836 5010
rect 38780 4956 38836 4958
rect 38332 4172 38388 4228
rect 37660 3612 37716 3668
rect 39788 6300 39844 6356
rect 39788 6076 39844 6132
rect 39900 5906 39956 5908
rect 39900 5854 39902 5906
rect 39902 5854 39954 5906
rect 39954 5854 39956 5906
rect 39900 5852 39956 5854
rect 39900 5292 39956 5348
rect 38892 3276 38948 3332
rect 39004 3388 39060 3444
rect 40236 7420 40292 7476
rect 40348 7362 40404 7364
rect 40348 7310 40350 7362
rect 40350 7310 40402 7362
rect 40402 7310 40404 7362
rect 40348 7308 40404 7310
rect 40236 6972 40292 7028
rect 40124 6578 40180 6580
rect 40124 6526 40126 6578
rect 40126 6526 40178 6578
rect 40178 6526 40180 6578
rect 40124 6524 40180 6526
rect 40236 6466 40292 6468
rect 40236 6414 40238 6466
rect 40238 6414 40290 6466
rect 40290 6414 40292 6466
rect 40236 6412 40292 6414
rect 40124 5906 40180 5908
rect 40124 5854 40126 5906
rect 40126 5854 40178 5906
rect 40178 5854 40180 5906
rect 40124 5852 40180 5854
rect 40124 5628 40180 5684
rect 41356 12236 41412 12292
rect 41356 11788 41412 11844
rect 41468 11564 41524 11620
rect 41916 12290 41972 12292
rect 41916 12238 41918 12290
rect 41918 12238 41970 12290
rect 41970 12238 41972 12290
rect 41916 12236 41972 12238
rect 41580 11900 41636 11956
rect 41468 11228 41524 11284
rect 43372 13580 43428 13636
rect 42700 13356 42756 13412
rect 43148 13468 43204 13524
rect 42700 13186 42756 13188
rect 42700 13134 42702 13186
rect 42702 13134 42754 13186
rect 42754 13134 42756 13186
rect 42700 13132 42756 13134
rect 42252 12684 42308 12740
rect 42812 12178 42868 12180
rect 42812 12126 42814 12178
rect 42814 12126 42866 12178
rect 42866 12126 42868 12178
rect 42812 12124 42868 12126
rect 44268 14530 44324 14532
rect 44268 14478 44270 14530
rect 44270 14478 44322 14530
rect 44322 14478 44324 14530
rect 44268 14476 44324 14478
rect 44156 14140 44212 14196
rect 43820 13356 43876 13412
rect 43260 12290 43316 12292
rect 43260 12238 43262 12290
rect 43262 12238 43314 12290
rect 43314 12238 43316 12290
rect 43260 12236 43316 12238
rect 44380 13468 44436 13524
rect 43932 12124 43988 12180
rect 45052 18844 45108 18900
rect 45612 20076 45668 20132
rect 44940 18060 44996 18116
rect 45612 18844 45668 18900
rect 44940 17836 44996 17892
rect 45276 18338 45332 18340
rect 45276 18286 45278 18338
rect 45278 18286 45330 18338
rect 45330 18286 45332 18338
rect 45276 18284 45332 18286
rect 45836 18562 45892 18564
rect 45836 18510 45838 18562
rect 45838 18510 45890 18562
rect 45890 18510 45892 18562
rect 45836 18508 45892 18510
rect 46060 18450 46116 18452
rect 46060 18398 46062 18450
rect 46062 18398 46114 18450
rect 46114 18398 46116 18450
rect 46060 18396 46116 18398
rect 47180 18674 47236 18676
rect 47180 18622 47182 18674
rect 47182 18622 47234 18674
rect 47234 18622 47236 18674
rect 47180 18620 47236 18622
rect 46620 18396 46676 18452
rect 45052 17388 45108 17444
rect 44828 17164 44884 17220
rect 44716 16156 44772 16212
rect 44604 14700 44660 14756
rect 42700 11564 42756 11620
rect 43596 11394 43652 11396
rect 43596 11342 43598 11394
rect 43598 11342 43650 11394
rect 43650 11342 43652 11394
rect 43596 11340 43652 11342
rect 42812 11282 42868 11284
rect 42812 11230 42814 11282
rect 42814 11230 42866 11282
rect 42866 11230 42868 11282
rect 42812 11228 42868 11230
rect 43372 10722 43428 10724
rect 43372 10670 43374 10722
rect 43374 10670 43426 10722
rect 43426 10670 43428 10722
rect 43372 10668 43428 10670
rect 43484 10610 43540 10612
rect 43484 10558 43486 10610
rect 43486 10558 43538 10610
rect 43538 10558 43540 10610
rect 43484 10556 43540 10558
rect 42252 10108 42308 10164
rect 42700 10220 42756 10276
rect 41916 9884 41972 9940
rect 41132 9212 41188 9268
rect 41916 9266 41972 9268
rect 41916 9214 41918 9266
rect 41918 9214 41970 9266
rect 41970 9214 41972 9266
rect 41916 9212 41972 9214
rect 41468 9042 41524 9044
rect 41468 8990 41470 9042
rect 41470 8990 41522 9042
rect 41522 8990 41524 9042
rect 41468 8988 41524 8990
rect 41356 8876 41412 8932
rect 41692 8764 41748 8820
rect 40572 6524 40628 6580
rect 41020 7250 41076 7252
rect 41020 7198 41022 7250
rect 41022 7198 41074 7250
rect 41074 7198 41076 7250
rect 41020 7196 41076 7198
rect 41244 7084 41300 7140
rect 41132 6860 41188 6916
rect 41020 5628 41076 5684
rect 40460 5180 40516 5236
rect 40348 5068 40404 5124
rect 40236 4562 40292 4564
rect 40236 4510 40238 4562
rect 40238 4510 40290 4562
rect 40290 4510 40292 4562
rect 40236 4508 40292 4510
rect 40796 3666 40852 3668
rect 40796 3614 40798 3666
rect 40798 3614 40850 3666
rect 40850 3614 40852 3666
rect 40796 3612 40852 3614
rect 41468 6748 41524 6804
rect 41356 6300 41412 6356
rect 41580 5068 41636 5124
rect 41244 3500 41300 3556
rect 41692 4844 41748 4900
rect 42476 8428 42532 8484
rect 41916 8146 41972 8148
rect 41916 8094 41918 8146
rect 41918 8094 41970 8146
rect 41970 8094 41972 8146
rect 41916 8092 41972 8094
rect 41916 7868 41972 7924
rect 42140 7868 42196 7924
rect 42364 7644 42420 7700
rect 43932 10780 43988 10836
rect 43484 9996 43540 10052
rect 42812 8930 42868 8932
rect 42812 8878 42814 8930
rect 42814 8878 42866 8930
rect 42866 8878 42868 8930
rect 42812 8876 42868 8878
rect 42812 7644 42868 7700
rect 42700 7532 42756 7588
rect 42476 6300 42532 6356
rect 42700 7308 42756 7364
rect 41804 4284 41860 4340
rect 41916 5740 41972 5796
rect 42028 5292 42084 5348
rect 42252 5852 42308 5908
rect 42924 7308 42980 7364
rect 42812 5740 42868 5796
rect 42140 4508 42196 4564
rect 42700 4956 42756 5012
rect 42028 4226 42084 4228
rect 42028 4174 42030 4226
rect 42030 4174 42082 4226
rect 42082 4174 42084 4226
rect 42028 4172 42084 4174
rect 42364 3612 42420 3668
rect 42924 5068 42980 5124
rect 43036 4396 43092 4452
rect 43148 8652 43204 8708
rect 44268 10722 44324 10724
rect 44268 10670 44270 10722
rect 44270 10670 44322 10722
rect 44322 10670 44324 10722
rect 44268 10668 44324 10670
rect 45500 16940 45556 16996
rect 46396 18338 46452 18340
rect 46396 18286 46398 18338
rect 46398 18286 46450 18338
rect 46450 18286 46452 18338
rect 46396 18284 46452 18286
rect 46060 17724 46116 17780
rect 44940 15708 44996 15764
rect 44940 14812 44996 14868
rect 44828 13356 44884 13412
rect 45164 13244 45220 13300
rect 44828 12962 44884 12964
rect 44828 12910 44830 12962
rect 44830 12910 44882 12962
rect 44882 12910 44884 12962
rect 44828 12908 44884 12910
rect 44940 12850 44996 12852
rect 44940 12798 44942 12850
rect 44942 12798 44994 12850
rect 44994 12798 44996 12850
rect 44940 12796 44996 12798
rect 44828 11394 44884 11396
rect 44828 11342 44830 11394
rect 44830 11342 44882 11394
rect 44882 11342 44884 11394
rect 44828 11340 44884 11342
rect 45612 16156 45668 16212
rect 46284 16940 46340 16996
rect 47964 20076 48020 20132
rect 48076 18956 48132 19012
rect 47852 18396 47908 18452
rect 47516 18172 47572 18228
rect 47628 18060 47684 18116
rect 46956 16994 47012 16996
rect 46956 16942 46958 16994
rect 46958 16942 47010 16994
rect 47010 16942 47012 16994
rect 46956 16940 47012 16942
rect 46172 16882 46228 16884
rect 46172 16830 46174 16882
rect 46174 16830 46226 16882
rect 46226 16830 46228 16882
rect 46172 16828 46228 16830
rect 46060 16716 46116 16772
rect 45948 15314 46004 15316
rect 45948 15262 45950 15314
rect 45950 15262 46002 15314
rect 46002 15262 46004 15314
rect 45948 15260 46004 15262
rect 46844 16770 46900 16772
rect 46844 16718 46846 16770
rect 46846 16718 46898 16770
rect 46898 16718 46900 16770
rect 46844 16716 46900 16718
rect 46396 16210 46452 16212
rect 46396 16158 46398 16210
rect 46398 16158 46450 16210
rect 46450 16158 46452 16210
rect 46396 16156 46452 16158
rect 47292 16882 47348 16884
rect 47292 16830 47294 16882
rect 47294 16830 47346 16882
rect 47346 16830 47348 16882
rect 47292 16828 47348 16830
rect 48188 17778 48244 17780
rect 48188 17726 48190 17778
rect 48190 17726 48242 17778
rect 48242 17726 48244 17778
rect 48188 17724 48244 17726
rect 48300 17276 48356 17332
rect 48076 16994 48132 16996
rect 48076 16942 48078 16994
rect 48078 16942 48130 16994
rect 48130 16942 48132 16994
rect 48076 16940 48132 16942
rect 47516 16156 47572 16212
rect 46732 15372 46788 15428
rect 47292 15260 47348 15316
rect 47404 15036 47460 15092
rect 47068 14588 47124 14644
rect 45836 14476 45892 14532
rect 46732 13746 46788 13748
rect 46732 13694 46734 13746
rect 46734 13694 46786 13746
rect 46786 13694 46788 13746
rect 46732 13692 46788 13694
rect 47404 13692 47460 13748
rect 45388 13244 45444 13300
rect 46060 12850 46116 12852
rect 46060 12798 46062 12850
rect 46062 12798 46114 12850
rect 46114 12798 46116 12850
rect 46060 12796 46116 12798
rect 47964 13468 48020 13524
rect 46508 12124 46564 12180
rect 45276 11340 45332 11396
rect 44716 10780 44772 10836
rect 44828 10610 44884 10612
rect 44828 10558 44830 10610
rect 44830 10558 44882 10610
rect 44882 10558 44884 10610
rect 44828 10556 44884 10558
rect 44156 9212 44212 9268
rect 43260 8316 43316 8372
rect 43484 7308 43540 7364
rect 43708 8818 43764 8820
rect 43708 8766 43710 8818
rect 43710 8766 43762 8818
rect 43762 8766 43764 8818
rect 43708 8764 43764 8766
rect 44156 8540 44212 8596
rect 44156 8370 44212 8372
rect 44156 8318 44158 8370
rect 44158 8318 44210 8370
rect 44210 8318 44212 8370
rect 44156 8316 44212 8318
rect 43708 7868 43764 7924
rect 43820 6860 43876 6916
rect 44156 8092 44212 8148
rect 43932 7980 43988 8036
rect 43820 6412 43876 6468
rect 43260 5180 43316 5236
rect 43708 4508 43764 4564
rect 44268 8034 44324 8036
rect 44268 7982 44270 8034
rect 44270 7982 44322 8034
rect 44322 7982 44324 8034
rect 44268 7980 44324 7982
rect 45052 9602 45108 9604
rect 45052 9550 45054 9602
rect 45054 9550 45106 9602
rect 45106 9550 45108 9602
rect 45052 9548 45108 9550
rect 44940 9212 44996 9268
rect 44716 9100 44772 9156
rect 45388 8988 45444 9044
rect 44940 8428 44996 8484
rect 45164 8540 45220 8596
rect 45388 8316 45444 8372
rect 44044 5740 44100 5796
rect 44156 6860 44212 6916
rect 43932 5068 43988 5124
rect 43932 4562 43988 4564
rect 43932 4510 43934 4562
rect 43934 4510 43986 4562
rect 43986 4510 43988 4562
rect 43932 4508 43988 4510
rect 44492 6524 44548 6580
rect 44268 5180 44324 5236
rect 44268 4956 44324 5012
rect 43148 3724 43204 3780
rect 43932 4284 43988 4340
rect 43708 3554 43764 3556
rect 43708 3502 43710 3554
rect 43710 3502 43762 3554
rect 43762 3502 43764 3554
rect 43708 3500 43764 3502
rect 45052 7196 45108 7252
rect 44828 6300 44884 6356
rect 44604 4732 44660 4788
rect 44716 6188 44772 6244
rect 44828 5682 44884 5684
rect 44828 5630 44830 5682
rect 44830 5630 44882 5682
rect 44882 5630 44884 5682
rect 44828 5628 44884 5630
rect 44716 5292 44772 5348
rect 44828 5404 44884 5460
rect 44604 3388 44660 3444
rect 44940 5068 44996 5124
rect 45836 10834 45892 10836
rect 45836 10782 45838 10834
rect 45838 10782 45890 10834
rect 45890 10782 45892 10834
rect 45836 10780 45892 10782
rect 46284 12066 46340 12068
rect 46284 12014 46286 12066
rect 46286 12014 46338 12066
rect 46338 12014 46340 12066
rect 46284 12012 46340 12014
rect 46844 11452 46900 11508
rect 47740 11506 47796 11508
rect 47740 11454 47742 11506
rect 47742 11454 47794 11506
rect 47794 11454 47796 11506
rect 47740 11452 47796 11454
rect 46172 10220 46228 10276
rect 47180 10220 47236 10276
rect 45948 10108 46004 10164
rect 45836 9042 45892 9044
rect 45836 8990 45838 9042
rect 45838 8990 45890 9042
rect 45890 8990 45892 9042
rect 45836 8988 45892 8990
rect 46844 10108 46900 10164
rect 46620 8204 46676 8260
rect 46396 7420 46452 7476
rect 45276 6524 45332 6580
rect 45164 4450 45220 4452
rect 45164 4398 45166 4450
rect 45166 4398 45218 4450
rect 45218 4398 45220 4450
rect 45164 4396 45220 4398
rect 46396 4956 46452 5012
rect 46508 5068 46564 5124
rect 45836 4898 45892 4900
rect 45836 4846 45838 4898
rect 45838 4846 45890 4898
rect 45890 4846 45892 4898
rect 45836 4844 45892 4846
rect 45276 3500 45332 3556
rect 46732 5740 46788 5796
rect 46620 4508 46676 4564
rect 46956 9548 47012 9604
rect 47180 9602 47236 9604
rect 47180 9550 47182 9602
rect 47182 9550 47234 9602
rect 47234 9550 47236 9602
rect 47180 9548 47236 9550
rect 47068 8876 47124 8932
rect 48188 10108 48244 10164
rect 47964 8988 48020 9044
rect 47964 8818 48020 8820
rect 47964 8766 47966 8818
rect 47966 8766 48018 8818
rect 48018 8766 48020 8818
rect 47964 8764 48020 8766
rect 47404 8540 47460 8596
rect 47964 8092 48020 8148
rect 48188 7980 48244 8036
rect 47964 7420 48020 7476
rect 47292 6018 47348 6020
rect 47292 5966 47294 6018
rect 47294 5966 47346 6018
rect 47346 5966 47348 6018
rect 47292 5964 47348 5966
rect 47068 5516 47124 5572
rect 47852 5404 47908 5460
rect 47964 5292 48020 5348
rect 47740 5180 47796 5236
rect 47404 4956 47460 5012
rect 46956 4060 47012 4116
rect 46732 3612 46788 3668
rect 47628 4562 47684 4564
rect 47628 4510 47630 4562
rect 47630 4510 47682 4562
rect 47682 4510 47684 4562
rect 47628 4508 47684 4510
rect 47852 4338 47908 4340
rect 47852 4286 47854 4338
rect 47854 4286 47906 4338
rect 47906 4286 47908 4338
rect 47852 4284 47908 4286
rect 47628 3724 47684 3780
rect 48076 3442 48132 3444
rect 48076 3390 48078 3442
rect 48078 3390 48130 3442
rect 48130 3390 48132 3442
rect 48076 3388 48132 3390
<< metal3 >>
rect 32946 46956 32956 47012
rect 33012 46956 36988 47012
rect 37044 46956 37054 47012
rect 49200 46452 50000 46480
rect 45266 46396 45276 46452
rect 45332 46396 50000 46452
rect 49200 46368 50000 46396
rect 4466 46228 4476 46284
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4740 46228 4750 46284
rect 35186 46228 35196 46284
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35460 46228 35470 46284
rect 26226 46060 26236 46116
rect 26292 46060 29372 46116
rect 29428 46060 29438 46116
rect 30258 46060 30268 46116
rect 30324 46060 33180 46116
rect 33236 46060 33246 46116
rect 10658 45948 10668 46004
rect 10724 45948 13916 46004
rect 13972 45948 13982 46004
rect 15250 45836 15260 45892
rect 15316 45836 16268 45892
rect 16324 45836 16334 45892
rect 37314 45836 37324 45892
rect 37380 45836 39788 45892
rect 39844 45836 39854 45892
rect 49200 45780 50000 45808
rect 24546 45724 24556 45780
rect 24612 45724 25340 45780
rect 25396 45724 25406 45780
rect 45042 45724 45052 45780
rect 45108 45724 50000 45780
rect 49200 45696 50000 45724
rect 7410 45612 7420 45668
rect 7476 45612 8092 45668
rect 8148 45612 11564 45668
rect 11620 45612 11630 45668
rect 18162 45612 18172 45668
rect 18228 45612 20076 45668
rect 20132 45612 20142 45668
rect 37874 45612 37884 45668
rect 37940 45612 38892 45668
rect 38948 45612 38958 45668
rect 19826 45444 19836 45500
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 20100 45444 20110 45500
rect 1698 45388 1708 45444
rect 1764 45388 1774 45444
rect 11106 45388 11116 45444
rect 11172 45388 12236 45444
rect 12292 45388 12302 45444
rect 17602 45388 17612 45444
rect 17668 45388 19292 45444
rect 19348 45388 19358 45444
rect 0 45108 800 45136
rect 1708 45108 1764 45388
rect 22978 45276 22988 45332
rect 23044 45276 25564 45332
rect 25620 45276 25630 45332
rect 35186 45276 35196 45332
rect 35252 45276 40796 45332
rect 40852 45276 40862 45332
rect 44370 45276 44380 45332
rect 44436 45276 46060 45332
rect 46116 45276 46126 45332
rect 23090 45164 23100 45220
rect 23156 45164 23884 45220
rect 23940 45164 25676 45220
rect 25732 45164 25742 45220
rect 37650 45164 37660 45220
rect 37716 45164 42028 45220
rect 42084 45164 42094 45220
rect 49200 45108 50000 45136
rect 0 45052 1764 45108
rect 10098 45052 10108 45108
rect 10164 45052 13692 45108
rect 13748 45052 17164 45108
rect 17220 45052 17230 45108
rect 22866 45052 22876 45108
rect 22932 45052 24444 45108
rect 24500 45052 25340 45108
rect 25396 45052 25406 45108
rect 27346 45052 27356 45108
rect 27412 45052 30380 45108
rect 30436 45052 30446 45108
rect 33954 45052 33964 45108
rect 34020 45052 36316 45108
rect 36372 45052 37100 45108
rect 37156 45052 37772 45108
rect 37828 45052 37838 45108
rect 38322 45052 38332 45108
rect 38388 45052 44604 45108
rect 44660 45052 44670 45108
rect 46834 45052 46844 45108
rect 46900 45052 50000 45108
rect 0 45024 800 45052
rect 49200 45024 50000 45052
rect 6178 44940 6188 44996
rect 6244 44940 7980 44996
rect 8036 44940 8046 44996
rect 8418 44940 8428 44996
rect 8484 44940 9660 44996
rect 9716 44940 11788 44996
rect 11844 44940 11854 44996
rect 19282 44940 19292 44996
rect 19348 44940 20412 44996
rect 20468 44940 20478 44996
rect 22642 44940 22652 44996
rect 22708 44940 23660 44996
rect 23716 44940 23726 44996
rect 44706 44940 44716 44996
rect 44772 44940 45052 44996
rect 45108 44940 45118 44996
rect 7980 44884 8036 44940
rect 7980 44828 8764 44884
rect 8820 44828 9548 44884
rect 9604 44828 10108 44884
rect 10164 44828 10174 44884
rect 35410 44828 35420 44884
rect 35476 44828 39004 44884
rect 39060 44828 39070 44884
rect 26562 44716 26572 44772
rect 26628 44716 28588 44772
rect 28644 44716 28654 44772
rect 4466 44660 4476 44716
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4740 44660 4750 44716
rect 35186 44660 35196 44716
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35460 44660 35470 44716
rect 18694 44492 18732 44548
rect 18788 44492 18798 44548
rect 26898 44492 26908 44548
rect 26964 44492 27692 44548
rect 27748 44492 27758 44548
rect 31714 44492 31724 44548
rect 31780 44492 34524 44548
rect 34580 44492 34590 44548
rect 39218 44492 39228 44548
rect 39284 44492 44940 44548
rect 44996 44492 45006 44548
rect 0 44436 800 44464
rect 49200 44436 50000 44464
rect 0 44380 21980 44436
rect 22036 44380 22046 44436
rect 31602 44380 31612 44436
rect 31668 44380 33068 44436
rect 33124 44380 33134 44436
rect 33282 44380 33292 44436
rect 33348 44380 37100 44436
rect 37156 44380 37166 44436
rect 40674 44380 40684 44436
rect 40740 44380 43260 44436
rect 43316 44380 45836 44436
rect 45892 44380 45902 44436
rect 47730 44380 47740 44436
rect 47796 44380 50000 44436
rect 0 44352 800 44380
rect 33292 44324 33348 44380
rect 49200 44352 50000 44380
rect 21858 44268 21868 44324
rect 21924 44268 28700 44324
rect 28756 44268 28766 44324
rect 29922 44268 29932 44324
rect 29988 44268 30380 44324
rect 30436 44268 33348 44324
rect 8418 44156 8428 44212
rect 8484 44156 12908 44212
rect 12964 44156 12974 44212
rect 33170 44156 33180 44212
rect 33236 44156 35980 44212
rect 36036 44156 36046 44212
rect 1474 44044 1484 44100
rect 1540 44044 7196 44100
rect 7252 44044 7262 44100
rect 8306 44044 8316 44100
rect 8372 44044 8988 44100
rect 9044 44044 9054 44100
rect 14588 44044 17052 44100
rect 17108 44044 17118 44100
rect 28354 44044 28364 44100
rect 28420 44044 29372 44100
rect 29428 44044 30268 44100
rect 30324 44044 30334 44100
rect 14588 43876 14644 44044
rect 40002 43932 40012 43988
rect 40068 43932 42028 43988
rect 42084 43932 45276 43988
rect 45332 43932 45342 43988
rect 19826 43876 19836 43932
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 20100 43876 20110 43932
rect 13682 43820 13692 43876
rect 13748 43820 14140 43876
rect 14196 43820 14644 43876
rect 19058 43820 19068 43876
rect 19124 43820 19572 43876
rect 38658 43820 38668 43876
rect 38724 43820 44716 43876
rect 44772 43820 44782 43876
rect 19516 43764 19572 43820
rect 49200 43764 50000 43792
rect 10994 43708 11004 43764
rect 11060 43708 11676 43764
rect 11732 43708 11742 43764
rect 11890 43708 11900 43764
rect 11956 43708 12572 43764
rect 12628 43708 12638 43764
rect 12898 43708 12908 43764
rect 12964 43708 14700 43764
rect 14756 43708 15988 43764
rect 18610 43708 18620 43764
rect 18676 43708 19292 43764
rect 19348 43708 19358 43764
rect 19516 43708 20412 43764
rect 20468 43708 20478 43764
rect 26114 43708 26124 43764
rect 26180 43708 26572 43764
rect 26628 43708 26638 43764
rect 29138 43708 29148 43764
rect 29204 43708 29820 43764
rect 29876 43708 29886 43764
rect 31938 43708 31948 43764
rect 32004 43708 34412 43764
rect 34468 43708 39564 43764
rect 39620 43708 39630 43764
rect 48290 43708 48300 43764
rect 48356 43708 50000 43764
rect 15932 43652 15988 43708
rect 49200 43680 50000 43708
rect 3938 43596 3948 43652
rect 4004 43596 4844 43652
rect 4900 43596 5628 43652
rect 5684 43596 6076 43652
rect 6132 43596 6142 43652
rect 9538 43596 9548 43652
rect 9604 43596 11452 43652
rect 11508 43596 11518 43652
rect 12338 43596 12348 43652
rect 12404 43596 12796 43652
rect 12852 43596 12862 43652
rect 14466 43596 14476 43652
rect 14532 43596 15596 43652
rect 15652 43596 15662 43652
rect 15932 43596 19012 43652
rect 30930 43596 30940 43652
rect 30996 43596 32172 43652
rect 32228 43596 32238 43652
rect 33954 43596 33964 43652
rect 34020 43596 36988 43652
rect 37044 43596 37054 43652
rect 38546 43596 38556 43652
rect 38612 43596 40908 43652
rect 40964 43596 40974 43652
rect 18956 43540 19012 43596
rect 10546 43484 10556 43540
rect 10612 43484 11564 43540
rect 11620 43484 11630 43540
rect 12674 43484 12684 43540
rect 12740 43484 13916 43540
rect 13972 43484 13982 43540
rect 14476 43484 15708 43540
rect 15764 43484 15774 43540
rect 18946 43484 18956 43540
rect 19012 43484 22428 43540
rect 22484 43484 22494 43540
rect 36754 43484 36764 43540
rect 36820 43484 39340 43540
rect 39396 43484 39406 43540
rect 41234 43484 41244 43540
rect 41300 43484 42924 43540
rect 42980 43484 42990 43540
rect 4834 43372 4844 43428
rect 4900 43372 5740 43428
rect 5796 43372 5806 43428
rect 13122 43372 13132 43428
rect 13188 43372 13692 43428
rect 13748 43372 13758 43428
rect 13794 43260 13804 43316
rect 13860 43260 14252 43316
rect 14308 43260 14318 43316
rect 14476 43204 14532 43484
rect 10882 43148 10892 43204
rect 10948 43148 14532 43204
rect 14700 43372 21084 43428
rect 21140 43372 22092 43428
rect 22148 43372 24892 43428
rect 24948 43372 24958 43428
rect 32274 43372 32284 43428
rect 32340 43372 34076 43428
rect 34132 43372 34142 43428
rect 4466 43092 4476 43148
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4740 43092 4750 43148
rect 11666 43036 11676 43092
rect 11732 43036 14028 43092
rect 14084 43036 14094 43092
rect 14700 42980 14756 43372
rect 6626 42924 6636 42980
rect 6692 42924 14756 42980
rect 15092 43260 16268 43316
rect 16324 43260 16334 43316
rect 15092 42868 15148 43260
rect 35186 43092 35196 43148
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35460 43092 35470 43148
rect 49200 43092 50000 43120
rect 48178 43036 48188 43092
rect 48244 43036 50000 43092
rect 49200 43008 50000 43036
rect 32498 42924 32508 42980
rect 32564 42924 34524 42980
rect 34580 42924 34590 42980
rect 36418 42924 36428 42980
rect 36484 42924 37212 42980
rect 37268 42924 37278 42980
rect 10098 42812 10108 42868
rect 10164 42812 10892 42868
rect 10948 42812 10958 42868
rect 14018 42812 14028 42868
rect 14084 42812 15148 42868
rect 10546 42700 10556 42756
rect 10612 42700 11340 42756
rect 11396 42700 12460 42756
rect 12516 42700 12526 42756
rect 19170 42700 19180 42756
rect 19236 42700 19740 42756
rect 19796 42700 23212 42756
rect 23268 42700 23278 42756
rect 28466 42700 28476 42756
rect 28532 42700 30268 42756
rect 30324 42700 31836 42756
rect 31892 42700 35084 42756
rect 35140 42700 35150 42756
rect 47394 42700 47404 42756
rect 47460 42700 48188 42756
rect 48244 42700 48254 42756
rect 6374 42588 6412 42644
rect 6468 42588 6478 42644
rect 9202 42588 9212 42644
rect 9268 42588 11452 42644
rect 11508 42588 15260 42644
rect 15316 42588 15326 42644
rect 17938 42588 17948 42644
rect 18004 42588 18620 42644
rect 18676 42588 19516 42644
rect 19572 42588 20636 42644
rect 20692 42588 20702 42644
rect 27346 42588 27356 42644
rect 27412 42588 29260 42644
rect 29316 42588 29326 42644
rect 42914 42588 42924 42644
rect 42980 42588 43820 42644
rect 43876 42588 43886 42644
rect 2146 42476 2156 42532
rect 2212 42476 3948 42532
rect 4004 42476 4014 42532
rect 8642 42476 8652 42532
rect 8708 42476 10220 42532
rect 10276 42476 10286 42532
rect 14018 42476 14028 42532
rect 14084 42476 14364 42532
rect 14420 42476 14430 42532
rect 14690 42476 14700 42532
rect 14756 42476 15036 42532
rect 15092 42476 15102 42532
rect 19058 42476 19068 42532
rect 19124 42476 19964 42532
rect 20020 42476 20030 42532
rect 25890 42476 25900 42532
rect 25956 42476 26572 42532
rect 26628 42476 26638 42532
rect 31602 42476 31612 42532
rect 31668 42476 34188 42532
rect 34244 42476 34254 42532
rect 49200 42420 50000 42448
rect 13794 42364 13804 42420
rect 13860 42364 19180 42420
rect 19236 42364 19246 42420
rect 48178 42364 48188 42420
rect 48244 42364 50000 42420
rect 19826 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20110 42364
rect 49200 42336 50000 42364
rect 6290 42252 6300 42308
rect 6356 42252 6636 42308
rect 6692 42252 6702 42308
rect 14690 42252 14700 42308
rect 14756 42252 15316 42308
rect 15260 42196 15316 42252
rect 7942 42140 7980 42196
rect 8036 42140 8046 42196
rect 8652 42140 9996 42196
rect 10052 42140 15148 42196
rect 15260 42140 15596 42196
rect 15652 42140 15662 42196
rect 16594 42140 16604 42196
rect 16660 42140 18340 42196
rect 20402 42140 20412 42196
rect 20468 42140 20916 42196
rect 45042 42140 45052 42196
rect 45108 42140 46844 42196
rect 46900 42140 46910 42196
rect 2258 42028 2268 42084
rect 2324 42028 2334 42084
rect 4246 42028 4284 42084
rect 4340 42028 4350 42084
rect 2268 41972 2324 42028
rect 8652 41972 8708 42140
rect 15092 42084 15148 42140
rect 18284 42084 18340 42140
rect 8866 42028 8876 42084
rect 8932 42028 10108 42084
rect 10164 42028 10174 42084
rect 11106 42028 11116 42084
rect 11172 42028 12348 42084
rect 12404 42028 12414 42084
rect 15092 42028 17500 42084
rect 17556 42028 17566 42084
rect 18274 42028 18284 42084
rect 18340 42028 19852 42084
rect 19908 42028 19918 42084
rect 1698 41916 1708 41972
rect 1764 41916 2324 41972
rect 3826 41916 3836 41972
rect 3892 41916 5404 41972
rect 5460 41916 5470 41972
rect 7410 41916 7420 41972
rect 7476 41916 8708 41972
rect 9426 41916 9436 41972
rect 9492 41916 9884 41972
rect 9940 41916 10668 41972
rect 10724 41916 10734 41972
rect 14018 41916 14028 41972
rect 14084 41916 17388 41972
rect 17444 41916 17454 41972
rect 18498 41916 18508 41972
rect 18564 41916 19964 41972
rect 20020 41916 20030 41972
rect 4946 41804 4956 41860
rect 5012 41804 6748 41860
rect 6804 41804 6814 41860
rect 9090 41804 9100 41860
rect 9156 41804 10108 41860
rect 10164 41804 12908 41860
rect 12964 41804 12974 41860
rect 13570 41804 13580 41860
rect 13636 41804 16156 41860
rect 16212 41804 16222 41860
rect 16482 41804 16492 41860
rect 16548 41804 18060 41860
rect 18116 41804 18126 41860
rect 20860 41748 20916 42140
rect 21970 41916 21980 41972
rect 22036 41916 25116 41972
rect 25172 41916 25182 41972
rect 32274 41916 32284 41972
rect 32340 41916 35868 41972
rect 35924 41916 35934 41972
rect 37538 41916 37548 41972
rect 37604 41916 39228 41972
rect 39284 41916 39294 41972
rect 39666 41916 39676 41972
rect 39732 41916 43596 41972
rect 43652 41916 43662 41972
rect 21634 41804 21644 41860
rect 21700 41804 23100 41860
rect 23156 41804 23166 41860
rect 24546 41804 24556 41860
rect 24612 41804 25340 41860
rect 25396 41804 25406 41860
rect 34626 41804 34636 41860
rect 34692 41804 35980 41860
rect 36036 41804 39900 41860
rect 39956 41804 39966 41860
rect 40114 41804 40124 41860
rect 40180 41804 41020 41860
rect 41076 41804 43932 41860
rect 43988 41804 44492 41860
rect 44548 41804 44558 41860
rect 45826 41804 45836 41860
rect 45892 41804 47740 41860
rect 47796 41804 47806 41860
rect 49200 41748 50000 41776
rect 12562 41692 12572 41748
rect 12628 41692 13356 41748
rect 13412 41692 13422 41748
rect 15092 41692 15260 41748
rect 15316 41692 15326 41748
rect 20850 41692 20860 41748
rect 20916 41692 20926 41748
rect 23538 41692 23548 41748
rect 23604 41692 23884 41748
rect 23940 41692 23950 41748
rect 24882 41692 24892 41748
rect 24948 41692 26348 41748
rect 26404 41692 26414 41748
rect 39218 41692 39228 41748
rect 39284 41692 44268 41748
rect 44324 41692 44334 41748
rect 47954 41692 47964 41748
rect 48020 41692 50000 41748
rect 15092 41636 15148 41692
rect 49200 41664 50000 41692
rect 12674 41580 12684 41636
rect 12740 41580 14924 41636
rect 14980 41580 15148 41636
rect 15362 41580 15372 41636
rect 15428 41580 16268 41636
rect 16324 41580 16334 41636
rect 4466 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4750 41580
rect 35186 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35470 41580
rect 12898 41468 12908 41524
rect 12964 41468 15820 41524
rect 15876 41468 15886 41524
rect 2258 41356 2268 41412
rect 2324 41356 8764 41412
rect 8820 41356 8830 41412
rect 14914 41356 14924 41412
rect 14980 41356 15708 41412
rect 15764 41356 16604 41412
rect 16660 41356 16670 41412
rect 36194 41356 36204 41412
rect 36260 41356 37212 41412
rect 37268 41356 37278 41412
rect 5842 41244 5852 41300
rect 5908 41244 6972 41300
rect 7028 41244 7038 41300
rect 13794 41244 13804 41300
rect 13860 41244 15036 41300
rect 15092 41244 15102 41300
rect 15250 41244 15260 41300
rect 15316 41244 16268 41300
rect 16324 41244 16334 41300
rect 31266 41244 31276 41300
rect 31332 41244 32284 41300
rect 32340 41244 32350 41300
rect 5730 41132 5740 41188
rect 5796 41132 8764 41188
rect 8820 41132 11900 41188
rect 11956 41132 11966 41188
rect 13570 41132 13580 41188
rect 13636 41132 13916 41188
rect 13972 41132 13982 41188
rect 15092 41132 22372 41188
rect 36194 41132 36204 41188
rect 36260 41132 38892 41188
rect 38948 41132 38958 41188
rect 44146 41132 44156 41188
rect 44212 41132 45724 41188
rect 45780 41132 45790 41188
rect 15092 41076 15148 41132
rect 22316 41076 22372 41132
rect 5058 41020 5068 41076
rect 5124 41020 7084 41076
rect 7140 41020 7150 41076
rect 7410 41020 7420 41076
rect 7476 41020 11004 41076
rect 11060 41020 15148 41076
rect 15922 41020 15932 41076
rect 15988 41020 15998 41076
rect 17378 41020 17388 41076
rect 17444 41020 18284 41076
rect 18340 41020 18900 41076
rect 22306 41020 22316 41076
rect 22372 41020 22382 41076
rect 33618 41020 33628 41076
rect 33684 41020 34300 41076
rect 34356 41020 34366 41076
rect 38210 41020 38220 41076
rect 38276 41020 39228 41076
rect 39284 41020 39294 41076
rect 39778 41020 39788 41076
rect 39844 41020 42364 41076
rect 42420 41020 42430 41076
rect 1810 40908 1820 40964
rect 1876 40908 2156 40964
rect 2212 40908 2222 40964
rect 13570 40908 13580 40964
rect 13636 40908 15596 40964
rect 15652 40908 15662 40964
rect 15932 40852 15988 41020
rect 18844 40964 18900 41020
rect 18844 40908 20636 40964
rect 20692 40908 20702 40964
rect 36418 40908 36428 40964
rect 36484 40908 37436 40964
rect 37492 40908 37502 40964
rect 41010 40908 41020 40964
rect 41076 40908 43708 40964
rect 43764 40908 43774 40964
rect 18844 40852 18900 40908
rect 12562 40796 12572 40852
rect 12628 40796 14028 40852
rect 14084 40796 15988 40852
rect 18834 40796 18844 40852
rect 18900 40796 18910 40852
rect 33506 40796 33516 40852
rect 33572 40796 34748 40852
rect 34804 40796 35196 40852
rect 35252 40796 42028 40852
rect 42084 40796 42700 40852
rect 42756 40796 42766 40852
rect 19826 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20110 40796
rect 8082 40684 8092 40740
rect 8148 40684 9772 40740
rect 9828 40684 10220 40740
rect 10276 40684 11228 40740
rect 11284 40684 11294 40740
rect 16034 40684 16044 40740
rect 16100 40684 17276 40740
rect 17332 40684 17342 40740
rect 38612 40684 39676 40740
rect 39732 40684 39742 40740
rect 38612 40628 38668 40684
rect 4834 40572 4844 40628
rect 4900 40572 7980 40628
rect 8036 40572 8046 40628
rect 15474 40572 15484 40628
rect 15540 40572 16156 40628
rect 16212 40572 16222 40628
rect 18050 40572 18060 40628
rect 18116 40572 18284 40628
rect 18340 40572 22876 40628
rect 22932 40572 26460 40628
rect 26516 40572 26526 40628
rect 34962 40572 34972 40628
rect 35028 40572 36316 40628
rect 36372 40572 38668 40628
rect 39330 40572 39340 40628
rect 39396 40572 41804 40628
rect 41860 40572 41870 40628
rect 5506 40460 5516 40516
rect 5572 40460 6300 40516
rect 6356 40460 6366 40516
rect 9762 40460 9772 40516
rect 9828 40460 11452 40516
rect 11508 40460 11518 40516
rect 12982 40460 13020 40516
rect 13076 40460 13086 40516
rect 16258 40460 16268 40516
rect 16324 40460 18620 40516
rect 18676 40460 18686 40516
rect 35634 40460 35644 40516
rect 35700 40460 37772 40516
rect 37828 40460 41692 40516
rect 41748 40460 44156 40516
rect 44212 40460 44222 40516
rect 0 40404 800 40432
rect 49200 40404 50000 40432
rect 0 40348 1596 40404
rect 1652 40348 1662 40404
rect 6178 40348 6188 40404
rect 6244 40348 11340 40404
rect 11396 40348 11406 40404
rect 13682 40348 13692 40404
rect 13748 40348 14252 40404
rect 14308 40348 14318 40404
rect 16706 40348 16716 40404
rect 16772 40348 18508 40404
rect 18564 40348 19180 40404
rect 19236 40348 19246 40404
rect 29138 40348 29148 40404
rect 29204 40348 29932 40404
rect 29988 40348 29998 40404
rect 38770 40348 38780 40404
rect 38836 40348 39788 40404
rect 39844 40348 39854 40404
rect 40226 40348 40236 40404
rect 40292 40348 44940 40404
rect 44996 40348 45006 40404
rect 46946 40348 46956 40404
rect 47012 40348 50000 40404
rect 0 40320 800 40348
rect 49200 40320 50000 40348
rect 2482 40236 2492 40292
rect 2548 40236 3724 40292
rect 3780 40236 3790 40292
rect 7522 40236 7532 40292
rect 7588 40236 9548 40292
rect 9604 40236 10108 40292
rect 10164 40236 10174 40292
rect 16034 40236 16044 40292
rect 16100 40236 20636 40292
rect 20692 40236 20702 40292
rect 20962 40236 20972 40292
rect 21028 40236 21756 40292
rect 21812 40236 21822 40292
rect 33954 40236 33964 40292
rect 34020 40236 35196 40292
rect 35252 40236 35262 40292
rect 2930 40124 2940 40180
rect 2996 40124 3388 40180
rect 3444 40124 3454 40180
rect 6626 40124 6636 40180
rect 6692 40124 8540 40180
rect 8596 40124 11788 40180
rect 11844 40124 13244 40180
rect 13300 40124 16268 40180
rect 16324 40124 16334 40180
rect 18162 40124 18172 40180
rect 18228 40124 19292 40180
rect 19348 40124 19852 40180
rect 19908 40124 19918 40180
rect 26002 40124 26012 40180
rect 26068 40124 28588 40180
rect 28644 40124 28654 40180
rect 34850 40124 34860 40180
rect 34916 40124 37324 40180
rect 37380 40124 37390 40180
rect 37762 40124 37772 40180
rect 37828 40124 41804 40180
rect 41860 40124 43484 40180
rect 43540 40124 43550 40180
rect 3490 40012 3500 40068
rect 3556 40012 4060 40068
rect 4116 40012 4126 40068
rect 23202 40012 23212 40068
rect 23268 40012 23660 40068
rect 23716 40012 33964 40068
rect 34020 40012 34030 40068
rect 41346 40012 41356 40068
rect 41412 40012 42028 40068
rect 42084 40012 45612 40068
rect 45668 40012 45678 40068
rect 4466 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4750 40012
rect 35186 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35470 40012
rect 2258 39788 2268 39844
rect 2324 39788 3164 39844
rect 3220 39788 3948 39844
rect 4004 39788 4014 39844
rect 8306 39788 8316 39844
rect 8372 39788 11564 39844
rect 11620 39788 12348 39844
rect 12404 39788 12414 39844
rect 12898 39788 12908 39844
rect 12964 39788 13468 39844
rect 13524 39788 13534 39844
rect 38658 39788 38668 39844
rect 38724 39788 42812 39844
rect 42868 39788 42878 39844
rect 43362 39788 43372 39844
rect 43428 39788 45500 39844
rect 45556 39788 45566 39844
rect 0 39732 800 39760
rect 49200 39732 50000 39760
rect 0 39676 2604 39732
rect 2660 39676 2996 39732
rect 3266 39676 3276 39732
rect 3332 39676 5964 39732
rect 6020 39676 6030 39732
rect 6748 39676 10892 39732
rect 10948 39676 10958 39732
rect 16006 39676 16044 39732
rect 16100 39676 16110 39732
rect 31938 39676 31948 39732
rect 32004 39676 32732 39732
rect 32788 39676 32798 39732
rect 35858 39676 35868 39732
rect 35924 39676 36428 39732
rect 36484 39676 37100 39732
rect 37156 39676 39004 39732
rect 39060 39676 40124 39732
rect 40180 39676 40190 39732
rect 45266 39676 45276 39732
rect 45332 39676 46060 39732
rect 46116 39676 46126 39732
rect 47842 39676 47852 39732
rect 47908 39676 50000 39732
rect 0 39648 800 39676
rect 2940 39620 2996 39676
rect 6748 39620 6804 39676
rect 49200 39648 50000 39676
rect 2940 39564 3500 39620
rect 3556 39564 3566 39620
rect 5842 39564 5852 39620
rect 5908 39564 5964 39620
rect 6020 39564 6030 39620
rect 6178 39564 6188 39620
rect 6244 39564 6748 39620
rect 6804 39564 6814 39620
rect 9986 39564 9996 39620
rect 10052 39564 14252 39620
rect 14308 39564 15820 39620
rect 15876 39564 17724 39620
rect 17780 39564 17790 39620
rect 24098 39564 24108 39620
rect 24164 39564 26124 39620
rect 26180 39564 26190 39620
rect 29250 39564 29260 39620
rect 29316 39564 30380 39620
rect 30436 39564 30446 39620
rect 2930 39452 2940 39508
rect 2996 39452 5404 39508
rect 5460 39452 6188 39508
rect 6244 39452 6254 39508
rect 10322 39452 10332 39508
rect 10388 39452 16996 39508
rect 17154 39452 17164 39508
rect 17220 39452 18844 39508
rect 18900 39452 18910 39508
rect 19058 39452 19068 39508
rect 19124 39452 19404 39508
rect 19460 39452 19470 39508
rect 24658 39452 24668 39508
rect 24724 39452 25228 39508
rect 25284 39452 25294 39508
rect 39890 39452 39900 39508
rect 39956 39452 40908 39508
rect 40964 39452 40974 39508
rect 16940 39396 16996 39452
rect 3490 39340 3500 39396
rect 3556 39340 6636 39396
rect 6692 39340 8540 39396
rect 8596 39340 8606 39396
rect 12226 39340 12236 39396
rect 12292 39340 12684 39396
rect 12740 39340 14588 39396
rect 14644 39340 14654 39396
rect 15222 39340 15260 39396
rect 15316 39340 15326 39396
rect 15586 39340 15596 39396
rect 15652 39340 16044 39396
rect 16100 39340 16110 39396
rect 16940 39340 20300 39396
rect 20356 39340 20366 39396
rect 26114 39340 26124 39396
rect 26180 39340 26796 39396
rect 26852 39340 27244 39396
rect 27300 39340 28476 39396
rect 28532 39340 29260 39396
rect 29316 39340 29326 39396
rect 3332 39228 6524 39284
rect 6580 39228 6590 39284
rect 6822 39228 6860 39284
rect 6916 39228 15148 39284
rect 15204 39228 17612 39284
rect 17668 39228 17678 39284
rect 27010 39228 27020 39284
rect 27076 39228 29036 39284
rect 29092 39228 29820 39284
rect 29876 39228 29886 39284
rect 3332 39172 3388 39228
rect 19826 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20110 39228
rect 1362 39116 1372 39172
rect 1428 39116 3388 39172
rect 4386 39116 4396 39172
rect 4452 39116 8652 39172
rect 8708 39116 8718 39172
rect 14690 39116 14700 39172
rect 14756 39116 14924 39172
rect 14980 39116 14990 39172
rect 15250 39116 15260 39172
rect 15316 39116 15820 39172
rect 15876 39116 15886 39172
rect 49200 39060 50000 39088
rect 3826 39004 3836 39060
rect 3892 39004 4284 39060
rect 4340 39004 4350 39060
rect 5282 39004 5292 39060
rect 5348 39004 5852 39060
rect 5908 39004 6748 39060
rect 6804 39004 6814 39060
rect 8530 39004 8540 39060
rect 8596 39004 8876 39060
rect 8932 39004 11788 39060
rect 11844 39004 12124 39060
rect 12180 39004 14476 39060
rect 14532 39004 14542 39060
rect 14914 39004 14924 39060
rect 14980 39004 15708 39060
rect 15764 39004 16492 39060
rect 16548 39004 16558 39060
rect 18610 39004 18620 39060
rect 18676 39004 22652 39060
rect 22708 39004 22718 39060
rect 30482 39004 30492 39060
rect 30548 39004 31836 39060
rect 31892 39004 34524 39060
rect 34580 39004 34590 39060
rect 38612 39004 39564 39060
rect 39620 39004 40012 39060
rect 40068 39004 40348 39060
rect 40404 39004 41692 39060
rect 41748 39004 47516 39060
rect 47572 39004 47582 39060
rect 47954 39004 47964 39060
rect 48020 39004 50000 39060
rect 38612 38948 38668 39004
rect 49200 38976 50000 39004
rect 3154 38892 3164 38948
rect 3220 38892 6020 38948
rect 6290 38892 6300 38948
rect 6356 38892 7084 38948
rect 7140 38892 9884 38948
rect 9940 38892 9950 38948
rect 19506 38892 19516 38948
rect 19572 38892 20188 38948
rect 20244 38892 20254 38948
rect 30034 38892 30044 38948
rect 30100 38892 31052 38948
rect 31108 38892 31118 38948
rect 38098 38892 38108 38948
rect 38164 38892 38668 38948
rect 4722 38780 4732 38836
rect 4788 38780 5740 38836
rect 5796 38780 5806 38836
rect 5964 38612 6020 38892
rect 11330 38780 11340 38836
rect 11396 38780 13356 38836
rect 13412 38780 16884 38836
rect 18050 38780 18060 38836
rect 18116 38780 18788 38836
rect 20290 38780 20300 38836
rect 20356 38780 22092 38836
rect 22148 38780 22158 38836
rect 33394 38780 33404 38836
rect 33460 38780 34076 38836
rect 34132 38780 34142 38836
rect 39890 38780 39900 38836
rect 39956 38780 45836 38836
rect 45892 38780 45902 38836
rect 16828 38724 16884 38780
rect 15474 38668 15484 38724
rect 15540 38668 15932 38724
rect 15988 38668 16380 38724
rect 16436 38668 16446 38724
rect 16818 38668 16828 38724
rect 16884 38668 17388 38724
rect 17444 38668 17454 38724
rect 4610 38556 4620 38612
rect 4676 38556 4956 38612
rect 5012 38556 5022 38612
rect 5954 38556 5964 38612
rect 6020 38556 6030 38612
rect 8306 38556 8316 38612
rect 8372 38556 8428 38612
rect 8484 38556 8494 38612
rect 15334 38556 15372 38612
rect 15428 38556 15438 38612
rect 18732 38500 18788 38780
rect 21532 38612 21588 38780
rect 27682 38668 27692 38724
rect 27748 38668 29484 38724
rect 29540 38668 29550 38724
rect 30370 38668 30380 38724
rect 30436 38668 32284 38724
rect 32340 38668 32350 38724
rect 37538 38668 37548 38724
rect 37604 38668 38668 38724
rect 38724 38668 40684 38724
rect 40740 38668 40750 38724
rect 21522 38556 21532 38612
rect 21588 38556 21598 38612
rect 21970 38556 21980 38612
rect 22036 38556 23324 38612
rect 23380 38556 23390 38612
rect 31378 38556 31388 38612
rect 31444 38556 32172 38612
rect 32228 38556 33292 38612
rect 33348 38556 33358 38612
rect 34402 38556 34412 38612
rect 34468 38556 35196 38612
rect 35252 38556 37772 38612
rect 37828 38556 37838 38612
rect 8530 38444 8540 38500
rect 8596 38444 9660 38500
rect 9716 38444 17724 38500
rect 17780 38444 17790 38500
rect 18722 38444 18732 38500
rect 18788 38444 18798 38500
rect 0 38388 800 38416
rect 4466 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4750 38444
rect 17724 38388 17780 38444
rect 35186 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35470 38444
rect 0 38332 1708 38388
rect 1764 38332 1774 38388
rect 7634 38332 7644 38388
rect 7700 38332 7756 38388
rect 7812 38332 9324 38388
rect 9380 38332 9390 38388
rect 11330 38332 11340 38388
rect 11396 38332 11406 38388
rect 17724 38332 22876 38388
rect 22932 38332 22942 38388
rect 0 38304 800 38332
rect 11340 38276 11396 38332
rect 3332 38220 11396 38276
rect 18498 38220 18508 38276
rect 18564 38220 19852 38276
rect 19908 38220 19918 38276
rect 3332 38164 3388 38220
rect 2258 38108 2268 38164
rect 2324 38108 3388 38164
rect 3490 38108 3500 38164
rect 3556 38108 4172 38164
rect 4228 38108 4238 38164
rect 6822 38108 6860 38164
rect 6916 38108 6926 38164
rect 7634 38108 7644 38164
rect 7700 38108 8316 38164
rect 8372 38108 8382 38164
rect 13906 38108 13916 38164
rect 13972 38108 18956 38164
rect 19012 38108 19404 38164
rect 19460 38108 19470 38164
rect 43138 38108 43148 38164
rect 43204 38108 44156 38164
rect 44212 38108 44940 38164
rect 44996 38108 45006 38164
rect 1698 37996 1708 38052
rect 1764 37996 3388 38052
rect 3444 37996 3454 38052
rect 4386 37996 4396 38052
rect 4452 37996 4956 38052
rect 5012 37996 5022 38052
rect 8978 37996 8988 38052
rect 9044 37996 9436 38052
rect 9492 37996 9502 38052
rect 11106 37996 11116 38052
rect 11172 37996 12348 38052
rect 12404 37996 13804 38052
rect 13860 37996 13870 38052
rect 15334 37996 15372 38052
rect 15428 37996 15438 38052
rect 15922 37996 15932 38052
rect 15988 37996 16268 38052
rect 16324 37996 16334 38052
rect 17154 37996 17164 38052
rect 17220 37996 17836 38052
rect 17892 37996 17902 38052
rect 22754 37996 22764 38052
rect 22820 37996 26012 38052
rect 26068 37996 26078 38052
rect 43362 37996 43372 38052
rect 43428 37996 48188 38052
rect 48244 37996 48254 38052
rect 0 37716 800 37744
rect 1708 37716 1764 37996
rect 2818 37884 2828 37940
rect 2884 37884 4508 37940
rect 4564 37884 4574 37940
rect 5170 37884 5180 37940
rect 5236 37884 6188 37940
rect 6244 37884 6254 37940
rect 11218 37884 11228 37940
rect 11284 37884 12460 37940
rect 12516 37884 14364 37940
rect 14420 37884 14430 37940
rect 17490 37884 17500 37940
rect 17556 37884 18060 37940
rect 18116 37884 18508 37940
rect 18564 37884 18574 37940
rect 20402 37884 20412 37940
rect 20468 37884 21644 37940
rect 21700 37884 21710 37940
rect 36194 37884 36204 37940
rect 36260 37884 37212 37940
rect 37268 37884 37278 37940
rect 41682 37884 41692 37940
rect 41748 37884 46060 37940
rect 46116 37884 46126 37940
rect 3602 37772 3612 37828
rect 3668 37772 6076 37828
rect 6132 37772 6142 37828
rect 10882 37772 10892 37828
rect 10948 37772 13804 37828
rect 13860 37772 13870 37828
rect 14018 37772 14028 37828
rect 14084 37772 16044 37828
rect 16100 37772 16110 37828
rect 17714 37772 17724 37828
rect 17780 37772 17790 37828
rect 22866 37772 22876 37828
rect 22932 37772 24220 37828
rect 24276 37772 24286 37828
rect 41458 37772 41468 37828
rect 41524 37772 43036 37828
rect 43092 37772 43102 37828
rect 17724 37716 17780 37772
rect 0 37660 1764 37716
rect 3798 37660 3836 37716
rect 3892 37660 3902 37716
rect 4162 37660 4172 37716
rect 4228 37660 6860 37716
rect 6916 37660 6926 37716
rect 12450 37660 12460 37716
rect 12516 37660 17780 37716
rect 0 37632 800 37660
rect 19826 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20110 37660
rect 2828 37548 3052 37604
rect 3108 37548 5068 37604
rect 5124 37548 5134 37604
rect 10210 37548 10220 37604
rect 10276 37548 15036 37604
rect 15092 37548 15102 37604
rect 15698 37548 15708 37604
rect 15764 37548 18732 37604
rect 18788 37548 18798 37604
rect 23734 37548 23772 37604
rect 23828 37548 23838 37604
rect 2828 37492 2884 37548
rect 2818 37436 2828 37492
rect 2884 37436 2894 37492
rect 3602 37436 3612 37492
rect 3668 37436 3948 37492
rect 4004 37436 4014 37492
rect 4918 37436 4956 37492
rect 5012 37436 5022 37492
rect 9650 37436 9660 37492
rect 9716 37436 13244 37492
rect 13300 37436 13310 37492
rect 15138 37436 15148 37492
rect 15204 37436 15820 37492
rect 15876 37436 17276 37492
rect 17332 37436 17342 37492
rect 19282 37436 19292 37492
rect 19348 37436 19358 37492
rect 19506 37436 19516 37492
rect 19572 37436 20188 37492
rect 20244 37436 20254 37492
rect 22754 37436 22764 37492
rect 22820 37436 23436 37492
rect 23492 37436 24668 37492
rect 24724 37436 24734 37492
rect 32162 37436 32172 37492
rect 32228 37436 35420 37492
rect 35476 37436 35486 37492
rect 39890 37436 39900 37492
rect 39956 37436 41020 37492
rect 41076 37436 42140 37492
rect 42196 37436 43708 37492
rect 19292 37380 19348 37436
rect 3042 37324 3052 37380
rect 3108 37324 8204 37380
rect 8260 37324 9996 37380
rect 10052 37324 10062 37380
rect 10322 37324 10332 37380
rect 10388 37324 11676 37380
rect 11732 37324 11742 37380
rect 14802 37324 14812 37380
rect 14868 37324 17724 37380
rect 17780 37324 19348 37380
rect 20850 37324 20860 37380
rect 20916 37324 21644 37380
rect 21700 37324 21710 37380
rect 22530 37324 22540 37380
rect 22596 37324 23548 37380
rect 23604 37324 25340 37380
rect 25396 37324 25406 37380
rect 43652 37268 43708 37436
rect 3500 37212 4172 37268
rect 4228 37212 4238 37268
rect 4722 37212 4732 37268
rect 4788 37212 8092 37268
rect 8148 37212 8158 37268
rect 9314 37212 9324 37268
rect 9380 37212 9884 37268
rect 9940 37212 9950 37268
rect 10658 37212 10668 37268
rect 10724 37212 11564 37268
rect 11620 37212 11630 37268
rect 12786 37212 12796 37268
rect 12852 37212 13580 37268
rect 13636 37212 13646 37268
rect 16342 37212 16380 37268
rect 16436 37212 16446 37268
rect 16594 37212 16604 37268
rect 16660 37212 17388 37268
rect 17444 37212 17454 37268
rect 20290 37212 20300 37268
rect 20356 37212 21084 37268
rect 21140 37212 21868 37268
rect 21924 37212 21934 37268
rect 23314 37212 23324 37268
rect 23380 37212 24332 37268
rect 24388 37212 24398 37268
rect 43652 37212 44940 37268
rect 44996 37212 45006 37268
rect 3500 37156 3556 37212
rect 3490 37100 3500 37156
rect 3556 37100 3566 37156
rect 3938 37100 3948 37156
rect 4004 37100 8204 37156
rect 8260 37100 8270 37156
rect 10098 37100 10108 37156
rect 10164 37100 10174 37156
rect 11106 37100 11116 37156
rect 11172 37100 17332 37156
rect 18722 37100 18732 37156
rect 18788 37100 21532 37156
rect 21588 37100 21598 37156
rect 23846 37100 23884 37156
rect 23940 37100 23950 37156
rect 42018 37100 42028 37156
rect 42084 37100 43932 37156
rect 43988 37100 43998 37156
rect 10108 37044 10164 37100
rect 2034 36988 2044 37044
rect 2100 36988 3388 37044
rect 3714 36988 3724 37044
rect 3780 36988 4732 37044
rect 4788 36988 4798 37044
rect 5618 36988 5628 37044
rect 5684 36988 5964 37044
rect 6020 36988 6030 37044
rect 7410 36988 7420 37044
rect 7476 36988 9660 37044
rect 9716 36988 9726 37044
rect 10108 36988 11004 37044
rect 11060 36988 11070 37044
rect 1698 36876 1708 36932
rect 1764 36876 2940 36932
rect 2996 36876 3006 36932
rect 3332 36708 3388 36988
rect 17276 36932 17332 37100
rect 17276 36876 19572 36932
rect 37090 36876 37100 36932
rect 37156 36876 39452 36932
rect 39508 36876 39518 36932
rect 4466 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4750 36876
rect 19516 36820 19572 36876
rect 35186 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35470 36876
rect 9986 36764 9996 36820
rect 10052 36764 10444 36820
rect 10500 36764 11116 36820
rect 11172 36764 11182 36820
rect 11442 36764 11452 36820
rect 11508 36764 12796 36820
rect 12852 36764 12862 36820
rect 18722 36764 18732 36820
rect 18788 36764 19180 36820
rect 19236 36764 19246 36820
rect 19506 36764 19516 36820
rect 19572 36764 19582 36820
rect 20738 36764 20748 36820
rect 20804 36764 22988 36820
rect 23044 36764 23054 36820
rect 29474 36764 29484 36820
rect 29540 36764 31276 36820
rect 31332 36764 31342 36820
rect 3332 36652 10500 36708
rect 11554 36652 11564 36708
rect 11620 36652 14140 36708
rect 14196 36652 14206 36708
rect 15092 36652 15932 36708
rect 15988 36652 15998 36708
rect 10444 36596 10500 36652
rect 15092 36596 15148 36652
rect 4162 36540 4172 36596
rect 4228 36540 4732 36596
rect 4788 36540 4844 36596
rect 4900 36540 4910 36596
rect 6402 36540 6412 36596
rect 6468 36540 7420 36596
rect 7476 36540 7486 36596
rect 10444 36540 11676 36596
rect 11732 36540 11742 36596
rect 12898 36540 12908 36596
rect 12964 36540 13692 36596
rect 13748 36540 13758 36596
rect 14578 36540 14588 36596
rect 14644 36540 15148 36596
rect 16818 36540 16828 36596
rect 16884 36540 18284 36596
rect 18340 36540 20412 36596
rect 20468 36540 20478 36596
rect 26852 36540 28028 36596
rect 28084 36540 29484 36596
rect 29540 36540 29820 36596
rect 29876 36540 29886 36596
rect 38210 36540 38220 36596
rect 38276 36540 39900 36596
rect 39956 36540 39966 36596
rect 26852 36484 26908 36540
rect 3332 36428 7308 36484
rect 7364 36428 7374 36484
rect 7522 36428 7532 36484
rect 7588 36428 7756 36484
rect 7812 36428 7822 36484
rect 24098 36428 24108 36484
rect 24164 36428 26908 36484
rect 29250 36428 29260 36484
rect 29316 36428 31612 36484
rect 31668 36428 31678 36484
rect 35298 36428 35308 36484
rect 35364 36428 36316 36484
rect 36372 36428 39004 36484
rect 39060 36428 42476 36484
rect 42532 36428 43148 36484
rect 43204 36428 43214 36484
rect 3332 36260 3388 36428
rect 6178 36316 6188 36372
rect 6244 36316 13356 36372
rect 13412 36316 13422 36372
rect 14886 36316 14924 36372
rect 14980 36316 14990 36372
rect 16594 36316 16604 36372
rect 16660 36316 17052 36372
rect 17108 36316 17118 36372
rect 44146 36316 44156 36372
rect 44212 36316 45052 36372
rect 45108 36316 45118 36372
rect 2258 36204 2268 36260
rect 2324 36204 3164 36260
rect 3220 36204 3388 36260
rect 7084 36204 9100 36260
rect 9156 36204 9772 36260
rect 9828 36204 9838 36260
rect 12338 36204 12348 36260
rect 12404 36204 13020 36260
rect 13076 36204 13804 36260
rect 13860 36204 14588 36260
rect 14644 36204 14654 36260
rect 15026 36204 15036 36260
rect 15092 36204 17164 36260
rect 17220 36204 17230 36260
rect 21858 36204 21868 36260
rect 21924 36204 22652 36260
rect 22708 36204 22718 36260
rect 26114 36204 26124 36260
rect 26180 36204 27244 36260
rect 27300 36204 27310 36260
rect 31378 36204 31388 36260
rect 31444 36204 34860 36260
rect 34916 36204 35756 36260
rect 35812 36204 35822 36260
rect 7084 36148 7140 36204
rect 12348 36148 12404 36204
rect 7074 36092 7084 36148
rect 7140 36092 7150 36148
rect 7606 36092 7644 36148
rect 7700 36092 7710 36148
rect 8194 36092 8204 36148
rect 8260 36092 8540 36148
rect 8596 36092 8606 36148
rect 9426 36092 9436 36148
rect 9492 36092 12404 36148
rect 16230 36092 16268 36148
rect 16324 36092 16334 36148
rect 19826 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20110 36092
rect 5842 35980 5852 36036
rect 5908 35980 5964 36036
rect 6020 35980 13580 36036
rect 13636 35980 13646 36036
rect 17602 35980 17612 36036
rect 17668 35980 18284 36036
rect 18340 35980 18350 36036
rect 18946 35980 18956 36036
rect 19012 35980 19068 36036
rect 19124 35980 19134 36036
rect 5394 35868 5404 35924
rect 5460 35868 5628 35924
rect 5684 35868 6636 35924
rect 6692 35868 6702 35924
rect 14690 35868 14700 35924
rect 14756 35868 19964 35924
rect 20020 35868 20030 35924
rect 23426 35868 23436 35924
rect 23492 35868 24332 35924
rect 24388 35868 24398 35924
rect 32610 35868 32620 35924
rect 32676 35868 33292 35924
rect 33348 35868 33358 35924
rect 40114 35868 40124 35924
rect 40180 35868 41692 35924
rect 41748 35868 41758 35924
rect 43652 35868 45612 35924
rect 45668 35868 45678 35924
rect 43652 35812 43708 35868
rect 5058 35756 5068 35812
rect 5124 35756 6860 35812
rect 6916 35756 6926 35812
rect 8082 35756 8092 35812
rect 8148 35756 8988 35812
rect 9044 35756 9884 35812
rect 9940 35756 9950 35812
rect 10882 35756 10892 35812
rect 10948 35756 11340 35812
rect 11396 35756 11406 35812
rect 16006 35756 16044 35812
rect 16100 35756 16604 35812
rect 16660 35756 16670 35812
rect 17686 35756 17724 35812
rect 17780 35756 18060 35812
rect 18116 35756 18126 35812
rect 19394 35756 19404 35812
rect 19460 35756 21532 35812
rect 21588 35756 21598 35812
rect 40226 35756 40236 35812
rect 40292 35756 43708 35812
rect 0 35700 800 35728
rect 10892 35700 10948 35756
rect 0 35644 1708 35700
rect 1764 35644 1774 35700
rect 3266 35644 3276 35700
rect 3332 35644 5740 35700
rect 5796 35644 5806 35700
rect 7858 35644 7868 35700
rect 7924 35644 8204 35700
rect 8260 35644 8428 35700
rect 8484 35644 8494 35700
rect 9650 35644 9660 35700
rect 9716 35644 10948 35700
rect 12348 35644 16828 35700
rect 16884 35644 16894 35700
rect 17798 35644 17836 35700
rect 17892 35644 17902 35700
rect 20850 35644 20860 35700
rect 20916 35644 23324 35700
rect 23380 35644 23390 35700
rect 30818 35644 30828 35700
rect 30884 35644 31612 35700
rect 31668 35644 32060 35700
rect 32116 35644 32126 35700
rect 44594 35644 44604 35700
rect 44660 35644 47068 35700
rect 47124 35644 47852 35700
rect 47908 35644 47918 35700
rect 0 35616 800 35644
rect 12348 35476 12404 35644
rect 16146 35532 16156 35588
rect 16212 35532 16380 35588
rect 16436 35532 16446 35588
rect 18274 35532 18284 35588
rect 18340 35532 25900 35588
rect 25956 35532 25966 35588
rect 16380 35476 16436 35532
rect 12338 35420 12348 35476
rect 12404 35420 12414 35476
rect 14578 35420 14588 35476
rect 14644 35420 15708 35476
rect 15764 35420 15774 35476
rect 16370 35420 16380 35476
rect 16436 35420 16446 35476
rect 10434 35308 10444 35364
rect 10500 35308 13244 35364
rect 13300 35308 13310 35364
rect 16230 35308 16268 35364
rect 16324 35308 16334 35364
rect 23734 35308 23772 35364
rect 23828 35308 23838 35364
rect 23986 35308 23996 35364
rect 24052 35308 24062 35364
rect 39778 35308 39788 35364
rect 39844 35308 42420 35364
rect 4466 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4750 35308
rect 23996 35252 24052 35308
rect 35186 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35470 35308
rect 1810 35196 1820 35252
rect 1876 35196 2156 35252
rect 2212 35196 2222 35252
rect 2706 35196 2716 35252
rect 2772 35196 4060 35252
rect 4116 35196 4126 35252
rect 5926 35196 5964 35252
rect 6020 35196 7420 35252
rect 7476 35196 7486 35252
rect 9538 35196 9548 35252
rect 9604 35196 9772 35252
rect 9828 35196 9838 35252
rect 11106 35196 11116 35252
rect 11172 35196 12236 35252
rect 12292 35196 12302 35252
rect 13570 35196 13580 35252
rect 13636 35196 17500 35252
rect 17556 35196 21532 35252
rect 21588 35196 21598 35252
rect 21746 35196 21756 35252
rect 21812 35196 22988 35252
rect 23044 35196 26124 35252
rect 26180 35196 26190 35252
rect 0 35028 800 35056
rect 1820 35028 1876 35196
rect 21532 35140 21588 35196
rect 42364 35140 42420 35308
rect 43260 35308 43708 35364
rect 43260 35252 43316 35308
rect 43652 35252 43708 35308
rect 43250 35196 43260 35252
rect 43316 35196 43326 35252
rect 43652 35196 44268 35252
rect 44324 35196 45836 35252
rect 45892 35196 45902 35252
rect 2258 35084 2268 35140
rect 2324 35084 8428 35140
rect 8484 35084 8764 35140
rect 8820 35084 8830 35140
rect 9426 35084 9436 35140
rect 9492 35084 10892 35140
rect 10948 35084 10958 35140
rect 11302 35084 11340 35140
rect 11396 35084 11406 35140
rect 14028 35084 15148 35140
rect 17938 35084 17948 35140
rect 18004 35084 18508 35140
rect 18564 35084 18574 35140
rect 19170 35084 19180 35140
rect 19236 35084 19740 35140
rect 19796 35084 19806 35140
rect 21532 35084 22540 35140
rect 22596 35084 22606 35140
rect 42364 35084 43316 35140
rect 43474 35084 43484 35140
rect 43540 35084 46228 35140
rect 14028 35028 14084 35084
rect 15092 35028 15148 35084
rect 43260 35028 43316 35084
rect 46172 35028 46228 35084
rect 49200 35028 50000 35056
rect 0 34972 1876 35028
rect 2044 34972 3612 35028
rect 3668 34972 3678 35028
rect 3826 34972 3836 35028
rect 3892 34972 3930 35028
rect 5030 34972 5068 35028
rect 5124 34972 5134 35028
rect 5954 34972 5964 35028
rect 6020 34972 6300 35028
rect 6356 34972 6366 35028
rect 6626 34972 6636 35028
rect 6692 34972 7196 35028
rect 7252 34972 7262 35028
rect 8866 34972 8876 35028
rect 8932 34972 10108 35028
rect 10164 34972 14084 35028
rect 14242 34972 14252 35028
rect 14308 34972 14924 35028
rect 14980 34972 14990 35028
rect 15092 34972 15260 35028
rect 15316 34972 15326 35028
rect 17714 34972 17724 35028
rect 17780 34972 18732 35028
rect 18788 34972 18798 35028
rect 18946 34972 18956 35028
rect 19012 34972 19292 35028
rect 19348 34972 19358 35028
rect 19628 34972 21308 35028
rect 21364 34972 21374 35028
rect 28018 34972 28028 35028
rect 28084 34972 29148 35028
rect 29204 34972 29214 35028
rect 41346 34972 41356 35028
rect 41412 34972 42252 35028
rect 42308 34972 42318 35028
rect 43260 34972 45052 35028
rect 45108 34972 45118 35028
rect 46172 34972 50000 35028
rect 0 34944 800 34972
rect 2044 34916 2100 34972
rect 19628 34916 19684 34972
rect 49200 34944 50000 34972
rect 1698 34860 1708 34916
rect 1764 34860 2100 34916
rect 2930 34860 2940 34916
rect 2996 34860 3500 34916
rect 3556 34860 3566 34916
rect 3714 34860 3724 34916
rect 3780 34860 6020 34916
rect 9426 34860 9436 34916
rect 9492 34860 10556 34916
rect 10612 34860 10622 34916
rect 12898 34860 12908 34916
rect 12964 34860 14028 34916
rect 14084 34860 14094 34916
rect 14438 34860 14476 34916
rect 14532 34860 14542 34916
rect 15026 34860 15036 34916
rect 15092 34860 15484 34916
rect 15540 34860 15550 34916
rect 17602 34860 17612 34916
rect 17668 34860 19628 34916
rect 19684 34860 19694 34916
rect 20066 34860 20076 34916
rect 20132 34860 22428 34916
rect 22484 34860 22494 34916
rect 22754 34860 22764 34916
rect 22820 34860 22876 34916
rect 22932 34860 23212 34916
rect 23268 34860 23548 34916
rect 31378 34860 31388 34916
rect 31444 34860 33460 34916
rect 41122 34860 41132 34916
rect 41188 34860 42812 34916
rect 42868 34860 42878 34916
rect 5964 34804 6020 34860
rect 3378 34748 3388 34804
rect 3444 34748 4396 34804
rect 4452 34748 4462 34804
rect 5954 34748 5964 34804
rect 6020 34748 6030 34804
rect 7522 34748 7532 34804
rect 7588 34748 8540 34804
rect 8596 34748 9884 34804
rect 9940 34748 9950 34804
rect 10098 34748 10108 34804
rect 10164 34748 10202 34804
rect 10434 34748 10444 34804
rect 10500 34748 11116 34804
rect 11172 34748 11182 34804
rect 11666 34748 11676 34804
rect 11732 34748 14140 34804
rect 14196 34748 14206 34804
rect 17938 34748 17948 34804
rect 18004 34748 18844 34804
rect 18900 34748 18910 34804
rect 19058 34748 19068 34804
rect 19124 34748 19134 34804
rect 19506 34748 19516 34804
rect 19572 34748 19852 34804
rect 19908 34748 19918 34804
rect 20178 34748 20188 34804
rect 20244 34748 22540 34804
rect 22596 34748 22606 34804
rect 19068 34692 19124 34748
rect 23492 34692 23548 34860
rect 33404 34804 33460 34860
rect 26450 34748 26460 34804
rect 26516 34748 28140 34804
rect 28196 34748 28206 34804
rect 29922 34748 29932 34804
rect 29988 34748 32060 34804
rect 32116 34748 32126 34804
rect 33394 34748 33404 34804
rect 33460 34748 35532 34804
rect 35588 34748 35598 34804
rect 42242 34748 42252 34804
rect 42308 34748 44940 34804
rect 44996 34748 45006 34804
rect 2930 34636 2940 34692
rect 2996 34636 3006 34692
rect 3602 34636 3612 34692
rect 3668 34636 11452 34692
rect 11508 34636 11518 34692
rect 14578 34636 14588 34692
rect 14644 34636 16380 34692
rect 16436 34636 16446 34692
rect 18498 34636 18508 34692
rect 18564 34636 18956 34692
rect 19012 34636 19124 34692
rect 19282 34636 19292 34692
rect 19348 34636 19740 34692
rect 19796 34636 19806 34692
rect 23492 34636 24108 34692
rect 24164 34636 24174 34692
rect 24630 34636 24668 34692
rect 24724 34636 24734 34692
rect 34850 34636 34860 34692
rect 34916 34636 36092 34692
rect 36148 34636 36158 34692
rect 37762 34636 37772 34692
rect 37828 34636 40908 34692
rect 40964 34636 42364 34692
rect 42420 34636 44604 34692
rect 44660 34636 45164 34692
rect 45220 34636 45230 34692
rect 1810 34524 1820 34580
rect 1876 34524 2604 34580
rect 2660 34524 2670 34580
rect 2940 34468 2996 34636
rect 3332 34524 16716 34580
rect 16772 34524 16782 34580
rect 22754 34524 22764 34580
rect 22820 34524 22830 34580
rect 41346 34524 41356 34580
rect 41412 34524 43820 34580
rect 43876 34524 43886 34580
rect 3332 34468 3388 34524
rect 19826 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20110 34524
rect 2940 34412 3388 34468
rect 3602 34412 3612 34468
rect 3668 34412 4284 34468
rect 4340 34412 4350 34468
rect 8166 34412 8204 34468
rect 8260 34412 8270 34468
rect 10770 34412 10780 34468
rect 10836 34412 12572 34468
rect 12628 34412 12638 34468
rect 13542 34412 13580 34468
rect 13636 34412 13646 34468
rect 14354 34412 14364 34468
rect 14420 34412 15596 34468
rect 15652 34412 15662 34468
rect 22764 34356 22820 34524
rect 49200 34356 50000 34384
rect 2594 34300 2604 34356
rect 2660 34300 2670 34356
rect 2930 34300 2940 34356
rect 2996 34300 3612 34356
rect 3668 34300 3836 34356
rect 3892 34300 3902 34356
rect 4722 34300 4732 34356
rect 4788 34300 5180 34356
rect 5236 34300 6188 34356
rect 6244 34300 6254 34356
rect 6402 34300 6412 34356
rect 6468 34300 6748 34356
rect 6804 34300 6814 34356
rect 8754 34300 8764 34356
rect 8820 34300 9436 34356
rect 9492 34300 9502 34356
rect 10546 34300 10556 34356
rect 10612 34300 11340 34356
rect 11396 34300 11406 34356
rect 16258 34300 16268 34356
rect 16324 34300 16940 34356
rect 16996 34300 17006 34356
rect 18722 34300 18732 34356
rect 18788 34300 19852 34356
rect 19908 34300 19918 34356
rect 21858 34300 21868 34356
rect 21924 34300 25340 34356
rect 25396 34300 25406 34356
rect 47954 34300 47964 34356
rect 48020 34300 50000 34356
rect 2604 34132 2660 34300
rect 2818 34188 2828 34244
rect 2884 34188 3388 34244
rect 3444 34188 3454 34244
rect 6850 34188 6860 34244
rect 6916 34188 8876 34244
rect 8932 34188 9212 34244
rect 9268 34188 9278 34244
rect 10322 34188 10332 34244
rect 10388 34188 10500 34244
rect 12450 34188 12460 34244
rect 12516 34188 12684 34244
rect 12740 34188 12750 34244
rect 15092 34188 15596 34244
rect 15652 34188 15662 34244
rect 18946 34188 18956 34244
rect 19012 34188 19628 34244
rect 19684 34188 19694 34244
rect 2604 34076 4396 34132
rect 4452 34076 10220 34132
rect 10276 34076 10286 34132
rect 10444 34020 10500 34188
rect 15092 34132 15148 34188
rect 22540 34132 22596 34300
rect 49200 34272 50000 34300
rect 28802 34188 28812 34244
rect 28868 34188 29932 34244
rect 29988 34188 29998 34244
rect 43138 34188 43148 34244
rect 43204 34188 44156 34244
rect 44212 34188 44222 34244
rect 12786 34076 12796 34132
rect 12852 34076 13020 34132
rect 13076 34076 13086 34132
rect 14578 34076 14588 34132
rect 14644 34076 15148 34132
rect 17938 34076 17948 34132
rect 18004 34076 19180 34132
rect 19236 34076 19246 34132
rect 22530 34076 22540 34132
rect 22596 34076 22606 34132
rect 22978 34076 22988 34132
rect 23044 34076 24668 34132
rect 24724 34076 25788 34132
rect 25844 34076 25854 34132
rect 6626 33964 6636 34020
rect 6692 33964 7308 34020
rect 7364 33964 8708 34020
rect 9314 33964 9324 34020
rect 9380 33964 10052 34020
rect 10434 33964 10444 34020
rect 10500 33964 10510 34020
rect 16706 33964 16716 34020
rect 16772 33964 17388 34020
rect 17444 33964 17454 34020
rect 24210 33964 24220 34020
rect 24276 33964 26012 34020
rect 26068 33964 26078 34020
rect 29250 33964 29260 34020
rect 29316 33964 30268 34020
rect 30324 33964 30334 34020
rect 33506 33964 33516 34020
rect 33572 33964 35756 34020
rect 35812 33964 35822 34020
rect 43810 33964 43820 34020
rect 43876 33964 44268 34020
rect 44324 33964 44334 34020
rect 8652 33908 8708 33964
rect 9996 33908 10052 33964
rect 1698 33852 1708 33908
rect 1764 33852 2044 33908
rect 2100 33852 2110 33908
rect 3378 33852 3388 33908
rect 3444 33852 7812 33908
rect 8642 33852 8652 33908
rect 8708 33852 9660 33908
rect 9716 33852 9726 33908
rect 9996 33852 10332 33908
rect 10388 33852 10398 33908
rect 15250 33852 15260 33908
rect 15316 33852 28364 33908
rect 28420 33852 28430 33908
rect 32050 33852 32060 33908
rect 32116 33852 33852 33908
rect 33908 33852 33918 33908
rect 35522 33852 35532 33908
rect 35588 33852 37100 33908
rect 37156 33852 37166 33908
rect 7756 33796 7812 33852
rect 7746 33740 7756 33796
rect 7812 33740 10052 33796
rect 11442 33740 11452 33796
rect 11508 33740 13468 33796
rect 13524 33740 13534 33796
rect 15698 33740 15708 33796
rect 15764 33740 17500 33796
rect 17556 33740 19516 33796
rect 19572 33740 19582 33796
rect 0 33684 800 33712
rect 4466 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4750 33740
rect 9996 33684 10052 33740
rect 35186 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35470 33740
rect 49200 33684 50000 33712
rect 0 33628 2604 33684
rect 2660 33628 2670 33684
rect 6402 33628 6412 33684
rect 6468 33628 6972 33684
rect 7028 33628 7420 33684
rect 7476 33628 7486 33684
rect 8530 33628 8540 33684
rect 8596 33628 9212 33684
rect 9268 33628 9278 33684
rect 9986 33628 9996 33684
rect 10052 33628 10556 33684
rect 10612 33628 10622 33684
rect 13122 33628 13132 33684
rect 13188 33628 13692 33684
rect 13748 33628 13758 33684
rect 17378 33628 17388 33684
rect 17444 33628 19292 33684
rect 19348 33628 19358 33684
rect 23090 33628 23100 33684
rect 23156 33628 23772 33684
rect 23828 33628 23838 33684
rect 24322 33628 24332 33684
rect 24388 33628 24892 33684
rect 24948 33628 24958 33684
rect 37426 33628 37436 33684
rect 37492 33628 39340 33684
rect 39396 33628 40908 33684
rect 40964 33628 40974 33684
rect 47394 33628 47404 33684
rect 47460 33628 50000 33684
rect 0 33600 800 33628
rect 49200 33600 50000 33628
rect 2818 33516 2828 33572
rect 2884 33516 3276 33572
rect 3332 33516 3836 33572
rect 3892 33516 3902 33572
rect 4834 33516 4844 33572
rect 4900 33516 5180 33572
rect 5236 33516 5246 33572
rect 8866 33516 8876 33572
rect 8932 33516 9100 33572
rect 9156 33516 9166 33572
rect 12086 33516 12124 33572
rect 12180 33516 12190 33572
rect 13794 33516 13804 33572
rect 13860 33516 21756 33572
rect 21812 33516 22316 33572
rect 22372 33516 22382 33572
rect 3574 33404 3612 33460
rect 3668 33404 3678 33460
rect 4162 33404 4172 33460
rect 4228 33404 10108 33460
rect 10164 33404 10174 33460
rect 11106 33404 11116 33460
rect 11172 33404 12012 33460
rect 12068 33404 12078 33460
rect 12310 33404 12348 33460
rect 12404 33404 12414 33460
rect 15362 33404 15372 33460
rect 15428 33404 20188 33460
rect 20244 33404 20254 33460
rect 32946 33404 32956 33460
rect 33012 33404 33404 33460
rect 33460 33404 37772 33460
rect 37828 33404 37838 33460
rect 45266 33404 45276 33460
rect 45332 33404 46060 33460
rect 46116 33404 46126 33460
rect 2146 33292 2156 33348
rect 2212 33292 6636 33348
rect 6692 33292 6702 33348
rect 9874 33292 9884 33348
rect 9940 33292 18508 33348
rect 18564 33292 18574 33348
rect 23090 33292 23100 33348
rect 23156 33292 23884 33348
rect 23940 33292 23950 33348
rect 28578 33292 28588 33348
rect 28644 33292 31164 33348
rect 31220 33292 31230 33348
rect 33954 33292 33964 33348
rect 34020 33292 35196 33348
rect 35252 33292 35262 33348
rect 1362 33180 1372 33236
rect 1428 33180 6300 33236
rect 6356 33180 6366 33236
rect 8418 33180 8428 33236
rect 8484 33180 9548 33236
rect 9604 33180 10668 33236
rect 10724 33180 10734 33236
rect 11452 33180 12908 33236
rect 12964 33180 12974 33236
rect 13234 33180 13244 33236
rect 13300 33180 15372 33236
rect 15428 33180 15438 33236
rect 15586 33180 15596 33236
rect 15652 33180 15662 33236
rect 15810 33180 15820 33236
rect 15876 33180 16828 33236
rect 16884 33180 16894 33236
rect 24210 33180 24220 33236
rect 24276 33180 25452 33236
rect 25508 33180 25518 33236
rect 35522 33180 35532 33236
rect 35588 33180 35980 33236
rect 36036 33180 38780 33236
rect 38836 33180 38846 33236
rect 43474 33180 43484 33236
rect 43540 33180 49364 33236
rect 11452 33124 11508 33180
rect 15596 33124 15652 33180
rect 3826 33068 3836 33124
rect 3892 33068 4508 33124
rect 4564 33068 4574 33124
rect 5954 33068 5964 33124
rect 6020 33068 8764 33124
rect 8820 33068 8830 33124
rect 11442 33068 11452 33124
rect 11508 33068 11518 33124
rect 11666 33068 11676 33124
rect 11732 33068 15652 33124
rect 22950 33068 22988 33124
rect 23044 33068 23054 33124
rect 23762 33068 23772 33124
rect 23828 33068 24444 33124
rect 24500 33068 25340 33124
rect 25396 33068 25406 33124
rect 28578 33068 28588 33124
rect 28644 33068 29372 33124
rect 29428 33068 37212 33124
rect 37268 33068 37278 33124
rect 38098 33068 38108 33124
rect 38164 33068 40460 33124
rect 40516 33068 40526 33124
rect 0 33012 800 33040
rect 0 32956 4844 33012
rect 4900 32956 4910 33012
rect 8838 32956 8876 33012
rect 8932 32956 8942 33012
rect 12114 32956 12124 33012
rect 12180 32956 12348 33012
rect 12404 32956 12414 33012
rect 13794 32956 13804 33012
rect 13860 32956 16044 33012
rect 16100 32956 16110 33012
rect 0 32928 800 32956
rect 19826 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20110 32956
rect 2258 32844 2268 32900
rect 2324 32844 9324 32900
rect 9380 32844 10332 32900
rect 10388 32844 10398 32900
rect 3042 32732 3052 32788
rect 3108 32732 3612 32788
rect 3668 32732 3678 32788
rect 4498 32732 4508 32788
rect 4564 32732 4844 32788
rect 4900 32732 5068 32788
rect 5124 32732 5134 32788
rect 15362 32732 15372 32788
rect 15428 32732 15708 32788
rect 15764 32732 16268 32788
rect 16324 32732 16828 32788
rect 16884 32732 16894 32788
rect 18918 32732 18956 32788
rect 19012 32732 19022 32788
rect 2930 32620 2940 32676
rect 2996 32620 3948 32676
rect 4004 32620 4014 32676
rect 9538 32620 9548 32676
rect 9604 32620 12796 32676
rect 12852 32620 15036 32676
rect 15092 32620 15102 32676
rect 15922 32620 15932 32676
rect 15988 32620 16940 32676
rect 16996 32620 19516 32676
rect 19572 32620 19582 32676
rect 21970 32620 21980 32676
rect 22036 32620 22316 32676
rect 22372 32620 22382 32676
rect 23874 32620 23884 32676
rect 23940 32620 24668 32676
rect 24724 32620 24734 32676
rect 32274 32620 32284 32676
rect 32340 32620 33964 32676
rect 34020 32620 34030 32676
rect 35746 32620 35756 32676
rect 35812 32620 41580 32676
rect 41636 32620 43708 32676
rect 43764 32620 43774 32676
rect 3332 32508 3388 32620
rect 22316 32564 22372 32620
rect 49308 32564 49364 33180
rect 3444 32508 3454 32564
rect 5394 32508 5404 32564
rect 5460 32508 6300 32564
rect 6356 32508 6366 32564
rect 7858 32508 7868 32564
rect 7924 32508 8316 32564
rect 8372 32508 9996 32564
rect 10052 32508 11788 32564
rect 11844 32508 11854 32564
rect 12450 32508 12460 32564
rect 12516 32508 15484 32564
rect 15540 32508 15550 32564
rect 22082 32508 22092 32564
rect 22148 32508 22158 32564
rect 22316 32508 23436 32564
rect 23492 32508 23502 32564
rect 40114 32508 40124 32564
rect 40180 32508 45612 32564
rect 45668 32508 45678 32564
rect 49084 32508 49364 32564
rect 22092 32452 22148 32508
rect 2258 32396 2268 32452
rect 2324 32396 5628 32452
rect 5684 32396 5694 32452
rect 6626 32396 6636 32452
rect 6692 32396 7308 32452
rect 7364 32396 8988 32452
rect 9044 32396 9156 32452
rect 9650 32396 9660 32452
rect 9716 32396 12012 32452
rect 12068 32396 12236 32452
rect 12292 32396 12302 32452
rect 15138 32396 15148 32452
rect 15204 32396 17164 32452
rect 17220 32396 17230 32452
rect 20178 32396 20188 32452
rect 20244 32396 20972 32452
rect 21028 32396 21038 32452
rect 22092 32396 23324 32452
rect 23380 32396 26236 32452
rect 26292 32396 26302 32452
rect 0 32340 800 32368
rect 6636 32340 6692 32396
rect 0 32284 1484 32340
rect 1540 32284 1550 32340
rect 4274 32284 4284 32340
rect 4340 32284 5180 32340
rect 5236 32284 6692 32340
rect 9100 32340 9156 32396
rect 49084 32340 49140 32508
rect 49200 32340 50000 32368
rect 9100 32284 11452 32340
rect 11508 32284 13916 32340
rect 13972 32284 13982 32340
rect 14690 32284 14700 32340
rect 14756 32284 17388 32340
rect 17444 32284 17454 32340
rect 22950 32284 22988 32340
rect 23044 32284 23054 32340
rect 41906 32284 41916 32340
rect 41972 32284 48188 32340
rect 48244 32284 48254 32340
rect 49084 32284 50000 32340
rect 0 32256 800 32284
rect 49200 32256 50000 32284
rect 8754 32172 8764 32228
rect 8820 32172 9772 32228
rect 9828 32172 9838 32228
rect 18834 32172 18844 32228
rect 18900 32172 21196 32228
rect 21252 32172 23660 32228
rect 23716 32172 24556 32228
rect 24612 32172 24622 32228
rect 4466 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4750 32172
rect 35186 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35470 32172
rect 6738 32060 6748 32116
rect 6804 32060 11116 32116
rect 11172 32060 11182 32116
rect 15026 32060 15036 32116
rect 15092 32060 16156 32116
rect 16212 32060 16222 32116
rect 17462 32060 17500 32116
rect 17556 32060 17566 32116
rect 39330 32060 39340 32116
rect 39396 32060 41020 32116
rect 41076 32060 41086 32116
rect 4498 31948 4508 32004
rect 4564 31948 5740 32004
rect 5796 31948 5806 32004
rect 7522 31948 7532 32004
rect 7588 31948 9100 32004
rect 9156 31948 9166 32004
rect 9650 31948 9660 32004
rect 9716 31948 10668 32004
rect 10724 31948 10734 32004
rect 11330 31948 11340 32004
rect 11396 31948 13580 32004
rect 13636 31948 13646 32004
rect 19282 31948 19292 32004
rect 19348 31948 19852 32004
rect 19908 31948 19918 32004
rect 39666 31948 39676 32004
rect 39732 31948 40180 32004
rect 40124 31892 40180 31948
rect 47012 31948 47180 32004
rect 47236 31948 47246 32004
rect 4162 31836 4172 31892
rect 4228 31836 5068 31892
rect 5124 31836 5134 31892
rect 6626 31836 6636 31892
rect 6692 31836 15148 31892
rect 21382 31836 21420 31892
rect 21476 31836 21486 31892
rect 21746 31836 21756 31892
rect 21812 31836 22428 31892
rect 22484 31836 22764 31892
rect 22820 31836 23100 31892
rect 23156 31836 23996 31892
rect 24052 31836 24062 31892
rect 24210 31836 24220 31892
rect 24276 31836 24892 31892
rect 24948 31836 24958 31892
rect 26562 31836 26572 31892
rect 26628 31836 27916 31892
rect 27972 31836 27982 31892
rect 31042 31836 31052 31892
rect 31108 31836 32060 31892
rect 32116 31836 32126 31892
rect 38658 31836 38668 31892
rect 38724 31836 39788 31892
rect 39844 31836 39854 31892
rect 40124 31836 41748 31892
rect 3154 31724 3164 31780
rect 3220 31724 4060 31780
rect 4116 31724 4126 31780
rect 5842 31724 5852 31780
rect 5908 31724 6972 31780
rect 7028 31724 7038 31780
rect 7970 31724 7980 31780
rect 8036 31724 8204 31780
rect 8260 31724 8270 31780
rect 8754 31724 8764 31780
rect 8820 31724 11004 31780
rect 11060 31724 11070 31780
rect 11554 31724 11564 31780
rect 11620 31724 12124 31780
rect 12180 31724 12190 31780
rect 0 31668 800 31696
rect 15092 31668 15148 31836
rect 41692 31780 41748 31836
rect 20290 31724 20300 31780
rect 20356 31724 25788 31780
rect 25844 31724 25854 31780
rect 28578 31724 28588 31780
rect 28644 31724 29148 31780
rect 29204 31724 32396 31780
rect 32452 31724 32462 31780
rect 41682 31724 41692 31780
rect 41748 31724 43148 31780
rect 43204 31724 43214 31780
rect 43810 31724 43820 31780
rect 43876 31724 45836 31780
rect 45892 31724 45902 31780
rect 47012 31668 47068 31948
rect 49200 31668 50000 31696
rect 0 31612 1820 31668
rect 1876 31612 1886 31668
rect 3266 31612 3276 31668
rect 0 31584 800 31612
rect 3332 31220 3388 31668
rect 3444 31612 3454 31668
rect 5506 31612 5516 31668
rect 5572 31612 7532 31668
rect 7588 31612 7598 31668
rect 8530 31612 8540 31668
rect 8596 31612 10108 31668
rect 10164 31612 10174 31668
rect 10742 31612 10780 31668
rect 10836 31612 10846 31668
rect 11442 31612 11452 31668
rect 11508 31612 12572 31668
rect 12628 31612 12796 31668
rect 12852 31612 12862 31668
rect 15092 31612 15484 31668
rect 15540 31612 15550 31668
rect 18610 31612 18620 31668
rect 18676 31612 22764 31668
rect 22820 31612 22830 31668
rect 34626 31612 34636 31668
rect 34692 31612 35308 31668
rect 35364 31612 42588 31668
rect 42644 31612 42654 31668
rect 47012 31612 50000 31668
rect 4050 31500 4060 31556
rect 4116 31500 6412 31556
rect 6468 31500 6478 31556
rect 6636 31332 6692 31612
rect 49200 31584 50000 31612
rect 10658 31500 10668 31556
rect 10724 31500 13020 31556
rect 13076 31500 15148 31556
rect 16146 31500 16156 31556
rect 16212 31500 19516 31556
rect 19572 31500 19582 31556
rect 23986 31500 23996 31556
rect 24052 31500 24556 31556
rect 24612 31500 26908 31556
rect 8754 31388 8764 31444
rect 8820 31388 9324 31444
rect 9380 31388 9390 31444
rect 9762 31388 9772 31444
rect 9828 31388 11116 31444
rect 11172 31388 11182 31444
rect 6626 31276 6636 31332
rect 6692 31276 6702 31332
rect 7644 31276 13244 31332
rect 13300 31276 13310 31332
rect 7644 31220 7700 31276
rect 15092 31220 15148 31500
rect 19826 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20110 31388
rect 3332 31164 7700 31220
rect 8726 31164 8764 31220
rect 8820 31164 8830 31220
rect 9538 31164 9548 31220
rect 9604 31164 14028 31220
rect 14084 31164 14094 31220
rect 15092 31164 20524 31220
rect 20580 31164 20590 31220
rect 26852 31108 26908 31500
rect 29586 31164 29596 31220
rect 29652 31164 30716 31220
rect 30772 31164 30782 31220
rect 38434 31164 38444 31220
rect 38500 31164 41132 31220
rect 41188 31164 41198 31220
rect 3332 31052 4844 31108
rect 4900 31052 9436 31108
rect 9492 31052 9502 31108
rect 9734 31052 9772 31108
rect 9828 31052 9838 31108
rect 18946 31052 18956 31108
rect 19012 31052 21308 31108
rect 21364 31052 21374 31108
rect 26852 31052 31388 31108
rect 31444 31052 34860 31108
rect 34916 31052 34926 31108
rect 0 30996 800 31024
rect 3332 30996 3388 31052
rect 49200 30996 50000 31024
rect 0 30940 1708 30996
rect 1764 30940 1774 30996
rect 2370 30940 2380 30996
rect 2436 30940 3388 30996
rect 3714 30940 3724 30996
rect 3780 30940 4956 30996
rect 5012 30940 5022 30996
rect 6514 30940 6524 30996
rect 6580 30940 8988 30996
rect 9044 30940 9548 30996
rect 9604 30940 9614 30996
rect 10098 30940 10108 30996
rect 10164 30940 11564 30996
rect 11620 30940 13356 30996
rect 13412 30940 13422 30996
rect 17826 30940 17836 30996
rect 17892 30940 20524 30996
rect 20580 30940 20590 30996
rect 24994 30940 25004 30996
rect 25060 30940 25340 30996
rect 25396 30940 25406 30996
rect 45266 30940 45276 30996
rect 45332 30940 50000 30996
rect 0 30912 800 30940
rect 49200 30912 50000 30940
rect 3938 30828 3948 30884
rect 4004 30828 5404 30884
rect 5460 30828 5470 30884
rect 6178 30828 6188 30884
rect 6244 30828 7084 30884
rect 7140 30828 7150 30884
rect 8194 30828 8204 30884
rect 8260 30828 14476 30884
rect 14532 30828 14542 30884
rect 19478 30828 19516 30884
rect 19572 30828 19582 30884
rect 19730 30828 19740 30884
rect 19796 30828 21532 30884
rect 21588 30828 22652 30884
rect 22708 30828 22876 30884
rect 22932 30828 22942 30884
rect 24770 30828 24780 30884
rect 24836 30828 26012 30884
rect 26068 30828 26078 30884
rect 37986 30828 37996 30884
rect 38052 30828 38780 30884
rect 38836 30828 38846 30884
rect 42802 30828 42812 30884
rect 42868 30828 43820 30884
rect 43876 30828 43886 30884
rect 6402 30716 6412 30772
rect 6468 30716 6972 30772
rect 7028 30716 7038 30772
rect 7746 30716 7756 30772
rect 7812 30716 9660 30772
rect 9716 30716 9726 30772
rect 13682 30716 13692 30772
rect 13748 30716 15372 30772
rect 15428 30716 15438 30772
rect 11106 30604 11116 30660
rect 11172 30604 12348 30660
rect 12404 30604 15708 30660
rect 15764 30604 15774 30660
rect 22194 30604 22204 30660
rect 22260 30604 23772 30660
rect 23828 30604 23838 30660
rect 4466 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4750 30604
rect 35186 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35470 30604
rect 10546 30492 10556 30548
rect 10612 30492 10780 30548
rect 10836 30492 10846 30548
rect 12450 30492 12460 30548
rect 12516 30492 15036 30548
rect 15092 30492 15102 30548
rect 20738 30492 20748 30548
rect 20804 30492 21308 30548
rect 21364 30492 21374 30548
rect 24098 30492 24108 30548
rect 24164 30492 26908 30548
rect 26964 30492 28140 30548
rect 28196 30492 28206 30548
rect 4274 30380 4284 30436
rect 4340 30380 5068 30436
rect 5124 30380 6300 30436
rect 6356 30380 6366 30436
rect 10658 30380 10668 30436
rect 10724 30380 11228 30436
rect 11284 30380 11294 30436
rect 12562 30380 12572 30436
rect 12628 30380 13580 30436
rect 13636 30380 13646 30436
rect 14242 30380 14252 30436
rect 14308 30380 19908 30436
rect 20290 30380 20300 30436
rect 20356 30380 23996 30436
rect 24052 30380 24062 30436
rect 0 30324 800 30352
rect 0 30268 1820 30324
rect 1876 30268 1886 30324
rect 4946 30268 4956 30324
rect 5012 30268 8204 30324
rect 8260 30268 8270 30324
rect 0 30240 800 30268
rect 11228 30212 11284 30380
rect 19852 30324 19908 30380
rect 49200 30324 50000 30352
rect 12898 30268 12908 30324
rect 12964 30268 14476 30324
rect 14532 30268 14542 30324
rect 14690 30268 14700 30324
rect 14756 30268 15036 30324
rect 15092 30268 15260 30324
rect 15316 30268 15326 30324
rect 18498 30268 18508 30324
rect 18564 30268 18956 30324
rect 19012 30268 19022 30324
rect 19170 30268 19180 30324
rect 19236 30268 19628 30324
rect 19684 30268 19694 30324
rect 19852 30268 20692 30324
rect 21746 30268 21756 30324
rect 21812 30268 24444 30324
rect 24500 30268 24510 30324
rect 25330 30268 25340 30324
rect 25396 30268 26908 30324
rect 46274 30268 46284 30324
rect 46340 30268 50000 30324
rect 1698 30156 1708 30212
rect 1764 30156 4172 30212
rect 4228 30156 4238 30212
rect 7858 30156 7868 30212
rect 7924 30156 8428 30212
rect 8484 30156 8494 30212
rect 10854 30156 10892 30212
rect 10948 30156 10958 30212
rect 11228 30156 14028 30212
rect 14084 30156 14094 30212
rect 14578 30156 14588 30212
rect 14644 30156 16268 30212
rect 16324 30156 16334 30212
rect 16594 30156 16604 30212
rect 16660 30156 17164 30212
rect 17220 30156 18060 30212
rect 18116 30156 18126 30212
rect 19394 30156 19404 30212
rect 19460 30156 19964 30212
rect 20020 30156 20030 30212
rect 20636 30100 20692 30268
rect 26852 30212 26908 30268
rect 49200 30240 50000 30268
rect 21970 30156 21980 30212
rect 22036 30156 22540 30212
rect 22596 30156 24556 30212
rect 24612 30156 24622 30212
rect 26852 30156 28588 30212
rect 28644 30156 28654 30212
rect 37202 30156 37212 30212
rect 37268 30156 38220 30212
rect 38276 30156 40684 30212
rect 40740 30156 40750 30212
rect 42690 30156 42700 30212
rect 42756 30156 45388 30212
rect 45444 30156 45454 30212
rect 4274 30044 4284 30100
rect 4340 30044 18284 30100
rect 18340 30044 18350 30100
rect 20626 30044 20636 30100
rect 20692 30044 20702 30100
rect 21410 30044 21420 30100
rect 21476 30044 21644 30100
rect 21700 30044 21710 30100
rect 31826 30044 31836 30100
rect 10434 29932 10444 29988
rect 10500 29932 11788 29988
rect 12786 29932 12796 29988
rect 12852 29932 13916 29988
rect 13972 29932 13982 29988
rect 15362 29932 15372 29988
rect 15428 29932 18508 29988
rect 18564 29932 18574 29988
rect 18946 29932 18956 29988
rect 19012 29932 19180 29988
rect 19236 29932 19404 29988
rect 19460 29932 19470 29988
rect 19628 29932 20356 29988
rect 20514 29932 20524 29988
rect 20580 29932 22652 29988
rect 22708 29932 22718 29988
rect 26226 29932 26236 29988
rect 26292 29932 26908 29988
rect 26964 29932 26974 29988
rect 27122 29932 27132 29988
rect 27188 29932 29260 29988
rect 29316 29932 29596 29988
rect 29652 29932 29662 29988
rect 11732 29876 11788 29932
rect 19628 29876 19684 29932
rect 11732 29820 12572 29876
rect 12628 29820 12638 29876
rect 13794 29820 13804 29876
rect 13860 29820 14588 29876
rect 14644 29820 14654 29876
rect 15092 29820 17836 29876
rect 17892 29820 19684 29876
rect 20300 29876 20356 29932
rect 20300 29820 25452 29876
rect 25508 29820 25518 29876
rect 15092 29764 15148 29820
rect 19826 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20110 29820
rect 31892 29764 31948 30100
rect 33170 29932 33180 29988
rect 33236 29932 34524 29988
rect 34580 29932 34590 29988
rect 43474 29932 43484 29988
rect 43540 29932 44044 29988
rect 44100 29932 44940 29988
rect 44996 29932 47404 29988
rect 47460 29932 47470 29988
rect 6402 29708 6412 29764
rect 6468 29708 15148 29764
rect 16482 29708 16492 29764
rect 16548 29708 19460 29764
rect 31892 29708 34076 29764
rect 34132 29708 35644 29764
rect 35700 29708 46060 29764
rect 46116 29708 46126 29764
rect 0 29652 800 29680
rect 19404 29652 19460 29708
rect 49200 29652 50000 29680
rect 0 29596 2492 29652
rect 2548 29596 2558 29652
rect 3332 29596 4284 29652
rect 4340 29596 7644 29652
rect 7700 29596 9660 29652
rect 9716 29596 10556 29652
rect 10612 29596 10622 29652
rect 16370 29596 16380 29652
rect 16436 29596 17052 29652
rect 17108 29596 17118 29652
rect 18050 29596 18060 29652
rect 18116 29596 18396 29652
rect 18452 29596 18462 29652
rect 19394 29596 19404 29652
rect 19460 29596 20412 29652
rect 20468 29596 20478 29652
rect 47058 29596 47068 29652
rect 47124 29596 50000 29652
rect 0 29568 800 29596
rect 3332 29540 3388 29596
rect 18060 29540 18116 29596
rect 49200 29568 50000 29596
rect 2706 29484 2716 29540
rect 2772 29484 3388 29540
rect 8306 29484 8316 29540
rect 8372 29484 10668 29540
rect 10724 29484 11116 29540
rect 11172 29484 11182 29540
rect 12982 29484 13020 29540
rect 13076 29484 13086 29540
rect 15362 29484 15372 29540
rect 15428 29484 16044 29540
rect 16100 29484 17276 29540
rect 17332 29484 18116 29540
rect 25890 29484 25900 29540
rect 25956 29484 27020 29540
rect 27076 29484 27086 29540
rect 27682 29484 27692 29540
rect 27748 29484 31276 29540
rect 31332 29484 31342 29540
rect 31892 29484 37212 29540
rect 37268 29484 37278 29540
rect 2482 29372 2492 29428
rect 2548 29372 2828 29428
rect 2884 29372 2894 29428
rect 3154 29372 3164 29428
rect 3220 29372 6748 29428
rect 6804 29372 6814 29428
rect 8988 29372 15820 29428
rect 15876 29372 20188 29428
rect 20244 29372 21308 29428
rect 21364 29372 21374 29428
rect 21746 29372 21756 29428
rect 21812 29372 22092 29428
rect 22148 29372 22158 29428
rect 28578 29372 28588 29428
rect 28644 29372 29484 29428
rect 29540 29372 29550 29428
rect 2492 29204 2548 29372
rect 2706 29260 2716 29316
rect 2772 29260 4396 29316
rect 4452 29260 4462 29316
rect 4946 29260 4956 29316
rect 5012 29260 6972 29316
rect 7028 29260 7038 29316
rect 8988 29204 9044 29372
rect 11778 29260 11788 29316
rect 11844 29260 13804 29316
rect 13860 29260 13870 29316
rect 14018 29260 14028 29316
rect 14084 29260 16268 29316
rect 16324 29260 16334 29316
rect 16594 29260 16604 29316
rect 16660 29260 18956 29316
rect 19012 29260 20076 29316
rect 20132 29260 20142 29316
rect 21074 29260 21084 29316
rect 21140 29260 24108 29316
rect 24164 29260 24174 29316
rect 20076 29204 20132 29260
rect 1810 29148 1820 29204
rect 1876 29148 3388 29204
rect 3490 29148 3500 29204
rect 3556 29148 9044 29204
rect 9762 29148 9772 29204
rect 9828 29148 10332 29204
rect 10388 29148 10398 29204
rect 10546 29148 10556 29204
rect 10612 29148 16716 29204
rect 16772 29148 16782 29204
rect 20076 29148 22652 29204
rect 22708 29148 22718 29204
rect 0 28980 800 29008
rect 0 28924 3052 28980
rect 3108 28924 3118 28980
rect 0 28896 800 28924
rect 3332 28868 3388 29148
rect 31892 29092 31948 29484
rect 35970 29372 35980 29428
rect 36036 29372 37324 29428
rect 37380 29372 41020 29428
rect 41076 29372 42700 29428
rect 42756 29372 42766 29428
rect 33394 29260 33404 29316
rect 33460 29260 35196 29316
rect 35252 29260 35262 29316
rect 35410 29260 35420 29316
rect 35476 29260 39340 29316
rect 39396 29260 39406 29316
rect 33058 29148 33068 29204
rect 33124 29148 34860 29204
rect 34916 29148 34926 29204
rect 8418 29036 8428 29092
rect 8484 29036 10108 29092
rect 10164 29036 10174 29092
rect 10434 29036 10444 29092
rect 10500 29036 11004 29092
rect 11060 29036 11070 29092
rect 20626 29036 20636 29092
rect 20692 29036 21308 29092
rect 21364 29036 21374 29092
rect 29586 29036 29596 29092
rect 29652 29036 30044 29092
rect 30100 29036 31948 29092
rect 4466 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4750 29036
rect 35186 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35470 29036
rect 49200 28980 50000 29008
rect 4834 28924 4844 28980
rect 4900 28924 12684 28980
rect 12740 28924 12750 28980
rect 19730 28924 19740 28980
rect 19796 28924 20412 28980
rect 20468 28924 23884 28980
rect 23940 28924 32732 28980
rect 32788 28924 32798 28980
rect 38322 28924 38332 28980
rect 38388 28924 39116 28980
rect 39172 28924 39900 28980
rect 39956 28924 42364 28980
rect 42420 28924 43484 28980
rect 43540 28924 43550 28980
rect 47730 28924 47740 28980
rect 47796 28924 50000 28980
rect 4844 28868 4900 28924
rect 49200 28896 50000 28924
rect 3332 28812 4900 28868
rect 5170 28812 5180 28868
rect 5236 28812 5740 28868
rect 5796 28812 6860 28868
rect 6916 28812 6926 28868
rect 8754 28812 8764 28868
rect 8820 28812 9436 28868
rect 9492 28812 9502 28868
rect 12114 28812 12124 28868
rect 12180 28812 15596 28868
rect 15652 28812 15662 28868
rect 16930 28812 16940 28868
rect 16996 28812 20188 28868
rect 20244 28812 20254 28868
rect 29698 28812 29708 28868
rect 29764 28812 30716 28868
rect 30772 28812 30782 28868
rect 41458 28812 41468 28868
rect 41524 28812 43820 28868
rect 43876 28812 43886 28868
rect 45602 28812 45612 28868
rect 45668 28812 45678 28868
rect 45612 28756 45668 28812
rect 2594 28700 2604 28756
rect 2660 28700 4396 28756
rect 4452 28700 10444 28756
rect 10500 28700 10510 28756
rect 12898 28700 12908 28756
rect 12964 28700 13468 28756
rect 13524 28700 13534 28756
rect 13682 28700 13692 28756
rect 13748 28700 13786 28756
rect 14242 28700 14252 28756
rect 14308 28700 17724 28756
rect 17780 28700 17790 28756
rect 30258 28700 30268 28756
rect 30324 28700 31836 28756
rect 31892 28700 31902 28756
rect 40460 28700 45668 28756
rect 3154 28588 3164 28644
rect 3220 28588 3836 28644
rect 3892 28588 3902 28644
rect 4610 28588 4620 28644
rect 4676 28588 5628 28644
rect 5684 28588 5694 28644
rect 7186 28588 7196 28644
rect 7252 28588 8092 28644
rect 8148 28588 8158 28644
rect 8530 28588 8540 28644
rect 8596 28588 9772 28644
rect 9828 28588 9838 28644
rect 10770 28588 10780 28644
rect 10836 28588 10892 28644
rect 10948 28588 10958 28644
rect 11218 28588 11228 28644
rect 11284 28588 12236 28644
rect 12292 28588 12302 28644
rect 13010 28588 13020 28644
rect 13076 28588 14028 28644
rect 14084 28588 14094 28644
rect 17938 28588 17948 28644
rect 18004 28588 18172 28644
rect 18228 28588 18956 28644
rect 19012 28588 19022 28644
rect 22978 28588 22988 28644
rect 23044 28588 23436 28644
rect 23492 28588 23502 28644
rect 23650 28588 23660 28644
rect 23716 28588 26236 28644
rect 26292 28588 26572 28644
rect 26628 28588 26638 28644
rect 40460 28532 40516 28700
rect 40674 28588 40684 28644
rect 40740 28588 41916 28644
rect 41972 28588 41982 28644
rect 43362 28588 43372 28644
rect 43428 28588 44884 28644
rect 8390 28476 8428 28532
rect 8484 28476 8494 28532
rect 15250 28476 15260 28532
rect 15316 28476 16044 28532
rect 16100 28476 21196 28532
rect 21252 28476 21262 28532
rect 22754 28476 22764 28532
rect 22820 28476 23996 28532
rect 24052 28476 24062 28532
rect 25778 28476 25788 28532
rect 25844 28476 26908 28532
rect 26964 28476 26974 28532
rect 27458 28476 27468 28532
rect 27524 28476 32844 28532
rect 32900 28476 32910 28532
rect 36194 28476 36204 28532
rect 36260 28476 36540 28532
rect 36596 28476 40516 28532
rect 41570 28476 41580 28532
rect 41636 28476 42252 28532
rect 42308 28476 42318 28532
rect 44828 28420 44884 28588
rect 5842 28364 5852 28420
rect 5908 28364 6412 28420
rect 6468 28364 6478 28420
rect 13346 28364 13356 28420
rect 13412 28364 17948 28420
rect 18004 28364 18014 28420
rect 44818 28364 44828 28420
rect 44884 28364 44894 28420
rect 0 28308 800 28336
rect 49200 28308 50000 28336
rect 0 28252 1708 28308
rect 1764 28252 1774 28308
rect 2258 28252 2268 28308
rect 2324 28252 11788 28308
rect 11844 28252 11854 28308
rect 13906 28252 13916 28308
rect 13972 28252 14476 28308
rect 14532 28252 14542 28308
rect 43250 28252 43260 28308
rect 43316 28252 45500 28308
rect 45556 28252 45566 28308
rect 47954 28252 47964 28308
rect 48020 28252 50000 28308
rect 0 28224 800 28252
rect 19826 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20110 28252
rect 49200 28224 50000 28252
rect 3332 28140 16492 28196
rect 16548 28140 16558 28196
rect 3332 28084 3388 28140
rect 2258 28028 2268 28084
rect 2324 28028 3388 28084
rect 5730 28028 5740 28084
rect 5796 28028 6300 28084
rect 6356 28028 6366 28084
rect 11554 28028 11564 28084
rect 11620 28028 11788 28084
rect 11844 28028 12684 28084
rect 12740 28028 12750 28084
rect 15026 28028 15036 28084
rect 15092 28028 15820 28084
rect 15876 28028 15886 28084
rect 17266 28028 17276 28084
rect 17332 28028 17836 28084
rect 17892 28028 19180 28084
rect 19236 28028 19246 28084
rect 45154 28028 45164 28084
rect 45220 28028 47628 28084
rect 47684 28028 47694 28084
rect 47842 28028 47852 28084
rect 47908 28028 47918 28084
rect 1362 27916 1372 27972
rect 1428 27916 6972 27972
rect 7028 27916 7038 27972
rect 8194 27916 8204 27972
rect 8260 27916 15036 27972
rect 15092 27916 15102 27972
rect 17714 27916 17724 27972
rect 17780 27916 22204 27972
rect 22260 27916 22270 27972
rect 23090 27916 23100 27972
rect 23156 27916 25788 27972
rect 25844 27916 25854 27972
rect 43922 27916 43932 27972
rect 43988 27916 46620 27972
rect 46676 27916 46686 27972
rect 47852 27860 47908 28028
rect 7186 27804 7196 27860
rect 7252 27804 10108 27860
rect 10164 27804 10332 27860
rect 10388 27804 10780 27860
rect 10836 27804 10846 27860
rect 12450 27804 12460 27860
rect 12516 27804 15260 27860
rect 15316 27804 15326 27860
rect 16818 27804 16828 27860
rect 16884 27804 18396 27860
rect 18452 27804 18462 27860
rect 21298 27804 21308 27860
rect 21364 27804 23436 27860
rect 23492 27804 23502 27860
rect 26674 27804 26684 27860
rect 26740 27804 27356 27860
rect 27412 27804 27422 27860
rect 47852 27804 48132 27860
rect 2482 27692 2492 27748
rect 2548 27692 5068 27748
rect 5124 27692 5134 27748
rect 7858 27692 7868 27748
rect 7924 27692 9772 27748
rect 9828 27692 9838 27748
rect 11218 27692 11228 27748
rect 11284 27692 11900 27748
rect 11956 27692 11966 27748
rect 14242 27692 14252 27748
rect 14308 27692 16044 27748
rect 16100 27692 16110 27748
rect 39666 27692 39676 27748
rect 39732 27692 40348 27748
rect 40404 27692 40414 27748
rect 0 27636 800 27664
rect 48076 27636 48132 27804
rect 49200 27636 50000 27664
rect 0 27580 3388 27636
rect 3444 27580 3454 27636
rect 3714 27580 3724 27636
rect 3780 27580 8820 27636
rect 8978 27580 8988 27636
rect 9044 27580 9548 27636
rect 9604 27580 9996 27636
rect 10052 27580 12908 27636
rect 12964 27580 16156 27636
rect 16212 27580 16222 27636
rect 48076 27580 50000 27636
rect 0 27552 800 27580
rect 8764 27524 8820 27580
rect 49200 27552 50000 27580
rect 8764 27468 10108 27524
rect 10164 27468 12012 27524
rect 12068 27468 12078 27524
rect 12562 27468 12572 27524
rect 12628 27468 13244 27524
rect 13300 27468 14812 27524
rect 14868 27468 14878 27524
rect 15026 27468 15036 27524
rect 15092 27468 16716 27524
rect 16772 27468 18060 27524
rect 18116 27468 18126 27524
rect 4466 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4750 27468
rect 11732 27412 11788 27468
rect 35186 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35470 27468
rect 6402 27356 6412 27412
rect 6468 27356 6860 27412
rect 6916 27356 6926 27412
rect 10658 27356 10668 27412
rect 10724 27356 11340 27412
rect 11396 27356 11406 27412
rect 11732 27356 15036 27412
rect 15092 27356 15102 27412
rect 4050 27244 4060 27300
rect 4116 27244 5964 27300
rect 6020 27244 6030 27300
rect 6514 27244 6524 27300
rect 6580 27244 8988 27300
rect 9044 27244 11900 27300
rect 11956 27244 11966 27300
rect 12226 27244 12236 27300
rect 12292 27244 14924 27300
rect 14980 27244 15148 27300
rect 21186 27244 21196 27300
rect 21252 27244 23996 27300
rect 24052 27244 24062 27300
rect 32386 27244 32396 27300
rect 32452 27244 45612 27300
rect 45668 27244 45678 27300
rect 3154 27132 3164 27188
rect 3220 27132 4956 27188
rect 5012 27132 5022 27188
rect 6748 27132 8764 27188
rect 8820 27132 9100 27188
rect 9156 27132 11116 27188
rect 11172 27132 11564 27188
rect 11620 27132 11630 27188
rect 11778 27132 11788 27188
rect 11844 27132 13356 27188
rect 13412 27132 13422 27188
rect 6748 27076 6804 27132
rect 15092 27076 15148 27244
rect 15698 27132 15708 27188
rect 15764 27132 20580 27188
rect 20738 27132 20748 27188
rect 20804 27132 22764 27188
rect 22820 27132 22830 27188
rect 26450 27132 26460 27188
rect 26516 27132 27132 27188
rect 27188 27132 27198 27188
rect 45266 27132 45276 27188
rect 45332 27132 46060 27188
rect 46116 27132 46126 27188
rect 20524 27076 20580 27132
rect 4732 27020 6804 27076
rect 6962 27020 6972 27076
rect 7028 27020 7196 27076
rect 7252 27020 7262 27076
rect 8082 27020 8092 27076
rect 8148 27020 8652 27076
rect 8708 27020 9324 27076
rect 9380 27020 9390 27076
rect 10770 27020 10780 27076
rect 10836 27020 11900 27076
rect 11956 27020 11966 27076
rect 15092 27020 15372 27076
rect 15428 27020 15438 27076
rect 15810 27020 15820 27076
rect 15876 27020 15886 27076
rect 20524 27020 22092 27076
rect 22148 27020 22158 27076
rect 22978 27020 22988 27076
rect 23044 27020 24444 27076
rect 24500 27020 31612 27076
rect 31668 27020 35868 27076
rect 35924 27020 37772 27076
rect 37828 27020 37838 27076
rect 0 26964 800 26992
rect 4732 26964 4788 27020
rect 15820 26964 15876 27020
rect 0 26908 2436 26964
rect 4722 26908 4732 26964
rect 4788 26908 4798 26964
rect 5740 26908 6524 26964
rect 6580 26908 6590 26964
rect 6962 26908 6972 26964
rect 7028 26908 7038 26964
rect 10546 26908 10556 26964
rect 10612 26908 12348 26964
rect 12404 26908 12414 26964
rect 13906 26908 13916 26964
rect 13972 26908 15876 26964
rect 16034 26908 16044 26964
rect 16100 26908 17388 26964
rect 17444 26908 17836 26964
rect 17892 26908 17902 26964
rect 23538 26908 23548 26964
rect 23604 26908 24556 26964
rect 24612 26908 24622 26964
rect 38322 26908 38332 26964
rect 38388 26908 39676 26964
rect 39732 26908 39742 26964
rect 0 26880 800 26908
rect 2380 26852 2436 26908
rect 5740 26852 5796 26908
rect 6972 26852 7028 26908
rect 2370 26796 2380 26852
rect 2436 26796 2446 26852
rect 2706 26796 2716 26852
rect 2772 26796 3612 26852
rect 3668 26796 3678 26852
rect 5618 26796 5628 26852
rect 5684 26796 5796 26852
rect 5964 26796 8316 26852
rect 8372 26796 8382 26852
rect 10322 26796 10332 26852
rect 10388 26796 10668 26852
rect 10724 26796 10734 26852
rect 11302 26796 11340 26852
rect 11396 26796 11406 26852
rect 11554 26796 11564 26852
rect 11620 26796 12124 26852
rect 12180 26796 12190 26852
rect 12348 26796 21308 26852
rect 21364 26796 21374 26852
rect 43362 26796 43372 26852
rect 43428 26796 44268 26852
rect 44324 26796 44334 26852
rect 5964 26740 6020 26796
rect 12348 26740 12404 26796
rect 2482 26684 2492 26740
rect 2548 26684 4620 26740
rect 4676 26684 4686 26740
rect 5170 26684 5180 26740
rect 5236 26684 5740 26740
rect 5796 26684 5806 26740
rect 5954 26684 5964 26740
rect 6020 26684 6030 26740
rect 6626 26684 6636 26740
rect 6692 26684 12404 26740
rect 13794 26684 13804 26740
rect 13860 26684 14588 26740
rect 14644 26684 14654 26740
rect 14802 26684 14812 26740
rect 14868 26684 15708 26740
rect 15764 26684 15774 26740
rect 16482 26684 16492 26740
rect 16548 26684 17164 26740
rect 17220 26684 17230 26740
rect 19826 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20110 26684
rect 2146 26572 2156 26628
rect 2212 26572 3500 26628
rect 3556 26572 4844 26628
rect 4900 26572 4910 26628
rect 5058 26572 5068 26628
rect 5124 26572 6748 26628
rect 6804 26572 6814 26628
rect 15362 26572 15372 26628
rect 15428 26572 16884 26628
rect 16828 26516 16884 26572
rect 2930 26460 2940 26516
rect 2996 26460 4396 26516
rect 4452 26460 5516 26516
rect 5572 26460 6636 26516
rect 6692 26460 6702 26516
rect 8978 26460 8988 26516
rect 9044 26460 10892 26516
rect 10948 26460 11452 26516
rect 11508 26460 11518 26516
rect 14018 26460 14028 26516
rect 14084 26460 16492 26516
rect 16548 26460 16558 26516
rect 16828 26460 21196 26516
rect 21252 26460 21262 26516
rect 38210 26460 38220 26516
rect 38276 26460 39676 26516
rect 39732 26460 39742 26516
rect 5058 26348 5068 26404
rect 5124 26348 11676 26404
rect 11732 26348 11742 26404
rect 12450 26348 12460 26404
rect 12516 26348 18284 26404
rect 18340 26348 18350 26404
rect 24434 26348 24444 26404
rect 24500 26348 26908 26404
rect 27794 26348 27804 26404
rect 27860 26348 28588 26404
rect 28644 26348 29484 26404
rect 29540 26348 29550 26404
rect 0 26292 800 26320
rect 26852 26292 26908 26348
rect 0 26236 1708 26292
rect 1764 26236 1774 26292
rect 6738 26236 6748 26292
rect 6804 26236 7196 26292
rect 7252 26236 7262 26292
rect 8082 26236 8092 26292
rect 8148 26236 8158 26292
rect 9986 26236 9996 26292
rect 10052 26236 16156 26292
rect 16212 26236 16222 26292
rect 16706 26236 16716 26292
rect 16772 26236 23772 26292
rect 23828 26236 23838 26292
rect 26852 26236 27468 26292
rect 27524 26236 27534 26292
rect 39218 26236 39228 26292
rect 39284 26236 44716 26292
rect 44772 26236 45388 26292
rect 45444 26236 45454 26292
rect 0 26208 800 26236
rect 8092 26180 8148 26236
rect 2930 26124 2940 26180
rect 2996 26124 5404 26180
rect 5460 26124 5470 26180
rect 7634 26124 7644 26180
rect 7700 26124 8036 26180
rect 8092 26124 10108 26180
rect 10164 26124 10174 26180
rect 11330 26124 11340 26180
rect 11396 26124 11900 26180
rect 11956 26124 11966 26180
rect 13682 26124 13692 26180
rect 13748 26124 15596 26180
rect 15652 26124 15662 26180
rect 18498 26124 18508 26180
rect 18564 26124 18844 26180
rect 18900 26124 18910 26180
rect 20178 26124 20188 26180
rect 20244 26124 22092 26180
rect 22148 26124 22158 26180
rect 36306 26124 36316 26180
rect 36372 26124 37548 26180
rect 37604 26124 37614 26180
rect 40114 26124 40124 26180
rect 40180 26124 40908 26180
rect 40964 26124 41916 26180
rect 41972 26124 43260 26180
rect 43316 26124 43326 26180
rect 7980 26068 8036 26124
rect 6290 26012 6300 26068
rect 6356 26012 6860 26068
rect 6916 26012 7756 26068
rect 7812 26012 7822 26068
rect 7980 26012 17276 26068
rect 17332 26012 17342 26068
rect 18386 26012 18396 26068
rect 18452 26012 27020 26068
rect 27076 26012 27086 26068
rect 7858 25900 7868 25956
rect 7924 25900 9884 25956
rect 9940 25900 13468 25956
rect 13524 25900 13534 25956
rect 22754 25900 22764 25956
rect 22820 25900 23212 25956
rect 23268 25900 23278 25956
rect 37314 25900 37324 25956
rect 37380 25900 45612 25956
rect 45668 25900 45678 25956
rect 4466 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4750 25900
rect 35186 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35470 25900
rect 1698 25788 1708 25844
rect 1764 25788 3052 25844
rect 3108 25788 3118 25844
rect 3826 25788 3836 25844
rect 3892 25788 3902 25844
rect 8194 25788 8204 25844
rect 8260 25788 8652 25844
rect 8708 25788 9548 25844
rect 9604 25788 9614 25844
rect 10098 25788 10108 25844
rect 10164 25788 14700 25844
rect 14756 25788 14766 25844
rect 19842 25788 19852 25844
rect 19908 25788 20412 25844
rect 20468 25788 20478 25844
rect 21410 25788 21420 25844
rect 21476 25788 22876 25844
rect 22932 25788 22942 25844
rect 3836 25732 3892 25788
rect 3836 25676 15148 25732
rect 18162 25676 18172 25732
rect 18228 25676 23772 25732
rect 23828 25676 23838 25732
rect 38322 25676 38332 25732
rect 38388 25676 39116 25732
rect 39172 25676 39788 25732
rect 39844 25676 39854 25732
rect 40338 25676 40348 25732
rect 40404 25676 41748 25732
rect 0 25620 800 25648
rect 0 25564 1708 25620
rect 1764 25564 2716 25620
rect 2772 25564 2782 25620
rect 4610 25564 4620 25620
rect 4676 25564 6972 25620
rect 7028 25564 7038 25620
rect 9314 25564 9324 25620
rect 9380 25564 13580 25620
rect 13636 25564 13646 25620
rect 0 25536 800 25564
rect 15092 25508 15148 25676
rect 15250 25564 15260 25620
rect 15316 25564 16380 25620
rect 16436 25564 16446 25620
rect 18050 25564 18060 25620
rect 18116 25564 18126 25620
rect 19282 25564 19292 25620
rect 19348 25564 22316 25620
rect 22372 25564 22382 25620
rect 24546 25564 24556 25620
rect 24612 25564 26124 25620
rect 26180 25564 26190 25620
rect 30370 25564 30380 25620
rect 30436 25564 32172 25620
rect 32228 25564 32238 25620
rect 38770 25564 38780 25620
rect 38836 25564 40572 25620
rect 40628 25564 40638 25620
rect 18060 25508 18116 25564
rect 41692 25508 41748 25676
rect 49200 25620 50000 25648
rect 43362 25564 43372 25620
rect 43428 25564 44044 25620
rect 44100 25564 44110 25620
rect 47954 25564 47964 25620
rect 48020 25564 50000 25620
rect 49200 25536 50000 25564
rect 6738 25452 6748 25508
rect 6804 25452 8092 25508
rect 8148 25452 8158 25508
rect 10406 25452 10444 25508
rect 10500 25452 10510 25508
rect 12674 25452 12684 25508
rect 12740 25452 13356 25508
rect 13412 25452 13422 25508
rect 15092 25452 15708 25508
rect 15764 25452 16716 25508
rect 16772 25452 16782 25508
rect 17266 25452 17276 25508
rect 17332 25452 17836 25508
rect 17892 25452 17902 25508
rect 18060 25452 18396 25508
rect 18452 25452 18462 25508
rect 19842 25452 19852 25508
rect 19908 25452 21420 25508
rect 21476 25452 21486 25508
rect 29362 25452 29372 25508
rect 29428 25452 33068 25508
rect 33124 25452 33134 25508
rect 39554 25452 39564 25508
rect 39620 25452 40460 25508
rect 40516 25452 41244 25508
rect 41300 25452 41310 25508
rect 41682 25452 41692 25508
rect 41748 25452 42364 25508
rect 42420 25452 42430 25508
rect 11330 25340 11340 25396
rect 11396 25340 12460 25396
rect 12516 25340 12526 25396
rect 15782 25340 15820 25396
rect 15876 25340 15886 25396
rect 16930 25340 16940 25396
rect 16996 25340 17500 25396
rect 17556 25340 18284 25396
rect 18340 25340 18732 25396
rect 18788 25340 18798 25396
rect 20178 25340 20188 25396
rect 20244 25340 20412 25396
rect 20468 25340 20478 25396
rect 37538 25340 37548 25396
rect 37604 25340 38780 25396
rect 38836 25340 38846 25396
rect 40562 25340 40572 25396
rect 40628 25340 43036 25396
rect 43092 25340 43102 25396
rect 44594 25340 44604 25396
rect 44660 25340 46060 25396
rect 46116 25340 46126 25396
rect 2482 25228 2492 25284
rect 2548 25228 3276 25284
rect 3332 25228 3342 25284
rect 12674 25228 12684 25284
rect 12740 25228 14476 25284
rect 14532 25228 14542 25284
rect 16678 25228 16716 25284
rect 16772 25228 16782 25284
rect 17042 25228 17052 25284
rect 17108 25228 17836 25284
rect 17892 25228 20300 25284
rect 20356 25228 22428 25284
rect 22484 25228 23212 25284
rect 23268 25228 23278 25284
rect 39330 25228 39340 25284
rect 39396 25228 39788 25284
rect 39844 25228 40796 25284
rect 40852 25228 40862 25284
rect 43138 25228 43148 25284
rect 43204 25228 43484 25284
rect 43540 25228 43550 25284
rect 2930 25116 2940 25172
rect 2996 25116 3388 25172
rect 5170 25116 5180 25172
rect 5236 25116 6972 25172
rect 7028 25116 9996 25172
rect 10052 25116 10668 25172
rect 10724 25116 10734 25172
rect 11078 25116 11116 25172
rect 11172 25116 11182 25172
rect 11414 25116 11452 25172
rect 11508 25116 11518 25172
rect 17602 25116 17612 25172
rect 17668 25116 18844 25172
rect 18900 25116 19404 25172
rect 19460 25116 19470 25172
rect 0 24948 800 24976
rect 3332 24948 3388 25116
rect 19826 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20110 25116
rect 11666 25004 11676 25060
rect 11732 25004 17276 25060
rect 17332 25004 17342 25060
rect 18274 25004 18284 25060
rect 18340 25004 18378 25060
rect 43698 25004 43708 25060
rect 43764 25004 45276 25060
rect 45332 25004 47404 25060
rect 47460 25004 47470 25060
rect 49200 24948 50000 24976
rect 0 24892 2436 24948
rect 3332 24892 13692 24948
rect 13748 24892 13758 24948
rect 16716 24892 17500 24948
rect 17556 24892 17566 24948
rect 30034 24892 30044 24948
rect 30100 24892 30940 24948
rect 30996 24892 31006 24948
rect 45154 24892 45164 24948
rect 45220 24892 50000 24948
rect 0 24864 800 24892
rect 2380 24724 2436 24892
rect 10770 24780 10780 24836
rect 10836 24780 11900 24836
rect 11956 24780 11966 24836
rect 15698 24780 15708 24836
rect 15764 24780 16156 24836
rect 16212 24780 16222 24836
rect 2370 24668 2380 24724
rect 2436 24668 2446 24724
rect 5590 24668 5628 24724
rect 5684 24668 9548 24724
rect 9604 24668 9614 24724
rect 10882 24668 10892 24724
rect 10948 24668 11228 24724
rect 11284 24668 11564 24724
rect 11620 24668 12012 24724
rect 12068 24668 13020 24724
rect 13076 24668 13086 24724
rect 2146 24556 2156 24612
rect 2212 24556 3388 24612
rect 3444 24556 3454 24612
rect 6738 24556 6748 24612
rect 6804 24556 8876 24612
rect 8932 24556 8942 24612
rect 6402 24444 6412 24500
rect 6468 24444 11340 24500
rect 11396 24444 11406 24500
rect 12338 24444 12348 24500
rect 12404 24444 13356 24500
rect 13412 24444 13916 24500
rect 13972 24444 13982 24500
rect 5058 24332 5068 24388
rect 5124 24332 15148 24388
rect 4466 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4750 24332
rect 15092 24276 15148 24332
rect 11106 24220 11116 24276
rect 11172 24220 11340 24276
rect 11396 24220 11406 24276
rect 13906 24220 13916 24276
rect 13972 24220 14476 24276
rect 14532 24220 14924 24276
rect 14980 24220 14990 24276
rect 15092 24220 15372 24276
rect 15428 24220 15438 24276
rect 16716 24164 16772 24892
rect 49200 24864 50000 24892
rect 41794 24780 41804 24836
rect 41860 24780 42700 24836
rect 42756 24780 43820 24836
rect 43876 24780 44940 24836
rect 44996 24780 45724 24836
rect 45780 24780 45790 24836
rect 16930 24668 16940 24724
rect 16996 24668 18060 24724
rect 18116 24668 18126 24724
rect 29250 24668 29260 24724
rect 29316 24668 30828 24724
rect 30884 24668 30894 24724
rect 41122 24668 41132 24724
rect 41188 24668 42476 24724
rect 42532 24668 42542 24724
rect 19842 24556 19852 24612
rect 19908 24556 20748 24612
rect 20804 24556 21868 24612
rect 21924 24556 21934 24612
rect 40002 24556 40012 24612
rect 40068 24556 41020 24612
rect 41076 24556 41086 24612
rect 38658 24444 38668 24500
rect 38724 24444 40348 24500
rect 40404 24444 40414 24500
rect 40674 24444 40684 24500
rect 40740 24444 42140 24500
rect 42196 24444 42206 24500
rect 37986 24332 37996 24388
rect 38052 24332 43036 24388
rect 43092 24332 43102 24388
rect 35186 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35470 24332
rect 49200 24276 50000 24304
rect 44034 24220 44044 24276
rect 44100 24220 50000 24276
rect 49200 24192 50000 24220
rect 2034 24108 2044 24164
rect 2100 24108 16772 24164
rect 4610 23996 4620 24052
rect 4676 23996 8204 24052
rect 8260 23996 8270 24052
rect 11778 23996 11788 24052
rect 11844 23996 16212 24052
rect 16930 23996 16940 24052
rect 16996 23996 17836 24052
rect 17892 23996 17902 24052
rect 26786 23996 26796 24052
rect 26852 23996 27804 24052
rect 27860 23996 27870 24052
rect 36306 23996 36316 24052
rect 36372 23996 37100 24052
rect 37156 23996 44940 24052
rect 44996 23996 45006 24052
rect 16156 23940 16212 23996
rect 6514 23884 6524 23940
rect 6580 23884 6748 23940
rect 6804 23884 6814 23940
rect 7186 23884 7196 23940
rect 7252 23884 11900 23940
rect 11956 23884 12460 23940
rect 12516 23884 12526 23940
rect 16156 23884 17276 23940
rect 17332 23884 17342 23940
rect 28578 23884 28588 23940
rect 28644 23884 29372 23940
rect 29428 23884 30828 23940
rect 30884 23884 30894 23940
rect 35970 23884 35980 23940
rect 36036 23884 45612 23940
rect 45668 23884 45678 23940
rect 6290 23772 6300 23828
rect 6356 23772 6860 23828
rect 6916 23772 6926 23828
rect 9202 23772 9212 23828
rect 9268 23772 10892 23828
rect 10948 23772 10958 23828
rect 12226 23772 12236 23828
rect 12292 23772 13580 23828
rect 13636 23772 13646 23828
rect 15362 23772 15372 23828
rect 15428 23772 15708 23828
rect 15764 23772 15774 23828
rect 16034 23772 16044 23828
rect 16100 23772 18284 23828
rect 18340 23772 18350 23828
rect 36418 23772 36428 23828
rect 36484 23772 40012 23828
rect 40068 23772 40078 23828
rect 41906 23772 41916 23828
rect 41972 23772 42588 23828
rect 42644 23772 42654 23828
rect 43138 23772 43148 23828
rect 43204 23772 43596 23828
rect 43652 23772 43662 23828
rect 6066 23660 6076 23716
rect 6132 23660 8652 23716
rect 8708 23660 8988 23716
rect 9044 23660 9054 23716
rect 9986 23660 9996 23716
rect 10052 23660 10556 23716
rect 10612 23660 10622 23716
rect 11666 23660 11676 23716
rect 11732 23660 14476 23716
rect 14532 23660 14542 23716
rect 17378 23660 17388 23716
rect 17444 23660 21700 23716
rect 35522 23660 35532 23716
rect 35588 23660 37436 23716
rect 37492 23660 37502 23716
rect 47394 23660 47404 23716
rect 47460 23660 48300 23716
rect 48356 23660 48366 23716
rect 0 23604 800 23632
rect 0 23548 1708 23604
rect 1764 23548 1774 23604
rect 6290 23548 6300 23604
rect 6356 23548 6972 23604
rect 7028 23548 7038 23604
rect 9202 23548 9212 23604
rect 9268 23548 10108 23604
rect 10164 23548 10174 23604
rect 10770 23548 10780 23604
rect 10836 23548 14252 23604
rect 14308 23548 14318 23604
rect 0 23520 800 23548
rect 11564 23492 11620 23548
rect 19826 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20110 23548
rect 11554 23436 11564 23492
rect 11620 23436 11630 23492
rect 21644 23380 21700 23660
rect 49200 23604 50000 23632
rect 23426 23548 23436 23604
rect 23492 23548 24332 23604
rect 24388 23548 28700 23604
rect 28756 23548 32732 23604
rect 32788 23548 32798 23604
rect 35858 23548 35868 23604
rect 35924 23548 38892 23604
rect 38948 23548 38958 23604
rect 47954 23548 47964 23604
rect 48020 23548 50000 23604
rect 38444 23492 38500 23548
rect 49200 23520 50000 23548
rect 22418 23436 22428 23492
rect 22484 23436 25228 23492
rect 25284 23436 25294 23492
rect 25442 23436 25452 23492
rect 25508 23436 29036 23492
rect 29092 23436 29102 23492
rect 30258 23436 30268 23492
rect 30324 23436 32060 23492
rect 32116 23436 32126 23492
rect 38434 23436 38444 23492
rect 38500 23436 38510 23492
rect 41794 23436 41804 23492
rect 41860 23436 42364 23492
rect 42420 23436 44044 23492
rect 44100 23436 44110 23492
rect 6626 23324 6636 23380
rect 6692 23324 9436 23380
rect 9492 23324 11788 23380
rect 11844 23324 11854 23380
rect 12562 23324 12572 23380
rect 12628 23324 17836 23380
rect 17892 23324 17902 23380
rect 21644 23324 26572 23380
rect 26628 23324 26638 23380
rect 29362 23324 29372 23380
rect 29428 23324 30940 23380
rect 30996 23324 31006 23380
rect 37426 23324 37436 23380
rect 37492 23324 37884 23380
rect 37940 23324 37950 23380
rect 40002 23324 40012 23380
rect 40068 23324 40796 23380
rect 40852 23324 40862 23380
rect 44370 23324 44380 23380
rect 44436 23324 46508 23380
rect 46564 23324 46574 23380
rect 6514 23212 6524 23268
rect 6580 23212 8652 23268
rect 8708 23212 10108 23268
rect 10164 23212 10174 23268
rect 15026 23212 15036 23268
rect 15092 23212 16156 23268
rect 16212 23212 16222 23268
rect 22866 23212 22876 23268
rect 22932 23212 24220 23268
rect 24276 23212 24286 23268
rect 25554 23212 25564 23268
rect 25620 23212 27580 23268
rect 27636 23212 29484 23268
rect 29540 23212 29550 23268
rect 31042 23212 31052 23268
rect 31108 23212 31500 23268
rect 31556 23212 31566 23268
rect 31938 23212 31948 23268
rect 32004 23212 33740 23268
rect 33796 23212 33806 23268
rect 40114 23212 40124 23268
rect 40180 23212 42924 23268
rect 42980 23212 45388 23268
rect 45444 23212 45454 23268
rect 46834 23212 46844 23268
rect 46900 23212 47180 23268
rect 47236 23212 48188 23268
rect 48244 23212 48254 23268
rect 7410 23100 7420 23156
rect 7476 23100 9660 23156
rect 9716 23100 9726 23156
rect 10518 23100 10556 23156
rect 10612 23100 10622 23156
rect 10882 23100 10892 23156
rect 10948 23100 13244 23156
rect 13300 23100 14924 23156
rect 14980 23100 14990 23156
rect 24322 23100 24332 23156
rect 24388 23100 25340 23156
rect 25396 23100 25676 23156
rect 25732 23100 25742 23156
rect 29670 23100 29708 23156
rect 29764 23100 29774 23156
rect 35522 23100 35532 23156
rect 35588 23100 42028 23156
rect 42084 23100 42094 23156
rect 42802 23100 42812 23156
rect 42868 23100 43484 23156
rect 43540 23100 43550 23156
rect 1810 22988 1820 23044
rect 1876 22988 3948 23044
rect 4004 22988 4844 23044
rect 4900 22988 4910 23044
rect 7634 22988 7644 23044
rect 7700 22988 14028 23044
rect 14084 22988 14094 23044
rect 36082 22988 36092 23044
rect 36148 22988 37996 23044
rect 38052 22988 39900 23044
rect 39956 22988 39966 23044
rect 49200 22932 50000 22960
rect 2034 22876 2044 22932
rect 2100 22876 4900 22932
rect 9426 22876 9436 22932
rect 9492 22876 9884 22932
rect 9940 22876 9950 22932
rect 16006 22876 16044 22932
rect 16100 22876 16110 22932
rect 18386 22876 18396 22932
rect 18452 22876 23660 22932
rect 23716 22876 23726 22932
rect 39666 22876 39676 22932
rect 39732 22876 40908 22932
rect 40964 22876 40974 22932
rect 41234 22876 41244 22932
rect 41300 22876 43148 22932
rect 43204 22876 43214 22932
rect 46946 22876 46956 22932
rect 47012 22876 50000 22932
rect 4466 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4750 22764
rect 4844 22596 4900 22876
rect 49200 22848 50000 22876
rect 5842 22764 5852 22820
rect 5908 22764 7196 22820
rect 7252 22764 7262 22820
rect 8754 22764 8764 22820
rect 8820 22764 10108 22820
rect 10164 22764 10332 22820
rect 10388 22764 10398 22820
rect 14466 22764 14476 22820
rect 14532 22764 15148 22820
rect 15204 22764 28364 22820
rect 28420 22764 28430 22820
rect 35186 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35470 22764
rect 8082 22652 8092 22708
rect 8148 22652 8428 22708
rect 8484 22652 8494 22708
rect 11330 22652 11340 22708
rect 11396 22652 12796 22708
rect 12852 22652 14140 22708
rect 14196 22652 14206 22708
rect 17826 22652 17836 22708
rect 17892 22652 23436 22708
rect 23492 22652 26348 22708
rect 26404 22652 26414 22708
rect 2482 22540 2492 22596
rect 2548 22540 3388 22596
rect 4844 22540 15372 22596
rect 15428 22540 19068 22596
rect 19124 22540 19134 22596
rect 26002 22540 26012 22596
rect 26068 22540 32508 22596
rect 32564 22540 32574 22596
rect 3332 22372 3388 22540
rect 4610 22428 4620 22484
rect 4676 22428 7308 22484
rect 7364 22428 9212 22484
rect 9268 22428 9278 22484
rect 9762 22428 9772 22484
rect 9828 22428 9838 22484
rect 10220 22428 15148 22484
rect 29586 22428 29596 22484
rect 29652 22428 30940 22484
rect 30996 22428 31006 22484
rect 44370 22428 44380 22484
rect 44436 22428 46284 22484
rect 46340 22428 47068 22484
rect 47124 22428 47134 22484
rect 9772 22372 9828 22428
rect 3332 22316 9828 22372
rect 6738 22204 6748 22260
rect 6804 22204 8708 22260
rect 8866 22204 8876 22260
rect 8932 22204 9324 22260
rect 9380 22204 9996 22260
rect 10052 22204 10062 22260
rect 8652 22148 8708 22204
rect 10220 22148 10276 22428
rect 15092 22372 15148 22428
rect 10434 22316 10444 22372
rect 10500 22316 14028 22372
rect 14084 22316 14094 22372
rect 15092 22316 21084 22372
rect 21140 22316 21150 22372
rect 30706 22316 30716 22372
rect 30772 22316 32060 22372
rect 32116 22316 32284 22372
rect 32340 22316 32350 22372
rect 37874 22316 37884 22372
rect 37940 22316 39844 22372
rect 40002 22316 40012 22372
rect 40068 22316 40572 22372
rect 40628 22316 40638 22372
rect 14028 22260 14084 22316
rect 39788 22260 39844 22316
rect 49200 22260 50000 22288
rect 13122 22204 13132 22260
rect 13188 22204 13468 22260
rect 13524 22204 13534 22260
rect 14028 22204 21756 22260
rect 21812 22204 21822 22260
rect 22530 22204 22540 22260
rect 22596 22204 22876 22260
rect 22932 22204 22942 22260
rect 37548 22204 39564 22260
rect 39620 22204 39630 22260
rect 39778 22204 39788 22260
rect 39844 22204 39854 22260
rect 40786 22204 40796 22260
rect 40852 22204 42252 22260
rect 42308 22204 42318 22260
rect 45266 22204 45276 22260
rect 45332 22204 46060 22260
rect 46116 22204 46126 22260
rect 47954 22204 47964 22260
rect 48020 22204 50000 22260
rect 37548 22148 37604 22204
rect 49200 22176 50000 22204
rect 6066 22092 6076 22148
rect 6132 22092 7756 22148
rect 7812 22092 7822 22148
rect 8652 22092 10276 22148
rect 12898 22092 12908 22148
rect 12964 22092 13692 22148
rect 13748 22092 13758 22148
rect 15586 22092 15596 22148
rect 15652 22092 20188 22148
rect 20244 22092 20254 22148
rect 37538 22092 37548 22148
rect 37604 22092 37614 22148
rect 38098 22092 38108 22148
rect 38164 22092 38174 22148
rect 38434 22092 38444 22148
rect 38500 22092 45612 22148
rect 45668 22092 45678 22148
rect 12114 21980 12124 22036
rect 12180 21980 12684 22036
rect 12740 21980 12750 22036
rect 19826 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20110 21980
rect 38108 21924 38164 22092
rect 38882 21980 38892 22036
rect 38948 21980 43484 22036
rect 43540 21980 43550 22036
rect 45378 21980 45388 22036
rect 45444 21980 46060 22036
rect 46116 21980 46126 22036
rect 7644 21868 8764 21924
rect 8820 21868 8830 21924
rect 10882 21868 10892 21924
rect 10948 21868 13244 21924
rect 13300 21868 14476 21924
rect 14532 21868 14542 21924
rect 29138 21868 29148 21924
rect 29204 21868 29708 21924
rect 29764 21868 31388 21924
rect 31444 21868 31454 21924
rect 38108 21868 40012 21924
rect 40068 21868 40078 21924
rect 7644 21812 7700 21868
rect 5618 21756 5628 21812
rect 5684 21756 6972 21812
rect 7028 21756 7700 21812
rect 7858 21756 7868 21812
rect 7924 21756 8652 21812
rect 8708 21756 20636 21812
rect 20692 21756 22988 21812
rect 23044 21756 23212 21812
rect 23268 21756 23278 21812
rect 29250 21756 29260 21812
rect 29316 21756 30828 21812
rect 30884 21756 30894 21812
rect 42130 21756 42140 21812
rect 42196 21756 42812 21812
rect 42868 21756 43260 21812
rect 43316 21756 43326 21812
rect 43586 21756 43596 21812
rect 43652 21756 45388 21812
rect 45444 21756 45454 21812
rect 6738 21644 6748 21700
rect 6804 21644 7644 21700
rect 7700 21644 8092 21700
rect 8148 21644 8158 21700
rect 11442 21644 11452 21700
rect 11508 21644 12124 21700
rect 12180 21644 12190 21700
rect 12898 21644 12908 21700
rect 12964 21644 13804 21700
rect 13860 21644 13870 21700
rect 37538 21644 37548 21700
rect 37604 21644 39004 21700
rect 39060 21644 39070 21700
rect 49200 21588 50000 21616
rect 5058 21532 5068 21588
rect 5124 21532 5852 21588
rect 5908 21532 12236 21588
rect 12292 21532 14812 21588
rect 14868 21532 15484 21588
rect 15540 21532 15550 21588
rect 20290 21532 20300 21588
rect 20356 21532 23100 21588
rect 23156 21532 23166 21588
rect 26786 21532 26796 21588
rect 26852 21532 27692 21588
rect 27748 21532 27758 21588
rect 30146 21532 30156 21588
rect 30212 21532 30492 21588
rect 30548 21532 30558 21588
rect 30818 21532 30828 21588
rect 30884 21532 32060 21588
rect 32116 21532 32126 21588
rect 44146 21532 44156 21588
rect 44212 21532 47516 21588
rect 47572 21532 47582 21588
rect 48290 21532 48300 21588
rect 48356 21532 50000 21588
rect 49200 21504 50000 21532
rect 5170 21420 5180 21476
rect 5236 21420 7420 21476
rect 7476 21420 7486 21476
rect 8978 21420 8988 21476
rect 9044 21420 11228 21476
rect 11284 21420 11788 21476
rect 11844 21420 11854 21476
rect 14690 21420 14700 21476
rect 14756 21420 16492 21476
rect 16548 21420 16558 21476
rect 36866 21420 36876 21476
rect 36932 21420 37660 21476
rect 37716 21420 37726 21476
rect 4610 21308 4620 21364
rect 4676 21308 10332 21364
rect 10388 21308 10398 21364
rect 21634 21308 21644 21364
rect 21700 21308 22428 21364
rect 22484 21308 23660 21364
rect 23716 21308 24220 21364
rect 24276 21308 28252 21364
rect 28308 21308 28318 21364
rect 34626 21308 34636 21364
rect 34692 21308 35196 21364
rect 35252 21308 38332 21364
rect 38388 21308 38398 21364
rect 45042 21308 45052 21364
rect 45108 21308 46956 21364
rect 47012 21308 47022 21364
rect 8418 21196 8428 21252
rect 8484 21196 13580 21252
rect 13636 21196 13646 21252
rect 41906 21196 41916 21252
rect 41972 21196 43260 21252
rect 43316 21196 43326 21252
rect 4466 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4750 21196
rect 35186 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35470 21196
rect 35970 20972 35980 21028
rect 36036 20972 37212 21028
rect 37268 20972 38444 21028
rect 38500 20972 38510 21028
rect 49200 20916 50000 20944
rect 10658 20860 10668 20916
rect 10724 20860 10892 20916
rect 10948 20860 10958 20916
rect 11302 20860 11340 20916
rect 11396 20860 11406 20916
rect 22978 20860 22988 20916
rect 23044 20860 23996 20916
rect 24052 20860 24062 20916
rect 31266 20860 31276 20916
rect 31332 20860 32172 20916
rect 32228 20860 32238 20916
rect 35746 20860 35756 20916
rect 35812 20860 36428 20916
rect 36484 20860 37660 20916
rect 37716 20860 42028 20916
rect 42084 20860 43148 20916
rect 43204 20860 43214 20916
rect 47506 20860 47516 20916
rect 47572 20860 50000 20916
rect 49200 20832 50000 20860
rect 6514 20748 6524 20804
rect 6580 20748 7868 20804
rect 7924 20748 8876 20804
rect 8932 20748 8942 20804
rect 10882 20748 10892 20804
rect 10948 20748 11564 20804
rect 11620 20748 11630 20804
rect 13906 20748 13916 20804
rect 13972 20748 18956 20804
rect 19012 20748 19022 20804
rect 21970 20748 21980 20804
rect 22036 20748 22764 20804
rect 22820 20748 23212 20804
rect 23268 20748 23278 20804
rect 30930 20748 30940 20804
rect 30996 20748 31500 20804
rect 31556 20748 34636 20804
rect 34692 20748 34702 20804
rect 40002 20748 40012 20804
rect 40068 20748 46620 20804
rect 46676 20748 46686 20804
rect 10546 20636 10556 20692
rect 10612 20636 14700 20692
rect 14756 20636 14766 20692
rect 15810 20636 15820 20692
rect 15876 20636 16604 20692
rect 16660 20636 16670 20692
rect 26562 20636 26572 20692
rect 26628 20636 31948 20692
rect 32004 20636 32014 20692
rect 42130 20636 42140 20692
rect 42196 20636 42924 20692
rect 42980 20636 42990 20692
rect 10882 20524 10892 20580
rect 10948 20524 11788 20580
rect 11844 20524 11854 20580
rect 12236 20468 12292 20636
rect 12646 20524 12684 20580
rect 12740 20524 12750 20580
rect 14102 20524 14140 20580
rect 14196 20524 14206 20580
rect 14578 20524 14588 20580
rect 14644 20524 16380 20580
rect 16436 20524 16446 20580
rect 16706 20524 16716 20580
rect 16772 20524 17276 20580
rect 17332 20524 18060 20580
rect 18116 20524 18126 20580
rect 27570 20524 27580 20580
rect 27636 20524 28364 20580
rect 28420 20524 31052 20580
rect 31108 20524 38668 20580
rect 12226 20412 12236 20468
rect 12292 20412 12302 20468
rect 15474 20412 15484 20468
rect 15540 20412 18284 20468
rect 18340 20412 18350 20468
rect 34402 20412 34412 20468
rect 34468 20412 35308 20468
rect 35364 20412 35374 20468
rect 38612 20412 38668 20524
rect 38724 20412 38734 20468
rect 19826 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20110 20412
rect 7410 20300 7420 20356
rect 7476 20300 9100 20356
rect 9156 20300 9166 20356
rect 10882 20300 10892 20356
rect 10948 20300 12124 20356
rect 12180 20300 12190 20356
rect 16370 20300 16380 20356
rect 16436 20300 16940 20356
rect 16996 20300 17006 20356
rect 49200 20244 50000 20272
rect 5404 20188 5740 20244
rect 5796 20188 6524 20244
rect 6580 20188 6590 20244
rect 7522 20188 7532 20244
rect 7588 20188 8204 20244
rect 8260 20188 8270 20244
rect 15698 20188 15708 20244
rect 15764 20188 16044 20244
rect 16100 20188 16110 20244
rect 23090 20188 23100 20244
rect 23156 20188 24108 20244
rect 24164 20188 24174 20244
rect 30370 20188 30380 20244
rect 30436 20188 31276 20244
rect 31332 20188 31342 20244
rect 32386 20188 32396 20244
rect 32452 20188 33292 20244
rect 33348 20188 34300 20244
rect 34356 20188 34366 20244
rect 44146 20188 44156 20244
rect 44212 20188 45052 20244
rect 45108 20188 45118 20244
rect 47964 20188 50000 20244
rect 5404 20132 5460 20188
rect 47964 20132 48020 20188
rect 49200 20160 50000 20188
rect 1698 20076 1708 20132
rect 1764 20076 3612 20132
rect 3668 20076 3678 20132
rect 4162 20076 4172 20132
rect 4228 20076 5460 20132
rect 5618 20076 5628 20132
rect 5684 20076 5964 20132
rect 6020 20076 6030 20132
rect 8642 20076 8652 20132
rect 8708 20076 9772 20132
rect 9828 20076 10556 20132
rect 10612 20076 10622 20132
rect 11106 20076 11116 20132
rect 11172 20076 13020 20132
rect 13076 20076 13086 20132
rect 13570 20076 13580 20132
rect 13636 20076 18956 20132
rect 19012 20076 19022 20132
rect 19730 20076 19740 20132
rect 19796 20076 20972 20132
rect 21028 20076 21038 20132
rect 30146 20076 30156 20132
rect 30212 20076 32284 20132
rect 32340 20076 32350 20132
rect 38994 20076 39004 20132
rect 39060 20076 41244 20132
rect 41300 20076 41310 20132
rect 43698 20076 43708 20132
rect 43764 20076 45612 20132
rect 45668 20076 45678 20132
rect 47954 20076 47964 20132
rect 48020 20076 48030 20132
rect 3490 19964 3500 20020
rect 3556 19964 4396 20020
rect 4452 19964 4462 20020
rect 6066 19964 6076 20020
rect 6132 19964 6860 20020
rect 6916 19964 6926 20020
rect 8530 19964 8540 20020
rect 8596 19964 9548 20020
rect 9604 19964 9614 20020
rect 11554 19964 11564 20020
rect 11620 19964 13916 20020
rect 13972 19964 13982 20020
rect 16034 19964 16044 20020
rect 16100 19964 16110 20020
rect 28018 19964 28028 20020
rect 28084 19964 28924 20020
rect 28980 19964 28990 20020
rect 40002 19964 40012 20020
rect 40068 19964 42476 20020
rect 42532 19964 42542 20020
rect 2482 19852 2492 19908
rect 2548 19852 4060 19908
rect 4116 19852 4126 19908
rect 4946 19852 4956 19908
rect 5012 19852 5740 19908
rect 5796 19852 5806 19908
rect 6402 19852 6412 19908
rect 6468 19852 7420 19908
rect 7476 19852 7486 19908
rect 9426 19852 9436 19908
rect 9492 19852 9772 19908
rect 9828 19852 10108 19908
rect 10164 19852 12908 19908
rect 12964 19852 12974 19908
rect 14018 19852 14028 19908
rect 14084 19852 15372 19908
rect 15428 19852 15438 19908
rect 16044 19796 16100 19964
rect 39218 19852 39228 19908
rect 39284 19852 41020 19908
rect 41076 19852 41086 19908
rect 4722 19740 4732 19796
rect 4788 19740 8764 19796
rect 8820 19740 8830 19796
rect 10210 19740 10220 19796
rect 10276 19740 11004 19796
rect 11060 19740 11070 19796
rect 13346 19740 13356 19796
rect 13412 19740 16100 19796
rect 20738 19740 20748 19796
rect 20804 19740 20814 19796
rect 27010 19740 27020 19796
rect 27076 19740 28812 19796
rect 28868 19740 28878 19796
rect 29250 19740 29260 19796
rect 29316 19740 36092 19796
rect 36148 19740 36158 19796
rect 39890 19740 39900 19796
rect 39956 19740 43372 19796
rect 43428 19740 43438 19796
rect 20748 19684 20804 19740
rect 14242 19628 14252 19684
rect 14308 19628 20804 19684
rect 41234 19628 41244 19684
rect 41300 19628 42700 19684
rect 42756 19628 43708 19684
rect 43764 19628 43774 19684
rect 4466 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4750 19628
rect 35186 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35470 19628
rect 6962 19516 6972 19572
rect 7028 19516 15820 19572
rect 15876 19516 15886 19572
rect 16818 19516 16828 19572
rect 16884 19516 16940 19572
rect 16996 19516 17006 19572
rect 4834 19404 4844 19460
rect 4900 19404 5180 19460
rect 5236 19404 5246 19460
rect 14466 19404 14476 19460
rect 14532 19404 17388 19460
rect 17444 19404 17454 19460
rect 27906 19404 27916 19460
rect 27972 19404 31836 19460
rect 31892 19404 31902 19460
rect 33170 19404 33180 19460
rect 33236 19404 35308 19460
rect 35364 19404 35374 19460
rect 2146 19292 2156 19348
rect 2212 19292 3500 19348
rect 3556 19292 5292 19348
rect 5348 19292 5358 19348
rect 15810 19292 15820 19348
rect 15876 19292 18844 19348
rect 18900 19292 18910 19348
rect 25554 19292 25564 19348
rect 25620 19292 25900 19348
rect 25956 19292 25966 19348
rect 29698 19292 29708 19348
rect 29764 19292 30156 19348
rect 30212 19292 30222 19348
rect 31266 19292 31276 19348
rect 31332 19292 33964 19348
rect 34020 19292 34030 19348
rect 39890 19292 39900 19348
rect 39956 19292 43036 19348
rect 43092 19292 43102 19348
rect 3602 19180 3612 19236
rect 3668 19180 3948 19236
rect 4004 19180 5068 19236
rect 5124 19180 5134 19236
rect 5394 19180 5404 19236
rect 5460 19180 8428 19236
rect 8484 19180 8494 19236
rect 10220 19180 10668 19236
rect 10724 19180 10734 19236
rect 12226 19180 12236 19236
rect 12292 19180 12908 19236
rect 12964 19180 12974 19236
rect 13682 19180 13692 19236
rect 13748 19180 14924 19236
rect 14980 19180 14990 19236
rect 20402 19180 20412 19236
rect 20468 19180 21308 19236
rect 21364 19180 21374 19236
rect 30258 19180 30268 19236
rect 30324 19180 33180 19236
rect 33236 19180 33246 19236
rect 41010 19180 41020 19236
rect 41076 19180 41692 19236
rect 41748 19180 42588 19236
rect 42644 19180 42654 19236
rect 10220 19124 10276 19180
rect 9314 19068 9324 19124
rect 9380 19068 9884 19124
rect 9940 19068 9950 19124
rect 10210 19068 10220 19124
rect 10276 19068 10286 19124
rect 10434 19068 10444 19124
rect 10500 19068 11116 19124
rect 11172 19068 11182 19124
rect 29250 19068 29260 19124
rect 29316 19068 29820 19124
rect 29876 19068 29886 19124
rect 32274 19068 32284 19124
rect 32340 19068 34188 19124
rect 34244 19068 34860 19124
rect 34916 19068 34926 19124
rect 35410 19068 35420 19124
rect 35476 19068 36764 19124
rect 36820 19068 36830 19124
rect 3826 18956 3836 19012
rect 3892 18956 4284 19012
rect 4340 18956 4350 19012
rect 5282 18956 5292 19012
rect 5348 18956 6076 19012
rect 6132 18956 7420 19012
rect 7476 18956 8204 19012
rect 8260 18956 8270 19012
rect 12114 18956 12124 19012
rect 12180 18956 13468 19012
rect 13524 18956 13534 19012
rect 16034 18956 16044 19012
rect 16100 18956 16716 19012
rect 16772 18956 16782 19012
rect 16930 18956 16940 19012
rect 16996 18956 17034 19012
rect 21970 18956 21980 19012
rect 22036 18956 28588 19012
rect 28644 18956 29708 19012
rect 29764 18956 30604 19012
rect 30660 18956 30670 19012
rect 30902 18956 30940 19012
rect 30996 18956 31006 19012
rect 31238 18956 31276 19012
rect 31332 18956 31342 19012
rect 32050 18956 32060 19012
rect 32116 18956 33516 19012
rect 33572 18956 33582 19012
rect 44258 18956 44268 19012
rect 44324 18956 48076 19012
rect 48132 18956 48142 19012
rect 29474 18844 29484 18900
rect 29540 18844 31164 18900
rect 31220 18844 31230 18900
rect 37650 18844 37660 18900
rect 37716 18844 45052 18900
rect 45108 18844 45612 18900
rect 45668 18844 45678 18900
rect 19826 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20110 18844
rect 9090 18732 9100 18788
rect 9156 18732 17276 18788
rect 17332 18732 17342 18788
rect 28690 18732 28700 18788
rect 28756 18732 30940 18788
rect 30996 18732 31006 18788
rect 31266 18732 31276 18788
rect 31332 18732 31612 18788
rect 31668 18732 31836 18788
rect 31892 18732 31902 18788
rect 33058 18732 33068 18788
rect 33124 18732 34300 18788
rect 34356 18732 36428 18788
rect 36484 18732 36494 18788
rect 10546 18620 10556 18676
rect 10612 18620 12796 18676
rect 12852 18620 12862 18676
rect 15922 18620 15932 18676
rect 15988 18620 16268 18676
rect 16324 18620 16334 18676
rect 19506 18620 19516 18676
rect 19572 18620 20748 18676
rect 20804 18620 23996 18676
rect 24052 18620 25452 18676
rect 25508 18620 25518 18676
rect 25890 18620 25900 18676
rect 25956 18620 26572 18676
rect 26628 18620 29036 18676
rect 29092 18620 29596 18676
rect 29652 18620 29662 18676
rect 30370 18620 30380 18676
rect 30436 18620 32508 18676
rect 32564 18620 32844 18676
rect 32900 18620 32910 18676
rect 40450 18620 40460 18676
rect 40516 18620 41356 18676
rect 41412 18620 41422 18676
rect 42438 18620 42476 18676
rect 42532 18620 42542 18676
rect 43474 18620 43484 18676
rect 43540 18620 47180 18676
rect 47236 18620 47246 18676
rect 42476 18564 42532 18620
rect 4834 18508 4844 18564
rect 4900 18508 5068 18564
rect 5124 18508 5134 18564
rect 8978 18508 8988 18564
rect 9044 18508 13244 18564
rect 13300 18508 13310 18564
rect 21756 18508 22652 18564
rect 22708 18508 25788 18564
rect 25844 18508 25854 18564
rect 28354 18508 28364 18564
rect 28420 18508 29932 18564
rect 29988 18508 29998 18564
rect 30146 18508 30156 18564
rect 30212 18508 31164 18564
rect 31220 18508 32956 18564
rect 33012 18508 33022 18564
rect 35298 18508 35308 18564
rect 35364 18508 36204 18564
rect 36260 18508 37212 18564
rect 37268 18508 37278 18564
rect 42242 18508 42252 18564
rect 42308 18508 42318 18564
rect 42476 18508 45836 18564
rect 45892 18508 45902 18564
rect 21756 18452 21812 18508
rect 30156 18452 30212 18508
rect 42252 18452 42308 18508
rect 1810 18396 1820 18452
rect 1876 18396 4060 18452
rect 4116 18396 4126 18452
rect 4610 18396 4620 18452
rect 4676 18396 9548 18452
rect 9604 18396 11900 18452
rect 11956 18396 11966 18452
rect 12562 18396 12572 18452
rect 12628 18396 14588 18452
rect 14644 18396 14654 18452
rect 21074 18396 21084 18452
rect 21140 18396 21812 18452
rect 23426 18396 23436 18452
rect 23492 18396 24220 18452
rect 24276 18396 24286 18452
rect 25666 18396 25676 18452
rect 25732 18396 26460 18452
rect 26516 18396 27244 18452
rect 27300 18396 27310 18452
rect 29810 18396 29820 18452
rect 29876 18396 30212 18452
rect 36642 18396 36652 18452
rect 36708 18396 37100 18452
rect 37156 18396 37166 18452
rect 38612 18396 39900 18452
rect 39956 18396 39966 18452
rect 40338 18396 40348 18452
rect 40404 18396 42308 18452
rect 42914 18396 42924 18452
rect 42980 18396 43260 18452
rect 43316 18396 43326 18452
rect 44706 18396 44716 18452
rect 44772 18396 46060 18452
rect 46116 18396 46126 18452
rect 46610 18396 46620 18452
rect 46676 18396 47852 18452
rect 47908 18396 47918 18452
rect 38612 18340 38668 18396
rect 2482 18284 2492 18340
rect 2548 18284 5180 18340
rect 5236 18284 5246 18340
rect 10322 18284 10332 18340
rect 10388 18284 11564 18340
rect 11620 18284 11630 18340
rect 21522 18284 21532 18340
rect 21588 18284 23884 18340
rect 23940 18284 23950 18340
rect 24322 18284 24332 18340
rect 24388 18284 25564 18340
rect 25620 18284 25630 18340
rect 27010 18284 27020 18340
rect 27076 18284 27086 18340
rect 31714 18284 31724 18340
rect 31780 18284 33068 18340
rect 33124 18284 33134 18340
rect 36418 18284 36428 18340
rect 36484 18284 38668 18340
rect 27020 18228 27076 18284
rect 42252 18228 42308 18396
rect 45266 18284 45276 18340
rect 45332 18284 46396 18340
rect 46452 18284 46462 18340
rect 4162 18172 4172 18228
rect 4228 18172 7084 18228
rect 7140 18172 7308 18228
rect 7364 18172 7374 18228
rect 10882 18172 10892 18228
rect 10948 18172 12236 18228
rect 12292 18172 13804 18228
rect 13860 18172 13870 18228
rect 14802 18172 14812 18228
rect 14868 18172 16268 18228
rect 16324 18172 16334 18228
rect 27020 18172 38444 18228
rect 38500 18172 38510 18228
rect 42130 18172 42140 18228
rect 42196 18172 42308 18228
rect 42662 18172 42700 18228
rect 42756 18172 42766 18228
rect 43474 18172 43484 18228
rect 43540 18172 47516 18228
rect 47572 18172 47582 18228
rect 6514 18060 6524 18116
rect 6580 18060 7868 18116
rect 7924 18060 10780 18116
rect 10836 18060 11788 18116
rect 11844 18060 11854 18116
rect 36194 18060 36204 18116
rect 36260 18060 37324 18116
rect 37380 18060 40572 18116
rect 40628 18060 40638 18116
rect 44930 18060 44940 18116
rect 44996 18060 47628 18116
rect 47684 18060 47694 18116
rect 4466 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4750 18060
rect 35186 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35470 18060
rect 5170 17948 5180 18004
rect 5236 17948 5740 18004
rect 5796 17948 5806 18004
rect 6860 17948 6972 18004
rect 7028 17948 7038 18004
rect 8194 17948 8204 18004
rect 8260 17948 12684 18004
rect 12740 17948 13580 18004
rect 13636 17948 21420 18004
rect 21476 17948 21486 18004
rect 30930 17948 30940 18004
rect 30996 17948 31836 18004
rect 31892 17948 34412 18004
rect 34468 17948 34478 18004
rect 44370 17948 44380 18004
rect 44436 17948 44446 18004
rect 6860 17892 6916 17948
rect 44380 17892 44436 17948
rect 3938 17836 3948 17892
rect 4004 17836 12572 17892
rect 12628 17836 12638 17892
rect 31266 17836 31276 17892
rect 31332 17836 40236 17892
rect 40292 17836 43708 17892
rect 43764 17836 44940 17892
rect 44996 17836 45006 17892
rect 1922 17724 1932 17780
rect 1988 17724 1998 17780
rect 5842 17724 5852 17780
rect 5908 17724 7084 17780
rect 7140 17724 7150 17780
rect 11106 17724 11116 17780
rect 11172 17724 11452 17780
rect 11508 17724 11518 17780
rect 16370 17724 16380 17780
rect 16436 17724 16828 17780
rect 16884 17724 16894 17780
rect 30146 17724 30156 17780
rect 30212 17724 30828 17780
rect 30884 17724 30894 17780
rect 42018 17724 42028 17780
rect 42084 17724 42700 17780
rect 42756 17724 42766 17780
rect 44034 17724 44044 17780
rect 44100 17724 44110 17780
rect 46050 17724 46060 17780
rect 46116 17724 48188 17780
rect 48244 17724 48254 17780
rect 0 17556 800 17584
rect 1932 17556 1988 17724
rect 5618 17612 5628 17668
rect 5684 17612 6300 17668
rect 6356 17612 7196 17668
rect 7252 17612 7262 17668
rect 14018 17612 14028 17668
rect 14084 17612 14588 17668
rect 14644 17612 17500 17668
rect 17556 17612 17566 17668
rect 19730 17612 19740 17668
rect 19796 17612 22092 17668
rect 22148 17612 22158 17668
rect 25218 17612 25228 17668
rect 25284 17612 31500 17668
rect 31556 17612 31836 17668
rect 31892 17612 31902 17668
rect 32274 17612 32284 17668
rect 32340 17612 32620 17668
rect 32676 17612 32686 17668
rect 40338 17612 40348 17668
rect 40404 17612 43708 17668
rect 43764 17612 43774 17668
rect 0 17500 1988 17556
rect 5954 17500 5964 17556
rect 6020 17500 6636 17556
rect 6692 17500 8652 17556
rect 8708 17500 8718 17556
rect 9090 17500 9100 17556
rect 9156 17500 16940 17556
rect 16996 17500 17836 17556
rect 17892 17500 21980 17556
rect 22036 17500 22046 17556
rect 32946 17500 32956 17556
rect 33012 17500 35644 17556
rect 35700 17500 35710 17556
rect 39218 17500 39228 17556
rect 39284 17500 40572 17556
rect 40628 17500 40638 17556
rect 42354 17500 42364 17556
rect 42420 17500 42700 17556
rect 42756 17500 42766 17556
rect 0 17472 800 17500
rect 44044 17444 44100 17724
rect 5058 17388 5068 17444
rect 5124 17388 5740 17444
rect 5796 17388 5806 17444
rect 7970 17388 7980 17444
rect 8036 17388 8540 17444
rect 8596 17388 8606 17444
rect 15810 17388 15820 17444
rect 15876 17388 16268 17444
rect 16324 17388 17500 17444
rect 17556 17388 17948 17444
rect 18004 17388 18284 17444
rect 18340 17388 22596 17444
rect 32050 17388 32060 17444
rect 32116 17388 34972 17444
rect 35028 17388 35532 17444
rect 35588 17388 35598 17444
rect 38434 17388 38444 17444
rect 38500 17388 40908 17444
rect 40964 17388 40974 17444
rect 44044 17388 44604 17444
rect 44660 17388 45052 17444
rect 45108 17388 45118 17444
rect 22540 17332 22596 17388
rect 3826 17276 3836 17332
rect 3892 17276 6748 17332
rect 6804 17276 8428 17332
rect 8484 17276 8494 17332
rect 11890 17276 11900 17332
rect 11956 17276 12684 17332
rect 12740 17276 14476 17332
rect 14532 17276 14542 17332
rect 22530 17276 22540 17332
rect 22596 17276 38668 17332
rect 38724 17276 40460 17332
rect 40516 17276 40526 17332
rect 44370 17276 44380 17332
rect 44436 17276 48300 17332
rect 48356 17276 48366 17332
rect 19826 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20110 17276
rect 11302 17164 11340 17220
rect 11396 17164 11406 17220
rect 17602 17164 17612 17220
rect 17668 17164 19292 17220
rect 19348 17164 19358 17220
rect 31490 17164 31500 17220
rect 31556 17164 32060 17220
rect 32116 17164 32126 17220
rect 36530 17164 36540 17220
rect 36596 17164 36606 17220
rect 37538 17164 37548 17220
rect 37604 17164 37884 17220
rect 37940 17164 37950 17220
rect 40226 17164 40236 17220
rect 40292 17164 41132 17220
rect 41188 17164 41198 17220
rect 42774 17164 42812 17220
rect 42868 17164 42878 17220
rect 44034 17164 44044 17220
rect 44100 17164 44828 17220
rect 44884 17164 44894 17220
rect 36540 17108 36596 17164
rect 3266 17052 3276 17108
rect 3332 17052 4172 17108
rect 4228 17052 5068 17108
rect 5124 17052 5134 17108
rect 14466 17052 14476 17108
rect 14532 17052 19628 17108
rect 19684 17052 19694 17108
rect 22082 17052 22092 17108
rect 22148 17052 23772 17108
rect 23828 17052 25228 17108
rect 25284 17052 25294 17108
rect 31826 17052 31836 17108
rect 31892 17052 33068 17108
rect 33124 17052 33134 17108
rect 34626 17052 34636 17108
rect 34692 17052 35420 17108
rect 35476 17052 41356 17108
rect 41412 17052 41422 17108
rect 42476 17052 43260 17108
rect 43316 17052 43326 17108
rect 43698 17052 43708 17108
rect 43764 17052 44492 17108
rect 44548 17052 44558 17108
rect 42476 16996 42532 17052
rect 5282 16940 5292 16996
rect 5348 16940 12236 16996
rect 12292 16940 12302 16996
rect 12460 16940 14924 16996
rect 14980 16940 14990 16996
rect 23314 16940 23324 16996
rect 23380 16940 28924 16996
rect 28980 16940 29260 16996
rect 29316 16940 29326 16996
rect 31714 16940 31724 16996
rect 31780 16940 31790 16996
rect 32834 16940 32844 16996
rect 32900 16940 33964 16996
rect 34020 16940 34972 16996
rect 35028 16940 35038 16996
rect 36530 16940 36540 16996
rect 36596 16940 38220 16996
rect 38276 16940 39004 16996
rect 39060 16940 39070 16996
rect 39442 16940 39452 16996
rect 39508 16940 39900 16996
rect 39956 16940 39966 16996
rect 40786 16940 40796 16996
rect 40852 16940 42532 16996
rect 42690 16940 42700 16996
rect 42756 16940 44268 16996
rect 44324 16940 44334 16996
rect 45490 16940 45500 16996
rect 45556 16940 46284 16996
rect 46340 16940 46956 16996
rect 47012 16940 48076 16996
rect 48132 16940 48142 16996
rect 12460 16884 12516 16940
rect 31724 16884 31780 16940
rect 2818 16828 2828 16884
rect 2884 16828 3500 16884
rect 3556 16828 3566 16884
rect 8082 16828 8092 16884
rect 8148 16828 8540 16884
rect 8596 16828 8606 16884
rect 10658 16828 10668 16884
rect 10724 16828 12124 16884
rect 12180 16828 12516 16884
rect 13458 16828 13468 16884
rect 13524 16828 13534 16884
rect 13794 16828 13804 16884
rect 13860 16828 15148 16884
rect 15204 16828 15214 16884
rect 16818 16828 16828 16884
rect 16884 16828 22316 16884
rect 22372 16828 22382 16884
rect 23874 16828 23884 16884
rect 23940 16828 24780 16884
rect 24836 16828 29484 16884
rect 29540 16828 29550 16884
rect 31724 16828 33516 16884
rect 33572 16828 34860 16884
rect 34916 16828 34926 16884
rect 39106 16828 39116 16884
rect 39172 16828 40908 16884
rect 40964 16828 40974 16884
rect 41122 16828 41132 16884
rect 41188 16828 41916 16884
rect 41972 16828 43484 16884
rect 43540 16828 43550 16884
rect 43810 16828 43820 16884
rect 43876 16828 44156 16884
rect 44212 16828 44222 16884
rect 46162 16828 46172 16884
rect 46228 16828 47292 16884
rect 47348 16828 47358 16884
rect 13468 16772 13524 16828
rect 1698 16716 1708 16772
rect 1764 16716 3164 16772
rect 3220 16716 3230 16772
rect 3378 16716 3388 16772
rect 3444 16716 5292 16772
rect 5348 16716 6076 16772
rect 6132 16716 6142 16772
rect 9762 16716 9772 16772
rect 9828 16716 10780 16772
rect 10836 16716 15372 16772
rect 15428 16716 16044 16772
rect 16100 16716 16110 16772
rect 16930 16716 16940 16772
rect 16996 16716 17500 16772
rect 17556 16716 21868 16772
rect 21924 16716 21934 16772
rect 22194 16716 22204 16772
rect 22260 16716 26236 16772
rect 26292 16716 26302 16772
rect 33842 16716 33852 16772
rect 33908 16716 34188 16772
rect 34244 16716 34254 16772
rect 38612 16716 40796 16772
rect 40852 16716 40862 16772
rect 46050 16716 46060 16772
rect 46116 16716 46844 16772
rect 46900 16716 46910 16772
rect 38612 16660 38668 16716
rect 4498 16604 4508 16660
rect 4564 16604 4956 16660
rect 5012 16604 5628 16660
rect 5684 16604 14140 16660
rect 14196 16604 14206 16660
rect 22866 16604 22876 16660
rect 22932 16604 23660 16660
rect 23716 16604 23726 16660
rect 33058 16604 33068 16660
rect 33124 16604 38668 16660
rect 39890 16604 39900 16660
rect 39956 16604 40684 16660
rect 40740 16604 41916 16660
rect 41972 16604 41982 16660
rect 5170 16492 5180 16548
rect 5236 16492 7420 16548
rect 7476 16492 7486 16548
rect 37538 16492 37548 16548
rect 37604 16492 42924 16548
rect 42980 16492 42990 16548
rect 4466 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4750 16492
rect 35186 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35470 16492
rect 6626 16380 6636 16436
rect 6692 16380 12796 16436
rect 12852 16380 16660 16436
rect 20738 16380 20748 16436
rect 20804 16380 22428 16436
rect 22484 16380 24780 16436
rect 24836 16380 27916 16436
rect 27972 16380 27982 16436
rect 39554 16380 39564 16436
rect 39620 16380 41580 16436
rect 41636 16380 42812 16436
rect 42868 16380 42878 16436
rect 16604 16324 16660 16380
rect 3602 16268 3612 16324
rect 3668 16268 5852 16324
rect 5908 16268 5918 16324
rect 12562 16268 12572 16324
rect 12628 16268 14476 16324
rect 14532 16268 14542 16324
rect 16604 16268 21812 16324
rect 33842 16268 33852 16324
rect 33908 16268 37212 16324
rect 37268 16268 37278 16324
rect 38098 16268 38108 16324
rect 38164 16268 38668 16324
rect 38724 16268 38734 16324
rect 40338 16268 40348 16324
rect 40404 16268 41020 16324
rect 41076 16268 41086 16324
rect 21756 16212 21812 16268
rect 4610 16156 4620 16212
rect 4676 16156 5068 16212
rect 5124 16156 6188 16212
rect 6244 16156 6254 16212
rect 7634 16156 7644 16212
rect 7700 16156 8428 16212
rect 8484 16156 10556 16212
rect 10612 16156 10622 16212
rect 17266 16156 17276 16212
rect 17332 16156 20748 16212
rect 20804 16156 20814 16212
rect 21746 16156 21756 16212
rect 21812 16156 28700 16212
rect 28756 16156 28766 16212
rect 40114 16156 40124 16212
rect 40180 16156 42028 16212
rect 42084 16156 42094 16212
rect 42998 16156 43036 16212
rect 43092 16156 43102 16212
rect 44706 16156 44716 16212
rect 44772 16156 45612 16212
rect 45668 16156 46396 16212
rect 46452 16156 47516 16212
rect 47572 16156 47582 16212
rect 7410 16044 7420 16100
rect 7476 16044 7486 16100
rect 8082 16044 8092 16100
rect 8148 16044 11004 16100
rect 11060 16044 11070 16100
rect 18274 16044 18284 16100
rect 18340 16044 22204 16100
rect 22260 16044 22270 16100
rect 23650 16044 23660 16100
rect 23716 16044 24668 16100
rect 24724 16044 24734 16100
rect 34290 16044 34300 16100
rect 34356 16044 34860 16100
rect 34916 16044 35196 16100
rect 35252 16044 37212 16100
rect 37268 16044 37278 16100
rect 7420 15988 7476 16044
rect 7420 15932 9884 15988
rect 9940 15932 10332 15988
rect 10388 15932 10398 15988
rect 12002 15932 12012 15988
rect 12068 15932 13692 15988
rect 13748 15932 17388 15988
rect 17444 15932 17454 15988
rect 19954 15932 19964 15988
rect 20020 15932 21644 15988
rect 21700 15932 21710 15988
rect 23202 15932 23212 15988
rect 23268 15932 23436 15988
rect 23492 15932 24332 15988
rect 24388 15932 24398 15988
rect 28578 15932 28588 15988
rect 28644 15932 30268 15988
rect 30324 15932 30334 15988
rect 31602 15932 31612 15988
rect 31668 15932 33068 15988
rect 33124 15932 33134 15988
rect 40002 15932 40012 15988
rect 40068 15932 41244 15988
rect 41300 15932 41310 15988
rect 41458 15932 41468 15988
rect 41524 15932 41562 15988
rect 12562 15820 12572 15876
rect 12628 15820 13244 15876
rect 13300 15820 13310 15876
rect 14018 15820 14028 15876
rect 14084 15820 16492 15876
rect 16548 15820 16558 15876
rect 21644 15764 21700 15932
rect 24098 15820 24108 15876
rect 24164 15820 27916 15876
rect 27972 15820 27982 15876
rect 31126 15820 31164 15876
rect 31220 15820 31230 15876
rect 34178 15820 34188 15876
rect 34244 15820 35868 15876
rect 35924 15820 38220 15876
rect 38276 15820 38444 15876
rect 38500 15820 38510 15876
rect 39778 15820 39788 15876
rect 39844 15820 40236 15876
rect 40292 15820 42252 15876
rect 42308 15820 42318 15876
rect 21644 15708 24444 15764
rect 24500 15708 25676 15764
rect 25732 15708 25742 15764
rect 40898 15708 40908 15764
rect 40964 15708 42476 15764
rect 42532 15708 44940 15764
rect 44996 15708 45006 15764
rect 19826 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20110 15708
rect 17266 15596 17276 15652
rect 17332 15596 18396 15652
rect 18452 15596 18462 15652
rect 20402 15596 20412 15652
rect 20468 15596 22764 15652
rect 22820 15596 22830 15652
rect 26012 15596 32900 15652
rect 34402 15596 34412 15652
rect 34468 15596 34972 15652
rect 35028 15596 35756 15652
rect 35812 15596 37996 15652
rect 38052 15596 43036 15652
rect 43092 15596 43102 15652
rect 18396 15540 18452 15596
rect 9874 15484 9884 15540
rect 9940 15484 11004 15540
rect 11060 15484 11900 15540
rect 11956 15484 11966 15540
rect 18396 15484 21084 15540
rect 21140 15484 21868 15540
rect 21924 15484 21934 15540
rect 26012 15428 26068 15596
rect 7074 15372 7084 15428
rect 7140 15372 9548 15428
rect 9604 15372 11340 15428
rect 11396 15372 16380 15428
rect 16436 15372 16446 15428
rect 17714 15372 17724 15428
rect 17780 15372 25340 15428
rect 25396 15372 26012 15428
rect 26068 15372 26078 15428
rect 26674 15372 26684 15428
rect 26740 15372 27692 15428
rect 27748 15372 27758 15428
rect 4946 15260 4956 15316
rect 5012 15260 5292 15316
rect 5348 15260 6860 15316
rect 6916 15260 7868 15316
rect 7924 15260 7934 15316
rect 11106 15260 11116 15316
rect 11172 15260 11788 15316
rect 11844 15260 11854 15316
rect 12114 15260 12124 15316
rect 12180 15260 12236 15316
rect 12292 15260 12302 15316
rect 17378 15260 17388 15316
rect 17444 15260 20412 15316
rect 20468 15260 20478 15316
rect 23958 15260 23996 15316
rect 24052 15260 24062 15316
rect 24210 15260 24220 15316
rect 24276 15260 26124 15316
rect 26180 15260 26190 15316
rect 26852 15260 27580 15316
rect 27636 15260 27646 15316
rect 26852 15204 26908 15260
rect 2482 15148 2492 15204
rect 2548 15148 4844 15204
rect 4900 15148 4910 15204
rect 10322 15148 10332 15204
rect 10388 15148 12684 15204
rect 12740 15148 14588 15204
rect 14644 15148 15820 15204
rect 15876 15148 15886 15204
rect 16930 15148 16940 15204
rect 16996 15148 18620 15204
rect 18676 15148 18686 15204
rect 23538 15148 23548 15204
rect 23604 15148 24108 15204
rect 24164 15148 24174 15204
rect 26002 15148 26012 15204
rect 26068 15148 26908 15204
rect 32844 15204 32900 15596
rect 33814 15484 33852 15540
rect 33908 15484 33918 15540
rect 34514 15484 34524 15540
rect 34580 15484 37324 15540
rect 37380 15484 37772 15540
rect 37828 15484 37838 15540
rect 38322 15484 38332 15540
rect 38388 15484 40012 15540
rect 40068 15484 40796 15540
rect 40852 15484 42140 15540
rect 42196 15484 42206 15540
rect 40338 15372 40348 15428
rect 40404 15372 42588 15428
rect 42644 15372 42654 15428
rect 43036 15372 46732 15428
rect 46788 15372 46798 15428
rect 43036 15316 43092 15372
rect 36082 15260 36092 15316
rect 36148 15260 36876 15316
rect 36932 15260 39676 15316
rect 39732 15260 39742 15316
rect 41570 15260 41580 15316
rect 41636 15260 43092 15316
rect 43810 15260 43820 15316
rect 43876 15260 45948 15316
rect 46004 15260 47292 15316
rect 47348 15260 47358 15316
rect 32844 15148 41020 15204
rect 41076 15148 42364 15204
rect 42420 15148 42430 15204
rect 44146 15036 44156 15092
rect 44212 15036 47404 15092
rect 47460 15036 47470 15092
rect 39106 14924 39116 14980
rect 39172 14924 40012 14980
rect 40068 14924 40078 14980
rect 4466 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4750 14924
rect 35186 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35470 14924
rect 35634 14812 35644 14868
rect 35700 14812 36540 14868
rect 36596 14812 36606 14868
rect 43138 14812 43148 14868
rect 43204 14812 44940 14868
rect 44996 14812 45006 14868
rect 25554 14700 25564 14756
rect 25620 14700 29932 14756
rect 29988 14700 30940 14756
rect 30996 14700 31006 14756
rect 34290 14700 34300 14756
rect 34356 14700 35756 14756
rect 35812 14700 35822 14756
rect 40114 14700 40124 14756
rect 40180 14700 43596 14756
rect 43652 14700 44604 14756
rect 44660 14700 44670 14756
rect 4610 14588 4620 14644
rect 4676 14588 6076 14644
rect 6132 14588 6142 14644
rect 9986 14588 9996 14644
rect 10052 14588 10780 14644
rect 10836 14588 10846 14644
rect 11554 14588 11564 14644
rect 11620 14588 12012 14644
rect 12068 14588 12908 14644
rect 12964 14588 13468 14644
rect 13524 14588 17724 14644
rect 17780 14588 17790 14644
rect 20626 14588 20636 14644
rect 20692 14588 21196 14644
rect 21252 14588 21262 14644
rect 23650 14588 23660 14644
rect 23716 14588 26236 14644
rect 26292 14588 26302 14644
rect 28466 14588 28476 14644
rect 28532 14588 39564 14644
rect 39620 14588 39630 14644
rect 40562 14588 40572 14644
rect 40628 14588 41804 14644
rect 41860 14588 41870 14644
rect 43474 14588 43484 14644
rect 43540 14588 47068 14644
rect 47124 14588 47134 14644
rect 8642 14476 8652 14532
rect 8708 14476 9660 14532
rect 9716 14476 10668 14532
rect 10724 14476 10734 14532
rect 16482 14476 16492 14532
rect 16548 14476 17500 14532
rect 17556 14476 21308 14532
rect 21364 14476 22540 14532
rect 22596 14476 24556 14532
rect 24612 14476 25340 14532
rect 25396 14476 25406 14532
rect 28690 14476 28700 14532
rect 28756 14476 29484 14532
rect 29540 14476 29820 14532
rect 29876 14476 30156 14532
rect 30212 14476 30222 14532
rect 36306 14476 36316 14532
rect 36372 14476 37548 14532
rect 37604 14476 39004 14532
rect 39060 14476 39340 14532
rect 39396 14476 39406 14532
rect 40002 14476 40012 14532
rect 40068 14476 41132 14532
rect 41188 14476 41198 14532
rect 41430 14476 41468 14532
rect 41524 14476 41534 14532
rect 41682 14476 41692 14532
rect 41748 14476 42700 14532
rect 42756 14476 42766 14532
rect 44258 14476 44268 14532
rect 44324 14476 45836 14532
rect 45892 14476 45902 14532
rect 27234 14364 27244 14420
rect 27300 14364 28028 14420
rect 28084 14364 28094 14420
rect 31238 14364 31276 14420
rect 31332 14364 31342 14420
rect 33282 14364 33292 14420
rect 33348 14364 37884 14420
rect 37940 14364 40852 14420
rect 42130 14364 42140 14420
rect 42196 14364 43484 14420
rect 43540 14364 43550 14420
rect 40796 14308 40852 14364
rect 12786 14252 12796 14308
rect 12852 14252 16716 14308
rect 16772 14252 16782 14308
rect 24546 14252 24556 14308
rect 24612 14252 27356 14308
rect 27412 14252 27422 14308
rect 30706 14252 30716 14308
rect 30772 14252 34636 14308
rect 34692 14252 34702 14308
rect 38434 14252 38444 14308
rect 38500 14252 38668 14308
rect 39666 14252 39676 14308
rect 39732 14252 40460 14308
rect 40516 14252 40526 14308
rect 40786 14252 40796 14308
rect 40852 14252 40862 14308
rect 42018 14252 42028 14308
rect 42084 14252 42700 14308
rect 42756 14252 42766 14308
rect 38612 14196 38668 14252
rect 24742 14140 24780 14196
rect 24836 14140 24846 14196
rect 26114 14140 26124 14196
rect 26180 14140 27244 14196
rect 27300 14140 27310 14196
rect 27458 14140 27468 14196
rect 27524 14140 29596 14196
rect 29652 14140 33180 14196
rect 33236 14140 33246 14196
rect 38612 14140 40684 14196
rect 40740 14140 41244 14196
rect 41300 14140 41310 14196
rect 42354 14140 42364 14196
rect 42420 14140 44156 14196
rect 44212 14140 44222 14196
rect 19826 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20110 14140
rect 5058 14028 5068 14084
rect 5124 14028 5852 14084
rect 5908 14028 6636 14084
rect 6692 14028 7196 14084
rect 7252 14028 9660 14084
rect 9716 14028 10220 14084
rect 10276 14028 10286 14084
rect 30370 14028 30380 14084
rect 30436 14028 30716 14084
rect 30772 14028 31724 14084
rect 31780 14028 39788 14084
rect 39844 14028 41020 14084
rect 41076 14028 41086 14084
rect 5394 13916 5404 13972
rect 5460 13916 10444 13972
rect 10500 13916 10510 13972
rect 12786 13916 12796 13972
rect 12852 13916 14140 13972
rect 14196 13916 14206 13972
rect 18722 13916 18732 13972
rect 18788 13916 20636 13972
rect 20692 13916 20702 13972
rect 33404 13916 35644 13972
rect 35700 13916 36092 13972
rect 36148 13916 36158 13972
rect 37874 13916 37884 13972
rect 37940 13916 40012 13972
rect 40068 13916 40078 13972
rect 9874 13804 9884 13860
rect 9940 13804 12236 13860
rect 12292 13804 12302 13860
rect 20066 13804 20076 13860
rect 20132 13804 23828 13860
rect 24434 13804 24444 13860
rect 24500 13804 25004 13860
rect 25060 13804 29260 13860
rect 29316 13804 29326 13860
rect 29474 13804 29484 13860
rect 29540 13804 31276 13860
rect 31332 13804 31342 13860
rect 23772 13748 23828 13804
rect 33404 13748 33460 13916
rect 41458 13804 41468 13860
rect 41524 13804 42252 13860
rect 42308 13804 42812 13860
rect 42868 13804 42878 13860
rect 11330 13692 11340 13748
rect 11396 13692 12684 13748
rect 12740 13692 12750 13748
rect 23762 13692 23772 13748
rect 23828 13692 29372 13748
rect 29428 13692 29438 13748
rect 31154 13692 31164 13748
rect 31220 13692 33404 13748
rect 33460 13692 33470 13748
rect 33954 13692 33964 13748
rect 34020 13692 34300 13748
rect 34356 13692 34366 13748
rect 36418 13692 36428 13748
rect 36484 13692 36876 13748
rect 36932 13692 36942 13748
rect 38546 13692 38556 13748
rect 38612 13692 39004 13748
rect 39060 13692 39070 13748
rect 40450 13692 40460 13748
rect 40516 13692 41580 13748
rect 41636 13692 41646 13748
rect 46722 13692 46732 13748
rect 46788 13692 47404 13748
rect 47460 13692 47470 13748
rect 2482 13580 2492 13636
rect 2548 13580 4732 13636
rect 4788 13580 4798 13636
rect 9202 13580 9212 13636
rect 9268 13580 10444 13636
rect 10500 13580 10510 13636
rect 19170 13580 19180 13636
rect 19236 13580 20076 13636
rect 20132 13580 21980 13636
rect 22036 13580 22046 13636
rect 23314 13580 23324 13636
rect 23380 13580 23660 13636
rect 23716 13580 23726 13636
rect 23986 13580 23996 13636
rect 24052 13580 25116 13636
rect 25172 13580 25182 13636
rect 28018 13580 28028 13636
rect 28084 13580 28476 13636
rect 28532 13580 28924 13636
rect 28980 13580 32284 13636
rect 32340 13580 32350 13636
rect 39666 13580 39676 13636
rect 39732 13580 42476 13636
rect 42532 13580 43372 13636
rect 43428 13580 43438 13636
rect 9426 13468 9436 13524
rect 9492 13468 10220 13524
rect 10276 13468 10286 13524
rect 16594 13468 16604 13524
rect 16660 13468 19068 13524
rect 19124 13468 19134 13524
rect 19394 13468 19404 13524
rect 19460 13468 20636 13524
rect 20692 13468 20702 13524
rect 31266 13468 31276 13524
rect 31332 13468 31500 13524
rect 31556 13468 31566 13524
rect 34626 13468 34636 13524
rect 34692 13468 35588 13524
rect 35858 13468 35868 13524
rect 35924 13468 43148 13524
rect 43204 13468 43214 13524
rect 44370 13468 44380 13524
rect 44436 13468 47964 13524
rect 48020 13468 48030 13524
rect 26338 13356 26348 13412
rect 26404 13356 27244 13412
rect 27300 13356 27310 13412
rect 31126 13356 31164 13412
rect 31220 13356 31230 13412
rect 4466 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4750 13356
rect 35186 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35470 13356
rect 35532 13300 35588 13468
rect 35970 13356 35980 13412
rect 36036 13356 37212 13412
rect 37268 13356 37660 13412
rect 37716 13356 37726 13412
rect 40898 13356 40908 13412
rect 40964 13356 42700 13412
rect 42756 13356 42766 13412
rect 43810 13356 43820 13412
rect 43876 13356 44828 13412
rect 44884 13356 44894 13412
rect 13122 13244 13132 13300
rect 13188 13244 23100 13300
rect 23156 13244 23166 13300
rect 23958 13244 23996 13300
rect 24052 13244 24062 13300
rect 35532 13244 45164 13300
rect 45220 13244 45388 13300
rect 45444 13244 45454 13300
rect 4722 13132 4732 13188
rect 4788 13132 5180 13188
rect 5236 13132 5246 13188
rect 35410 13132 35420 13188
rect 35476 13132 42140 13188
rect 42196 13132 42700 13188
rect 42756 13132 42766 13188
rect 5282 13020 5292 13076
rect 5348 13020 10444 13076
rect 10500 13020 10510 13076
rect 12002 13020 12012 13076
rect 12068 13020 13468 13076
rect 13524 13020 13534 13076
rect 16258 13020 16268 13076
rect 16324 13020 18172 13076
rect 18228 13020 18238 13076
rect 19618 13020 19628 13076
rect 19684 13020 21868 13076
rect 21924 13020 21934 13076
rect 23538 13020 23548 13076
rect 23604 13020 24332 13076
rect 24388 13020 26908 13076
rect 26964 13020 26974 13076
rect 28690 13020 28700 13076
rect 28756 13020 30380 13076
rect 30436 13020 36764 13076
rect 36820 13020 36830 13076
rect 39442 13020 39452 13076
rect 39508 13020 41132 13076
rect 41188 13020 41692 13076
rect 41748 13020 41758 13076
rect 17714 12908 17724 12964
rect 17780 12908 17790 12964
rect 26226 12908 26236 12964
rect 26292 12908 27468 12964
rect 27524 12908 28252 12964
rect 28308 12908 28318 12964
rect 41458 12908 41468 12964
rect 41524 12908 44828 12964
rect 44884 12908 44894 12964
rect 17724 12852 17780 12908
rect 4610 12796 4620 12852
rect 4676 12796 5068 12852
rect 5124 12796 5852 12852
rect 5908 12796 5918 12852
rect 14466 12796 14476 12852
rect 14532 12796 15036 12852
rect 15092 12796 15372 12852
rect 15428 12796 15438 12852
rect 16706 12796 16716 12852
rect 16772 12796 29596 12852
rect 29652 12796 29662 12852
rect 29810 12796 29820 12852
rect 29876 12796 30268 12852
rect 30324 12796 30334 12852
rect 34402 12796 34412 12852
rect 34468 12796 34972 12852
rect 35028 12796 40012 12852
rect 40068 12796 40078 12852
rect 44930 12796 44940 12852
rect 44996 12796 46060 12852
rect 46116 12796 46126 12852
rect 5730 12684 5740 12740
rect 5796 12684 8876 12740
rect 8932 12684 8942 12740
rect 14018 12684 14028 12740
rect 14084 12684 15148 12740
rect 15204 12684 15214 12740
rect 19170 12684 19180 12740
rect 19236 12684 20188 12740
rect 20244 12684 20254 12740
rect 26852 12684 37772 12740
rect 37828 12684 37838 12740
rect 41458 12684 41468 12740
rect 41524 12684 42252 12740
rect 42308 12684 42318 12740
rect 26852 12628 26908 12684
rect 20626 12572 20636 12628
rect 20692 12572 22764 12628
rect 22820 12572 26908 12628
rect 28028 12572 37996 12628
rect 38052 12572 38062 12628
rect 19826 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20110 12572
rect 8866 12460 8876 12516
rect 8932 12460 9996 12516
rect 10052 12460 10062 12516
rect 26852 12460 27300 12516
rect 3154 12348 3164 12404
rect 3220 12348 4284 12404
rect 4340 12348 4350 12404
rect 10434 12348 10444 12404
rect 10500 12348 11116 12404
rect 11172 12348 11182 12404
rect 18722 12348 18732 12404
rect 18788 12348 20076 12404
rect 20132 12348 20142 12404
rect 22754 12348 22764 12404
rect 22820 12348 24220 12404
rect 24276 12348 24286 12404
rect 26786 12348 26796 12404
rect 26852 12348 26908 12460
rect 27244 12404 27300 12460
rect 27234 12348 27244 12404
rect 27300 12348 27310 12404
rect 28028 12292 28084 12572
rect 28242 12460 28252 12516
rect 28308 12460 29260 12516
rect 29316 12460 29326 12516
rect 30156 12460 33292 12516
rect 33348 12460 33358 12516
rect 30156 12404 30212 12460
rect 29362 12348 29372 12404
rect 29428 12348 30212 12404
rect 30370 12348 30380 12404
rect 30436 12348 31724 12404
rect 31780 12348 31790 12404
rect 3602 12236 3612 12292
rect 3668 12236 4732 12292
rect 4788 12236 4798 12292
rect 8978 12236 8988 12292
rect 9044 12236 9996 12292
rect 10052 12236 11228 12292
rect 11284 12236 11294 12292
rect 21970 12236 21980 12292
rect 22036 12236 23436 12292
rect 23492 12236 28084 12292
rect 30258 12236 30268 12292
rect 30324 12236 31836 12292
rect 31892 12236 31902 12292
rect 37090 12236 37100 12292
rect 37156 12236 38780 12292
rect 38836 12236 38846 12292
rect 41346 12236 41356 12292
rect 41412 12236 41916 12292
rect 41972 12236 43260 12292
rect 43316 12236 43326 12292
rect 3826 12124 3836 12180
rect 3892 12124 4508 12180
rect 4564 12124 5292 12180
rect 5348 12124 5358 12180
rect 8530 12124 8540 12180
rect 8596 12124 15932 12180
rect 15988 12124 18172 12180
rect 18228 12124 18238 12180
rect 26114 12124 26124 12180
rect 26180 12124 28252 12180
rect 28308 12124 28318 12180
rect 30034 12124 30044 12180
rect 30100 12124 30940 12180
rect 30996 12124 31006 12180
rect 34738 12124 34748 12180
rect 34804 12124 35532 12180
rect 35588 12124 35598 12180
rect 37314 12124 37324 12180
rect 37380 12124 39340 12180
rect 39396 12124 39406 12180
rect 42802 12124 42812 12180
rect 42868 12124 43932 12180
rect 43988 12124 46508 12180
rect 46564 12124 46574 12180
rect 2482 12012 2492 12068
rect 2548 12012 3276 12068
rect 3332 12012 3342 12068
rect 10098 12012 10108 12068
rect 10164 12012 10668 12068
rect 10724 12012 14028 12068
rect 14084 12012 14094 12068
rect 15698 12012 15708 12068
rect 15764 12012 16604 12068
rect 16660 12012 16670 12068
rect 18498 12012 18508 12068
rect 18564 12012 19516 12068
rect 19572 12012 19582 12068
rect 25330 12012 25340 12068
rect 25396 12012 27244 12068
rect 27300 12012 27310 12068
rect 32386 12012 32396 12068
rect 32452 12012 33292 12068
rect 33348 12012 33740 12068
rect 33796 12012 35084 12068
rect 35140 12012 36316 12068
rect 36372 12012 36382 12068
rect 37762 12012 37772 12068
rect 37828 12012 38668 12068
rect 38882 12012 38892 12068
rect 38948 12012 46284 12068
rect 46340 12012 46350 12068
rect 38612 11956 38668 12012
rect 15138 11900 15148 11956
rect 15204 11900 16492 11956
rect 16548 11900 18956 11956
rect 19012 11900 19022 11956
rect 31154 11900 31164 11956
rect 31220 11900 31948 11956
rect 32004 11900 32014 11956
rect 32162 11900 32172 11956
rect 32228 11900 35644 11956
rect 35700 11900 38332 11956
rect 38388 11900 38398 11956
rect 38612 11900 41580 11956
rect 41636 11900 41646 11956
rect 20178 11788 20188 11844
rect 20244 11788 21924 11844
rect 37426 11788 37436 11844
rect 37492 11788 37996 11844
rect 38052 11788 41356 11844
rect 41412 11788 41422 11844
rect 4466 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4750 11788
rect 21868 11732 21924 11788
rect 35186 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35470 11788
rect 7746 11676 7756 11732
rect 7812 11676 8764 11732
rect 8820 11676 9884 11732
rect 9940 11676 13692 11732
rect 13748 11676 13758 11732
rect 21868 11676 35028 11732
rect 36194 11676 36204 11732
rect 36260 11676 36540 11732
rect 36596 11676 40236 11732
rect 40292 11676 40302 11732
rect 34972 11620 35028 11676
rect 3378 11564 3388 11620
rect 3444 11564 4732 11620
rect 4788 11564 4798 11620
rect 9314 11564 9324 11620
rect 9380 11564 11004 11620
rect 11060 11564 11676 11620
rect 11732 11564 11742 11620
rect 31042 11564 31052 11620
rect 31108 11564 32508 11620
rect 32564 11564 32574 11620
rect 34972 11564 36988 11620
rect 37044 11564 40908 11620
rect 40964 11564 41468 11620
rect 41524 11564 42700 11620
rect 42756 11564 42766 11620
rect 4610 11452 4620 11508
rect 4676 11452 5628 11508
rect 5684 11452 5694 11508
rect 8306 11452 8316 11508
rect 8372 11452 10668 11508
rect 10724 11452 10734 11508
rect 12450 11452 12460 11508
rect 12516 11452 13020 11508
rect 13076 11452 13086 11508
rect 28130 11452 28140 11508
rect 28196 11452 29036 11508
rect 29092 11452 29102 11508
rect 35074 11452 35084 11508
rect 35140 11452 36204 11508
rect 36260 11452 36270 11508
rect 38434 11452 38444 11508
rect 38500 11452 39788 11508
rect 39844 11452 40236 11508
rect 40292 11452 40684 11508
rect 40740 11452 40750 11508
rect 46834 11452 46844 11508
rect 46900 11452 47740 11508
rect 47796 11452 47806 11508
rect 9874 11340 9884 11396
rect 9940 11340 10220 11396
rect 10276 11340 11228 11396
rect 11284 11340 12236 11396
rect 12292 11340 12302 11396
rect 12786 11340 12796 11396
rect 12852 11340 13468 11396
rect 13524 11340 13534 11396
rect 19506 11340 19516 11396
rect 19572 11340 20748 11396
rect 20804 11340 28476 11396
rect 28532 11340 29372 11396
rect 29428 11340 29438 11396
rect 30818 11340 30828 11396
rect 30884 11340 31836 11396
rect 31892 11340 31902 11396
rect 38210 11340 38220 11396
rect 38276 11340 39228 11396
rect 39284 11340 39676 11396
rect 39732 11340 39742 11396
rect 43586 11340 43596 11396
rect 43652 11340 44828 11396
rect 44884 11340 45276 11396
rect 45332 11340 45342 11396
rect 5058 11228 5068 11284
rect 5124 11228 5964 11284
rect 6020 11228 6524 11284
rect 6580 11228 12684 11284
rect 12740 11228 12750 11284
rect 29698 11228 29708 11284
rect 29764 11228 30604 11284
rect 30660 11228 30670 11284
rect 36978 11228 36988 11284
rect 37044 11228 37548 11284
rect 37604 11228 37614 11284
rect 38612 11228 39004 11284
rect 39060 11228 39070 11284
rect 41458 11228 41468 11284
rect 41524 11228 42812 11284
rect 42868 11228 42878 11284
rect 38612 11172 38668 11228
rect 6626 11116 6636 11172
rect 6692 11116 7868 11172
rect 7924 11116 7934 11172
rect 8194 11116 8204 11172
rect 8260 11116 9660 11172
rect 9716 11116 9726 11172
rect 12002 11116 12012 11172
rect 12068 11116 12460 11172
rect 12516 11116 12526 11172
rect 30818 11116 30828 11172
rect 30884 11116 33852 11172
rect 33908 11116 33918 11172
rect 35522 11116 35532 11172
rect 35588 11116 35980 11172
rect 36036 11116 38668 11172
rect 25106 11004 25116 11060
rect 25172 11004 30604 11060
rect 30660 11004 30670 11060
rect 19826 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20110 11004
rect 8194 10780 8204 10836
rect 8260 10780 8988 10836
rect 9044 10780 10556 10836
rect 10612 10780 10622 10836
rect 29362 10780 29372 10836
rect 29428 10780 31164 10836
rect 31220 10780 31724 10836
rect 31780 10780 31790 10836
rect 43922 10780 43932 10836
rect 43988 10780 44716 10836
rect 44772 10780 45836 10836
rect 45892 10780 45902 10836
rect 10742 10668 10780 10724
rect 10836 10668 10846 10724
rect 24882 10668 24892 10724
rect 24948 10668 26012 10724
rect 26068 10668 26078 10724
rect 37090 10668 37100 10724
rect 37156 10668 37996 10724
rect 38052 10668 38062 10724
rect 43362 10668 43372 10724
rect 43428 10668 44268 10724
rect 44324 10668 44334 10724
rect 4946 10556 4956 10612
rect 5012 10556 5292 10612
rect 5348 10556 5358 10612
rect 9762 10556 9772 10612
rect 9828 10556 10892 10612
rect 10948 10556 10958 10612
rect 28018 10556 28028 10612
rect 28084 10556 28700 10612
rect 28756 10556 28766 10612
rect 29474 10556 29484 10612
rect 29540 10556 30268 10612
rect 30324 10556 31164 10612
rect 31220 10556 31230 10612
rect 31378 10556 31388 10612
rect 31444 10556 31482 10612
rect 32050 10556 32060 10612
rect 32116 10556 33180 10612
rect 33236 10556 34076 10612
rect 34132 10556 34142 10612
rect 43474 10556 43484 10612
rect 43540 10556 44828 10612
rect 44884 10556 44894 10612
rect 8866 10444 8876 10500
rect 8932 10444 10780 10500
rect 10836 10444 10846 10500
rect 22418 10444 22428 10500
rect 22484 10444 22988 10500
rect 23044 10444 24668 10500
rect 24724 10444 25228 10500
rect 25284 10444 25294 10500
rect 27794 10444 27804 10500
rect 27860 10444 28588 10500
rect 28644 10444 28654 10500
rect 30146 10444 30156 10500
rect 30212 10444 33852 10500
rect 33908 10444 36652 10500
rect 36708 10444 36718 10500
rect 10546 10332 10556 10388
rect 10612 10332 11116 10388
rect 11172 10332 11182 10388
rect 28018 10332 28028 10388
rect 28084 10332 29932 10388
rect 29988 10332 29998 10388
rect 31042 10332 31052 10388
rect 31108 10332 31724 10388
rect 31780 10332 31790 10388
rect 23202 10220 23212 10276
rect 23268 10220 24444 10276
rect 24500 10220 24510 10276
rect 27458 10220 27468 10276
rect 27524 10220 29596 10276
rect 29652 10220 30156 10276
rect 30212 10220 30222 10276
rect 35858 10220 35868 10276
rect 35924 10220 42700 10276
rect 42756 10220 42766 10276
rect 45948 10220 46172 10276
rect 46228 10220 47180 10276
rect 47236 10220 47246 10276
rect 4466 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4750 10220
rect 35186 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35470 10220
rect 45948 10164 46004 10220
rect 15474 10108 15484 10164
rect 15540 10108 16772 10164
rect 39890 10108 39900 10164
rect 39956 10108 42252 10164
rect 42308 10108 42318 10164
rect 45938 10108 45948 10164
rect 46004 10108 46014 10164
rect 46834 10108 46844 10164
rect 46900 10108 48188 10164
rect 48244 10108 48254 10164
rect 16716 10052 16772 10108
rect 5282 9996 5292 10052
rect 5348 9996 6188 10052
rect 6244 9996 6972 10052
rect 7028 9996 7038 10052
rect 16716 9996 17724 10052
rect 17780 9996 17790 10052
rect 27682 9996 27692 10052
rect 27748 9996 30156 10052
rect 30212 9996 30222 10052
rect 30818 9996 30828 10052
rect 30884 9996 33740 10052
rect 33796 9996 36092 10052
rect 36148 9996 36158 10052
rect 38098 9996 38108 10052
rect 38164 9996 43484 10052
rect 43540 9996 43550 10052
rect 1698 9884 1708 9940
rect 1764 9884 5404 9940
rect 5460 9884 6076 9940
rect 6132 9884 6142 9940
rect 11890 9884 11900 9940
rect 11956 9884 12908 9940
rect 12964 9884 20188 9940
rect 20244 9884 20254 9940
rect 25666 9884 25676 9940
rect 25732 9884 26908 9940
rect 9986 9772 9996 9828
rect 10052 9772 10668 9828
rect 10724 9772 11452 9828
rect 11508 9772 11518 9828
rect 11666 9660 11676 9716
rect 11732 9660 17612 9716
rect 17668 9660 17678 9716
rect 21186 9660 21196 9716
rect 21252 9660 26236 9716
rect 26292 9660 26302 9716
rect 26852 9604 26908 9884
rect 38612 9884 38892 9940
rect 38948 9884 38958 9940
rect 40674 9884 40684 9940
rect 40740 9884 41916 9940
rect 41972 9884 41982 9940
rect 28578 9772 28588 9828
rect 28644 9772 29148 9828
rect 29204 9772 30716 9828
rect 30772 9772 30782 9828
rect 38612 9716 38668 9884
rect 30146 9660 30156 9716
rect 30212 9660 34636 9716
rect 34692 9660 36876 9716
rect 36932 9660 38668 9716
rect 5506 9548 5516 9604
rect 5572 9548 6524 9604
rect 6580 9548 6590 9604
rect 7074 9548 7084 9604
rect 7140 9548 7756 9604
rect 7812 9548 8988 9604
rect 9044 9548 9054 9604
rect 12674 9548 12684 9604
rect 12740 9548 13692 9604
rect 13748 9548 13758 9604
rect 16930 9548 16940 9604
rect 16996 9548 17948 9604
rect 18004 9548 19628 9604
rect 19684 9548 20188 9604
rect 20244 9548 21420 9604
rect 21476 9548 22092 9604
rect 22148 9548 22158 9604
rect 26852 9548 27580 9604
rect 27636 9548 29260 9604
rect 29316 9548 29326 9604
rect 45042 9548 45052 9604
rect 45108 9548 46956 9604
rect 47012 9548 47022 9604
rect 47170 9548 47180 9604
rect 47236 9548 47246 9604
rect 47180 9492 47236 9548
rect 49200 9492 50000 9520
rect 12226 9436 12236 9492
rect 12292 9436 12572 9492
rect 12628 9436 12638 9492
rect 47180 9436 50000 9492
rect 19826 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20110 9436
rect 49200 9408 50000 9436
rect 14914 9324 14924 9380
rect 14980 9324 15932 9380
rect 15988 9324 19348 9380
rect 33282 9324 33292 9380
rect 33348 9324 35196 9380
rect 35252 9324 35262 9380
rect 19292 9268 19348 9324
rect 2482 9212 2492 9268
rect 2548 9212 3836 9268
rect 3892 9212 3902 9268
rect 4050 9212 4060 9268
rect 4116 9212 4956 9268
rect 5012 9212 5022 9268
rect 14354 9212 14364 9268
rect 14420 9212 15036 9268
rect 15092 9212 15102 9268
rect 16034 9212 16044 9268
rect 16100 9212 16716 9268
rect 16772 9212 16782 9268
rect 17714 9212 17724 9268
rect 17780 9212 18844 9268
rect 18900 9212 18910 9268
rect 19292 9212 34300 9268
rect 34356 9212 34366 9268
rect 38770 9212 38780 9268
rect 38836 9212 41132 9268
rect 41188 9212 41916 9268
rect 41972 9212 41982 9268
rect 44146 9212 44156 9268
rect 44212 9212 44940 9268
rect 44996 9212 45006 9268
rect 4610 9100 4620 9156
rect 4676 9100 5180 9156
rect 5236 9100 5740 9156
rect 5796 9100 5806 9156
rect 14466 9100 14476 9156
rect 14532 9100 14812 9156
rect 14868 9100 18396 9156
rect 18452 9100 18462 9156
rect 34300 9044 34356 9212
rect 37314 9100 37324 9156
rect 37380 9100 44716 9156
rect 44772 9100 44782 9156
rect 3938 8988 3948 9044
rect 4004 8988 4956 9044
rect 5012 8988 7980 9044
rect 8036 8988 10668 9044
rect 10724 8988 10892 9044
rect 10948 8988 10958 9044
rect 15698 8988 15708 9044
rect 15764 8988 16492 9044
rect 16548 8988 16558 9044
rect 20178 8988 20188 9044
rect 20244 8988 21196 9044
rect 21252 8988 21644 9044
rect 21700 8988 21710 9044
rect 34300 8988 41468 9044
rect 41524 8988 41534 9044
rect 45378 8988 45388 9044
rect 45444 8988 45836 9044
rect 45892 8988 47964 9044
rect 48020 8988 48030 9044
rect 9986 8876 9996 8932
rect 10052 8876 10444 8932
rect 10500 8876 11900 8932
rect 11956 8876 11966 8932
rect 29922 8876 29932 8932
rect 29988 8876 34524 8932
rect 34580 8876 34590 8932
rect 34748 8876 39004 8932
rect 39060 8876 39900 8932
rect 39956 8876 39966 8932
rect 40338 8876 40348 8932
rect 40404 8876 41356 8932
rect 41412 8876 41422 8932
rect 42802 8876 42812 8932
rect 42868 8876 47068 8932
rect 47124 8876 47134 8932
rect 34748 8820 34804 8876
rect 49200 8820 50000 8848
rect 4386 8764 4396 8820
rect 4452 8764 5236 8820
rect 12562 8764 12572 8820
rect 12628 8764 16268 8820
rect 16324 8764 17948 8820
rect 18004 8764 18014 8820
rect 32274 8764 32284 8820
rect 32340 8764 32508 8820
rect 32564 8764 34804 8820
rect 35186 8764 35196 8820
rect 35252 8764 35588 8820
rect 39554 8764 39564 8820
rect 39620 8764 41692 8820
rect 41748 8764 43708 8820
rect 43764 8764 43774 8820
rect 47954 8764 47964 8820
rect 48020 8764 50000 8820
rect 4466 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4750 8652
rect 5180 8596 5236 8764
rect 35532 8708 35588 8764
rect 49200 8736 50000 8764
rect 8978 8652 8988 8708
rect 9044 8652 28252 8708
rect 28308 8652 28700 8708
rect 28756 8652 28766 8708
rect 35532 8652 35644 8708
rect 35700 8652 35710 8708
rect 40002 8652 40012 8708
rect 40068 8652 43148 8708
rect 43204 8652 43214 8708
rect 35186 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35470 8652
rect 5170 8540 5180 8596
rect 5236 8540 15148 8596
rect 15204 8540 15214 8596
rect 16482 8540 16492 8596
rect 16548 8540 27468 8596
rect 27524 8540 27534 8596
rect 38434 8540 38444 8596
rect 38500 8540 44156 8596
rect 44212 8540 44222 8596
rect 45154 8540 45164 8596
rect 45220 8540 47404 8596
rect 47460 8540 47470 8596
rect 10742 8428 10780 8484
rect 10836 8428 10846 8484
rect 16492 8372 16548 8540
rect 21522 8428 21532 8484
rect 21588 8428 22092 8484
rect 22148 8428 22428 8484
rect 22484 8428 22494 8484
rect 28476 8428 29932 8484
rect 29988 8428 29998 8484
rect 31266 8428 31276 8484
rect 31332 8428 31342 8484
rect 32498 8428 32508 8484
rect 32564 8428 32574 8484
rect 42466 8428 42476 8484
rect 42532 8428 44940 8484
rect 44996 8428 45006 8484
rect 28476 8372 28532 8428
rect 31276 8372 31332 8428
rect 32508 8372 32564 8428
rect 3332 8316 5852 8372
rect 5908 8316 7084 8372
rect 7140 8316 7150 8372
rect 13010 8316 13020 8372
rect 13076 8316 13468 8372
rect 13524 8316 16548 8372
rect 17826 8316 17836 8372
rect 17892 8316 17902 8372
rect 27906 8316 27916 8372
rect 27972 8316 28532 8372
rect 28690 8316 28700 8372
rect 28756 8316 33964 8372
rect 34020 8316 35980 8372
rect 36036 8316 36046 8372
rect 36530 8316 36540 8372
rect 36596 8316 40460 8372
rect 40516 8316 40526 8372
rect 43250 8316 43260 8372
rect 43316 8316 43326 8372
rect 44146 8316 44156 8372
rect 44212 8316 45388 8372
rect 45444 8316 45454 8372
rect 1810 8204 1820 8260
rect 1876 8204 3276 8260
rect 3332 8204 3388 8316
rect 17836 8260 17892 8316
rect 43260 8260 43316 8316
rect 9426 8204 9436 8260
rect 9492 8204 10780 8260
rect 10836 8204 12908 8260
rect 12964 8204 12974 8260
rect 13570 8204 13580 8260
rect 13636 8204 16268 8260
rect 16324 8204 17892 8260
rect 21970 8204 21980 8260
rect 22036 8204 30044 8260
rect 30100 8204 30110 8260
rect 31378 8204 31388 8260
rect 31444 8204 31612 8260
rect 31668 8204 31678 8260
rect 34514 8204 34524 8260
rect 34580 8204 38668 8260
rect 43260 8204 46620 8260
rect 46676 8204 46686 8260
rect 38612 8148 38668 8204
rect 49200 8148 50000 8176
rect 5506 8092 5516 8148
rect 5572 8092 6636 8148
rect 6692 8092 14028 8148
rect 14084 8092 14094 8148
rect 15586 8092 15596 8148
rect 15652 8092 16604 8148
rect 16660 8092 17388 8148
rect 17444 8092 17454 8148
rect 18722 8092 18732 8148
rect 18788 8092 27132 8148
rect 27188 8092 27580 8148
rect 27636 8092 29372 8148
rect 29428 8092 29438 8148
rect 35858 8092 35868 8148
rect 35924 8092 37324 8148
rect 37380 8092 38220 8148
rect 38276 8092 38286 8148
rect 38612 8092 41748 8148
rect 41906 8092 41916 8148
rect 41972 8092 44156 8148
rect 44212 8092 44222 8148
rect 47954 8092 47964 8148
rect 48020 8092 50000 8148
rect 8978 7980 8988 8036
rect 9044 7980 9772 8036
rect 9828 7980 9838 8036
rect 11890 7980 11900 8036
rect 11956 7980 18844 8036
rect 18900 7980 18910 8036
rect 14578 7868 14588 7924
rect 14644 7868 15596 7924
rect 15652 7868 15662 7924
rect 19404 7812 19460 8092
rect 41692 8036 41748 8092
rect 49200 8064 50000 8092
rect 26002 7980 26012 8036
rect 26068 7980 26908 8036
rect 29810 7980 29820 8036
rect 29876 7980 30716 8036
rect 30772 7980 30782 8036
rect 32582 7980 32620 8036
rect 32676 7980 32686 8036
rect 38098 7980 38108 8036
rect 38164 7980 39452 8036
rect 39508 7980 39518 8036
rect 41692 7980 43932 8036
rect 43988 7980 43998 8036
rect 44258 7980 44268 8036
rect 44324 7980 48188 8036
rect 48244 7980 48254 8036
rect 26852 7924 26908 7980
rect 26852 7868 27468 7924
rect 27524 7868 29596 7924
rect 29652 7868 30044 7924
rect 30100 7868 30110 7924
rect 31042 7868 31052 7924
rect 31108 7868 32732 7924
rect 32788 7868 41916 7924
rect 41972 7868 41982 7924
rect 42130 7868 42140 7924
rect 42196 7868 43708 7924
rect 43764 7868 43774 7924
rect 19826 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20110 7868
rect 13122 7756 13132 7812
rect 13188 7756 16828 7812
rect 16884 7756 17500 7812
rect 17556 7756 17566 7812
rect 19394 7756 19404 7812
rect 19460 7756 19470 7812
rect 11442 7644 11452 7700
rect 11508 7644 14252 7700
rect 14308 7644 14924 7700
rect 14980 7644 14990 7700
rect 17042 7644 17052 7700
rect 17108 7644 18396 7700
rect 18452 7644 26012 7700
rect 26068 7644 26078 7700
rect 35970 7644 35980 7700
rect 36036 7644 37212 7700
rect 37268 7644 38108 7700
rect 38164 7644 38174 7700
rect 42354 7644 42364 7700
rect 42420 7644 42812 7700
rect 42868 7644 42878 7700
rect 11554 7532 11564 7588
rect 11620 7532 12572 7588
rect 12628 7532 12638 7588
rect 19058 7532 19068 7588
rect 19124 7532 19740 7588
rect 19796 7532 21420 7588
rect 21476 7532 21486 7588
rect 25442 7532 25452 7588
rect 25508 7532 27132 7588
rect 27188 7532 31388 7588
rect 31444 7532 31454 7588
rect 38770 7532 38780 7588
rect 38836 7532 39900 7588
rect 39956 7532 39966 7588
rect 42690 7532 42700 7588
rect 42756 7532 43820 7588
rect 43876 7532 43886 7588
rect 49200 7476 50000 7504
rect 28914 7420 28924 7476
rect 28980 7420 29820 7476
rect 29876 7420 29886 7476
rect 33394 7420 33404 7476
rect 33460 7420 35420 7476
rect 35476 7420 35486 7476
rect 40226 7420 40236 7476
rect 40292 7420 46396 7476
rect 46452 7420 46462 7476
rect 47954 7420 47964 7476
rect 48020 7420 50000 7476
rect 49200 7392 50000 7420
rect 17938 7308 17948 7364
rect 18004 7308 18956 7364
rect 19012 7308 19022 7364
rect 23426 7308 23436 7364
rect 23492 7308 24444 7364
rect 24500 7308 24510 7364
rect 40338 7308 40348 7364
rect 40404 7308 42700 7364
rect 42756 7308 42766 7364
rect 42914 7308 42924 7364
rect 42980 7308 43484 7364
rect 43540 7308 43550 7364
rect 41010 7196 41020 7252
rect 41076 7196 45052 7252
rect 45108 7196 45118 7252
rect 5282 7084 5292 7140
rect 5348 7084 6524 7140
rect 6580 7084 8988 7140
rect 9044 7084 9054 7140
rect 38994 7084 39004 7140
rect 39060 7084 41244 7140
rect 41300 7084 41310 7140
rect 4466 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4750 7084
rect 35186 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35470 7084
rect 9090 6972 9100 7028
rect 9156 6972 12572 7028
rect 12628 6972 12638 7028
rect 28140 6972 30380 7028
rect 30436 6972 30446 7028
rect 40198 6972 40236 7028
rect 40292 6972 40302 7028
rect 9762 6860 9772 6916
rect 9828 6860 10332 6916
rect 10388 6860 10398 6916
rect 11666 6860 11676 6916
rect 11732 6860 12124 6916
rect 12180 6860 12190 6916
rect 12338 6860 12348 6916
rect 12404 6860 13020 6916
rect 13076 6860 13086 6916
rect 18396 6860 27916 6916
rect 27972 6860 27982 6916
rect 9874 6748 9884 6804
rect 9940 6748 10668 6804
rect 10724 6748 11452 6804
rect 11508 6748 13580 6804
rect 13636 6748 13646 6804
rect 12898 6636 12908 6692
rect 12964 6636 13692 6692
rect 13748 6636 13758 6692
rect 18396 6580 18452 6860
rect 28140 6804 28196 6972
rect 32274 6860 32284 6916
rect 32340 6860 33068 6916
rect 33124 6860 33134 6916
rect 35298 6860 35308 6916
rect 35364 6860 36428 6916
rect 36484 6860 36494 6916
rect 39890 6860 39900 6916
rect 39956 6860 41132 6916
rect 41188 6860 41198 6916
rect 43810 6860 43820 6916
rect 43876 6860 44156 6916
rect 44212 6860 44222 6916
rect 22876 6748 28196 6804
rect 29484 6748 29988 6804
rect 32162 6748 32172 6804
rect 32228 6748 32956 6804
rect 33012 6748 33022 6804
rect 35718 6748 35756 6804
rect 35812 6748 35822 6804
rect 36988 6748 37660 6804
rect 37716 6748 37884 6804
rect 37940 6748 39340 6804
rect 39396 6748 39406 6804
rect 39554 6748 39564 6804
rect 39620 6748 41468 6804
rect 41524 6748 43764 6804
rect 22876 6692 22932 6748
rect 29484 6692 29540 6748
rect 29932 6692 29988 6748
rect 36988 6692 37044 6748
rect 21970 6636 21980 6692
rect 22036 6636 22932 6692
rect 23090 6636 23100 6692
rect 23156 6636 29540 6692
rect 29698 6636 29708 6692
rect 29764 6636 29774 6692
rect 29932 6636 34468 6692
rect 34626 6636 34636 6692
rect 34692 6636 36652 6692
rect 36708 6636 36718 6692
rect 36876 6636 37044 6692
rect 37986 6636 37996 6692
rect 38052 6636 38556 6692
rect 38612 6636 38622 6692
rect 8082 6524 8092 6580
rect 8148 6524 11004 6580
rect 11060 6524 11070 6580
rect 12562 6524 12572 6580
rect 12628 6524 16268 6580
rect 16324 6524 18452 6580
rect 23650 6524 23660 6580
rect 23716 6524 24332 6580
rect 24388 6524 24398 6580
rect 29708 6468 29764 6636
rect 34412 6580 34468 6636
rect 36876 6580 36932 6636
rect 43708 6580 43764 6748
rect 31714 6524 31724 6580
rect 31780 6524 33740 6580
rect 33796 6524 33806 6580
rect 34412 6524 36932 6580
rect 37090 6524 37100 6580
rect 37156 6524 37772 6580
rect 37828 6524 37838 6580
rect 39442 6524 39452 6580
rect 39508 6524 40124 6580
rect 40180 6524 40572 6580
rect 40628 6524 40638 6580
rect 43708 6524 44492 6580
rect 44548 6524 45276 6580
rect 45332 6524 45342 6580
rect 12674 6412 12684 6468
rect 12740 6412 13132 6468
rect 13188 6412 13198 6468
rect 13682 6412 13692 6468
rect 13748 6412 14700 6468
rect 14756 6412 14766 6468
rect 17714 6412 17724 6468
rect 17780 6412 22596 6468
rect 22978 6412 22988 6468
rect 23044 6412 23996 6468
rect 24052 6412 24062 6468
rect 24668 6412 26348 6468
rect 26404 6412 26684 6468
rect 26740 6412 29764 6468
rect 34850 6412 34860 6468
rect 34916 6412 34926 6468
rect 36642 6412 36652 6468
rect 36708 6412 37996 6468
rect 38052 6412 38062 6468
rect 40226 6412 40236 6468
rect 40292 6412 43820 6468
rect 43876 6412 43886 6468
rect 22540 6356 22596 6412
rect 8642 6300 8652 6356
rect 8708 6300 9772 6356
rect 9828 6300 17556 6356
rect 21298 6300 21308 6356
rect 21364 6300 22204 6356
rect 22260 6300 22270 6356
rect 22540 6300 22820 6356
rect 6514 6188 6524 6244
rect 6580 6188 7644 6244
rect 7700 6188 11452 6244
rect 11508 6188 15148 6244
rect 15092 6132 15148 6188
rect 6290 6076 6300 6132
rect 6356 6076 7420 6132
rect 7476 6076 10108 6132
rect 10164 6076 10174 6132
rect 12450 6076 12460 6132
rect 12516 6076 12908 6132
rect 12964 6076 12974 6132
rect 13234 6076 13244 6132
rect 13300 6076 14700 6132
rect 14756 6076 14766 6132
rect 15092 6076 15484 6132
rect 15540 6076 15550 6132
rect 17500 6020 17556 6300
rect 19826 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20110 6300
rect 22204 6132 22260 6300
rect 22764 6244 22820 6300
rect 22754 6188 22764 6244
rect 22820 6188 22830 6244
rect 24668 6132 24724 6412
rect 34860 6356 34916 6412
rect 29474 6300 29484 6356
rect 29540 6300 30716 6356
rect 30772 6300 32060 6356
rect 32116 6300 32126 6356
rect 34860 6300 38668 6356
rect 39778 6300 39788 6356
rect 39844 6300 41356 6356
rect 41412 6300 41422 6356
rect 42466 6300 42476 6356
rect 42532 6300 44828 6356
rect 44884 6300 44894 6356
rect 38612 6244 38668 6300
rect 25666 6188 25676 6244
rect 25732 6188 26572 6244
rect 26628 6188 35196 6244
rect 35252 6188 35262 6244
rect 38612 6188 44716 6244
rect 44772 6188 44782 6244
rect 22204 6076 24724 6132
rect 29698 6076 29708 6132
rect 29764 6076 33180 6132
rect 33236 6076 35756 6132
rect 35812 6076 35822 6132
rect 36754 6076 36764 6132
rect 36820 6076 37324 6132
rect 37380 6076 39788 6132
rect 39844 6076 39854 6132
rect 10770 5964 10780 6020
rect 10836 5964 11228 6020
rect 11284 5964 11900 6020
rect 11956 5964 13132 6020
rect 13188 5964 13198 6020
rect 17490 5964 17500 6020
rect 17556 5964 20804 6020
rect 21410 5964 21420 6020
rect 21476 5964 23100 6020
rect 23156 5964 23166 6020
rect 23314 5964 23324 6020
rect 23380 5964 28084 6020
rect 28690 5964 28700 6020
rect 28756 5964 30940 6020
rect 30996 5964 31164 6020
rect 31220 5964 31230 6020
rect 31378 5964 31388 6020
rect 31444 5964 32060 6020
rect 32116 5964 32126 6020
rect 38882 5964 38892 6020
rect 38948 5964 47292 6020
rect 47348 5964 47358 6020
rect 20748 5908 20804 5964
rect 28028 5908 28084 5964
rect 31388 5908 31444 5964
rect 7074 5852 7084 5908
rect 7140 5852 8540 5908
rect 8596 5852 8606 5908
rect 8754 5852 8764 5908
rect 8820 5852 9996 5908
rect 10052 5852 10444 5908
rect 10500 5852 11116 5908
rect 11172 5852 11182 5908
rect 19842 5852 19852 5908
rect 19908 5852 20524 5908
rect 20580 5852 20590 5908
rect 20748 5852 21980 5908
rect 22036 5852 22046 5908
rect 22754 5852 22764 5908
rect 22820 5852 26236 5908
rect 26292 5852 26302 5908
rect 26786 5852 26796 5908
rect 26852 5852 27580 5908
rect 27636 5852 27646 5908
rect 28018 5852 28028 5908
rect 28084 5852 28588 5908
rect 28644 5852 31444 5908
rect 33842 5852 33852 5908
rect 33908 5852 33918 5908
rect 34514 5852 34524 5908
rect 34580 5852 35308 5908
rect 35364 5852 35374 5908
rect 39330 5852 39340 5908
rect 39396 5852 39900 5908
rect 39956 5852 39966 5908
rect 40114 5852 40124 5908
rect 40180 5852 42252 5908
rect 42308 5852 42318 5908
rect 33852 5796 33908 5852
rect 6738 5740 6748 5796
rect 6804 5740 7420 5796
rect 7476 5740 7486 5796
rect 8866 5740 8876 5796
rect 8932 5740 12236 5796
rect 12292 5740 12684 5796
rect 12740 5740 12750 5796
rect 13906 5740 13916 5796
rect 13972 5740 14924 5796
rect 14980 5740 16604 5796
rect 16660 5740 19572 5796
rect 20738 5740 20748 5796
rect 20804 5740 21532 5796
rect 21588 5740 23548 5796
rect 23604 5740 24444 5796
rect 24500 5740 24780 5796
rect 24836 5740 26908 5796
rect 26964 5740 26974 5796
rect 29036 5740 29372 5796
rect 29428 5740 31724 5796
rect 31780 5740 31790 5796
rect 32396 5740 33908 5796
rect 38546 5740 38556 5796
rect 38612 5740 41916 5796
rect 41972 5740 41982 5796
rect 42802 5740 42812 5796
rect 42868 5740 44044 5796
rect 44100 5740 46732 5796
rect 46788 5740 46798 5796
rect 19516 5684 19572 5740
rect 29036 5684 29092 5740
rect 11890 5628 11900 5684
rect 11956 5628 13468 5684
rect 13524 5628 13534 5684
rect 16930 5628 16940 5684
rect 16996 5628 18396 5684
rect 18452 5628 18462 5684
rect 19506 5628 19516 5684
rect 19572 5628 23324 5684
rect 23380 5628 23390 5684
rect 24210 5628 24220 5684
rect 24276 5628 25228 5684
rect 25284 5628 25294 5684
rect 26226 5628 26236 5684
rect 26292 5628 29092 5684
rect 29250 5628 29260 5684
rect 29316 5628 30380 5684
rect 30436 5628 30446 5684
rect 32396 5572 32452 5740
rect 32610 5628 32620 5684
rect 32676 5628 34860 5684
rect 34916 5628 34926 5684
rect 36642 5628 36652 5684
rect 36708 5628 38668 5684
rect 38724 5628 38734 5684
rect 40114 5628 40124 5684
rect 40180 5628 40236 5684
rect 40292 5628 40302 5684
rect 41010 5628 41020 5684
rect 41076 5628 44828 5684
rect 44884 5628 44894 5684
rect 16828 5516 22316 5572
rect 22372 5516 23100 5572
rect 23156 5516 23166 5572
rect 25442 5516 25452 5572
rect 25508 5516 25676 5572
rect 25732 5516 25742 5572
rect 26674 5516 26684 5572
rect 26740 5516 27020 5572
rect 27076 5516 27086 5572
rect 31826 5516 31836 5572
rect 31892 5516 32452 5572
rect 36082 5516 36092 5572
rect 36148 5516 47068 5572
rect 47124 5516 47134 5572
rect 0 5460 800 5488
rect 4466 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4750 5516
rect 0 5404 1708 5460
rect 1764 5404 1774 5460
rect 0 5376 800 5404
rect 16828 5348 16884 5516
rect 35186 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35470 5516
rect 29138 5404 29148 5460
rect 29204 5404 29820 5460
rect 29876 5404 29886 5460
rect 43810 5404 43820 5460
rect 43876 5404 44828 5460
rect 44884 5404 47852 5460
rect 47908 5404 47918 5460
rect 6738 5292 6748 5348
rect 6804 5292 7756 5348
rect 7812 5292 11004 5348
rect 11060 5292 13580 5348
rect 13636 5292 13804 5348
rect 13860 5292 13870 5348
rect 15026 5292 15036 5348
rect 15092 5292 16884 5348
rect 17714 5292 17724 5348
rect 17780 5292 19068 5348
rect 19124 5292 19134 5348
rect 21522 5292 21532 5348
rect 21588 5292 23772 5348
rect 23828 5292 23838 5348
rect 24770 5292 24780 5348
rect 24836 5292 28140 5348
rect 28196 5292 28206 5348
rect 33842 5292 33852 5348
rect 33908 5292 35644 5348
rect 35700 5292 35710 5348
rect 36530 5292 36540 5348
rect 36596 5292 37436 5348
rect 37492 5292 37502 5348
rect 37650 5292 37660 5348
rect 37716 5292 37726 5348
rect 39890 5292 39900 5348
rect 39956 5292 42028 5348
rect 42084 5292 42094 5348
rect 44706 5292 44716 5348
rect 44772 5292 47964 5348
rect 48020 5292 48030 5348
rect 8530 5180 8540 5236
rect 8596 5180 11788 5236
rect 11844 5180 11854 5236
rect 14466 5180 14476 5236
rect 14532 5180 15148 5236
rect 15204 5180 15214 5236
rect 16828 5124 16884 5292
rect 37660 5236 37716 5292
rect 17042 5180 17052 5236
rect 17108 5180 18732 5236
rect 18788 5180 20748 5236
rect 20804 5180 20814 5236
rect 20962 5180 20972 5236
rect 21028 5180 22764 5236
rect 22820 5180 22830 5236
rect 24882 5180 24892 5236
rect 24948 5180 26796 5236
rect 26852 5180 26862 5236
rect 35308 5180 37716 5236
rect 40450 5180 40460 5236
rect 40516 5180 43260 5236
rect 43316 5180 43326 5236
rect 44258 5180 44268 5236
rect 44324 5180 47740 5236
rect 47796 5180 47806 5236
rect 6738 5068 6748 5124
rect 6804 5068 8204 5124
rect 8260 5068 8270 5124
rect 8418 5068 8428 5124
rect 8484 5068 12572 5124
rect 12628 5068 12638 5124
rect 16828 5068 17836 5124
rect 17892 5068 17902 5124
rect 18050 5068 18060 5124
rect 18116 5068 18508 5124
rect 18564 5068 18574 5124
rect 18834 5068 18844 5124
rect 18900 5068 20412 5124
rect 20468 5068 20478 5124
rect 22418 5068 22428 5124
rect 22484 5068 23436 5124
rect 23492 5068 23502 5124
rect 24658 5068 24668 5124
rect 24724 5068 26684 5124
rect 26740 5068 26750 5124
rect 26852 5068 27804 5124
rect 27860 5068 29484 5124
rect 29540 5068 29550 5124
rect 31602 5068 31612 5124
rect 31668 5068 34692 5124
rect 19740 5012 19796 5068
rect 26852 5012 26908 5068
rect 34636 5012 34692 5068
rect 35308 5012 35364 5180
rect 35858 5068 35868 5124
rect 35924 5068 38108 5124
rect 38164 5068 38174 5124
rect 40338 5068 40348 5124
rect 40404 5068 41580 5124
rect 41636 5068 41646 5124
rect 42914 5068 42924 5124
rect 42980 5068 43932 5124
rect 43988 5068 43998 5124
rect 44930 5068 44940 5124
rect 44996 5068 46508 5124
rect 46564 5068 46574 5124
rect 4050 4956 4060 5012
rect 4116 4956 5068 5012
rect 5124 4956 5134 5012
rect 10882 4956 10892 5012
rect 10948 4956 11788 5012
rect 11844 4956 12684 5012
rect 12740 4956 13916 5012
rect 13972 4956 13982 5012
rect 19730 4956 19740 5012
rect 19796 4956 19806 5012
rect 22316 4956 22876 5012
rect 22932 4956 25676 5012
rect 25732 4956 26908 5012
rect 30370 4956 30380 5012
rect 30436 4956 33068 5012
rect 33124 4956 33134 5012
rect 34626 4956 34636 5012
rect 34692 4956 34702 5012
rect 35298 4956 35308 5012
rect 35364 4956 35374 5012
rect 38770 4956 38780 5012
rect 38836 4956 42700 5012
rect 42756 4956 44268 5012
rect 44324 4956 44334 5012
rect 46386 4956 46396 5012
rect 46452 4956 47404 5012
rect 47460 4956 47470 5012
rect 5068 4900 5124 4956
rect 22316 4900 22372 4956
rect 1698 4844 1708 4900
rect 1764 4844 1774 4900
rect 5068 4844 6300 4900
rect 6356 4844 6366 4900
rect 8866 4844 8876 4900
rect 8932 4844 14140 4900
rect 14196 4844 14206 4900
rect 22306 4844 22316 4900
rect 22372 4844 22382 4900
rect 25778 4844 25788 4900
rect 25844 4844 31276 4900
rect 31332 4844 31836 4900
rect 31892 4844 31902 4900
rect 41682 4844 41692 4900
rect 41748 4844 45836 4900
rect 45892 4844 45902 4900
rect 0 4788 800 4816
rect 1708 4788 1764 4844
rect 49200 4788 50000 4816
rect 0 4732 1764 4788
rect 11554 4732 11564 4788
rect 11620 4732 12908 4788
rect 12964 4732 12974 4788
rect 23986 4732 23996 4788
rect 24052 4732 24556 4788
rect 24612 4732 31500 4788
rect 31556 4732 31566 4788
rect 31714 4732 31724 4788
rect 31780 4732 34972 4788
rect 35028 4732 35756 4788
rect 35812 4732 35822 4788
rect 44594 4732 44604 4788
rect 44660 4732 50000 4788
rect 0 4704 800 4732
rect 19826 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20110 4732
rect 31500 4676 31556 4732
rect 49200 4704 50000 4732
rect 22194 4620 22204 4676
rect 22260 4620 25788 4676
rect 25844 4620 25854 4676
rect 31500 4620 34188 4676
rect 34244 4620 35196 4676
rect 35252 4620 35262 4676
rect 7522 4508 7532 4564
rect 7588 4508 9772 4564
rect 9828 4508 9838 4564
rect 15474 4508 15484 4564
rect 15540 4508 17948 4564
rect 18004 4508 18014 4564
rect 20178 4508 20188 4564
rect 20244 4508 22092 4564
rect 22148 4508 22158 4564
rect 30258 4508 30268 4564
rect 30324 4508 34076 4564
rect 34132 4508 36092 4564
rect 36148 4508 36158 4564
rect 40226 4508 40236 4564
rect 40292 4508 42140 4564
rect 42196 4508 43708 4564
rect 43764 4508 43932 4564
rect 43988 4508 43998 4564
rect 46610 4508 46620 4564
rect 46676 4508 47628 4564
rect 47684 4508 47694 4564
rect 6514 4396 6524 4452
rect 6580 4396 10780 4452
rect 10836 4396 10846 4452
rect 22754 4396 22764 4452
rect 22820 4396 23884 4452
rect 23940 4396 23950 4452
rect 32386 4396 32396 4452
rect 32452 4396 33964 4452
rect 34020 4396 35980 4452
rect 36036 4396 36046 4452
rect 43026 4396 43036 4452
rect 43092 4396 45164 4452
rect 45220 4396 45230 4452
rect 5842 4284 5852 4340
rect 5908 4284 7084 4340
rect 7140 4284 7150 4340
rect 7410 4284 7420 4340
rect 7476 4284 7486 4340
rect 41794 4284 41804 4340
rect 41860 4284 43932 4340
rect 43988 4284 47852 4340
rect 47908 4284 47918 4340
rect 7420 4228 7476 4284
rect 6178 4172 6188 4228
rect 6244 4172 7476 4228
rect 8978 4172 8988 4228
rect 9044 4172 13692 4228
rect 13748 4172 13758 4228
rect 14242 4172 14252 4228
rect 14308 4172 15820 4228
rect 15876 4172 16716 4228
rect 16772 4172 16782 4228
rect 24546 4172 24556 4228
rect 24612 4172 25228 4228
rect 25284 4172 25294 4228
rect 38322 4172 38332 4228
rect 38388 4172 42028 4228
rect 42084 4172 42094 4228
rect 0 4116 800 4144
rect 49200 4116 50000 4144
rect 0 4060 1708 4116
rect 1764 4060 1774 4116
rect 5506 4060 5516 4116
rect 5572 4060 6748 4116
rect 6804 4060 6814 4116
rect 9426 4060 9436 4116
rect 9492 4060 10668 4116
rect 10724 4060 10734 4116
rect 46946 4060 46956 4116
rect 47012 4060 50000 4116
rect 0 4032 800 4060
rect 49200 4032 50000 4060
rect 4466 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4750 3948
rect 35186 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35470 3948
rect 5058 3836 5068 3892
rect 5124 3836 9548 3892
rect 9604 3836 10780 3892
rect 10836 3836 10846 3892
rect 7970 3724 7980 3780
rect 8036 3724 9324 3780
rect 9380 3724 9390 3780
rect 29586 3724 29596 3780
rect 29652 3724 30940 3780
rect 30996 3724 31006 3780
rect 43138 3724 43148 3780
rect 43204 3724 47628 3780
rect 47684 3724 47694 3780
rect 4610 3612 4620 3668
rect 4676 3612 8428 3668
rect 8484 3612 10108 3668
rect 10164 3612 10174 3668
rect 17490 3612 17500 3668
rect 17556 3612 18620 3668
rect 18676 3612 18686 3668
rect 20850 3612 20860 3668
rect 20916 3612 22092 3668
rect 22148 3612 22158 3668
rect 26226 3612 26236 3668
rect 26292 3612 29372 3668
rect 29428 3612 29438 3668
rect 32946 3612 32956 3668
rect 33012 3612 33852 3668
rect 33908 3612 33918 3668
rect 37650 3612 37660 3668
rect 37716 3612 40796 3668
rect 40852 3612 40862 3668
rect 42354 3612 42364 3668
rect 42420 3612 46732 3668
rect 46788 3612 46798 3668
rect 4162 3500 4172 3556
rect 4228 3500 7420 3556
rect 7476 3500 7868 3556
rect 7924 3500 7934 3556
rect 12114 3500 12124 3556
rect 12180 3500 13468 3556
rect 13524 3500 14140 3556
rect 14196 3500 14206 3556
rect 20290 3500 20300 3556
rect 20356 3500 21084 3556
rect 21140 3500 21150 3556
rect 25890 3500 25900 3556
rect 25956 3500 28588 3556
rect 28644 3500 28654 3556
rect 30258 3500 30268 3556
rect 30324 3500 32284 3556
rect 32340 3500 32620 3556
rect 32676 3500 32686 3556
rect 33618 3500 33628 3556
rect 33684 3500 35084 3556
rect 35140 3500 36204 3556
rect 36260 3500 36270 3556
rect 41234 3500 41244 3556
rect 41300 3500 43708 3556
rect 43764 3500 43774 3556
rect 45266 3500 45276 3556
rect 45332 3500 48356 3556
rect 0 3444 800 3472
rect 48300 3444 48356 3500
rect 49200 3444 50000 3472
rect 0 3388 1708 3444
rect 1764 3388 1774 3444
rect 6066 3388 6076 3444
rect 6132 3388 6972 3444
rect 7028 3388 7038 3444
rect 30902 3388 30940 3444
rect 30996 3388 31006 3444
rect 38994 3388 39004 3444
rect 39060 3388 44604 3444
rect 44660 3388 44670 3444
rect 45836 3388 48076 3444
rect 48132 3388 48142 3444
rect 48300 3388 50000 3444
rect 0 3360 800 3388
rect 45836 3332 45892 3388
rect 49200 3360 50000 3388
rect 38882 3276 38892 3332
rect 38948 3276 45892 3332
rect 19826 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20110 3164
rect 0 2772 800 2800
rect 0 2716 2156 2772
rect 2212 2716 2222 2772
rect 0 2688 800 2716
<< via3 >>
rect 4476 46228 4532 46284
rect 4580 46228 4636 46284
rect 4684 46228 4740 46284
rect 35196 46228 35252 46284
rect 35300 46228 35356 46284
rect 35404 46228 35460 46284
rect 19836 45444 19892 45500
rect 19940 45444 19996 45500
rect 20044 45444 20100 45500
rect 4476 44660 4532 44716
rect 4580 44660 4636 44716
rect 4684 44660 4740 44716
rect 35196 44660 35252 44716
rect 35300 44660 35356 44716
rect 35404 44660 35460 44716
rect 18732 44492 18788 44548
rect 19836 43876 19892 43932
rect 19940 43876 19996 43932
rect 20044 43876 20100 43932
rect 10556 43484 10612 43540
rect 10892 43148 10948 43204
rect 4476 43092 4532 43148
rect 4580 43092 4636 43148
rect 4684 43092 4740 43148
rect 35196 43092 35252 43148
rect 35300 43092 35356 43148
rect 35404 43092 35460 43148
rect 19180 42700 19236 42756
rect 6412 42588 6468 42644
rect 19180 42364 19236 42420
rect 19836 42308 19892 42364
rect 19940 42308 19996 42364
rect 20044 42308 20100 42364
rect 7980 42140 8036 42196
rect 4284 42028 4340 42084
rect 5404 41916 5460 41972
rect 23884 41692 23940 41748
rect 4476 41524 4532 41580
rect 4580 41524 4636 41580
rect 4684 41524 4740 41580
rect 35196 41524 35252 41580
rect 35300 41524 35356 41580
rect 35404 41524 35460 41580
rect 19836 40740 19892 40796
rect 19940 40740 19996 40796
rect 20044 40740 20100 40796
rect 4844 40572 4900 40628
rect 5516 40460 5572 40516
rect 13020 40460 13076 40516
rect 4476 39956 4532 40012
rect 4580 39956 4636 40012
rect 4684 39956 4740 40012
rect 35196 39956 35252 40012
rect 35300 39956 35356 40012
rect 35404 39956 35460 40012
rect 16044 39676 16100 39732
rect 5964 39564 6020 39620
rect 6188 39564 6244 39620
rect 15260 39340 15316 39396
rect 6860 39228 6916 39284
rect 19836 39172 19892 39228
rect 19940 39172 19996 39228
rect 20044 39172 20100 39228
rect 14924 39116 14980 39172
rect 3836 39004 3892 39060
rect 13356 38780 13412 38836
rect 4956 38556 5012 38612
rect 8428 38556 8484 38612
rect 15372 38556 15428 38612
rect 17724 38444 17780 38500
rect 4476 38388 4532 38444
rect 4580 38388 4636 38444
rect 4684 38388 4740 38444
rect 35196 38388 35252 38444
rect 35300 38388 35356 38444
rect 35404 38388 35460 38444
rect 7644 38332 7700 38388
rect 6860 38108 6916 38164
rect 15372 37996 15428 38052
rect 17836 37996 17892 38052
rect 6188 37884 6244 37940
rect 3836 37660 3892 37716
rect 19836 37604 19892 37660
rect 19940 37604 19996 37660
rect 20044 37604 20100 37660
rect 23772 37548 23828 37604
rect 4956 37436 5012 37492
rect 16380 37212 16436 37268
rect 23884 37100 23940 37156
rect 5628 36988 5684 37044
rect 4476 36820 4532 36876
rect 4580 36820 4636 36876
rect 4684 36820 4740 36876
rect 35196 36820 35252 36876
rect 35300 36820 35356 36876
rect 35404 36820 35460 36876
rect 18732 36764 18788 36820
rect 4844 36540 4900 36596
rect 6412 36540 6468 36596
rect 14924 36316 14980 36372
rect 7644 36092 7700 36148
rect 8204 36092 8260 36148
rect 16268 36092 16324 36148
rect 19836 36036 19892 36092
rect 19940 36036 19996 36092
rect 20044 36036 20100 36092
rect 5964 35980 6020 36036
rect 19068 35980 19124 36036
rect 5404 35868 5460 35924
rect 16044 35756 16100 35812
rect 17724 35756 17780 35812
rect 17836 35644 17892 35700
rect 16380 35532 16436 35588
rect 10444 35308 10500 35364
rect 16268 35308 16324 35364
rect 23772 35308 23828 35364
rect 4476 35252 4532 35308
rect 4580 35252 4636 35308
rect 4684 35252 4740 35308
rect 35196 35252 35252 35308
rect 35300 35252 35356 35308
rect 35404 35252 35460 35308
rect 5964 35196 6020 35252
rect 9772 35196 9828 35252
rect 17500 35196 17556 35252
rect 8764 35084 8820 35140
rect 11340 35084 11396 35140
rect 3836 34972 3892 35028
rect 5068 34972 5124 35028
rect 15260 34972 15316 35028
rect 14476 34860 14532 34916
rect 22764 34860 22820 34916
rect 5964 34748 6020 34804
rect 10108 34748 10164 34804
rect 19068 34748 19124 34804
rect 19516 34748 19572 34804
rect 24668 34636 24724 34692
rect 19836 34468 19892 34524
rect 19940 34468 19996 34524
rect 20044 34468 20100 34524
rect 4284 34412 4340 34468
rect 8204 34412 8260 34468
rect 10780 34412 10836 34468
rect 13580 34412 13636 34468
rect 3612 34300 3668 34356
rect 3388 34188 3444 34244
rect 16716 33964 16772 34020
rect 3388 33852 3444 33908
rect 4476 33684 4532 33740
rect 4580 33684 4636 33740
rect 4684 33684 4740 33740
rect 35196 33684 35252 33740
rect 35300 33684 35356 33740
rect 35404 33684 35460 33740
rect 13692 33628 13748 33684
rect 8876 33516 8932 33572
rect 12124 33516 12180 33572
rect 3612 33404 3668 33460
rect 12348 33404 12404 33460
rect 15372 33404 15428 33460
rect 15372 33180 15428 33236
rect 11452 33068 11508 33124
rect 22988 33068 23044 33124
rect 8876 32956 8932 33012
rect 12124 32956 12180 33012
rect 19836 32900 19892 32956
rect 19940 32900 19996 32956
rect 20044 32900 20100 32956
rect 5068 32732 5124 32788
rect 18956 32732 19012 32788
rect 24668 32620 24724 32676
rect 3388 32508 3444 32564
rect 11452 32284 11508 32340
rect 22988 32284 23044 32340
rect 8764 32172 8820 32228
rect 4476 32116 4532 32172
rect 4580 32116 4636 32172
rect 4684 32116 4740 32172
rect 35196 32116 35252 32172
rect 35300 32116 35356 32172
rect 35404 32116 35460 32172
rect 17500 32060 17556 32116
rect 21420 31836 21476 31892
rect 7980 31724 8036 31780
rect 3388 31612 3444 31668
rect 5516 31612 5572 31668
rect 10780 31612 10836 31668
rect 22764 31612 22820 31668
rect 19836 31332 19892 31388
rect 19940 31332 19996 31388
rect 20044 31332 20100 31388
rect 8764 31164 8820 31220
rect 9772 31052 9828 31108
rect 19516 30828 19572 30884
rect 12348 30604 12404 30660
rect 4476 30548 4532 30604
rect 4580 30548 4636 30604
rect 4684 30548 4740 30604
rect 35196 30548 35252 30604
rect 35300 30548 35356 30604
rect 35404 30548 35460 30604
rect 10780 30492 10836 30548
rect 4284 30380 4340 30436
rect 13580 30380 13636 30436
rect 14700 30268 14756 30324
rect 10892 30156 10948 30212
rect 14028 30156 14084 30212
rect 21420 30044 21476 30100
rect 18956 29932 19012 29988
rect 19836 29764 19892 29820
rect 19940 29764 19996 29820
rect 20044 29764 20100 29820
rect 13020 29484 13076 29540
rect 15820 29372 15876 29428
rect 14028 29260 14084 29316
rect 8428 29036 8484 29092
rect 4476 28980 4532 29036
rect 4580 28980 4636 29036
rect 4684 28980 4740 29036
rect 35196 28980 35252 29036
rect 35300 28980 35356 29036
rect 35404 28980 35460 29036
rect 13692 28700 13748 28756
rect 3836 28588 3892 28644
rect 10780 28588 10836 28644
rect 8428 28476 8484 28532
rect 19836 28196 19892 28252
rect 19940 28196 19996 28252
rect 20044 28196 20100 28252
rect 6972 27916 7028 27972
rect 15036 27916 15092 27972
rect 15036 27468 15092 27524
rect 4476 27412 4532 27468
rect 4580 27412 4636 27468
rect 4684 27412 4740 27468
rect 35196 27412 35252 27468
rect 35300 27412 35356 27468
rect 35404 27412 35460 27468
rect 10668 27356 10724 27412
rect 5964 27244 6020 27300
rect 6972 27020 7028 27076
rect 11340 26796 11396 26852
rect 19836 26628 19892 26684
rect 19940 26628 19996 26684
rect 20044 26628 20100 26684
rect 4476 25844 4532 25900
rect 4580 25844 4636 25900
rect 4684 25844 4740 25900
rect 35196 25844 35252 25900
rect 35300 25844 35356 25900
rect 35404 25844 35460 25900
rect 14700 25788 14756 25844
rect 10444 25452 10500 25508
rect 15820 25340 15876 25396
rect 18284 25340 18340 25396
rect 16716 25228 16772 25284
rect 10668 25116 10724 25172
rect 11116 25116 11172 25172
rect 11452 25116 11508 25172
rect 19836 25060 19892 25116
rect 19940 25060 19996 25116
rect 20044 25060 20100 25116
rect 18284 25004 18340 25060
rect 5628 24668 5684 24724
rect 13356 24444 13412 24500
rect 4476 24276 4532 24332
rect 4580 24276 4636 24332
rect 4684 24276 4740 24332
rect 11116 24220 11172 24276
rect 14476 24220 14532 24276
rect 35196 24276 35252 24332
rect 35300 24276 35356 24332
rect 35404 24276 35460 24332
rect 6972 23548 7028 23604
rect 19836 23492 19892 23548
rect 19940 23492 19996 23548
rect 20044 23492 20100 23548
rect 10556 23100 10612 23156
rect 10892 23100 10948 23156
rect 29708 23100 29764 23156
rect 16044 22876 16100 22932
rect 4476 22708 4532 22764
rect 4580 22708 4636 22764
rect 4684 22708 4740 22764
rect 10108 22764 10164 22820
rect 35196 22708 35252 22764
rect 35300 22708 35356 22764
rect 35404 22708 35460 22764
rect 30940 22428 30996 22484
rect 12684 21980 12740 22036
rect 19836 21924 19892 21980
rect 19940 21924 19996 21980
rect 20044 21924 20100 21980
rect 4476 21140 4532 21196
rect 4580 21140 4636 21196
rect 4684 21140 4740 21196
rect 35196 21140 35252 21196
rect 35300 21140 35356 21196
rect 35404 21140 35460 21196
rect 10892 20860 10948 20916
rect 11340 20860 11396 20916
rect 12684 20524 12740 20580
rect 14140 20524 14196 20580
rect 19836 20356 19892 20412
rect 19940 20356 19996 20412
rect 20044 20356 20100 20412
rect 16044 20188 16100 20244
rect 31276 20188 31332 20244
rect 4476 19572 4532 19628
rect 4580 19572 4636 19628
rect 4684 19572 4740 19628
rect 35196 19572 35252 19628
rect 35300 19572 35356 19628
rect 35404 19572 35460 19628
rect 6972 19516 7028 19572
rect 15820 19516 15876 19572
rect 16940 19516 16996 19572
rect 15820 19292 15876 19348
rect 29708 19292 29764 19348
rect 43036 19292 43092 19348
rect 10668 19180 10724 19236
rect 16940 18956 16996 19012
rect 30940 18956 30996 19012
rect 31276 18956 31332 19012
rect 19836 18788 19892 18844
rect 19940 18788 19996 18844
rect 20044 18788 20100 18844
rect 42476 18620 42532 18676
rect 42924 18396 42980 18452
rect 42700 18172 42756 18228
rect 4476 18004 4532 18060
rect 4580 18004 4636 18060
rect 4684 18004 4740 18060
rect 35196 18004 35252 18060
rect 35300 18004 35356 18060
rect 35404 18004 35460 18060
rect 19836 17220 19892 17276
rect 19940 17220 19996 17276
rect 20044 17220 20100 17276
rect 11340 17164 11396 17220
rect 42812 17164 42868 17220
rect 12124 16828 12180 16884
rect 24780 16828 24836 16884
rect 42924 16492 42980 16548
rect 4476 16436 4532 16492
rect 4580 16436 4636 16492
rect 4684 16436 4740 16492
rect 35196 16436 35252 16492
rect 35300 16436 35356 16492
rect 35404 16436 35460 16492
rect 42812 16380 42868 16436
rect 43036 16156 43092 16212
rect 41468 15932 41524 15988
rect 31164 15820 31220 15876
rect 42476 15708 42532 15764
rect 19836 15652 19892 15708
rect 19940 15652 19996 15708
rect 20044 15652 20100 15708
rect 12124 15260 12180 15316
rect 23996 15260 24052 15316
rect 33852 15484 33908 15540
rect 4476 14868 4532 14924
rect 4580 14868 4636 14924
rect 4684 14868 4740 14924
rect 35196 14868 35252 14924
rect 35300 14868 35356 14924
rect 35404 14868 35460 14924
rect 41468 14476 41524 14532
rect 42700 14476 42756 14532
rect 31276 14364 31332 14420
rect 24780 14140 24836 14196
rect 19836 14084 19892 14140
rect 19940 14084 19996 14140
rect 20044 14084 20100 14140
rect 14140 13916 14196 13972
rect 31276 13468 31332 13524
rect 31164 13356 31220 13412
rect 4476 13300 4532 13356
rect 4580 13300 4636 13356
rect 4684 13300 4740 13356
rect 35196 13300 35252 13356
rect 35300 13300 35356 13356
rect 35404 13300 35460 13356
rect 23996 13244 24052 13300
rect 19836 12516 19892 12572
rect 19940 12516 19996 12572
rect 20044 12516 20100 12572
rect 10668 12012 10724 12068
rect 4476 11732 4532 11788
rect 4580 11732 4636 11788
rect 4684 11732 4740 11788
rect 35196 11732 35252 11788
rect 35300 11732 35356 11788
rect 35404 11732 35460 11788
rect 19836 10948 19892 11004
rect 19940 10948 19996 11004
rect 20044 10948 20100 11004
rect 10780 10668 10836 10724
rect 31388 10556 31444 10612
rect 33852 10444 33908 10500
rect 4476 10164 4532 10220
rect 4580 10164 4636 10220
rect 4684 10164 4740 10220
rect 35196 10164 35252 10220
rect 35300 10164 35356 10220
rect 35404 10164 35460 10220
rect 19836 9380 19892 9436
rect 19940 9380 19996 9436
rect 20044 9380 20100 9436
rect 4476 8596 4532 8652
rect 4580 8596 4636 8652
rect 4684 8596 4740 8652
rect 35196 8596 35252 8652
rect 35300 8596 35356 8652
rect 35404 8596 35460 8652
rect 10780 8428 10836 8484
rect 31388 8204 31444 8260
rect 32620 7980 32676 8036
rect 19836 7812 19892 7868
rect 19940 7812 19996 7868
rect 20044 7812 20100 7868
rect 43820 7532 43876 7588
rect 4476 7028 4532 7084
rect 4580 7028 4636 7084
rect 4684 7028 4740 7084
rect 35196 7028 35252 7084
rect 35300 7028 35356 7084
rect 35404 7028 35460 7084
rect 40236 6972 40292 7028
rect 35756 6748 35812 6804
rect 19836 6244 19892 6300
rect 19940 6244 19996 6300
rect 20044 6244 20100 6300
rect 30940 5964 30996 6020
rect 40236 5628 40292 5684
rect 4476 5460 4532 5516
rect 4580 5460 4636 5516
rect 4684 5460 4740 5516
rect 35196 5460 35252 5516
rect 35300 5460 35356 5516
rect 35404 5460 35460 5516
rect 43820 5404 43876 5460
rect 35756 4732 35812 4788
rect 19836 4676 19892 4732
rect 19940 4676 19996 4732
rect 20044 4676 20100 4732
rect 4476 3892 4532 3948
rect 4580 3892 4636 3948
rect 4684 3892 4740 3948
rect 35196 3892 35252 3948
rect 35300 3892 35356 3948
rect 35404 3892 35460 3948
rect 32620 3500 32676 3556
rect 30940 3388 30996 3444
rect 19836 3108 19892 3164
rect 19940 3108 19996 3164
rect 20044 3108 20100 3164
<< metal4 >>
rect 4448 46284 4768 46316
rect 4448 46228 4476 46284
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4740 46228 4768 46284
rect 4448 44716 4768 46228
rect 4448 44660 4476 44716
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4740 44660 4768 44716
rect 4448 43148 4768 44660
rect 19808 45500 20128 46316
rect 19808 45444 19836 45500
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 20100 45444 20128 45500
rect 18732 44548 18788 44558
rect 4448 43092 4476 43148
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4740 43092 4768 43148
rect 4284 42084 4340 42094
rect 3836 39060 3892 39070
rect 3836 37716 3892 39004
rect 3836 37650 3892 37660
rect 3836 35028 3892 35038
rect 3612 34356 3668 34366
rect 3388 34244 3444 34254
rect 3388 33908 3444 34188
rect 3388 33842 3444 33852
rect 3612 33460 3668 34300
rect 3612 33394 3668 33404
rect 3388 32564 3444 32574
rect 3388 31668 3444 32508
rect 3388 31602 3444 31612
rect 3836 28644 3892 34972
rect 4284 34468 4340 42028
rect 4284 30436 4340 34412
rect 4284 30370 4340 30380
rect 4448 41580 4768 43092
rect 10556 43540 10612 43550
rect 6412 42644 6468 42654
rect 4448 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4768 41580
rect 4448 40012 4768 41524
rect 5404 41972 5460 41982
rect 4448 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4768 40012
rect 4448 38444 4768 39956
rect 4448 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4768 38444
rect 4448 36876 4768 38388
rect 4448 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4768 36876
rect 4448 35308 4768 36820
rect 4844 40628 4900 40638
rect 4844 36596 4900 40572
rect 4956 38612 5012 38622
rect 4956 37492 5012 38556
rect 4956 37426 5012 37436
rect 4844 36530 4900 36540
rect 5404 35924 5460 41916
rect 5404 35858 5460 35868
rect 5516 40516 5572 40526
rect 4448 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4768 35308
rect 4448 33740 4768 35252
rect 4448 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4768 33740
rect 4448 32172 4768 33684
rect 5068 35028 5124 35038
rect 5068 32788 5124 34972
rect 5068 32722 5124 32732
rect 4448 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4768 32172
rect 4448 30604 4768 32116
rect 5516 31668 5572 40460
rect 5964 39620 6020 39630
rect 5516 31602 5572 31612
rect 5628 37044 5684 37054
rect 4448 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4768 30604
rect 3836 28578 3892 28588
rect 4448 29036 4768 30548
rect 4448 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4768 29036
rect 4448 27468 4768 28980
rect 4448 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4768 27468
rect 4448 25900 4768 27412
rect 4448 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4768 25900
rect 4448 24332 4768 25844
rect 5628 24724 5684 36988
rect 5964 36036 6020 39564
rect 6188 39620 6244 39630
rect 6188 37940 6244 39564
rect 6188 37874 6244 37884
rect 6412 36596 6468 42588
rect 7980 42196 8036 42206
rect 6860 39284 6916 39294
rect 6860 38164 6916 39228
rect 6860 38098 6916 38108
rect 7644 38388 7700 38398
rect 6412 36530 6468 36540
rect 7644 36148 7700 38332
rect 7644 36082 7700 36092
rect 5964 35970 6020 35980
rect 5964 35252 6020 35262
rect 5964 34804 6020 35196
rect 5964 27300 6020 34748
rect 7980 31780 8036 42140
rect 8428 38612 8484 38622
rect 8204 36148 8260 36158
rect 8204 34468 8260 36092
rect 8204 34402 8260 34412
rect 7980 31714 8036 31724
rect 8428 29092 8484 38556
rect 10444 35364 10500 35374
rect 9772 35252 9828 35262
rect 8764 35140 8820 35150
rect 8764 32228 8820 35084
rect 8876 33572 8932 33582
rect 8876 33012 8932 33516
rect 8876 32946 8932 32956
rect 8764 31220 8820 32172
rect 8764 31154 8820 31164
rect 9772 31108 9828 35196
rect 9772 31042 9828 31052
rect 10108 34804 10164 34814
rect 8428 28532 8484 29036
rect 8428 28466 8484 28476
rect 5964 27234 6020 27244
rect 6972 27972 7028 27982
rect 5628 24658 5684 24668
rect 6972 27076 7028 27916
rect 4448 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4768 24332
rect 4448 22764 4768 24276
rect 4448 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4768 22764
rect 4448 21196 4768 22708
rect 4448 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4768 21196
rect 4448 19628 4768 21140
rect 4448 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4768 19628
rect 4448 18060 4768 19572
rect 6972 23604 7028 27020
rect 6972 19572 7028 23548
rect 10108 22820 10164 34748
rect 10444 25508 10500 35308
rect 10444 25442 10500 25452
rect 10556 23156 10612 43484
rect 10892 43204 10948 43214
rect 10780 34468 10836 34478
rect 10780 31668 10836 34412
rect 10780 31602 10836 31612
rect 10780 30548 10836 30558
rect 10780 28644 10836 30492
rect 10892 30212 10948 43148
rect 13020 40516 13076 40526
rect 10892 30146 10948 30156
rect 11340 35140 11396 35150
rect 10780 28578 10836 28588
rect 10668 27412 10724 27422
rect 10668 25172 10724 27356
rect 11340 26852 11396 35084
rect 12124 33572 12180 33582
rect 11340 26786 11396 26796
rect 11452 33124 11508 33134
rect 11452 32340 11508 33068
rect 12124 33012 12180 33516
rect 12124 32946 12180 32956
rect 12348 33460 12404 33470
rect 10668 25106 10724 25116
rect 11116 25172 11172 25182
rect 11116 24276 11172 25116
rect 11452 25172 11508 32284
rect 12348 30660 12404 33404
rect 12348 30594 12404 30604
rect 13020 29540 13076 40460
rect 16044 39732 16100 39742
rect 15260 39396 15316 39406
rect 14924 39172 14980 39182
rect 13020 29474 13076 29484
rect 13356 38836 13412 38846
rect 11452 25106 11508 25116
rect 13356 24500 13412 38780
rect 14924 36372 14980 39116
rect 14924 36306 14980 36316
rect 15260 35028 15316 39340
rect 15372 38612 15428 38622
rect 15372 38052 15428 38556
rect 15372 37986 15428 37996
rect 16044 35812 16100 39676
rect 17724 38500 17780 38510
rect 16380 37268 16436 37278
rect 16044 35746 16100 35756
rect 16268 36148 16324 36158
rect 16268 35364 16324 36092
rect 16380 35588 16436 37212
rect 17724 35812 17780 38444
rect 17724 35746 17780 35756
rect 17836 38052 17892 38062
rect 17836 35700 17892 37996
rect 18732 36820 18788 44492
rect 19808 43932 20128 45444
rect 19808 43876 19836 43932
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 20100 43876 20128 43932
rect 19180 42756 19236 42766
rect 19180 42420 19236 42700
rect 19180 42354 19236 42364
rect 19808 42364 20128 43876
rect 18732 36754 18788 36764
rect 19808 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20128 42364
rect 19808 40796 20128 42308
rect 35168 46284 35488 46316
rect 35168 46228 35196 46284
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35460 46228 35488 46284
rect 35168 44716 35488 46228
rect 35168 44660 35196 44716
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35460 44660 35488 44716
rect 35168 43148 35488 44660
rect 35168 43092 35196 43148
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35460 43092 35488 43148
rect 19808 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20128 40796
rect 19808 39228 20128 40740
rect 19808 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20128 39228
rect 19808 37660 20128 39172
rect 19808 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20128 37660
rect 23884 41748 23940 41758
rect 19808 36092 20128 37604
rect 17836 35634 17892 35644
rect 19068 36036 19124 36046
rect 16380 35522 16436 35532
rect 16268 35298 16324 35308
rect 15260 34962 15316 34972
rect 17500 35252 17556 35262
rect 14476 34916 14532 34926
rect 13580 34468 13636 34478
rect 13580 30436 13636 34412
rect 13580 30370 13636 30380
rect 13692 33684 13748 33694
rect 13692 28756 13748 33628
rect 14028 30212 14084 30222
rect 14028 29316 14084 30156
rect 14028 29250 14084 29260
rect 13692 28690 13748 28700
rect 13356 24434 13412 24444
rect 11116 24210 11172 24220
rect 14476 24276 14532 34860
rect 16716 34020 16772 34030
rect 15372 33460 15428 33470
rect 15372 33236 15428 33404
rect 15372 33170 15428 33180
rect 14700 30324 14756 30334
rect 14700 25844 14756 30268
rect 15820 29428 15876 29438
rect 15036 27972 15092 27982
rect 15036 27524 15092 27916
rect 15036 27458 15092 27468
rect 14700 25778 14756 25788
rect 15820 25396 15876 29372
rect 15820 25330 15876 25340
rect 16716 25284 16772 33964
rect 17500 32116 17556 35196
rect 19068 34804 19124 35980
rect 19808 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20128 36092
rect 19068 34738 19124 34748
rect 19516 34804 19572 34814
rect 17500 32050 17556 32060
rect 18956 32788 19012 32798
rect 18956 29988 19012 32732
rect 19516 30884 19572 34748
rect 19516 30818 19572 30828
rect 19808 34524 20128 36036
rect 23772 37604 23828 37614
rect 23772 35364 23828 37548
rect 23884 37156 23940 41692
rect 23884 37090 23940 37100
rect 35168 41580 35488 43092
rect 35168 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35488 41580
rect 35168 40012 35488 41524
rect 35168 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35488 40012
rect 35168 38444 35488 39956
rect 35168 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35488 38444
rect 23772 35298 23828 35308
rect 35168 36876 35488 38388
rect 35168 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35488 36876
rect 35168 35308 35488 36820
rect 35168 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35488 35308
rect 19808 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20128 34524
rect 19808 32956 20128 34468
rect 19808 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20128 32956
rect 19808 31388 20128 32900
rect 22764 34916 22820 34926
rect 19808 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20128 31388
rect 18956 29922 19012 29932
rect 19808 29820 20128 31332
rect 21420 31892 21476 31902
rect 21420 30100 21476 31836
rect 22764 31668 22820 34860
rect 24668 34692 24724 34702
rect 22988 33124 23044 33134
rect 22988 32340 23044 33068
rect 24668 32676 24724 34636
rect 24668 32610 24724 32620
rect 35168 33740 35488 35252
rect 35168 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35488 33740
rect 22988 32274 23044 32284
rect 22764 31602 22820 31612
rect 35168 32172 35488 33684
rect 35168 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35488 32172
rect 21420 30034 21476 30044
rect 35168 30604 35488 32116
rect 35168 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35488 30604
rect 19808 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20128 29820
rect 19808 28252 20128 29764
rect 19808 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20128 28252
rect 19808 26684 20128 28196
rect 19808 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20128 26684
rect 16716 25218 16772 25228
rect 18284 25396 18340 25406
rect 18284 25060 18340 25340
rect 18284 24994 18340 25004
rect 19808 25116 20128 26628
rect 19808 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20128 25116
rect 14476 24210 14532 24220
rect 19808 23548 20128 25060
rect 19808 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20128 23548
rect 10556 23090 10612 23100
rect 10892 23156 10948 23166
rect 10108 22754 10164 22764
rect 10892 20916 10948 23100
rect 16044 22932 16100 22942
rect 12684 22036 12740 22046
rect 10892 20850 10948 20860
rect 11340 20916 11396 20926
rect 6972 19506 7028 19516
rect 4448 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4768 18060
rect 4448 16492 4768 18004
rect 4448 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4768 16492
rect 4448 14924 4768 16436
rect 4448 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4768 14924
rect 4448 13356 4768 14868
rect 4448 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4768 13356
rect 4448 11788 4768 13300
rect 10668 19236 10724 19246
rect 10668 12068 10724 19180
rect 11340 17220 11396 20860
rect 12684 20580 12740 21980
rect 12684 20514 12740 20524
rect 14140 20580 14196 20590
rect 11340 17154 11396 17164
rect 12124 16884 12180 16894
rect 12124 15316 12180 16828
rect 12124 15250 12180 15260
rect 14140 13972 14196 20524
rect 16044 20244 16100 22876
rect 16044 20178 16100 20188
rect 19808 21980 20128 23492
rect 35168 29036 35488 30548
rect 35168 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35488 29036
rect 35168 27468 35488 28980
rect 35168 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35488 27468
rect 35168 25900 35488 27412
rect 35168 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35488 25900
rect 35168 24332 35488 25844
rect 35168 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35488 24332
rect 19808 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20128 21980
rect 19808 20412 20128 21924
rect 19808 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20128 20412
rect 15820 19572 15876 19582
rect 15820 19348 15876 19516
rect 15820 19282 15876 19292
rect 16940 19572 16996 19582
rect 16940 19012 16996 19516
rect 16940 18946 16996 18956
rect 14140 13906 14196 13916
rect 19808 18844 20128 20356
rect 29708 23156 29764 23166
rect 29708 19348 29764 23100
rect 35168 22764 35488 24276
rect 35168 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35488 22764
rect 29708 19282 29764 19292
rect 30940 22484 30996 22494
rect 30940 19012 30996 22428
rect 35168 21196 35488 22708
rect 35168 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35488 21196
rect 30940 18946 30996 18956
rect 31276 20244 31332 20254
rect 31276 19012 31332 20188
rect 31276 18946 31332 18956
rect 35168 19628 35488 21140
rect 35168 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35488 19628
rect 19808 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20128 18844
rect 19808 17276 20128 18788
rect 19808 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20128 17276
rect 19808 15708 20128 17220
rect 35168 18060 35488 19572
rect 43036 19348 43092 19358
rect 35168 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35488 18060
rect 19808 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20128 15708
rect 19808 14140 20128 15652
rect 24780 16884 24836 16894
rect 19808 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20128 14140
rect 10668 12002 10724 12012
rect 19808 12572 20128 14084
rect 23996 15316 24052 15326
rect 23996 13300 24052 15260
rect 24780 14196 24836 16828
rect 35168 16492 35488 18004
rect 35168 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35488 16492
rect 24780 14130 24836 14140
rect 31164 15876 31220 15886
rect 31164 13412 31220 15820
rect 33852 15540 33908 15550
rect 31276 14420 31332 14430
rect 31276 13524 31332 14364
rect 31276 13458 31332 13468
rect 31164 13346 31220 13356
rect 23996 13234 24052 13244
rect 19808 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20128 12572
rect 4448 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4768 11788
rect 4448 10220 4768 11732
rect 19808 11004 20128 12516
rect 19808 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20128 11004
rect 4448 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4768 10220
rect 4448 8652 4768 10164
rect 4448 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4768 8652
rect 4448 7084 4768 8596
rect 10780 10724 10836 10734
rect 10780 8484 10836 10668
rect 10780 8418 10836 8428
rect 19808 9436 20128 10948
rect 19808 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20128 9436
rect 4448 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4768 7084
rect 4448 5516 4768 7028
rect 4448 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4768 5516
rect 4448 3948 4768 5460
rect 4448 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4768 3948
rect 4448 3076 4768 3892
rect 19808 7868 20128 9380
rect 31388 10612 31444 10622
rect 31388 8260 31444 10556
rect 33852 10500 33908 15484
rect 33852 10434 33908 10444
rect 35168 14924 35488 16436
rect 42476 18676 42532 18686
rect 35168 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35488 14924
rect 35168 13356 35488 14868
rect 41468 15988 41524 15998
rect 41468 14532 41524 15932
rect 42476 15764 42532 18620
rect 42924 18452 42980 18462
rect 42476 15698 42532 15708
rect 42700 18228 42756 18238
rect 41468 14466 41524 14476
rect 42700 14532 42756 18172
rect 42812 17220 42868 17230
rect 42812 16436 42868 17164
rect 42924 16548 42980 18396
rect 42924 16482 42980 16492
rect 42812 16370 42868 16380
rect 43036 16212 43092 19292
rect 43036 16146 43092 16156
rect 42700 14466 42756 14476
rect 35168 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35488 13356
rect 35168 11788 35488 13300
rect 35168 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35488 11788
rect 31388 8194 31444 8204
rect 35168 10220 35488 11732
rect 35168 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35488 10220
rect 35168 8652 35488 10164
rect 35168 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35488 8652
rect 19808 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20128 7868
rect 19808 6300 20128 7812
rect 19808 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20128 6300
rect 19808 4732 20128 6244
rect 32620 8036 32676 8046
rect 19808 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20128 4732
rect 19808 3164 20128 4676
rect 30940 6020 30996 6030
rect 30940 3444 30996 5964
rect 32620 3556 32676 7980
rect 32620 3490 32676 3500
rect 35168 7084 35488 8596
rect 35168 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35488 7084
rect 43820 7588 43876 7598
rect 35168 5516 35488 7028
rect 40236 7028 40292 7038
rect 35168 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35488 5516
rect 35168 3948 35488 5460
rect 35756 6804 35812 6814
rect 35756 4788 35812 6748
rect 40236 5684 40292 6972
rect 40236 5618 40292 5628
rect 43820 5460 43876 7532
rect 43820 5394 43876 5404
rect 35756 4722 35812 4732
rect 35168 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35488 3948
rect 30940 3378 30996 3388
rect 19808 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20128 3164
rect 19808 3076 20128 3108
rect 35168 3076 35488 3892
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1031_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 24304 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_2  _1032_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 22176 0 -1 29792
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1033_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 14672 0 1 26656
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1034_
timestamp 1698431365
transform 1 0 4816 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1035_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5824 0 1 37632
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1036_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 7168 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1037_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 12432 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1038_
timestamp 1698431365
transform -1 0 14672 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1039_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 4144 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1040_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 3472 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1041_
timestamp 1698431365
transform 1 0 11872 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1042_
timestamp 1698431365
transform -1 0 11872 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1043_
timestamp 1698431365
transform -1 0 11088 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1044_
timestamp 1698431365
transform -1 0 3136 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1045_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 2576 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1046_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 9856 0 -1 34496
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _1047_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 9968 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1048_
timestamp 1698431365
transform -1 0 26544 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1049_
timestamp 1698431365
transform -1 0 23520 0 -1 34496
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1050_
timestamp 1698431365
transform 1 0 21168 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1051_
timestamp 1698431365
transform -1 0 20720 0 1 34496
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1052_
timestamp 1698431365
transform -1 0 11200 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1053_
timestamp 1698431365
transform 1 0 4368 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1054_
timestamp 1698431365
transform -1 0 9856 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1055_
timestamp 1698431365
transform 1 0 8848 0 1 34496
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1056_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5600 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1057_
timestamp 1698431365
transform -1 0 7280 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1058_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 6272 0 -1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1059_
timestamp 1698431365
transform 1 0 15120 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1060_
timestamp 1698431365
transform -1 0 14896 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1061_
timestamp 1698431365
transform -1 0 13104 0 1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1062_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 9856 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1063_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 2016 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1064_
timestamp 1698431365
transform -1 0 13104 0 1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1065_
timestamp 1698431365
transform -1 0 18816 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1066_
timestamp 1698431365
transform 1 0 17248 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1067_
timestamp 1698431365
transform -1 0 18256 0 1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1068_
timestamp 1698431365
transform 1 0 16576 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1069_
timestamp 1698431365
transform -1 0 16016 0 -1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1070_
timestamp 1698431365
transform 1 0 8512 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1071_
timestamp 1698431365
transform 1 0 11648 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1072_
timestamp 1698431365
transform 1 0 11648 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1073_
timestamp 1698431365
transform -1 0 12544 0 1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1074_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 13104 0 1 31360
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _1075_
timestamp 1698431365
transform 1 0 10192 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  _1076_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 15904 0 1 32928
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1077_
timestamp 1698431365
transform 1 0 19600 0 1 26656
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _1078_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 19600 0 -1 25088
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1079_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 23184 0 -1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1080_
timestamp 1698431365
transform 1 0 6944 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1081_
timestamp 1698431365
transform 1 0 12208 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1082_
timestamp 1698431365
transform 1 0 12320 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1083_
timestamp 1698431365
transform -1 0 11984 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1084_
timestamp 1698431365
transform 1 0 10416 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1085_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 11312 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1086_
timestamp 1698431365
transform 1 0 15792 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1087_
timestamp 1698431365
transform 1 0 6048 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1088_
timestamp 1698431365
transform -1 0 15456 0 1 40768
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _1089_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 11200 0 -1 40768
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _1090_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 12320 0 -1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1091_
timestamp 1698431365
transform -1 0 5040 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1092_
timestamp 1698431365
transform 1 0 5488 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1093_
timestamp 1698431365
transform -1 0 7280 0 1 31360
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1094_
timestamp 1698431365
transform -1 0 26768 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1095_
timestamp 1698431365
transform -1 0 23184 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1096_
timestamp 1698431365
transform 1 0 18816 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1097_
timestamp 1698431365
transform 1 0 19712 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1098_
timestamp 1698431365
transform -1 0 19600 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1099_
timestamp 1698431365
transform -1 0 18144 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1100_
timestamp 1698431365
transform -1 0 20048 0 1 31360
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1101_
timestamp 1698431365
transform -1 0 19712 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1102_
timestamp 1698431365
transform -1 0 15904 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1103_
timestamp 1698431365
transform 1 0 15904 0 1 29792
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1104_
timestamp 1698431365
transform -1 0 19488 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1105_
timestamp 1698431365
transform -1 0 15232 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1106_
timestamp 1698431365
transform 1 0 13552 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1107_
timestamp 1698431365
transform 1 0 16128 0 1 37632
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _1108_
timestamp 1698431365
transform 1 0 15232 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1109_
timestamp 1698431365
transform -1 0 10528 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1110_
timestamp 1698431365
transform -1 0 27776 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1111_
timestamp 1698431365
transform -1 0 23856 0 1 34496
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_4  _1112_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 15344 0 -1 32928
box -86 -86 4902 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1113_
timestamp 1698431365
transform -1 0 7056 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1114_
timestamp 1698431365
transform -1 0 6608 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1115_
timestamp 1698431365
transform 1 0 8400 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_4  _1116_
timestamp 1698431365
transform 1 0 16128 0 1 32928
box -86 -86 4902 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1117_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 19040 0 1 31360
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1118_
timestamp 1698431365
transform 1 0 14224 0 1 29792
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1119_
timestamp 1698431365
transform -1 0 18816 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1120_
timestamp 1698431365
transform -1 0 6160 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1121_
timestamp 1698431365
transform 1 0 13104 0 -1 26656
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1122_
timestamp 1698431365
transform -1 0 17696 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _1123_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 14896 0 1 31360
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1124_
timestamp 1698431365
transform 1 0 11760 0 1 34496
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1125_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 15904 0 1 34496
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _1126_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 13440 0 1 34496
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1127_
timestamp 1698431365
transform 1 0 3136 0 1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _1128_
timestamp 1698431365
transform 1 0 11088 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1129_
timestamp 1698431365
transform 1 0 8624 0 -1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _1130_
timestamp 1698431365
transform 1 0 10080 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1131_
timestamp 1698431365
transform 1 0 12880 0 -1 34496
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1132_
timestamp 1698431365
transform 1 0 8624 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1133_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 10528 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1134_
timestamp 1698431365
transform -1 0 9408 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1135_
timestamp 1698431365
transform -1 0 6720 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1136_
timestamp 1698431365
transform -1 0 8512 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1137_
timestamp 1698431365
transform 1 0 7616 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _1138_
timestamp 1698431365
transform -1 0 9072 0 1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _1139_
timestamp 1698431365
transform -1 0 27776 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1140_
timestamp 1698431365
transform -1 0 23072 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _1141_
timestamp 1698431365
transform 1 0 17248 0 -1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1142_
timestamp 1698431365
transform -1 0 10304 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _1143_
timestamp 1698431365
transform 1 0 9520 0 1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1144_
timestamp 1698431365
transform -1 0 11200 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _1145_
timestamp 1698431365
transform 1 0 7056 0 1 39200
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1146_
timestamp 1698431365
transform 1 0 8288 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1147_
timestamp 1698431365
transform -1 0 17024 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _1148_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 10752 0 1 28224
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__or4_2  _1149_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 10976 0 -1 29792
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1150_
timestamp 1698431365
transform -1 0 16912 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1151_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 5264 0 1 28224
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1152_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 2240 0 -1 29792
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1153_
timestamp 1698431365
transform -1 0 13104 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1154_
timestamp 1698431365
transform -1 0 5488 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1155_
timestamp 1698431365
transform -1 0 7392 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1156_
timestamp 1698431365
transform 1 0 7280 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or4_2  _1157_
timestamp 1698431365
transform -1 0 8960 0 -1 40768
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _1158_
timestamp 1698431365
transform 1 0 3024 0 -1 36064
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1159_
timestamp 1698431365
transform -1 0 4480 0 1 31360
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1160_
timestamp 1698431365
transform 1 0 2576 0 -1 32928
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1161_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 9408 0 -1 28224
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1162_
timestamp 1698431365
transform -1 0 9184 0 -1 42336
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1163_
timestamp 1698431365
transform -1 0 9184 0 1 29792
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1164_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1568 0 -1 31360
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_4  _1165_
timestamp 1698431365
transform 1 0 3360 0 -1 29792
box -86 -86 4902 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1166_
timestamp 1698431365
transform 1 0 5488 0 1 29792
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1167_
timestamp 1698431365
transform -1 0 27104 0 1 34496
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1168_
timestamp 1698431365
transform -1 0 20608 0 1 40768
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1169_
timestamp 1698431365
transform -1 0 17920 0 -1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1170_
timestamp 1698431365
transform -1 0 16912 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1171_
timestamp 1698431365
transform -1 0 21168 0 -1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1172_
timestamp 1698431365
transform 1 0 16464 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _1173_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 17024 0 -1 40768
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1174_
timestamp 1698431365
transform -1 0 14112 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1175_
timestamp 1698431365
transform -1 0 16800 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1176_
timestamp 1698431365
transform -1 0 16576 0 -1 36064
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1177_
timestamp 1698431365
transform 1 0 8064 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1178_
timestamp 1698431365
transform 1 0 13328 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1179_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 16464 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _1180_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 10416 0 -1 31360
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _1181_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 13552 0 -1 31360
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1182_
timestamp 1698431365
transform -1 0 8400 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1183_
timestamp 1698431365
transform -1 0 22848 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1184_
timestamp 1698431365
transform 1 0 8960 0 1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _1185_
timestamp 1698431365
transform -1 0 10752 0 -1 40768
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1186_
timestamp 1698431365
transform 1 0 8512 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _1187_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 9072 0 1 40768
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1188_
timestamp 1698431365
transform -1 0 8288 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1189_
timestamp 1698431365
transform 1 0 5824 0 1 32928
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1190_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 7504 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1191_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 8288 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_2  _1192_
timestamp 1698431365
transform 1 0 11312 0 -1 31360
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _1193_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 8736 0 1 31360
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _1194_
timestamp 1698431365
transform -1 0 8624 0 -1 31360
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1195_
timestamp 1698431365
transform 1 0 4816 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1196_
timestamp 1698431365
transform -1 0 5712 0 -1 37632
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1197_
timestamp 1698431365
transform -1 0 12544 0 1 39200
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1198_
timestamp 1698431365
transform -1 0 6384 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1199_
timestamp 1698431365
transform 1 0 5488 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1200_
timestamp 1698431365
transform 1 0 8288 0 1 26656
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1201_
timestamp 1698431365
transform -1 0 13776 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1202_
timestamp 1698431365
transform -1 0 11648 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1203_
timestamp 1698431365
transform 1 0 6832 0 -1 26656
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1204_
timestamp 1698431365
transform -1 0 11760 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1205_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 9184 0 -1 25088
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _1206_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5712 0 -1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _1207_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5824 0 1 25088
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1208_
timestamp 1698431365
transform -1 0 7168 0 1 36064
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _1209_
timestamp 1698431365
transform 1 0 10080 0 -1 42336
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1210_
timestamp 1698431365
transform 1 0 10640 0 1 36064
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1211_
timestamp 1698431365
transform 1 0 18032 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _1212_
timestamp 1698431365
transform -1 0 16128 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _1213_
timestamp 1698431365
transform -1 0 14112 0 -1 39200
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1214_
timestamp 1698431365
transform 1 0 11648 0 1 37632
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1215_
timestamp 1698431365
transform -1 0 11648 0 1 37632
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1216_
timestamp 1698431365
transform 1 0 9184 0 1 37632
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1217_
timestamp 1698431365
transform 1 0 11424 0 -1 37632
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1218_
timestamp 1698431365
transform -1 0 11424 0 -1 37632
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1219_
timestamp 1698431365
transform 1 0 18144 0 -1 34496
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1220_
timestamp 1698431365
transform -1 0 22288 0 -1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1221_
timestamp 1698431365
transform -1 0 22512 0 1 32928
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1222_
timestamp 1698431365
transform -1 0 24864 0 -1 29792
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1223_
timestamp 1698431365
transform -1 0 25312 0 1 28224
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _1224_
timestamp 1698431365
transform 1 0 20720 0 -1 34496
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1225_
timestamp 1698431365
transform -1 0 20720 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1226_
timestamp 1698431365
transform 1 0 17472 0 -1 39200
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1227_
timestamp 1698431365
transform 1 0 14224 0 1 36064
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1228_
timestamp 1698431365
transform 1 0 16800 0 1 36064
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1229_
timestamp 1698431365
transform 1 0 19264 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1230_
timestamp 1698431365
transform 1 0 19936 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1231_
timestamp 1698431365
transform -1 0 22848 0 -1 37632
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _1232_
timestamp 1698431365
transform 1 0 19712 0 1 37632
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1233_
timestamp 1698431365
transform 1 0 19712 0 -1 37632
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1234_
timestamp 1698431365
transform -1 0 23744 0 -1 32928
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1235_
timestamp 1698431365
transform -1 0 22176 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1236_
timestamp 1698431365
transform -1 0 23632 0 1 36064
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _1237_
timestamp 1698431365
transform -1 0 24080 0 -1 36064
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _1238_
timestamp 1698431365
transform -1 0 15456 0 -1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1239_
timestamp 1698431365
transform -1 0 10752 0 1 23520
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1240_
timestamp 1698431365
transform -1 0 8176 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1241_
timestamp 1698431365
transform -1 0 20384 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1242_
timestamp 1698431365
transform 1 0 19600 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1243_
timestamp 1698431365
transform -1 0 21168 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1244_
timestamp 1698431365
transform -1 0 8848 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1245_
timestamp 1698431365
transform -1 0 47040 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1246_
timestamp 1698431365
transform -1 0 48048 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _1247_
timestamp 1698431365
transform 1 0 34384 0 1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _1248_
timestamp 1698431365
transform -1 0 44464 0 1 12544
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1249_
timestamp 1698431365
transform 1 0 35280 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1250_
timestamp 1698431365
transform -1 0 47040 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_4  _1251_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 37184 0 1 12544
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1252_
timestamp 1698431365
transform -1 0 48160 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_4  _1253_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 43008 0 -1 14112
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1254_
timestamp 1698431365
transform 1 0 34160 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1255_
timestamp 1698431365
transform -1 0 34160 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1256_
timestamp 1698431365
transform 1 0 34944 0 1 14112
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1257_
timestamp 1698431365
transform 1 0 35056 0 -1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _1258_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 45696 0 -1 12544
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1259_
timestamp 1698431365
transform -1 0 40544 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1260_
timestamp 1698431365
transform -1 0 42448 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1261_
timestamp 1698431365
transform -1 0 39984 0 -1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _1262_
timestamp 1698431365
transform -1 0 48160 0 -1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1263_
timestamp 1698431365
transform 1 0 34160 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _1264_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 44464 0 1 14112
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1265_
timestamp 1698431365
transform -1 0 30576 0 -1 12544
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1266_
timestamp 1698431365
transform 1 0 40768 0 -1 14112
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1267_
timestamp 1698431365
transform -1 0 20384 0 1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _1268_
timestamp 1698431365
transform -1 0 19824 0 -1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1269_
timestamp 1698431365
transform 1 0 21168 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1270_
timestamp 1698431365
transform 1 0 5488 0 1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1271_
timestamp 1698431365
transform -1 0 5264 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1272_
timestamp 1698431365
transform -1 0 8288 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1273_
timestamp 1698431365
transform 1 0 4592 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1274_
timestamp 1698431365
transform -1 0 5600 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1275_
timestamp 1698431365
transform 1 0 21168 0 1 14112
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1276_
timestamp 1698431365
transform 1 0 16800 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1277_
timestamp 1698431365
transform -1 0 8176 0 -1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1278_
timestamp 1698431365
transform -1 0 8288 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1279_
timestamp 1698431365
transform -1 0 5264 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1280_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 5152 0 -1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1281_
timestamp 1698431365
transform 1 0 10528 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1282_
timestamp 1698431365
transform -1 0 20944 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1283_
timestamp 1698431365
transform -1 0 12208 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1284_
timestamp 1698431365
transform -1 0 9856 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1285_
timestamp 1698431365
transform 1 0 17248 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1286_
timestamp 1698431365
transform -1 0 18144 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1287_
timestamp 1698431365
transform 1 0 9968 0 1 7840
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _1288_
timestamp 1698431365
transform 1 0 11200 0 -1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1289_
timestamp 1698431365
transform 1 0 6720 0 1 20384
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1290_
timestamp 1698431365
transform 1 0 12432 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1291_
timestamp 1698431365
transform 1 0 12208 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1292_
timestamp 1698431365
transform -1 0 5152 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1293_
timestamp 1698431365
transform -1 0 40544 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1294_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 39648 0 1 10976
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _1295_
timestamp 1698431365
transform -1 0 38640 0 -1 12544
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1296_
timestamp 1698431365
transform 1 0 36848 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1297_
timestamp 1698431365
transform 1 0 38640 0 -1 12544
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1298_
timestamp 1698431365
transform -1 0 23856 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1299_
timestamp 1698431365
transform -1 0 22176 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _1300_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 7280 0 -1 20384
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1301_
timestamp 1698431365
transform 1 0 3024 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1302_
timestamp 1698431365
transform -1 0 5936 0 -1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1303_
timestamp 1698431365
transform 1 0 5488 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1304_
timestamp 1698431365
transform 1 0 21616 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1305_
timestamp 1698431365
transform -1 0 23968 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1306_
timestamp 1698431365
transform -1 0 22736 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1307_
timestamp 1698431365
transform 1 0 9072 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1308_
timestamp 1698431365
transform 1 0 11536 0 1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1309_
timestamp 1698431365
transform 1 0 12096 0 1 10976
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1310_
timestamp 1698431365
transform 1 0 13328 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1311_
timestamp 1698431365
transform -1 0 11760 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1312_
timestamp 1698431365
transform -1 0 11312 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1313_
timestamp 1698431365
transform 1 0 5600 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1314_
timestamp 1698431365
transform 1 0 3472 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1315_
timestamp 1698431365
transform 1 0 8736 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1316_
timestamp 1698431365
transform -1 0 10080 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1317_
timestamp 1698431365
transform 1 0 8512 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1318_
timestamp 1698431365
transform -1 0 10304 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _1319_
timestamp 1698431365
transform 1 0 6160 0 -1 25088
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _1320_
timestamp 1698431365
transform 1 0 7840 0 1 18816
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _1321_
timestamp 1698431365
transform -1 0 5264 0 -1 20384
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1322_
timestamp 1698431365
transform -1 0 5264 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1323_
timestamp 1698431365
transform -1 0 4032 0 -1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1324_
timestamp 1698431365
transform -1 0 7616 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _1325_
timestamp 1698431365
transform 1 0 3360 0 1 18816
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1326_
timestamp 1698431365
transform 1 0 17248 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1327_
timestamp 1698431365
transform 1 0 17360 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1328_
timestamp 1698431365
transform -1 0 9520 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1329_
timestamp 1698431365
transform 1 0 10752 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1330_
timestamp 1698431365
transform 1 0 11088 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1331_
timestamp 1698431365
transform -1 0 9184 0 -1 20384
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _1332_
timestamp 1698431365
transform -1 0 8736 0 1 17248
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1333_
timestamp 1698431365
transform -1 0 8288 0 -1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1334_
timestamp 1698431365
transform -1 0 11424 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1335_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 10752 0 1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1336_
timestamp 1698431365
transform -1 0 5488 0 -1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _1337_
timestamp 1698431365
transform 1 0 3472 0 -1 17248
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1338_
timestamp 1698431365
transform -1 0 11424 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1339_
timestamp 1698431365
transform 1 0 10080 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1340_
timestamp 1698431365
transform -1 0 10192 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1341_
timestamp 1698431365
transform -1 0 11536 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _1342_
timestamp 1698431365
transform 1 0 7056 0 1 15680
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1343_
timestamp 1698431365
transform -1 0 7728 0 -1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1344_
timestamp 1698431365
transform -1 0 44016 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1345_
timestamp 1698431365
transform 1 0 35056 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1346_
timestamp 1698431365
transform 1 0 36848 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1347_
timestamp 1698431365
transform -1 0 38416 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1348_
timestamp 1698431365
transform 1 0 37744 0 1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1349_
timestamp 1698431365
transform 1 0 38416 0 -1 7840
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1350_
timestamp 1698431365
transform -1 0 43008 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1351_
timestamp 1698431365
transform 1 0 36288 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1352_
timestamp 1698431365
transform 1 0 37184 0 1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1353_
timestamp 1698431365
transform 1 0 38304 0 1 6272
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1354_
timestamp 1698431365
transform 1 0 25984 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or4_2  _1355_
timestamp 1698431365
transform 1 0 26656 0 1 12544
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1356_
timestamp 1698431365
transform 1 0 34496 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1357_
timestamp 1698431365
transform 1 0 37072 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1358_
timestamp 1698431365
transform -1 0 39312 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1359_
timestamp 1698431365
transform 1 0 35504 0 1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1360_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 34944 0 1 9408
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1361_
timestamp 1698431365
transform -1 0 36624 0 1 7840
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1362_
timestamp 1698431365
transform 1 0 39648 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1363_
timestamp 1698431365
transform 1 0 38976 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1364_
timestamp 1698431365
transform 1 0 39984 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1365_
timestamp 1698431365
transform 1 0 40320 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1366_
timestamp 1698431365
transform 1 0 40768 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1367_
timestamp 1698431365
transform 1 0 44016 0 -1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _1368_
timestamp 1698431365
transform 1 0 36064 0 -1 9408
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1369_
timestamp 1698431365
transform 1 0 44576 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1370_
timestamp 1698431365
transform -1 0 47712 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1371_
timestamp 1698431365
transform -1 0 46144 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1372_
timestamp 1698431365
transform 1 0 44800 0 1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1373_
timestamp 1698431365
transform 1 0 44576 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1374_
timestamp 1698431365
transform 1 0 44800 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1375_
timestamp 1698431365
transform -1 0 48160 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1376_
timestamp 1698431365
transform -1 0 35392 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1377_
timestamp 1698431365
transform 1 0 34048 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1378_
timestamp 1698431365
transform 1 0 35392 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1379_
timestamp 1698431365
transform -1 0 35392 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_2  _1380_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 32928 0 -1 17248
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1381_
timestamp 1698431365
transform -1 0 33712 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1382_
timestamp 1698431365
transform 1 0 32928 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1383_
timestamp 1698431365
transform 1 0 16576 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1384_
timestamp 1698431365
transform -1 0 33600 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1385_
timestamp 1698431365
transform 1 0 18816 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1386_
timestamp 1698431365
transform -1 0 19936 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1387_
timestamp 1698431365
transform -1 0 26880 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1388_
timestamp 1698431365
transform 1 0 22064 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1389_
timestamp 1698431365
transform -1 0 32480 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1390_
timestamp 1698431365
transform -1 0 34832 0 1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1391_
timestamp 1698431365
transform -1 0 34272 0 1 6272
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1392_
timestamp 1698431365
transform -1 0 35504 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1393_
timestamp 1698431365
transform -1 0 32144 0 -1 17248
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1394_
timestamp 1698431365
transform -1 0 30576 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1395_
timestamp 1698431365
transform -1 0 22176 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1396_
timestamp 1698431365
transform 1 0 20608 0 -1 7840
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1397_
timestamp 1698431365
transform 1 0 20272 0 -1 6272
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1398_
timestamp 1698431365
transform 1 0 19600 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1399_
timestamp 1698431365
transform -1 0 33600 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1400_
timestamp 1698431365
transform -1 0 32144 0 1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1401_
timestamp 1698431365
transform -1 0 31920 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1402_
timestamp 1698431365
transform 1 0 26992 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1403_
timestamp 1698431365
transform -1 0 28000 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1404_
timestamp 1698431365
transform -1 0 27888 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1405_
timestamp 1698431365
transform 1 0 26096 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1406_
timestamp 1698431365
transform 1 0 25648 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1407_
timestamp 1698431365
transform -1 0 32144 0 -1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1408_
timestamp 1698431365
transform -1 0 31248 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1409_
timestamp 1698431365
transform 1 0 29680 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1410_
timestamp 1698431365
transform -1 0 31248 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1411_
timestamp 1698431365
transform -1 0 30576 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1412_
timestamp 1698431365
transform 1 0 29232 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1413_
timestamp 1698431365
transform 1 0 28784 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1414_
timestamp 1698431365
transform -1 0 35728 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1415_
timestamp 1698431365
transform 1 0 25648 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1416_
timestamp 1698431365
transform -1 0 24304 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1417_
timestamp 1698431365
transform 1 0 22736 0 1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _1418_
timestamp 1698431365
transform -1 0 27776 0 -1 29792
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1419_
timestamp 1698431365
transform -1 0 35168 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1420_
timestamp 1698431365
transform 1 0 27104 0 1 43904
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1421_
timestamp 1698431365
transform -1 0 30688 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1422_
timestamp 1698431365
transform 1 0 37072 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1423_
timestamp 1698431365
transform -1 0 35952 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1424_
timestamp 1698431365
transform 1 0 29232 0 -1 39200
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1425_
timestamp 1698431365
transform -1 0 27888 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1426_
timestamp 1698431365
transform -1 0 41664 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1427_
timestamp 1698431365
transform -1 0 40544 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1428_
timestamp 1698431365
transform 1 0 38640 0 1 40768
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1429_
timestamp 1698431365
transform 1 0 35952 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1430_
timestamp 1698431365
transform -1 0 42336 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1431_
timestamp 1698431365
transform 1 0 41104 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1432_
timestamp 1698431365
transform 1 0 42672 0 1 42336
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1433_
timestamp 1698431365
transform -1 0 41440 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1434_
timestamp 1698431365
transform 1 0 44800 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1435_
timestamp 1698431365
transform 1 0 35616 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1436_
timestamp 1698431365
transform -1 0 44464 0 1 36064
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1437_
timestamp 1698431365
transform -1 0 45360 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1438_
timestamp 1698431365
transform -1 0 44464 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1439_
timestamp 1698431365
transform 1 0 41104 0 1 36064
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1440_
timestamp 1698431365
transform -1 0 40880 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1441_
timestamp 1698431365
transform -1 0 38080 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1442_
timestamp 1698431365
transform 1 0 34384 0 -1 36064
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1443_
timestamp 1698431365
transform -1 0 34272 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1444_
timestamp 1698431365
transform -1 0 39872 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1445_
timestamp 1698431365
transform 1 0 37632 0 -1 36064
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1446_
timestamp 1698431365
transform 1 0 37296 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1447_
timestamp 1698431365
transform 1 0 25088 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1448_
timestamp 1698431365
transform -1 0 44464 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1449_
timestamp 1698431365
transform 1 0 45808 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1450_
timestamp 1698431365
transform -1 0 48160 0 -1 15680
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1451_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 43120 0 -1 17248
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1452_
timestamp 1698431365
transform -1 0 37072 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_4  _1453_
timestamp 1698431365
transform 1 0 36512 0 -1 14112
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1454_
timestamp 1698431365
transform -1 0 38416 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1455_
timestamp 1698431365
transform 1 0 36848 0 1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1456_
timestamp 1698431365
transform -1 0 44016 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1457_
timestamp 1698431365
transform -1 0 43904 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1458_
timestamp 1698431365
transform -1 0 45248 0 -1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1459_
timestamp 1698431365
transform 1 0 42560 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1460_
timestamp 1698431365
transform -1 0 38304 0 -1 18816
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1461_
timestamp 1698431365
transform -1 0 39424 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1462_
timestamp 1698431365
transform 1 0 34048 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1463_
timestamp 1698431365
transform 1 0 37408 0 -1 15680
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1464_
timestamp 1698431365
transform 1 0 37744 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1465_
timestamp 1698431365
transform -1 0 41104 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_4  _1466_
timestamp 1698431365
transform 1 0 36848 0 1 17248
box -86 -86 4902 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1467_
timestamp 1698431365
transform -1 0 27776 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1468_
timestamp 1698431365
transform -1 0 26096 0 -1 18816
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1469_
timestamp 1698431365
transform -1 0 24528 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _1470_
timestamp 1698431365
transform -1 0 27552 0 1 28224
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1471_
timestamp 1698431365
transform 1 0 32928 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1472_
timestamp 1698431365
transform 1 0 33936 0 1 42336
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1473_
timestamp 1698431365
transform -1 0 31808 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1474_
timestamp 1698431365
transform 1 0 34048 0 1 40768
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1475_
timestamp 1698431365
transform 1 0 33376 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1476_
timestamp 1698431365
transform 1 0 41216 0 1 40768
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1477_
timestamp 1698431365
transform 1 0 40544 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1478_
timestamp 1698431365
transform -1 0 44128 0 -1 40768
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1479_
timestamp 1698431365
transform -1 0 44464 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1480_
timestamp 1698431365
transform 1 0 32928 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1481_
timestamp 1698431365
transform 1 0 42784 0 1 37632
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1482_
timestamp 1698431365
transform 1 0 41216 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1483_
timestamp 1698431365
transform -1 0 42560 0 -1 32928
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1484_
timestamp 1698431365
transform 1 0 44800 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1485_
timestamp 1698431365
transform 1 0 32256 0 1 34496
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1486_
timestamp 1698431365
transform -1 0 32592 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1487_
timestamp 1698431365
transform 1 0 34608 0 1 32928
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1488_
timestamp 1698431365
transform 1 0 34384 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1489_
timestamp 1698431365
transform 1 0 40768 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1490_
timestamp 1698431365
transform -1 0 39200 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1491_
timestamp 1698431365
transform -1 0 27104 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1492_
timestamp 1698431365
transform -1 0 26208 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1493_
timestamp 1698431365
transform -1 0 28560 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1494_
timestamp 1698431365
transform -1 0 28672 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _1495_
timestamp 1698431365
transform -1 0 27104 0 -1 17248
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1496_
timestamp 1698431365
transform 1 0 28672 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1497_
timestamp 1698431365
transform 1 0 28112 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1498_
timestamp 1698431365
transform 1 0 43904 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1499_
timestamp 1698431365
transform -1 0 36176 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1500_
timestamp 1698431365
transform 1 0 29456 0 1 17248
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1501_
timestamp 1698431365
transform 1 0 29904 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1502_
timestamp 1698431365
transform 1 0 29008 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1503_
timestamp 1698431365
transform -1 0 31248 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1504_
timestamp 1698431365
transform -1 0 31024 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1505_
timestamp 1698431365
transform 1 0 29344 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1506_
timestamp 1698431365
transform 1 0 29792 0 -1 18816
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1507_
timestamp 1698431365
transform -1 0 30688 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1508_
timestamp 1698431365
transform 1 0 29120 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1509_
timestamp 1698431365
transform 1 0 31920 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1510_
timestamp 1698431365
transform 1 0 31024 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1511_
timestamp 1698431365
transform 1 0 24976 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1512_
timestamp 1698431365
transform -1 0 36624 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1513_
timestamp 1698431365
transform 1 0 29008 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1514_
timestamp 1698431365
transform -1 0 34048 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1515_
timestamp 1698431365
transform 1 0 35952 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1516_
timestamp 1698431365
transform 1 0 32704 0 1 18816
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1517_
timestamp 1698431365
transform -1 0 30464 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1518_
timestamp 1698431365
transform 1 0 29008 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1519_
timestamp 1698431365
transform -1 0 32256 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1520_
timestamp 1698431365
transform 1 0 30800 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1521_
timestamp 1698431365
transform -1 0 34832 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1522_
timestamp 1698431365
transform 1 0 29904 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1523_
timestamp 1698431365
transform -1 0 34720 0 1 18816
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1524_
timestamp 1698431365
transform -1 0 31360 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1525_
timestamp 1698431365
transform 1 0 29008 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1526_
timestamp 1698431365
transform 1 0 30128 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1527_
timestamp 1698431365
transform 1 0 30688 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1528_
timestamp 1698431365
transform -1 0 33152 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1529_
timestamp 1698431365
transform 1 0 31584 0 -1 18816
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1530_
timestamp 1698431365
transform -1 0 32592 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1531_
timestamp 1698431365
transform 1 0 25312 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1532_
timestamp 1698431365
transform -1 0 28224 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1533_
timestamp 1698431365
transform 1 0 25984 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1534_
timestamp 1698431365
transform 1 0 31024 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1535_
timestamp 1698431365
transform 1 0 31696 0 1 18816
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1536_
timestamp 1698431365
transform -1 0 32368 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1537_
timestamp 1698431365
transform 1 0 25872 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1538_
timestamp 1698431365
transform -1 0 29120 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1539_
timestamp 1698431365
transform 1 0 26208 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1540_
timestamp 1698431365
transform -1 0 42560 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1541_
timestamp 1698431365
transform -1 0 40432 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1542_
timestamp 1698431365
transform -1 0 42560 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1543_
timestamp 1698431365
transform -1 0 40544 0 -1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1544_
timestamp 1698431365
transform 1 0 38864 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1545_
timestamp 1698431365
transform 1 0 40768 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1546_
timestamp 1698431365
transform -1 0 40544 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _1547_
timestamp 1698431365
transform 1 0 40544 0 1 15680
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1548_
timestamp 1698431365
transform 1 0 40320 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1549_
timestamp 1698431365
transform -1 0 43008 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1550_
timestamp 1698431365
transform -1 0 45808 0 1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1551_
timestamp 1698431365
transform -1 0 42560 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1552_
timestamp 1698431365
transform 1 0 42112 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1553_
timestamp 1698431365
transform 1 0 41104 0 -1 18816
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1554_
timestamp 1698431365
transform 1 0 42448 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _1555_
timestamp 1698431365
transform -1 0 41888 0 1 14112
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1556_
timestamp 1698431365
transform -1 0 41664 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1557_
timestamp 1698431365
transform -1 0 39984 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1558_
timestamp 1698431365
transform 1 0 41104 0 1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1559_
timestamp 1698431365
transform 1 0 44688 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1560_
timestamp 1698431365
transform -1 0 39872 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1561_
timestamp 1698431365
transform -1 0 39200 0 -1 9408
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1562_
timestamp 1698431365
transform 1 0 22400 0 -1 21952
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1563_
timestamp 1698431365
transform 1 0 21280 0 -1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1564_
timestamp 1698431365
transform -1 0 22960 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1565_
timestamp 1698431365
transform -1 0 6944 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1566_
timestamp 1698431365
transform 1 0 21280 0 1 43904
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1567_
timestamp 1698431365
transform -1 0 21952 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1568_
timestamp 1698431365
transform 1 0 25088 0 -1 42336
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1569_
timestamp 1698431365
transform -1 0 24752 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1570_
timestamp 1698431365
transform 1 0 22288 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1571_
timestamp 1698431365
transform 1 0 37632 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1572_
timestamp 1698431365
transform 1 0 37968 0 -1 29792
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1573_
timestamp 1698431365
transform 1 0 37296 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1574_
timestamp 1698431365
transform -1 0 44464 0 1 28224
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1575_
timestamp 1698431365
transform -1 0 45360 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1576_
timestamp 1698431365
transform 1 0 46704 0 -1 21952
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1577_
timestamp 1698431365
transform 1 0 44800 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1578_
timestamp 1698431365
transform 1 0 46592 0 -1 31360
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1579_
timestamp 1698431365
transform -1 0 46592 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1580_
timestamp 1698431365
transform 1 0 30800 0 1 26656
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1581_
timestamp 1698431365
transform -1 0 30800 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1582_
timestamp 1698431365
transform 1 0 34832 0 1 28224
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1583_
timestamp 1698431365
transform -1 0 34944 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1584_
timestamp 1698431365
transform 1 0 22400 0 1 21952
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1585_
timestamp 1698431365
transform 1 0 22960 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1586_
timestamp 1698431365
transform -1 0 23744 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1587_
timestamp 1698431365
transform 1 0 25088 0 -1 45472
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1588_
timestamp 1698431365
transform 1 0 24416 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1589_
timestamp 1698431365
transform 1 0 25648 0 -1 40768
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1590_
timestamp 1698431365
transform -1 0 25760 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1591_
timestamp 1698431365
transform -1 0 23744 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1592_
timestamp 1698431365
transform 1 0 34944 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1593_
timestamp 1698431365
transform 1 0 36960 0 1 40768
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1594_
timestamp 1698431365
transform 1 0 35952 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1595_
timestamp 1698431365
transform 1 0 44688 0 1 43904
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1596_
timestamp 1698431365
transform -1 0 39424 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1597_
timestamp 1698431365
transform 1 0 42784 0 1 39200
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1598_
timestamp 1698431365
transform 1 0 43008 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1599_
timestamp 1698431365
transform 1 0 40768 0 -1 40768
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1600_
timestamp 1698431365
transform -1 0 41440 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1601_
timestamp 1698431365
transform 1 0 33824 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1602_
timestamp 1698431365
transform 1 0 33824 0 -1 39200
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1603_
timestamp 1698431365
transform -1 0 33600 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1604_
timestamp 1698431365
transform 1 0 36960 0 1 37632
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1605_
timestamp 1698431365
transform 1 0 35952 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1606_
timestamp 1698431365
transform 1 0 31024 0 -1 45472
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1607_
timestamp 1698431365
transform -1 0 31808 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1608_
timestamp 1698431365
transform 1 0 38752 0 -1 43904
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1609_
timestamp 1698431365
transform -1 0 35616 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1610_
timestamp 1698431365
transform 1 0 23184 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1611_
timestamp 1698431365
transform -1 0 42560 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1612_
timestamp 1698431365
transform -1 0 40544 0 -1 39200
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1613_
timestamp 1698431365
transform 1 0 44800 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1614_
timestamp 1698431365
transform -1 0 38976 0 1 39200
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1615_
timestamp 1698431365
transform -1 0 43232 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1616_
timestamp 1698431365
transform 1 0 46592 0 1 43904
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1617_
timestamp 1698431365
transform 1 0 44800 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1618_
timestamp 1698431365
transform 1 0 46480 0 -1 39200
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1619_
timestamp 1698431365
transform -1 0 46480 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1620_
timestamp 1698431365
transform -1 0 33152 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1621_
timestamp 1698431365
transform 1 0 31024 0 -1 36064
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1622_
timestamp 1698431365
transform -1 0 29680 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1623_
timestamp 1698431365
transform 1 0 30912 0 -1 32928
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1624_
timestamp 1698431365
transform 1 0 28336 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1625_
timestamp 1698431365
transform 1 0 30688 0 -1 40768
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1626_
timestamp 1698431365
transform -1 0 30912 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1627_
timestamp 1698431365
transform 1 0 30800 0 -1 37632
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1628_
timestamp 1698431365
transform -1 0 31584 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1629_
timestamp 1698431365
transform -1 0 44912 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1630_
timestamp 1698431365
transform -1 0 40544 0 -1 32928
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1631_
timestamp 1698431365
transform -1 0 40992 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1632_
timestamp 1698431365
transform 1 0 40880 0 -1 31360
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1633_
timestamp 1698431365
transform 1 0 38192 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1634_
timestamp 1698431365
transform -1 0 44464 0 1 31360
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1635_
timestamp 1698431365
transform 1 0 44688 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1636_
timestamp 1698431365
transform 1 0 42560 0 1 34496
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1637_
timestamp 1698431365
transform 1 0 40992 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1638_
timestamp 1698431365
transform 1 0 23408 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1639_
timestamp 1698431365
transform 1 0 30464 0 -1 31360
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1640_
timestamp 1698431365
transform 1 0 29344 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1641_
timestamp 1698431365
transform 1 0 34048 0 -1 31360
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1642_
timestamp 1698431365
transform -1 0 33936 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1643_
timestamp 1698431365
transform 1 0 4816 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1644_
timestamp 1698431365
transform 1 0 12208 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1645_
timestamp 1698431365
transform -1 0 19600 0 1 7840
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1646_
timestamp 1698431365
transform 1 0 10192 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1647_
timestamp 1698431365
transform -1 0 16576 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1648_
timestamp 1698431365
transform -1 0 10752 0 1 17248
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1649_
timestamp 1698431365
transform -1 0 11088 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1650_
timestamp 1698431365
transform 1 0 5488 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1651_
timestamp 1698431365
transform 1 0 8848 0 1 12544
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1652_
timestamp 1698431365
transform -1 0 11200 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1653_
timestamp 1698431365
transform 1 0 9632 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _1654_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 10080 0 1 9408
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1655_
timestamp 1698431365
transform 1 0 11200 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1656_
timestamp 1698431365
transform 1 0 4816 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1657_
timestamp 1698431365
transform 1 0 16128 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1658_
timestamp 1698431365
transform -1 0 37296 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1659_
timestamp 1698431365
transform 1 0 14784 0 -1 9408
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1660_
timestamp 1698431365
transform 1 0 6384 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1661_
timestamp 1698431365
transform 1 0 12432 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1662_
timestamp 1698431365
transform -1 0 14448 0 1 7840
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1663_
timestamp 1698431365
transform 1 0 27888 0 -1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1664_
timestamp 1698431365
transform 1 0 29232 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1665_
timestamp 1698431365
transform -1 0 29568 0 1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1666_
timestamp 1698431365
transform -1 0 29904 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1667_
timestamp 1698431365
transform 1 0 28336 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1668_
timestamp 1698431365
transform -1 0 13104 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1669_
timestamp 1698431365
transform -1 0 16800 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1670_
timestamp 1698431365
transform 1 0 17696 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1671_
timestamp 1698431365
transform 1 0 18592 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and3_2  _1672_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 9856 0 -1 14112
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1673_
timestamp 1698431365
transform -1 0 12432 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1674_
timestamp 1698431365
transform 1 0 11312 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1675_
timestamp 1698431365
transform 1 0 10192 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1676_
timestamp 1698431365
transform -1 0 11872 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1677_
timestamp 1698431365
transform 1 0 10192 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _1678_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 14560 0 -1 25088
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _1679_
timestamp 1698431365
transform 1 0 13328 0 1 20384
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _1680_
timestamp 1698431365
transform -1 0 14672 0 -1 17248
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1681_
timestamp 1698431365
transform 1 0 19488 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1682_
timestamp 1698431365
transform 1 0 18368 0 -1 18816
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1683_
timestamp 1698431365
transform -1 0 18928 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1684_
timestamp 1698431365
transform 1 0 9520 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1685_
timestamp 1698431365
transform 1 0 10416 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_1  _1686_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 12544 0 1 20384
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1687_
timestamp 1698431365
transform -1 0 13888 0 -1 18816
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1688_
timestamp 1698431365
transform 1 0 13552 0 -1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1689_
timestamp 1698431365
transform 1 0 16352 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1690_
timestamp 1698431365
transform 1 0 15904 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1691_
timestamp 1698431365
transform 1 0 16128 0 1 18816
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1692_
timestamp 1698431365
transform 1 0 17136 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1693_
timestamp 1698431365
transform 1 0 18704 0 1 15680
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1694_
timestamp 1698431365
transform 1 0 18816 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1695_
timestamp 1698431365
transform -1 0 13104 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai222_2  _1696_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 10528 0 -1 20384
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1697_
timestamp 1698431365
transform -1 0 17024 0 -1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1698_
timestamp 1698431365
transform 1 0 16464 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1699_
timestamp 1698431365
transform 1 0 18032 0 -1 15680
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1700_
timestamp 1698431365
transform -1 0 18480 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1701_
timestamp 1698431365
transform -1 0 11872 0 1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _1702_
timestamp 1698431365
transform -1 0 15904 0 1 23520
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1703_
timestamp 1698431365
transform -1 0 16912 0 1 20384
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _1704_
timestamp 1698431365
transform -1 0 14560 0 1 18816
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1705_
timestamp 1698431365
transform 1 0 20160 0 -1 20384
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1706_
timestamp 1698431365
transform 1 0 21168 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1707_
timestamp 1698431365
transform -1 0 15568 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1708_
timestamp 1698431365
transform 1 0 15008 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1709_
timestamp 1698431365
transform 1 0 15904 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1710_
timestamp 1698431365
transform 1 0 14224 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1711_
timestamp 1698431365
transform 1 0 14336 0 1 20384
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1712_
timestamp 1698431365
transform 1 0 11200 0 -1 26656
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _1713_
timestamp 1698431365
transform 1 0 15904 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1714_
timestamp 1698431365
transform 1 0 22176 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1715_
timestamp 1698431365
transform 1 0 26208 0 -1 23520
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1716_
timestamp 1698431365
transform 1 0 26320 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1717_
timestamp 1698431365
transform 1 0 14560 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _1718_
timestamp 1698431365
transform 1 0 10528 0 1 25088
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1719_
timestamp 1698431365
transform -1 0 18928 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1720_
timestamp 1698431365
transform -1 0 18704 0 -1 26656
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1721_
timestamp 1698431365
transform 1 0 26432 0 -1 26656
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1722_
timestamp 1698431365
transform -1 0 27664 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1723_
timestamp 1698431365
transform 1 0 16464 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_2  _1724_
timestamp 1698431365
transform 1 0 10752 0 -1 23520
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1725_
timestamp 1698431365
transform 1 0 17696 0 1 23520
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1726_
timestamp 1698431365
transform 1 0 23072 0 -1 23520
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1727_
timestamp 1698431365
transform -1 0 23520 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1728_
timestamp 1698431365
transform 1 0 17360 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _1729_
timestamp 1698431365
transform 1 0 9408 0 -1 25088
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1730_
timestamp 1698431365
transform 1 0 17808 0 1 25088
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1731_
timestamp 1698431365
transform 1 0 23184 0 -1 26656
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1732_
timestamp 1698431365
transform -1 0 24752 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1733_
timestamp 1698431365
transform 1 0 13328 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1734_
timestamp 1698431365
transform 1 0 16352 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1735_
timestamp 1698431365
transform 1 0 15008 0 -1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1736_
timestamp 1698431365
transform -1 0 16800 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1737_
timestamp 1698431365
transform -1 0 15008 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1738_
timestamp 1698431365
transform 1 0 19152 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1739_
timestamp 1698431365
transform -1 0 19152 0 -1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1740_
timestamp 1698431365
transform 1 0 26320 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1741_
timestamp 1698431365
transform 1 0 26656 0 1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1742_
timestamp 1698431365
transform 1 0 29008 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1743_
timestamp 1698431365
transform 1 0 29008 0 1 42336
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1744_
timestamp 1698431365
transform -1 0 27552 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1745_
timestamp 1698431365
transform 1 0 28000 0 -1 40768
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1746_
timestamp 1698431365
transform 1 0 27216 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1747_
timestamp 1698431365
transform 1 0 37408 0 1 31360
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1748_
timestamp 1698431365
transform -1 0 37520 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1749_
timestamp 1698431365
transform 1 0 40880 0 1 28224
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1750_
timestamp 1698431365
transform 1 0 41104 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1751_
timestamp 1698431365
transform 1 0 29456 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1752_
timestamp 1698431365
transform 1 0 46256 0 -1 23520
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1753_
timestamp 1698431365
transform 1 0 44128 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1754_
timestamp 1698431365
transform -1 0 47936 0 -1 28224
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1755_
timestamp 1698431365
transform 1 0 44800 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1756_
timestamp 1698431365
transform 1 0 30464 0 1 28224
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1757_
timestamp 1698431365
transform -1 0 29904 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1758_
timestamp 1698431365
transform 1 0 34272 0 1 29792
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1759_
timestamp 1698431365
transform 1 0 32928 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1760_
timestamp 1698431365
transform 1 0 12656 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1761_
timestamp 1698431365
transform -1 0 22288 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1762_
timestamp 1698431365
transform -1 0 14224 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1763_
timestamp 1698431365
transform 1 0 17024 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1764_
timestamp 1698431365
transform 1 0 16464 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1765_
timestamp 1698431365
transform -1 0 9184 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1766_
timestamp 1698431365
transform -1 0 23184 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1767_
timestamp 1698431365
transform -1 0 15120 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1768_
timestamp 1698431365
transform -1 0 10528 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1769_
timestamp 1698431365
transform 1 0 7168 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _1770_
timestamp 1698431365
transform -1 0 10752 0 -1 23520
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1771_
timestamp 1698431365
transform -1 0 24864 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1772_
timestamp 1698431365
transform -1 0 6608 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1773_
timestamp 1698431365
transform 1 0 5936 0 1 21952
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1774_
timestamp 1698431365
transform 1 0 18816 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1775_
timestamp 1698431365
transform -1 0 28336 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1776_
timestamp 1698431365
transform 1 0 22624 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1777_
timestamp 1698431365
transform 1 0 23856 0 1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1778_
timestamp 1698431365
transform 1 0 22736 0 1 6272
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1779_
timestamp 1698431365
transform 1 0 10976 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1780_
timestamp 1698431365
transform -1 0 10304 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1781_
timestamp 1698431365
transform -1 0 18256 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1782_
timestamp 1698431365
transform -1 0 17808 0 -1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1783_
timestamp 1698431365
transform -1 0 18368 0 -1 4704
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1784_
timestamp 1698431365
transform -1 0 18704 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1785_
timestamp 1698431365
transform -1 0 14112 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1786_
timestamp 1698431365
transform 1 0 6832 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1787_
timestamp 1698431365
transform 1 0 8400 0 -1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1788_
timestamp 1698431365
transform 1 0 7280 0 -1 6272
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1789_
timestamp 1698431365
transform -1 0 7728 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1790_
timestamp 1698431365
transform 1 0 5936 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1791_
timestamp 1698431365
transform 1 0 7280 0 -1 4704
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1792_
timestamp 1698431365
transform 1 0 6160 0 1 4704
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1793_
timestamp 1698431365
transform 1 0 5488 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1794_
timestamp 1698431365
transform 1 0 10304 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1795_
timestamp 1698431365
transform -1 0 12320 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1796_
timestamp 1698431365
transform 1 0 7840 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1797_
timestamp 1698431365
transform 1 0 10864 0 1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1798_
timestamp 1698431365
transform 1 0 10528 0 1 4704
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1799_
timestamp 1698431365
transform 1 0 6384 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1800_
timestamp 1698431365
transform 1 0 8288 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1801_
timestamp 1698431365
transform 1 0 11648 0 -1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1802_
timestamp 1698431365
transform -1 0 14448 0 1 4704
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1803_
timestamp 1698431365
transform 1 0 8736 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1804_
timestamp 1698431365
transform -1 0 16912 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1805_
timestamp 1698431365
transform 1 0 12096 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1806_
timestamp 1698431365
transform -1 0 13440 0 -1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1807_
timestamp 1698431365
transform -1 0 13104 0 1 6272
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1808_
timestamp 1698431365
transform -1 0 11872 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1809_
timestamp 1698431365
transform -1 0 15792 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1810_
timestamp 1698431365
transform 1 0 12992 0 -1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1811_
timestamp 1698431365
transform -1 0 15680 0 1 4704
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1812_
timestamp 1698431365
transform 1 0 42560 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1813_
timestamp 1698431365
transform -1 0 44464 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1814_
timestamp 1698431365
transform 1 0 39872 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1815_
timestamp 1698431365
transform 1 0 39984 0 -1 4704
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1816_
timestamp 1698431365
transform 1 0 42448 0 1 4704
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1817_
timestamp 1698431365
transform -1 0 40544 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1818_
timestamp 1698431365
transform -1 0 45136 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1819_
timestamp 1698431365
transform -1 0 42672 0 1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1820_
timestamp 1698431365
transform -1 0 44464 0 1 6272
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1821_
timestamp 1698431365
transform -1 0 43120 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1822_
timestamp 1698431365
transform 1 0 43120 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1823_
timestamp 1698431365
transform 1 0 43680 0 -1 4704
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1824_
timestamp 1698431365
transform -1 0 44464 0 1 7840
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1825_
timestamp 1698431365
transform 1 0 45248 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1826_
timestamp 1698431365
transform 1 0 31920 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1827_
timestamp 1698431365
transform -1 0 48384 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1828_
timestamp 1698431365
transform 1 0 38640 0 1 4704
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1829_
timestamp 1698431365
transform 1 0 46592 0 -1 6272
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1830_
timestamp 1698431365
transform 1 0 42672 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1831_
timestamp 1698431365
transform -1 0 30800 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1832_
timestamp 1698431365
transform 1 0 30800 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1833_
timestamp 1698431365
transform 1 0 31472 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1834_
timestamp 1698431365
transform 1 0 33600 0 -1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1835_
timestamp 1698431365
transform -1 0 36624 0 1 4704
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1836_
timestamp 1698431365
transform 1 0 36176 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1837_
timestamp 1698431365
transform 1 0 31136 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1838_
timestamp 1698431365
transform -1 0 37968 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1839_
timestamp 1698431365
transform -1 0 35504 0 1 4704
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1840_
timestamp 1698431365
transform -1 0 36512 0 -1 4704
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1841_
timestamp 1698431365
transform 1 0 37968 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1842_
timestamp 1698431365
transform -1 0 35616 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1843_
timestamp 1698431365
transform -1 0 34720 0 -1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1844_
timestamp 1698431365
transform -1 0 34496 0 -1 4704
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1845_
timestamp 1698431365
transform -1 0 35168 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1846_
timestamp 1698431365
transform 1 0 21280 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1847_
timestamp 1698431365
transform 1 0 23632 0 -1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1848_
timestamp 1698431365
transform 1 0 21840 0 -1 4704
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1849_
timestamp 1698431365
transform -1 0 20384 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1850_
timestamp 1698431365
transform -1 0 26992 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1851_
timestamp 1698431365
transform -1 0 24864 0 -1 4704
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1852_
timestamp 1698431365
transform -1 0 26208 0 -1 4704
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1853_
timestamp 1698431365
transform -1 0 25536 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1854_
timestamp 1698431365
transform -1 0 33376 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1855_
timestamp 1698431365
transform -1 0 30688 0 -1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1856_
timestamp 1698431365
transform -1 0 30128 0 1 4704
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1857_
timestamp 1698431365
transform -1 0 28784 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1858_
timestamp 1698431365
transform -1 0 22960 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1859_
timestamp 1698431365
transform 1 0 21728 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _1860_
timestamp 1698431365
transform 1 0 21952 0 -1 6272
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1861_
timestamp 1698431365
transform -1 0 41776 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1862_
timestamp 1698431365
transform -1 0 35840 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1863_
timestamp 1698431365
transform 1 0 34944 0 -1 23520
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1864_
timestamp 1698431365
transform 1 0 35392 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _1865_
timestamp 1698431365
transform 1 0 36064 0 -1 17248
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1866_
timestamp 1698431365
transform 1 0 38192 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1867_
timestamp 1698431365
transform 1 0 34272 0 -1 25088
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1868_
timestamp 1698431365
transform -1 0 34272 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1869_
timestamp 1698431365
transform 1 0 34608 0 1 21952
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1870_
timestamp 1698431365
transform 1 0 34496 0 1 20384
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1871_
timestamp 1698431365
transform 1 0 33824 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1872_
timestamp 1698431365
transform 1 0 38192 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1873_
timestamp 1698431365
transform 1 0 34720 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1874_
timestamp 1698431365
transform 1 0 36848 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _1875_
timestamp 1698431365
transform 1 0 37744 0 -1 21952
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1876_
timestamp 1698431365
transform 1 0 38864 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1877_
timestamp 1698431365
transform 1 0 39536 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1878_
timestamp 1698431365
transform 1 0 38640 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1879_
timestamp 1698431365
transform -1 0 43008 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1880_
timestamp 1698431365
transform 1 0 41440 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _1881_
timestamp 1698431365
transform 1 0 41664 0 1 20384
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1882_
timestamp 1698431365
transform 1 0 40768 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1883_
timestamp 1698431365
transform -1 0 43904 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1884_
timestamp 1698431365
transform 1 0 42336 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1885_
timestamp 1698431365
transform -1 0 43008 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _1886_
timestamp 1698431365
transform -1 0 42112 0 1 21952
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1887_
timestamp 1698431365
transform 1 0 37520 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1888_
timestamp 1698431365
transform 1 0 43456 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1889_
timestamp 1698431365
transform 1 0 42560 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1890_
timestamp 1698431365
transform -1 0 42896 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _1891_
timestamp 1698431365
transform -1 0 42000 0 1 23520
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1892_
timestamp 1698431365
transform 1 0 42896 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1893_
timestamp 1698431365
transform 1 0 43008 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1894_
timestamp 1698431365
transform 1 0 40768 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _1895_
timestamp 1698431365
transform -1 0 43008 0 1 25088
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1896_
timestamp 1698431365
transform -1 0 37968 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1897_
timestamp 1698431365
transform -1 0 38864 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1898_
timestamp 1698431365
transform 1 0 38528 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _1899_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 40432 0 1 25088
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1900_
timestamp 1698431365
transform 1 0 39536 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1901_
timestamp 1698431365
transform 1 0 39424 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1902_
timestamp 1698431365
transform 1 0 22176 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1903_
timestamp 1698431365
transform 1 0 24528 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1904_
timestamp 1698431365
transform -1 0 31360 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1905_
timestamp 1698431365
transform 1 0 31360 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1906_
timestamp 1698431365
transform 1 0 30128 0 1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1907_
timestamp 1698431365
transform 1 0 29792 0 1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1908_
timestamp 1698431365
transform 1 0 30800 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1909_
timestamp 1698431365
transform -1 0 28672 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1910_
timestamp 1698431365
transform 1 0 25536 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1911_
timestamp 1698431365
transform 1 0 27440 0 -1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1912_
timestamp 1698431365
transform 1 0 22736 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1913_
timestamp 1698431365
transform -1 0 24528 0 1 15680
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1914_
timestamp 1698431365
transform -1 0 30800 0 -1 14112
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1915_
timestamp 1698431365
transform -1 0 24416 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1916_
timestamp 1698431365
transform -1 0 27440 0 -1 15680
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1917_
timestamp 1698431365
transform 1 0 23856 0 -1 15680
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1918_
timestamp 1698431365
transform 1 0 24640 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1919_
timestamp 1698431365
transform -1 0 26768 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1920_
timestamp 1698431365
transform 1 0 22848 0 1 14112
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1921_
timestamp 1698431365
transform 1 0 23184 0 -1 14112
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1922_
timestamp 1698431365
transform -1 0 23184 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _1923_
timestamp 1698431365
transform 1 0 26544 0 -1 14112
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1924_
timestamp 1698431365
transform -1 0 27664 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1925_
timestamp 1698431365
transform 1 0 24192 0 1 14112
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1926_
timestamp 1698431365
transform -1 0 24864 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1927_
timestamp 1698431365
transform -1 0 46368 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1928_
timestamp 1698431365
transform -1 0 44464 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1929_
timestamp 1698431365
transform 1 0 44688 0 1 18816
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1930_
timestamp 1698431365
transform -1 0 47824 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1931_
timestamp 1698431365
transform -1 0 46256 0 -1 18816
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1932_
timestamp 1698431365
transform 1 0 30016 0 1 14112
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1933_
timestamp 1698431365
transform 1 0 45696 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1934_
timestamp 1698431365
transform -1 0 40880 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1935_
timestamp 1698431365
transform 1 0 41888 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1936_
timestamp 1698431365
transform -1 0 38528 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _1937_
timestamp 1698431365
transform 1 0 38528 0 1 15680
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _1938_
timestamp 1698431365
transform 1 0 39312 0 -1 18816
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1939_
timestamp 1698431365
transform -1 0 42112 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1940_
timestamp 1698431365
transform 1 0 41104 0 -1 15680
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1941_
timestamp 1698431365
transform 1 0 46592 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1942_
timestamp 1698431365
transform 1 0 9184 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1943_
timestamp 1698431365
transform 1 0 9408 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1944_
timestamp 1698431365
transform 1 0 7616 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1945_
timestamp 1698431365
transform -1 0 6832 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1946_
timestamp 1698431365
transform -1 0 5600 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1947_
timestamp 1698431365
transform -1 0 4816 0 -1 9408
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1948_
timestamp 1698431365
transform -1 0 6832 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1949_
timestamp 1698431365
transform -1 0 5936 0 -1 9408
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1950_
timestamp 1698431365
transform 1 0 8064 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1951_
timestamp 1698431365
transform 1 0 6832 0 1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1952_
timestamp 1698431365
transform 1 0 7392 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1953_
timestamp 1698431365
transform 1 0 43232 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1954_
timestamp 1698431365
transform 1 0 44128 0 -1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1955_
timestamp 1698431365
transform 1 0 41328 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1956_
timestamp 1698431365
transform 1 0 31696 0 -1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1957_
timestamp 1698431365
transform 1 0 29008 0 1 10976
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1958_
timestamp 1698431365
transform 1 0 30576 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1959_
timestamp 1698431365
transform 1 0 28336 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1960_
timestamp 1698431365
transform 1 0 29232 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1961_
timestamp 1698431365
transform 1 0 30800 0 -1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1962_
timestamp 1698431365
transform 1 0 31024 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1963_
timestamp 1698431365
transform -1 0 17248 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1964_
timestamp 1698431365
transform 1 0 19824 0 1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1965_
timestamp 1698431365
transform 1 0 19264 0 1 25088
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1966_
timestamp 1698431365
transform 1 0 18928 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1967_
timestamp 1698431365
transform 1 0 19264 0 1 23520
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1968_
timestamp 1698431365
transform -1 0 19264 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1969_
timestamp 1698431365
transform 1 0 21952 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1970_
timestamp 1698431365
transform -1 0 23856 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1971_
timestamp 1698431365
transform 1 0 23744 0 -1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1972_
timestamp 1698431365
transform -1 0 16576 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1973_
timestamp 1698431365
transform -1 0 18256 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1974_
timestamp 1698431365
transform 1 0 21616 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1975_
timestamp 1698431365
transform 1 0 16352 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1976_
timestamp 1698431365
transform -1 0 18256 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1977_
timestamp 1698431365
transform -1 0 22960 0 1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1978_
timestamp 1698431365
transform 1 0 21280 0 1 29792
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1979_
timestamp 1698431365
transform 1 0 24304 0 -1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1980_
timestamp 1698431365
transform 1 0 18144 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1981_
timestamp 1698431365
transform -1 0 22512 0 -1 31360
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1982_
timestamp 1698431365
transform 1 0 17360 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1983_
timestamp 1698431365
transform -1 0 19824 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1984_
timestamp 1698431365
transform -1 0 20944 0 1 29792
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1985_
timestamp 1698431365
transform 1 0 20048 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1986_
timestamp 1698431365
transform 1 0 17248 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1987_
timestamp 1698431365
transform 1 0 22624 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1988_
timestamp 1698431365
transform 1 0 18256 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1989_
timestamp 1698431365
transform 1 0 22848 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1990_
timestamp 1698431365
transform -1 0 24640 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1991_
timestamp 1698431365
transform 1 0 24528 0 1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1992_
timestamp 1698431365
transform 1 0 23968 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1993_
timestamp 1698431365
transform 1 0 18256 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1994_
timestamp 1698431365
transform 1 0 22512 0 1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1995_
timestamp 1698431365
transform -1 0 23968 0 -1 37632
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1996_
timestamp 1698431365
transform -1 0 24528 0 -1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1997_
timestamp 1698431365
transform 1 0 24080 0 -1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1998_
timestamp 1698431365
transform 1 0 18256 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1999_
timestamp 1698431365
transform -1 0 18480 0 1 34496
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2000_
timestamp 1698431365
transform 1 0 17472 0 -1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2001_
timestamp 1698431365
transform -1 0 19376 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2002_
timestamp 1698431365
transform -1 0 23184 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2003_
timestamp 1698431365
transform 1 0 18816 0 -1 43904
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2004_
timestamp 1698431365
transform 1 0 18816 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2005_
timestamp 1698431365
transform -1 0 22064 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2006_
timestamp 1698431365
transform 1 0 21168 0 1 34496
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2007_
timestamp 1698431365
transform -1 0 22176 0 -1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2008_
timestamp 1698431365
transform 1 0 21056 0 -1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2009_
timestamp 1698431365
transform -1 0 20608 0 1 39200
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2010_
timestamp 1698431365
transform 1 0 18368 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2011_
timestamp 1698431365
transform -1 0 19264 0 1 39200
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2012_
timestamp 1698431365
transform 1 0 18144 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2013_
timestamp 1698431365
transform -1 0 18368 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2014_
timestamp 1698431365
transform 1 0 15568 0 1 39200
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2015_
timestamp 1698431365
transform 1 0 15568 0 1 40768
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2016_
timestamp 1698431365
transform -1 0 17584 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2017_
timestamp 1698431365
transform -1 0 18144 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2018_
timestamp 1698431365
transform 1 0 14448 0 -1 39200
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2019_
timestamp 1698431365
transform 1 0 15568 0 -1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2020_
timestamp 1698431365
transform 1 0 13440 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2021_
timestamp 1698431365
transform -1 0 14896 0 1 43904
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2022_
timestamp 1698431365
transform 1 0 13440 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2023_
timestamp 1698431365
transform -1 0 14448 0 1 39200
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2024_
timestamp 1698431365
transform 1 0 11984 0 1 40768
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2025_
timestamp 1698431365
transform -1 0 14112 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2026_
timestamp 1698431365
transform 1 0 9520 0 1 36064
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2027_
timestamp 1698431365
transform 1 0 9520 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2028_
timestamp 1698431365
transform -1 0 13104 0 1 43904
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2029_
timestamp 1698431365
transform 1 0 11200 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2030_
timestamp 1698431365
transform -1 0 6496 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2031_
timestamp 1698431365
transform -1 0 4704 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2032_
timestamp 1698431365
transform -1 0 8512 0 -1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2033_
timestamp 1698431365
transform -1 0 7952 0 1 34496
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2034_
timestamp 1698431365
transform 1 0 7168 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2035_
timestamp 1698431365
transform 1 0 2688 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2036_
timestamp 1698431365
transform -1 0 7952 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2037_
timestamp 1698431365
transform 1 0 7952 0 -1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _2038_
timestamp 1698431365
transform 1 0 7952 0 1 37632
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2039_
timestamp 1698431365
transform -1 0 4592 0 1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2040_
timestamp 1698431365
transform 1 0 3136 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2041_
timestamp 1698431365
transform -1 0 7168 0 -1 39200
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2042_
timestamp 1698431365
transform 1 0 5824 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2043_
timestamp 1698431365
transform -1 0 4144 0 -1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2044_
timestamp 1698431365
transform -1 0 4368 0 1 37632
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2045_
timestamp 1698431365
transform -1 0 7168 0 -1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2046_
timestamp 1698431365
transform 1 0 5488 0 -1 36064
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2047_
timestamp 1698431365
transform 1 0 2464 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2048_
timestamp 1698431365
transform 1 0 3696 0 -1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2049_
timestamp 1698431365
transform 1 0 4256 0 -1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2050_
timestamp 1698431365
transform 1 0 3248 0 -1 34496
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2051_
timestamp 1698431365
transform 1 0 2128 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2052_
timestamp 1698431365
transform -1 0 24752 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2053_
timestamp 1698431365
transform 1 0 10304 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2054_
timestamp 1698431365
transform 1 0 14672 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _2055_
timestamp 1698431365
transform -1 0 12432 0 1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2056_
timestamp 1698431365
transform -1 0 5264 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2057_
timestamp 1698431365
transform 1 0 3360 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2058_
timestamp 1698431365
transform -1 0 10304 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2059_
timestamp 1698431365
transform 1 0 15568 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2060_
timestamp 1698431365
transform 1 0 15232 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2061_
timestamp 1698431365
transform -1 0 15568 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2062_
timestamp 1698431365
transform 1 0 6608 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2063_
timestamp 1698431365
transform 1 0 5488 0 1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2064_
timestamp 1698431365
transform 1 0 4368 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2065_
timestamp 1698431365
transform 1 0 16688 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2066_
timestamp 1698431365
transform 1 0 10528 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2067_
timestamp 1698431365
transform -1 0 16688 0 1 43904
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _2068_
timestamp 1698431365
transform -1 0 16688 0 -1 43904
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2069_
timestamp 1698431365
transform 1 0 8176 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2070_
timestamp 1698431365
transform -1 0 8400 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2071_
timestamp 1698431365
transform 1 0 6048 0 1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2072_
timestamp 1698431365
transform 1 0 4816 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2073_
timestamp 1698431365
transform 1 0 4144 0 -1 31360
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2074_
timestamp 1698431365
transform -1 0 5040 0 1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2075_
timestamp 1698431365
transform -1 0 6608 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2076_
timestamp 1698431365
transform -1 0 8624 0 1 43904
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2077_
timestamp 1698431365
transform 1 0 7056 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _2078_
timestamp 1698431365
transform 1 0 43120 0 -1 18816
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2079_
timestamp 1698431365
transform 1 0 44128 0 -1 18816
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2080_
timestamp 1698431365
transform 1 0 46256 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2081_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 30016 0 -1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2082_
timestamp 1698431365
transform 1 0 25984 0 -1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2083_
timestamp 1698431365
transform 1 0 36512 0 -1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2084_
timestamp 1698431365
transform 1 0 37632 0 1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2085_
timestamp 1698431365
transform -1 0 45136 0 -1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2086_
timestamp 1698431365
transform 1 0 39088 0 1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2087_
timestamp 1698431365
transform 1 0 32368 0 1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2088_
timestamp 1698431365
transform 1 0 36848 0 1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2089_
timestamp 1698431365
transform 1 0 22512 0 1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2090_
timestamp 1698431365
transform 1 0 29456 0 -1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2091_
timestamp 1698431365
transform 1 0 32928 0 -1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2092_
timestamp 1698431365
transform -1 0 44688 0 -1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2093_
timestamp 1698431365
transform -1 0 44912 0 -1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2094_
timestamp 1698431365
transform 1 0 45136 0 1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2095_
timestamp 1698431365
transform 1 0 45136 0 1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2096_
timestamp 1698431365
transform 1 0 29008 0 1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2097_
timestamp 1698431365
transform -1 0 37072 0 -1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2098_
timestamp 1698431365
transform 1 0 25536 0 1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2099_
timestamp 1698431365
transform 1 0 29008 0 1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2100_
timestamp 1698431365
transform 1 0 31248 0 1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2101_
timestamp 1698431365
transform 1 0 30688 0 1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2102_
timestamp 1698431365
transform 1 0 29120 0 1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2103_
timestamp 1698431365
transform 1 0 25088 0 1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2104_
timestamp 1698431365
transform 1 0 25312 0 -1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2105_
timestamp 1698431365
transform 1 0 45136 0 1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2106_
timestamp 1698431365
transform 1 0 37968 0 1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2107_
timestamp 1698431365
transform 1 0 20608 0 -1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2108_
timestamp 1698431365
transform 1 0 23072 0 1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2109_
timestamp 1698431365
transform 1 0 36848 0 1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2110_
timestamp 1698431365
transform 1 0 42448 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2111_
timestamp 1698431365
transform 1 0 45136 0 1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2112_
timestamp 1698431365
transform 1 0 45136 0 1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2113_
timestamp 1698431365
transform 1 0 29344 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2114_
timestamp 1698431365
transform 1 0 33488 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2115_
timestamp 1698431365
transform -1 0 26208 0 1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2116_
timestamp 1698431365
transform 1 0 23744 0 1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2117_
timestamp 1698431365
transform 1 0 36176 0 -1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2118_
timestamp 1698431365
transform 1 0 36960 0 -1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2119_
timestamp 1698431365
transform 1 0 42336 0 -1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2120_
timestamp 1698431365
transform 1 0 38976 0 1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2121_
timestamp 1698431365
transform 1 0 31808 0 1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2122_
timestamp 1698431365
transform 1 0 35616 0 -1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2123_
timestamp 1698431365
transform 1 0 30128 0 1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2124_
timestamp 1698431365
transform 1 0 33712 0 -1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2125_
timestamp 1698431365
transform 1 0 44688 0 -1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2126_
timestamp 1698431365
transform 1 0 41664 0 -1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2127_
timestamp 1698431365
transform 1 0 45136 0 1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2128_
timestamp 1698431365
transform 1 0 44800 0 -1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2129_
timestamp 1698431365
transform 1 0 27776 0 -1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2130_
timestamp 1698431365
transform 1 0 29008 0 1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2131_
timestamp 1698431365
transform 1 0 29232 0 1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2132_
timestamp 1698431365
transform 1 0 29120 0 1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2133_
timestamp 1698431365
transform 1 0 37184 0 -1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2134_
timestamp 1698431365
transform 1 0 39088 0 1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2135_
timestamp 1698431365
transform -1 0 45920 0 -1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2136_
timestamp 1698431365
transform 1 0 40768 0 -1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2137_
timestamp 1698431365
transform 1 0 29008 0 1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2138_
timestamp 1698431365
transform 1 0 32256 0 1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2139_
timestamp 1698431365
transform 1 0 13552 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2140_
timestamp 1698431365
transform 1 0 16688 0 1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2141_
timestamp 1698431365
transform 1 0 13440 0 1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2142_
timestamp 1698431365
transform -1 0 14784 0 -1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2143_
timestamp 1698431365
transform -1 0 28784 0 1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2144_
timestamp 1698431365
transform 1 0 17696 0 1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2145_
timestamp 1698431365
transform 1 0 18592 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2146_
timestamp 1698431365
transform 1 0 17024 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2147_
timestamp 1698431365
transform 1 0 20832 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2148_
timestamp 1698431365
transform -1 0 28784 0 1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2149_
timestamp 1698431365
transform 1 0 25536 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2150_
timestamp 1698431365
transform 1 0 22288 0 1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2151_
timestamp 1698431365
transform 1 0 23072 0 1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2152_
timestamp 1698431365
transform 1 0 14672 0 1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2153_
timestamp 1698431365
transform 1 0 13776 0 1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2154_
timestamp 1698431365
transform 1 0 17696 0 1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2155_
timestamp 1698431365
transform 1 0 25648 0 -1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2156_
timestamp 1698431365
transform -1 0 28784 0 1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2157_
timestamp 1698431365
transform 1 0 35728 0 -1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2158_
timestamp 1698431365
transform 1 0 40768 0 -1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2159_
timestamp 1698431365
transform 1 0 45136 0 1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2160_
timestamp 1698431365
transform 1 0 45136 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2161_
timestamp 1698431365
transform 1 0 28224 0 -1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2162_
timestamp 1698431365
transform -1 0 36176 0 -1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2163_
timestamp 1698431365
transform 1 0 11984 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2164_
timestamp 1698431365
transform 1 0 1568 0 1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2165_
timestamp 1698431365
transform 1 0 4592 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _2166_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 36288 0 -1 7840
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _2167_
timestamp 1698431365
transform 1 0 19376 0 -1 9408
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _2168_
timestamp 1698431365
transform 1 0 24640 0 1 6272
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffnq_1  _2169_
timestamp 1698431365
transform 1 0 28112 0 -1 7840
box -86 -86 3446 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2170_
timestamp 1698431365
transform 1 0 22624 0 1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2171_
timestamp 1698431365
transform 1 0 16016 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2172_
timestamp 1698431365
transform 1 0 6272 0 1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _2173_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 7280 0 -1 4704
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2174_
timestamp 1698431365
transform 1 0 7280 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2175_
timestamp 1698431365
transform 1 0 12768 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2176_
timestamp 1698431365
transform 1 0 9744 0 -1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2177_
timestamp 1698431365
transform 1 0 13552 0 -1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2178_
timestamp 1698431365
transform 1 0 39200 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2179_
timestamp 1698431365
transform 1 0 41216 0 -1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2180_
timestamp 1698431365
transform 1 0 45136 0 1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2181_
timestamp 1698431365
transform 1 0 44240 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2182_
timestamp 1698431365
transform 1 0 35616 0 -1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2183_
timestamp 1698431365
transform -1 0 39760 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2184_
timestamp 1698431365
transform 1 0 31696 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2185_
timestamp 1698431365
transform 1 0 18480 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2186_
timestamp 1698431365
transform 1 0 23296 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2187_
timestamp 1698431365
transform 1 0 26544 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2188_
timestamp 1698431365
transform 1 0 1568 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2189_
timestamp 1698431365
transform 1 0 12320 0 -1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2190_
timestamp 1698431365
transform 1 0 1568 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2191_
timestamp 1698431365
transform -1 0 14784 0 -1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2192_
timestamp 1698431365
transform 1 0 1568 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2193_
timestamp 1698431365
transform -1 0 4816 0 1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2194_
timestamp 1698431365
transform 1 0 6944 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2195_
timestamp 1698431365
transform -1 0 4816 0 1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2196_
timestamp 1698431365
transform 1 0 1568 0 1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2197_
timestamp 1698431365
transform 1 0 5936 0 -1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2198_
timestamp 1698431365
transform -1 0 4816 0 1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2199_
timestamp 1698431365
transform 1 0 1568 0 1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2200_
timestamp 1698431365
transform 1 0 5600 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2201_
timestamp 1698431365
transform 1 0 16800 0 1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2202_
timestamp 1698431365
transform 1 0 36176 0 -1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2203_
timestamp 1698431365
transform -1 0 43792 0 1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2204_
timestamp 1698431365
transform 1 0 32928 0 -1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2205_
timestamp 1698431365
transform 1 0 34384 0 -1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2206_
timestamp 1698431365
transform 1 0 38192 0 1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2207_
timestamp 1698431365
transform -1 0 46368 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2208_
timestamp 1698431365
transform 1 0 42672 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2209_
timestamp 1698431365
transform -1 0 45024 0 -1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2210_
timestamp 1698431365
transform -1 0 39424 0 -1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2211_
timestamp 1698431365
transform 1 0 37296 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2212_
timestamp 1698431365
transform 1 0 17248 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _2213_
timestamp 1698431365
transform 1 0 14672 0 1 21952
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2214_
timestamp 1698431365
transform 1 0 20272 0 -1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2215_
timestamp 1698431365
transform 1 0 30576 0 1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2216_
timestamp 1698431365
transform 1 0 31584 0 1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2217_
timestamp 1698431365
transform 1 0 23184 0 1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2218_
timestamp 1698431365
transform 1 0 25088 0 -1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _2219_
timestamp 1698431365
transform 1 0 21168 0 1 12544
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2220_
timestamp 1698431365
transform 1 0 22288 0 1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2221_
timestamp 1698431365
transform 1 0 45136 0 1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2222_
timestamp 1698431365
transform 1 0 45136 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2223_
timestamp 1698431365
transform 1 0 1568 0 1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2224_
timestamp 1698431365
transform 1 0 3136 0 -1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2225_
timestamp 1698431365
transform 1 0 5936 0 -1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2226_
timestamp 1698431365
transform 1 0 44688 0 1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2227_
timestamp 1698431365
transform 1 0 41216 0 1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2228_
timestamp 1698431365
transform 1 0 32928 0 -1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2229_
timestamp 1698431365
transform 1 0 30688 0 1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2230_
timestamp 1698431365
transform 1 0 19040 0 -1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2231_
timestamp 1698431365
transform 1 0 17920 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2232_
timestamp 1698431365
transform 1 0 25088 0 -1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2233_
timestamp 1698431365
transform 1 0 24864 0 1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2234_
timestamp 1698431365
transform 1 0 25088 0 -1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2235_
timestamp 1698431365
transform 1 0 23856 0 1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2236_
timestamp 1698431365
transform 1 0 17584 0 1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2237_
timestamp 1698431365
transform -1 0 24080 0 -1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2238_
timestamp 1698431365
transform 1 0 17360 0 -1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2239_
timestamp 1698431365
transform -1 0 18816 0 1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2240_
timestamp 1698431365
transform 1 0 12208 0 -1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2241_
timestamp 1698431365
transform -1 0 13552 0 -1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2242_
timestamp 1698431365
transform 1 0 8624 0 1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _2243_
timestamp 1698431365
transform 1 0 5488 0 1 42336
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2244_
timestamp 1698431365
transform 1 0 2016 0 1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2245_
timestamp 1698431365
transform 1 0 1568 0 -1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _2246_
timestamp 1698431365
transform 1 0 1568 0 -1 39200
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2247_
timestamp 1698431365
transform 1 0 1568 0 1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2248_
timestamp 1698431365
transform 1 0 1568 0 1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2249_
timestamp 1698431365
transform -1 0 17360 0 1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2250_
timestamp 1698431365
transform 1 0 1568 0 1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _2251_
timestamp 1698431365
transform 1 0 13552 0 -1 45472
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2252_
timestamp 1698431365
transform 1 0 1568 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2253_
timestamp 1698431365
transform 1 0 5936 0 -1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _2254_
timestamp 1698431365
transform 1 0 45136 0 -1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2271_
timestamp 1698431365
transform 1 0 36848 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2272_
timestamp 1698431365
transform 1 0 35504 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2273_
timestamp 1698431365
transform 1 0 37968 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2274_
timestamp 1698431365
transform 1 0 43232 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2275_
timestamp 1698431365
transform 1 0 38528 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2276_
timestamp 1698431365
transform 1 0 39200 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1032__A2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 20272 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1035__A2
timestamp 1698431365
transform -1 0 5936 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1046__B2
timestamp 1698431365
transform 1 0 7728 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1047__A1
timestamp 1698431365
transform 1 0 8848 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1047__A2
timestamp 1698431365
transform -1 0 9968 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1049__A2
timestamp 1698431365
transform 1 0 23744 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1051__A2
timestamp 1698431365
transform 1 0 19040 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1054__I
timestamp 1698431365
transform 1 0 7280 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1057__I
timestamp 1698431365
transform -1 0 7056 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1064__A2
timestamp 1698431365
transform 1 0 8960 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1066__I
timestamp 1698431365
transform 1 0 16800 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1073__A1
timestamp 1698431365
transform 1 0 9632 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1073__A2
timestamp 1698431365
transform 1 0 8624 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1077__A2
timestamp 1698431365
transform 1 0 19376 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1078__A2
timestamp 1698431365
transform 1 0 21840 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1083__I
timestamp 1698431365
transform 1 0 8512 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1085__A1
timestamp 1698431365
transform 1 0 10304 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1086__I
timestamp 1698431365
transform 1 0 15792 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1089__A2
timestamp 1698431365
transform -1 0 11200 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1093__B2
timestamp 1698431365
transform -1 0 5712 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1096__I
timestamp 1698431365
transform 1 0 17136 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1102__I
timestamp 1698431365
transform 1 0 11088 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1103__A2
timestamp 1698431365
transform -1 0 18144 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1107__A2
timestamp 1698431365
transform 1 0 11312 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1107__B2
timestamp 1698431365
transform -1 0 13104 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1111__A2
timestamp 1698431365
transform 1 0 24080 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1112__B2
timestamp 1698431365
transform 1 0 7280 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1115__B2
timestamp 1698431365
transform 1 0 6608 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1125__A2
timestamp 1698431365
transform 1 0 12320 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1125__B
timestamp 1698431365
transform -1 0 15344 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1132__I
timestamp 1698431365
transform -1 0 5712 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1134__A1
timestamp 1698431365
transform -1 0 9856 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1145__A2
timestamp 1698431365
transform 1 0 8400 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1151__B
timestamp 1698431365
transform -1 0 2016 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1152__A1
timestamp 1698431365
transform 1 0 2800 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1155__I
timestamp 1698431365
transform 1 0 7392 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1159__B
timestamp 1698431365
transform 1 0 5040 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1162__A2
timestamp 1698431365
transform 1 0 9632 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1175__B
timestamp 1698431365
transform 1 0 13664 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1176__A1
timestamp 1698431365
transform 1 0 16016 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1179__A1
timestamp 1698431365
transform -1 0 15568 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1184__A2
timestamp 1698431365
transform -1 0 9184 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1187__A1
timestamp 1698431365
transform -1 0 12208 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1189__A2
timestamp 1698431365
transform -1 0 7168 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1193__B2
timestamp 1698431365
transform 1 0 8848 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1207__A1
timestamp 1698431365
transform -1 0 5936 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1208__B
timestamp 1698431365
transform -1 0 5488 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1212__A2
timestamp 1698431365
transform 1 0 10416 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1222__A3
timestamp 1698431365
transform 1 0 20048 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1226__A2
timestamp 1698431365
transform 1 0 17920 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1227__A2
timestamp 1698431365
transform -1 0 9520 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1229__I
timestamp 1698431365
transform 1 0 19712 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1236__A1
timestamp 1698431365
transform 1 0 23632 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1237__A1
timestamp 1698431365
transform -1 0 18368 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1239__A4
timestamp 1698431365
transform -1 0 10976 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1267__A2
timestamp 1698431365
transform 1 0 19152 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1268__A1
timestamp 1698431365
transform 1 0 19600 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1268__A2
timestamp 1698431365
transform 1 0 20608 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1270__C
timestamp 1698431365
transform 1 0 6608 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1275__A1
timestamp 1698431365
transform 1 0 23408 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1275__A2
timestamp 1698431365
transform 1 0 22960 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1277__C
timestamp 1698431365
transform -1 0 5264 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1287__A2
timestamp 1698431365
transform -1 0 9520 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1288__A2
timestamp 1698431365
transform 1 0 11984 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1295__A3
timestamp 1698431365
transform 1 0 41888 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1295__A4
timestamp 1698431365
transform -1 0 37968 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1296__I
timestamp 1698431365
transform 1 0 37520 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1298__I
timestamp 1698431365
transform -1 0 24304 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1300__B
timestamp 1698431365
transform 1 0 7392 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1306__I
timestamp 1698431365
transform 1 0 20720 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1308__A1
timestamp 1698431365
transform 1 0 12096 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1309__A2
timestamp 1698431365
transform 1 0 13104 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1315__I
timestamp 1698431365
transform 1 0 8512 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1318__A1
timestamp 1698431365
transform 1 0 12208 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1319__A4
timestamp 1698431365
transform -1 0 5264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1325__A3
timestamp 1698431365
transform -1 0 2240 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1327__I
timestamp 1698431365
transform 1 0 18256 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1328__A1
timestamp 1698431365
transform -1 0 9184 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1332__A1
timestamp 1698431365
transform -1 0 6832 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1337__A3
timestamp 1698431365
transform -1 0 5936 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1353__A1
timestamp 1698431365
transform 1 0 32480 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1383__I
timestamp 1698431365
transform 1 0 17472 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1384__A1
timestamp 1698431365
transform 1 0 35728 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1389__A1
timestamp 1698431365
transform 1 0 32144 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1402__A1
timestamp 1698431365
transform 1 0 25984 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1403__A1
timestamp 1698431365
transform 1 0 27104 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1409__A1
timestamp 1698431365
transform 1 0 29456 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1410__A1
timestamp 1698431365
transform 1 0 29456 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1420__S
timestamp 1698431365
transform -1 0 29456 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1423__I
timestamp 1698431365
transform 1 0 36176 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1424__S
timestamp 1698431365
transform 1 0 31808 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1428__S
timestamp 1698431365
transform 1 0 39648 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1432__S
timestamp 1698431365
transform 1 0 36288 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1436__I0
timestamp 1698431365
transform 1 0 44912 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1465__A1
timestamp 1698431365
transform 1 0 42672 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1466__A1
timestamp 1698431365
transform 1 0 38640 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1481__I0
timestamp 1698431365
transform -1 0 45136 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1491__B
timestamp 1698431365
transform -1 0 26208 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1492__A2
timestamp 1698431365
transform 1 0 25312 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1497__I
timestamp 1698431365
transform 1 0 27888 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1500__A2
timestamp 1698431365
transform 1 0 31248 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1502__A2
timestamp 1698431365
transform 1 0 28784 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1506__A2
timestamp 1698431365
transform 1 0 30800 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1508__A2
timestamp 1698431365
transform 1 0 28896 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1511__I
timestamp 1698431365
transform 1 0 24752 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1513__A1
timestamp 1698431365
transform -1 0 29792 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1517__B
timestamp 1698431365
transform 1 0 28560 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1524__B
timestamp 1698431365
transform -1 0 30912 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1555__A1
timestamp 1698431365
transform 1 0 42336 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1556__I
timestamp 1698431365
transform 1 0 42672 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1563__A2
timestamp 1698431365
transform 1 0 22400 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1565__I
timestamp 1698431365
transform 1 0 5488 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1566__S
timestamp 1698431365
transform 1 0 21056 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1568__S
timestamp 1698431365
transform 1 0 24864 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1572__S
timestamp 1698431365
transform 1 0 39872 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1574__S
timestamp 1698431365
transform 1 0 42224 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1576__S
timestamp 1698431365
transform -1 0 45136 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1578__S
timestamp 1698431365
transform 1 0 44912 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1611__I
timestamp 1698431365
transform -1 0 40992 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1612__S
timestamp 1698431365
transform 1 0 41664 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1614__S
timestamp 1698431365
transform 1 0 39984 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1616__S
timestamp 1698431365
transform 1 0 41216 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1618__S
timestamp 1698431365
transform 1 0 40320 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1620__I
timestamp 1698431365
transform 1 0 33376 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1629__I
timestamp 1698431365
transform 1 0 45136 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1634__I0
timestamp 1698431365
transform -1 0 42784 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1644__A1
timestamp 1698431365
transform 1 0 13552 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1646__I
timestamp 1698431365
transform 1 0 9968 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1647__I
timestamp 1698431365
transform -1 0 17024 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1654__A2
timestamp 1698431365
transform -1 0 10080 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1657__A2
timestamp 1698431365
transform 1 0 17920 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1659__A2
timestamp 1698431365
transform 1 0 15120 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1659__C
timestamp 1698431365
transform -1 0 16352 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1661__A2
timestamp 1698431365
transform 1 0 12208 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1662__A2
timestamp 1698431365
transform 1 0 11424 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1662__C
timestamp 1698431365
transform -1 0 13104 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1663__A1
timestamp 1698431365
transform 1 0 28672 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1664__I
timestamp 1698431365
transform 1 0 28560 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1666__I
timestamp 1698431365
transform 1 0 30128 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1668__A2
timestamp 1698431365
transform -1 0 13104 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1671__A1
timestamp 1698431365
transform 1 0 21392 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1678__A1
timestamp 1698431365
transform -1 0 11984 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1678__B2
timestamp 1698431365
transform -1 0 12432 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1680__C
timestamp 1698431365
transform 1 0 14896 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1685__A1
timestamp 1698431365
transform 1 0 10192 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1685__A2
timestamp 1698431365
transform 1 0 11760 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1686__A1
timestamp 1698431365
transform -1 0 10192 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1686__C2
timestamp 1698431365
transform 1 0 12768 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1690__A2
timestamp 1698431365
transform -1 0 15904 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1691__A1
timestamp 1698431365
transform -1 0 16128 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1695__A2
timestamp 1698431365
transform -1 0 13552 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1696__C2
timestamp 1698431365
transform -1 0 13104 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1697__A1
timestamp 1698431365
transform -1 0 15904 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1702__B2
timestamp 1698431365
transform -1 0 14000 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1703__A1
timestamp 1698431365
transform 1 0 15904 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1703__B2
timestamp 1698431365
transform -1 0 17360 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1709__A1
timestamp 1698431365
transform -1 0 16240 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1710__I
timestamp 1698431365
transform 1 0 14000 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1711__A2
timestamp 1698431365
transform -1 0 16576 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1718__A1
timestamp 1698431365
transform -1 0 13104 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1719__A1
timestamp 1698431365
transform -1 0 19152 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1724__A1
timestamp 1698431365
transform 1 0 14896 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1724__B2
timestamp 1698431365
transform -1 0 9968 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1724__C2
timestamp 1698431365
transform -1 0 10416 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1728__A1
timestamp 1698431365
transform -1 0 17696 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1729__A1
timestamp 1698431365
transform -1 0 6608 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1729__B2
timestamp 1698431365
transform -1 0 5712 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1739__A1
timestamp 1698431365
transform 1 0 20048 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1743__S
timestamp 1698431365
transform 1 0 30016 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1745__S
timestamp 1698431365
transform 1 0 29904 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1747__S
timestamp 1698431365
transform 1 0 37184 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1749__S
timestamp 1698431365
transform 1 0 40656 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1752__I0
timestamp 1698431365
transform 1 0 48160 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1752__S
timestamp 1698431365
transform -1 0 44464 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1754__S
timestamp 1698431365
transform 1 0 46032 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1756__S
timestamp 1698431365
transform 1 0 30240 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1758__S
timestamp 1698431365
transform 1 0 34048 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1760__I
timestamp 1698431365
transform 1 0 11312 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1765__I
timestamp 1698431365
transform -1 0 6160 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1768__B
timestamp 1698431365
transform -1 0 8848 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1770__A2
timestamp 1698431365
transform -1 0 7056 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1770__A3
timestamp 1698431365
transform -1 0 10192 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1773__A2
timestamp 1698431365
transform -1 0 7168 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1775__I
timestamp 1698431365
transform 1 0 28560 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1783__A2
timestamp 1698431365
transform 1 0 18368 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1785__I
timestamp 1698431365
transform -1 0 14448 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1788__A2
timestamp 1698431365
transform -1 0 6384 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1792__A2
timestamp 1698431365
transform 1 0 5040 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1804__I
timestamp 1698431365
transform 1 0 18368 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1807__B
timestamp 1698431365
transform -1 0 9184 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1809__I
timestamp 1698431365
transform 1 0 14672 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1815__A1
timestamp 1698431365
transform 1 0 30352 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1816__B
timestamp 1698431365
transform 1 0 27888 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1819__A1
timestamp 1698431365
transform 1 0 30800 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1820__B
timestamp 1698431365
transform 1 0 29904 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1823__A1
timestamp 1698431365
transform -1 0 32704 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1824__B
timestamp 1698431365
transform -1 0 34384 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1826__I
timestamp 1698431365
transform 1 0 31696 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1859__A2
timestamp 1698431365
transform -1 0 22064 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1861__A1
timestamp 1698431365
transform -1 0 37520 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1861__A2
timestamp 1698431365
transform 1 0 42784 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1865__C
timestamp 1698431365
transform 1 0 33824 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1870__I0
timestamp 1698431365
transform 1 0 36400 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1875__A1
timestamp 1698431365
transform 1 0 37520 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1881__A1
timestamp 1698431365
transform 1 0 43344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1881__B2
timestamp 1698431365
transform 1 0 42896 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1886__A1
timestamp 1698431365
transform 1 0 37072 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1891__A1
timestamp 1698431365
transform 1 0 37968 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1891__A2
timestamp 1698431365
transform 1 0 40992 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1895__A1
timestamp 1698431365
transform 1 0 40208 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1898__A2
timestamp 1698431365
transform -1 0 38528 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1899__A1
timestamp 1698431365
transform 1 0 39648 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1902__A2
timestamp 1698431365
transform 1 0 22512 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1906__A1
timestamp 1698431365
transform -1 0 28784 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1909__A1
timestamp 1698431365
transform 1 0 28896 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1910__A1
timestamp 1698431365
transform 1 0 26096 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1924__A1
timestamp 1698431365
transform -1 0 28112 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1928__B
timestamp 1698431365
transform 1 0 44912 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1932__A2
timestamp 1698431365
transform 1 0 29792 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1933__B
timestamp 1698431365
transform 1 0 46928 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1941__A1
timestamp 1698431365
transform 1 0 48048 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1951__A1
timestamp 1698431365
transform -1 0 7616 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1954__B
timestamp 1698431365
transform 1 0 34608 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1955__A2
timestamp 1698431365
transform 1 0 34272 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1957__A3
timestamp 1698431365
transform 1 0 28112 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1964__A1
timestamp 1698431365
transform 1 0 19600 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1964__A2
timestamp 1698431365
transform -1 0 19824 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1965__I1
timestamp 1698431365
transform 1 0 17584 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1967__I1
timestamp 1698431365
transform 1 0 19040 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1974__I
timestamp 1698431365
transform 1 0 21392 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1978__A1
timestamp 1698431365
transform 1 0 21392 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1978__A2
timestamp 1698431365
transform -1 0 21056 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1978__B
timestamp 1698431365
transform 1 0 24528 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1983__A1
timestamp 1698431365
transform 1 0 18928 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1989__B
timestamp 1698431365
transform 1 0 24528 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1990__A1
timestamp 1698431365
transform 1 0 23744 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1990__A2
timestamp 1698431365
transform 1 0 25312 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1992__A1
timestamp 1698431365
transform 1 0 24864 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1994__A1
timestamp 1698431365
transform 1 0 24080 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1995__A1
timestamp 1698431365
transform 1 0 22288 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1995__A2
timestamp 1698431365
transform 1 0 24080 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1995__B
timestamp 1698431365
transform -1 0 24752 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2000__A1
timestamp 1698431365
transform 1 0 18368 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2001__A1
timestamp 1698431365
transform 1 0 19376 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2004__A1
timestamp 1698431365
transform 1 0 19712 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2005__B
timestamp 1698431365
transform 1 0 21392 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2006__A1
timestamp 1698431365
transform 1 0 25312 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2006__A2
timestamp 1698431365
transform 1 0 18592 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2006__B
timestamp 1698431365
transform 1 0 25312 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2010__A1
timestamp 1698431365
transform -1 0 18144 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2013__I
timestamp 1698431365
transform 1 0 16800 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2014__A1
timestamp 1698431365
transform -1 0 18032 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2015__A1
timestamp 1698431365
transform -1 0 17136 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2015__A2
timestamp 1698431365
transform -1 0 15568 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2019__A1
timestamp 1698431365
transform -1 0 17696 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2020__A1
timestamp 1698431365
transform 1 0 10864 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2022__A1
timestamp 1698431365
transform -1 0 14672 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2023__A1
timestamp 1698431365
transform 1 0 9968 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2024__A1
timestamp 1698431365
transform -1 0 13776 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2024__A2
timestamp 1698431365
transform -1 0 12656 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2026__A1
timestamp 1698431365
transform 1 0 8960 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2029__A1
timestamp 1698431365
transform -1 0 11760 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2030__I
timestamp 1698431365
transform -1 0 6496 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2031__I
timestamp 1698431365
transform -1 0 4592 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2032__A1
timestamp 1698431365
transform -1 0 8624 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2035__I
timestamp 1698431365
transform -1 0 3584 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2037__A1
timestamp 1698431365
transform -1 0 3136 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2038__A1
timestamp 1698431365
transform -1 0 9856 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2041__A1
timestamp 1698431365
transform -1 0 5936 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2042__A1
timestamp 1698431365
transform -1 0 6944 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2042__A2
timestamp 1698431365
transform 1 0 4816 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2045__A1
timestamp 1698431365
transform 1 0 6832 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2046__A1
timestamp 1698431365
transform -1 0 6048 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2046__A2
timestamp 1698431365
transform -1 0 3920 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2049__A1
timestamp 1698431365
transform -1 0 3584 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2050__A1
timestamp 1698431365
transform -1 0 4368 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2050__A2
timestamp 1698431365
transform -1 0 3248 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2054__A1
timestamp 1698431365
transform 1 0 10192 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2055__A1
timestamp 1698431365
transform -1 0 12656 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2057__A1
timestamp 1698431365
transform -1 0 3920 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2057__A2
timestamp 1698431365
transform -1 0 2240 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2058__B
timestamp 1698431365
transform 1 0 8064 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2059__A1
timestamp 1698431365
transform -1 0 17696 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2060__A1
timestamp 1698431365
transform -1 0 15120 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2061__A1
timestamp 1698431365
transform -1 0 15792 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2062__B
timestamp 1698431365
transform -1 0 6160 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2063__A1
timestamp 1698431365
transform -1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2064__A2
timestamp 1698431365
transform 1 0 4144 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2065__A2
timestamp 1698431365
transform 1 0 17472 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2066__B
timestamp 1698431365
transform -1 0 10864 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2068__A1
timestamp 1698431365
transform 1 0 14112 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2068__A3
timestamp 1698431365
transform 1 0 15792 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2070__B
timestamp 1698431365
transform -1 0 7840 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2071__A1
timestamp 1698431365
transform 1 0 5040 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2071__A2
timestamp 1698431365
transform 1 0 5824 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2071__B
timestamp 1698431365
transform 1 0 7504 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2072__A2
timestamp 1698431365
transform 1 0 5040 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2074__A1
timestamp 1698431365
transform 1 0 5040 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2075__A1
timestamp 1698431365
transform -1 0 4816 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2075__A2
timestamp 1698431365
transform -1 0 4816 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2077__A1
timestamp 1698431365
transform -1 0 8176 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2080__A1
timestamp 1698431365
transform 1 0 45472 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2081__CLK
timestamp 1698431365
transform 1 0 29904 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2082__CLK
timestamp 1698431365
transform 1 0 29232 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2083__CLK
timestamp 1698431365
transform 1 0 40096 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2084__CLK
timestamp 1698431365
transform 1 0 39872 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2085__CLK
timestamp 1698431365
transform 1 0 40992 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2086__CLK
timestamp 1698431365
transform 1 0 42560 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2087__CLK
timestamp 1698431365
transform -1 0 33376 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2088__CLK
timestamp 1698431365
transform 1 0 40096 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2090__CLK
timestamp 1698431365
transform -1 0 33376 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2091__CLK
timestamp 1698431365
transform 1 0 32480 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2092__CLK
timestamp 1698431365
transform 1 0 43904 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2093__CLK
timestamp 1698431365
transform -1 0 41664 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2094__CLK
timestamp 1698431365
transform 1 0 44576 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2105__CLK
timestamp 1698431365
transform 1 0 43008 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2106__CLK
timestamp 1698431365
transform 1 0 38304 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2107__CLK
timestamp 1698431365
transform -1 0 19488 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2108__CLK
timestamp 1698431365
transform 1 0 26544 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2115__CLK
timestamp 1698431365
transform 1 0 26432 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2116__CLK
timestamp 1698431365
transform 1 0 27216 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2117__CLK
timestamp 1698431365
transform 1 0 40992 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2118__CLK
timestamp 1698431365
transform 1 0 39424 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2119__CLK
timestamp 1698431365
transform 1 0 42112 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2120__CLK
timestamp 1698431365
transform 1 0 42448 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2121__CLK
timestamp 1698431365
transform 1 0 31584 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2122__CLK
timestamp 1698431365
transform 1 0 38864 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2123__CLK
timestamp 1698431365
transform 1 0 37072 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2124__CLK
timestamp 1698431365
transform -1 0 41216 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2125__CLK
timestamp 1698431365
transform 1 0 41664 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2126__CLK
timestamp 1698431365
transform 1 0 36400 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2127__CLK
timestamp 1698431365
transform 1 0 37072 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2128__CLK
timestamp 1698431365
transform -1 0 45136 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2131__CLK
timestamp 1698431365
transform 1 0 32704 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2132__CLK
timestamp 1698431365
transform 1 0 32592 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2139__CLK
timestamp 1698431365
transform 1 0 18144 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2140__CLK
timestamp 1698431365
transform 1 0 20160 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2141__CLK
timestamp 1698431365
transform 1 0 17472 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2142__CLK
timestamp 1698431365
transform 1 0 15456 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2143__CLK
timestamp 1698431365
transform 1 0 29120 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2152__CLK
timestamp 1698431365
transform 1 0 14448 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2153__CLK
timestamp 1698431365
transform 1 0 17472 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2154__CLK
timestamp 1698431365
transform 1 0 21392 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2155__CLK
timestamp 1698431365
transform 1 0 29120 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2156__CLK
timestamp 1698431365
transform 1 0 28784 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2163__CLK
timestamp 1698431365
transform 1 0 15456 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2164__CLK
timestamp 1698431365
transform -1 0 5936 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2165__CLK
timestamp 1698431365
transform 1 0 5040 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2166__CLKN
timestamp 1698431365
transform 1 0 37184 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2167__CLKN
timestamp 1698431365
transform 1 0 22960 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2168__CLKN
timestamp 1698431365
transform 1 0 24416 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2169__CLKN
timestamp 1698431365
transform 1 0 32144 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2170__CLK
timestamp 1698431365
transform 1 0 22400 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2171__CLK
timestamp 1698431365
transform 1 0 10640 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2172__CLK
timestamp 1698431365
transform 1 0 8848 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2173__CLK
timestamp 1698431365
transform -1 0 5936 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2174__CLK
timestamp 1698431365
transform 1 0 6608 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2175__CLK
timestamp 1698431365
transform 1 0 18816 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2176__CLK
timestamp 1698431365
transform 1 0 9744 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2177__CLK
timestamp 1698431365
transform 1 0 17920 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2178__CLK
timestamp 1698431365
transform 1 0 33712 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2179__CLK
timestamp 1698431365
transform 1 0 31248 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2180__CLK
timestamp 1698431365
transform -1 0 28784 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2181__CLK
timestamp 1698431365
transform 1 0 33264 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2182__CLK
timestamp 1698431365
transform 1 0 33936 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2183__CLK
timestamp 1698431365
transform 1 0 32480 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2184__CLK
timestamp 1698431365
transform 1 0 34384 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2185__CLK
timestamp 1698431365
transform 1 0 21392 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2186__CLK
timestamp 1698431365
transform 1 0 20720 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2187__CLK
timestamp 1698431365
transform 1 0 27216 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2188__CLK
timestamp 1698431365
transform 1 0 5040 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2189__CLK
timestamp 1698431365
transform 1 0 15792 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2190__CLK
timestamp 1698431365
transform -1 0 6384 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2191__CLK
timestamp 1698431365
transform 1 0 15008 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2192__CLK
timestamp 1698431365
transform 1 0 5040 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2193__CLK
timestamp 1698431365
transform 1 0 5040 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2194__CLK
timestamp 1698431365
transform 1 0 10192 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2195__CLK
timestamp 1698431365
transform 1 0 6160 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2196__CLK
timestamp 1698431365
transform 1 0 6608 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2197__CLK
timestamp 1698431365
transform 1 0 9632 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2198__CLK
timestamp 1698431365
transform 1 0 6160 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2199__CLK
timestamp 1698431365
transform 1 0 6384 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2200__CLK
timestamp 1698431365
transform 1 0 9632 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2201__CLK
timestamp 1698431365
transform 1 0 20720 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2202__CLK
timestamp 1698431365
transform 1 0 39424 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2203__CLK
timestamp 1698431365
transform 1 0 40320 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2213__CLK
timestamp 1698431365
transform 1 0 14448 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2215__CLK
timestamp 1698431365
transform 1 0 34048 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2216__CLK
timestamp 1698431365
transform 1 0 35056 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2217__CLK
timestamp 1698431365
transform 1 0 22960 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2218__CLK
timestamp 1698431365
transform 1 0 24640 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2220__CLK
timestamp 1698431365
transform 1 0 22064 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2222__CLK
timestamp 1698431365
transform 1 0 44912 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2223__CLK
timestamp 1698431365
transform 1 0 5712 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2224__CLK
timestamp 1698431365
transform 1 0 7056 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2225__CLK
timestamp 1698431365
transform 1 0 9184 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2226__CLK
timestamp 1698431365
transform 1 0 35056 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2227__CLK
timestamp 1698431365
transform 1 0 38192 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2228__CLK
timestamp 1698431365
transform 1 0 36176 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2229__CLK
timestamp 1698431365
transform 1 0 34160 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2230__CLK
timestamp 1698431365
transform 1 0 22288 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2235__CLK
timestamp 1698431365
transform 1 0 28000 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2236__CLK
timestamp 1698431365
transform 1 0 20608 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2237__CLK
timestamp 1698431365
transform 1 0 24080 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2238__CLK
timestamp 1698431365
transform -1 0 21056 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2239__CLK
timestamp 1698431365
transform 1 0 17920 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2240__CLK
timestamp 1698431365
transform 1 0 17360 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2241__CLK
timestamp 1698431365
transform -1 0 13552 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2242__CLK
timestamp 1698431365
transform 1 0 10080 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2243__CLK
timestamp 1698431365
transform 1 0 7952 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2244__CLK
timestamp 1698431365
transform 1 0 3920 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2245__CLK
timestamp 1698431365
transform 1 0 4816 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2246__CLK
timestamp 1698431365
transform 1 0 1792 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2247__CLK
timestamp 1698431365
transform 1 0 3920 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2248__CLK
timestamp 1698431365
transform 1 0 5040 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2250__CLK
timestamp 1698431365
transform 1 0 3920 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2251__CLK
timestamp 1698431365
transform -1 0 17248 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2252__CLK
timestamp 1698431365
transform 1 0 4592 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2253__CLK
timestamp 1698431365
transform -1 0 9632 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_clk_I
timestamp 1698431365
transform 1 0 24640 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_0_0_clk_I
timestamp 1698431365
transform 1 0 17472 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_1_0_clk_I
timestamp 1698431365
transform 1 0 16464 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_2_0_clk_I
timestamp 1698431365
transform 1 0 25312 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_3_0_clk_I
timestamp 1698431365
transform 1 0 24192 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_4_0_clk_I
timestamp 1698431365
transform -1 0 11312 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_5_0_clk_I
timestamp 1698431365
transform 1 0 15008 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_6_0_clk_I
timestamp 1698431365
transform 1 0 23408 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_7_0_clk_I
timestamp 1698431365
transform 1 0 21280 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_8_0_clk_I
timestamp 1698431365
transform 1 0 33152 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_9_0_clk_I
timestamp 1698431365
transform 1 0 32704 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_10_0_clk_I
timestamp 1698431365
transform 1 0 36400 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_11_0_clk_I
timestamp 1698431365
transform 1 0 37184 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_12_0_clk_I
timestamp 1698431365
transform 1 0 28560 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_13_0_clk_I
timestamp 1698431365
transform 1 0 29232 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_14_0_clk_I
timestamp 1698431365
transform 1 0 37184 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_15_0_clk_I
timestamp 1698431365
transform 1 0 37072 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input1_I
timestamp 1698431365
transform 1 0 2912 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input2_I
timestamp 1698431365
transform -1 0 10752 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input3_I
timestamp 1698431365
transform 1 0 2240 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input4_I
timestamp 1698431365
transform 1 0 2912 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input5_I
timestamp 1698431365
transform 1 0 4816 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input6_I
timestamp 1698431365
transform 1 0 2464 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input7_I
timestamp 1698431365
transform 1 0 1792 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input8_I
timestamp 1698431365
transform 1 0 4368 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input9_I
timestamp 1698431365
transform 1 0 4816 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input10_I
timestamp 1698431365
transform 1 0 2464 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input11_I
timestamp 1698431365
transform 1 0 2464 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input12_I
timestamp 1698431365
transform 1 0 2912 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input13_I
timestamp 1698431365
transform 1 0 5040 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input14_I
timestamp 1698431365
transform 1 0 4368 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input15_I
timestamp 1698431365
transform 1 0 1904 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input16_I
timestamp 1698431365
transform 1 0 1792 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input17_I
timestamp 1698431365
transform -1 0 2688 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input18_I
timestamp 1698431365
transform 1 0 2800 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input19_I
timestamp 1698431365
transform -1 0 2240 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input20_I
timestamp 1698431365
transform 1 0 25312 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input21_I
timestamp 1698431365
transform -1 0 17808 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input22_I
timestamp 1698431365
transform -1 0 18256 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input23_I
timestamp 1698431365
transform 1 0 3360 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input24_I
timestamp 1698431365
transform 1 0 16240 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input25_I
timestamp 1698431365
transform -1 0 35056 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input26_I
timestamp 1698431365
transform -1 0 41216 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input27_I
timestamp 1698431365
transform -1 0 35952 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input28_I
timestamp 1698431365
transform -1 0 5152 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input29_I
timestamp 1698431365
transform -1 0 11536 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input30_I
timestamp 1698431365
transform -1 0 8736 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input31_I
timestamp 1698431365
transform -1 0 12096 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input32_I
timestamp 1698431365
transform 1 0 24416 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input33_I
timestamp 1698431365
transform -1 0 5936 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input34_I
timestamp 1698431365
transform -1 0 4256 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input35_I
timestamp 1698431365
transform 1 0 18368 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input36_I
timestamp 1698431365
transform 1 0 28112 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input37_I
timestamp 1698431365
transform -1 0 23632 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input38_I
timestamp 1698431365
transform 1 0 32592 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input39_I
timestamp 1698431365
transform 1 0 37744 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input40_I
timestamp 1698431365
transform 1 0 35728 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input41_I
timestamp 1698431365
transform -1 0 40096 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input42_I
timestamp 1698431365
transform -1 0 37968 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input43_I
timestamp 1698431365
transform -1 0 28784 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input44_I
timestamp 1698431365
transform -1 0 34944 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input45_I
timestamp 1698431365
transform -1 0 4704 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input46_I
timestamp 1698431365
transform -1 0 20944 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input47_I
timestamp 1698431365
transform -1 0 45136 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input48_I
timestamp 1698431365
transform -1 0 41888 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input49_I
timestamp 1698431365
transform -1 0 44464 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input50_I
timestamp 1698431365
transform -1 0 43568 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input51_I
timestamp 1698431365
transform 1 0 20272 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input52_I
timestamp 1698431365
transform 1 0 3248 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output59_I
timestamp 1698431365
transform 1 0 17472 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output61_I
timestamp 1698431365
transform 1 0 2800 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_clk dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 25088 0 -1 25088
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_0_0_clk dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 16464 0 1 14112
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_1_0_clk
timestamp 1698431365
transform 1 0 13328 0 1 15680
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_2_0_clk
timestamp 1698431365
transform -1 0 22736 0 -1 14112
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_3_0_clk
timestamp 1698431365
transform 1 0 20608 0 -1 15680
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_4_0_clk
timestamp 1698431365
transform 1 0 11760 0 -1 28224
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_5_0_clk
timestamp 1698431365
transform -1 0 16240 0 1 28224
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_6_0_clk
timestamp 1698431365
transform -1 0 22064 0 -1 28224
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_7_0_clk
timestamp 1698431365
transform 1 0 18256 0 -1 31360
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_8_0_clk
timestamp 1698431365
transform -1 0 35840 0 -1 18816
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_9_0_clk
timestamp 1698431365
transform 1 0 32928 0 -1 21952
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_10_0_clk
timestamp 1698431365
transform 1 0 37408 0 1 18816
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_11_0_clk
timestamp 1698431365
transform 1 0 37632 0 -1 20384
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_12_0_clk
timestamp 1698431365
transform 1 0 29008 0 -1 34496
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_13_0_clk
timestamp 1698431365
transform -1 0 32368 0 1 36064
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_14_0_clk
timestamp 1698431365
transform 1 0 37408 0 1 32928
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_15_0_clk
timestamp 1698431365
transform 1 0 37296 0 1 34496
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_10 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 2464 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_18 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 3360 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_22 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 3808 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_26
timestamp 1698431365
transform 1 0 4256 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_30
timestamp 1698431365
transform 1 0 4704 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_36
timestamp 1698431365
transform 1 0 5376 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_38 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5600 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_61
timestamp 1698431365
transform 1 0 8176 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_172
timestamp 1698431365
transform 1 0 20608 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_174
timestamp 1698431365
transform 1 0 20832 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_201
timestamp 1698431365
transform 1 0 23856 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_203
timestamp 1698431365
transform 1 0 24080 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_6 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 2016 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_72
timestamp 1698431365
transform 1 0 9408 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_99
timestamp 1698431365
transform 1 0 12432 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_101
timestamp 1698431365
transform 1 0 12656 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_139
timestamp 1698431365
transform 1 0 16912 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_152
timestamp 1698431365
transform 1 0 18368 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_182
timestamp 1698431365
transform 1 0 21728 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_222
timestamp 1698431365
transform 1 0 26208 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_224
timestamp 1698431365
transform 1 0 26432 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_302
timestamp 1698431365
transform 1 0 35168 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_343
timestamp 1698431365
transform 1 0 39760 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_418
timestamp 1698431365
transform 1 0 48160 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_6
timestamp 1698431365
transform 1 0 2016 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_22
timestamp 1698431365
transform 1 0 3808 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_30
timestamp 1698431365
transform 1 0 4704 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_32
timestamp 1698431365
transform 1 0 4928 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_41
timestamp 1698431365
transform 1 0 5936 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_98
timestamp 1698431365
transform 1 0 12320 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_117
timestamp 1698431365
transform 1 0 14448 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_128
timestamp 1698431365
transform 1 0 15680 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_130
timestamp 1698431365
transform 1 0 15904 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_170
timestamp 1698431365
transform 1 0 20384 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_172
timestamp 1698431365
transform 1 0 20608 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_177
timestamp 1698431365
transform 1 0 21168 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_229
timestamp 1698431365
transform 1 0 26992 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_233
timestamp 1698431365
transform 1 0 27440 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_269
timestamp 1698431365
transform 1 0 31472 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_331
timestamp 1698431365
transform 1 0 38416 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_419
timestamp 1698431365
transform 1 0 48272 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_3_6 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 2016 0 -1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_38
timestamp 1698431365
transform 1 0 5600 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_41
timestamp 1698431365
transform 1 0 5936 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_45
timestamp 1698431365
transform 1 0 6384 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_68
timestamp 1698431365
transform 1 0 8960 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_72
timestamp 1698431365
transform 1 0 9408 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_155
timestamp 1698431365
transform 1 0 18704 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_162
timestamp 1698431365
transform 1 0 19488 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_204
timestamp 1698431365
transform 1 0 24192 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_208
timestamp 1698431365
transform 1 0 24640 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_216
timestamp 1698431365
transform 1 0 25536 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_237
timestamp 1698431365
transform 1 0 27888 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_241
timestamp 1698431365
transform 1 0 28336 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_262
timestamp 1698431365
transform 1 0 30688 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_264
timestamp 1698431365
transform 1 0 30912 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_271
timestamp 1698431365
transform 1 0 31696 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_279
timestamp 1698431365
transform 1 0 32592 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_335
timestamp 1698431365
transform 1 0 38864 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_2
timestamp 1698431365
transform 1 0 1568 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_34
timestamp 1698431365
transform 1 0 5152 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_37
timestamp 1698431365
transform 1 0 5488 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_41
timestamp 1698431365
transform 1 0 5936 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_43
timestamp 1698431365
transform 1 0 6160 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_81
timestamp 1698431365
transform 1 0 10416 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_94
timestamp 1698431365
transform 1 0 11872 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_107
timestamp 1698431365
transform 1 0 13328 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_135
timestamp 1698431365
transform 1 0 16464 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_137
timestamp 1698431365
transform 1 0 16688 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_167
timestamp 1698431365
transform 1 0 20048 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_171
timestamp 1698431365
transform 1 0 20496 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_177
timestamp 1698431365
transform 1 0 21168 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_181
timestamp 1698431365
transform 1 0 21616 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_206
timestamp 1698431365
transform 1 0 24416 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_238
timestamp 1698431365
transform 1 0 28000 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_242
timestamp 1698431365
transform 1 0 28448 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_247
timestamp 1698431365
transform 1 0 29008 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_267
timestamp 1698431365
transform 1 0 31248 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_269
timestamp 1698431365
transform 1 0 31472 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_278
timestamp 1698431365
transform 1 0 32480 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_299
timestamp 1698431365
transform 1 0 34832 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_305
timestamp 1698431365
transform 1 0 35504 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_309
timestamp 1698431365
transform 1 0 35952 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_317
timestamp 1698431365
transform 1 0 36848 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_319
timestamp 1698431365
transform 1 0 37072 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_2
timestamp 1698431365
transform 1 0 1568 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_10
timestamp 1698431365
transform 1 0 2464 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_14
timestamp 1698431365
transform 1 0 2912 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_49
timestamp 1698431365
transform 1 0 6832 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_57
timestamp 1698431365
transform 1 0 7728 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_61
timestamp 1698431365
transform 1 0 8176 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_63
timestamp 1698431365
transform 1 0 8400 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_66
timestamp 1698431365
transform 1 0 8736 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_72
timestamp 1698431365
transform 1 0 9408 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_74
timestamp 1698431365
transform 1 0 9632 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_138
timestamp 1698431365
transform 1 0 16800 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_150
timestamp 1698431365
transform 1 0 18144 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_154
timestamp 1698431365
transform 1 0 18592 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_170
timestamp 1698431365
transform 1 0 20384 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_187
timestamp 1698431365
transform 1 0 22288 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_193
timestamp 1698431365
transform 1 0 22960 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_199
timestamp 1698431365
transform 1 0 23632 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_203
timestamp 1698431365
transform 1 0 24080 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_205
timestamp 1698431365
transform 1 0 24304 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_208
timestamp 1698431365
transform 1 0 24640 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_212
timestamp 1698431365
transform 1 0 25088 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_228
timestamp 1698431365
transform 1 0 26880 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_235
timestamp 1698431365
transform 1 0 27664 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_273
timestamp 1698431365
transform 1 0 31920 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_277
timestamp 1698431365
transform 1 0 32368 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_279
timestamp 1698431365
transform 1 0 32592 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_318
timestamp 1698431365
transform 1 0 36960 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_322
timestamp 1698431365
transform 1 0 37408 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_385
timestamp 1698431365
transform 1 0 44464 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_37
timestamp 1698431365
transform 1 0 5488 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_41
timestamp 1698431365
transform 1 0 5936 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_57
timestamp 1698431365
transform 1 0 7728 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_65
timestamp 1698431365
transform 1 0 8624 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_69
timestamp 1698431365
transform 1 0 9072 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_73
timestamp 1698431365
transform 1 0 9520 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_87
timestamp 1698431365
transform 1 0 11088 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_89
timestamp 1698431365
transform 1 0 11312 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_92
timestamp 1698431365
transform 1 0 11648 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_100
timestamp 1698431365
transform 1 0 12544 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_102
timestamp 1698431365
transform 1 0 12768 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_117
timestamp 1698431365
transform 1 0 14448 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_121
timestamp 1698431365
transform 1 0 14896 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_129
timestamp 1698431365
transform 1 0 15792 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_131
timestamp 1698431365
transform 1 0 16016 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_134
timestamp 1698431365
transform 1 0 16352 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_142
timestamp 1698431365
transform 1 0 17248 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_146
timestamp 1698431365
transform 1 0 17696 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_150
timestamp 1698431365
transform 1 0 18144 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_171
timestamp 1698431365
transform 1 0 20496 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_177
timestamp 1698431365
transform 1 0 21168 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_179
timestamp 1698431365
transform 1 0 21392 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_186
timestamp 1698431365
transform 1 0 22176 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_219
timestamp 1698431365
transform 1 0 25872 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_227
timestamp 1698431365
transform 1 0 26768 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_229
timestamp 1698431365
transform 1 0 26992 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_238
timestamp 1698431365
transform 1 0 28000 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_242
timestamp 1698431365
transform 1 0 28448 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_247
timestamp 1698431365
transform 1 0 29008 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_259
timestamp 1698431365
transform 1 0 30352 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_273
timestamp 1698431365
transform 1 0 31920 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_277
timestamp 1698431365
transform 1 0 32368 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_281
timestamp 1698431365
transform 1 0 32816 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_288
timestamp 1698431365
transform 1 0 33600 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_290
timestamp 1698431365
transform 1 0 33824 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_293
timestamp 1698431365
transform 1 0 34160 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_297
timestamp 1698431365
transform 1 0 34608 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_323
timestamp 1698431365
transform 1 0 37520 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_327
timestamp 1698431365
transform 1 0 37968 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_329
timestamp 1698431365
transform 1 0 38192 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_373
timestamp 1698431365
transform 1 0 43120 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_387
timestamp 1698431365
transform 1 0 44688 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_2
timestamp 1698431365
transform 1 0 1568 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_18
timestamp 1698431365
transform 1 0 3360 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_20
timestamp 1698431365
transform 1 0 3584 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_72
timestamp 1698431365
transform 1 0 9408 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_76
timestamp 1698431365
transform 1 0 9856 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_85
timestamp 1698431365
transform 1 0 10864 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_130
timestamp 1698431365
transform 1 0 15904 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_138
timestamp 1698431365
transform 1 0 16800 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_142
timestamp 1698431365
transform 1 0 17248 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_146
timestamp 1698431365
transform 1 0 17696 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_150
timestamp 1698431365
transform 1 0 18144 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_154
timestamp 1698431365
transform 1 0 18592 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_158
timestamp 1698431365
transform 1 0 19040 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_160
timestamp 1698431365
transform 1 0 19264 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_191
timestamp 1698431365
transform 1 0 22736 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_195
timestamp 1698431365
transform 1 0 23184 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_203
timestamp 1698431365
transform 1 0 24080 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_207
timestamp 1698431365
transform 1 0 24528 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_209
timestamp 1698431365
transform 1 0 24752 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_212
timestamp 1698431365
transform 1 0 25088 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_220
timestamp 1698431365
transform 1 0 25984 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_242
timestamp 1698431365
transform 1 0 28448 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_246
timestamp 1698431365
transform 1 0 28896 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_250
timestamp 1698431365
transform 1 0 29344 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_254
timestamp 1698431365
transform 1 0 29792 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_257
timestamp 1698431365
transform 1 0 30128 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_261
timestamp 1698431365
transform 1 0 30576 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_265
timestamp 1698431365
transform 1 0 31024 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_269
timestamp 1698431365
transform 1 0 31472 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_273
timestamp 1698431365
transform 1 0 31920 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_277
timestamp 1698431365
transform 1 0 32368 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_282
timestamp 1698431365
transform 1 0 32928 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_289
timestamp 1698431365
transform 1 0 33712 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_293
timestamp 1698431365
transform 1 0 34160 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_304
timestamp 1698431365
transform 1 0 35392 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_306
timestamp 1698431365
transform 1 0 35616 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_309
timestamp 1698431365
transform 1 0 35952 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_322
timestamp 1698431365
transform 1 0 37408 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_324
timestamp 1698431365
transform 1 0 37632 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_327
timestamp 1698431365
transform 1 0 37968 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_338
timestamp 1698431365
transform 1 0 39200 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_342
timestamp 1698431365
transform 1 0 39648 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_346
timestamp 1698431365
transform 1 0 40096 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_352
timestamp 1698431365
transform 1 0 40768 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_356
timestamp 1698431365
transform 1 0 41216 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_31
timestamp 1698431365
transform 1 0 4816 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_37
timestamp 1698431365
transform 1 0 5488 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_62
timestamp 1698431365
transform 1 0 8288 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_72
timestamp 1698431365
transform 1 0 9408 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_94
timestamp 1698431365
transform 1 0 11872 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_96
timestamp 1698431365
transform 1 0 12096 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_107
timestamp 1698431365
transform 1 0 13328 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_166
timestamp 1698431365
transform 1 0 19936 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_170
timestamp 1698431365
transform 1 0 20384 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_174
timestamp 1698431365
transform 1 0 20832 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_177
timestamp 1698431365
transform 1 0 21168 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_252
timestamp 1698431365
transform 1 0 29568 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_254
timestamp 1698431365
transform 1 0 29792 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_290
timestamp 1698431365
transform 1 0 33824 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_294
timestamp 1698431365
transform 1 0 34272 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_317
timestamp 1698431365
transform 1 0 36848 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_323
timestamp 1698431365
transform 1 0 37520 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_387
timestamp 1698431365
transform 1 0 44688 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_393
timestamp 1698431365
transform 1 0 45360 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_9_2
timestamp 1698431365
transform 1 0 1568 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_18
timestamp 1698431365
transform 1 0 3360 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_26
timestamp 1698431365
transform 1 0 4256 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_38
timestamp 1698431365
transform 1 0 5600 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_42
timestamp 1698431365
transform 1 0 6048 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_49
timestamp 1698431365
transform 1 0 6832 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_53
timestamp 1698431365
transform 1 0 7280 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_56
timestamp 1698431365
transform 1 0 7616 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_68
timestamp 1698431365
transform 1 0 8960 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_88
timestamp 1698431365
transform 1 0 11200 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_90
timestamp 1698431365
transform 1 0 11424 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_120
timestamp 1698431365
transform 1 0 14784 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_124
timestamp 1698431365
transform 1 0 15232 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_136
timestamp 1698431365
transform 1 0 16576 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_142
timestamp 1698431365
transform 1 0 17248 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_9_146
timestamp 1698431365
transform 1 0 17696 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_162
timestamp 1698431365
transform 1 0 19488 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_166
timestamp 1698431365
transform 1 0 19936 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_168
timestamp 1698431365
transform 1 0 20160 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_198
timestamp 1698431365
transform 1 0 23520 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_206
timestamp 1698431365
transform 1 0 24416 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_255
timestamp 1698431365
transform 1 0 29904 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_259
timestamp 1698431365
transform 1 0 30352 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_274
timestamp 1698431365
transform 1 0 32032 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_344
timestamp 1698431365
transform 1 0 39872 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_352
timestamp 1698431365
transform 1 0 40768 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_367
timestamp 1698431365
transform 1 0 42448 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_371
timestamp 1698431365
transform 1 0 42896 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_373
timestamp 1698431365
transform 1 0 43120 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_418
timestamp 1698431365
transform 1 0 48160 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_43
timestamp 1698431365
transform 1 0 6160 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_47
timestamp 1698431365
transform 1 0 6608 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_55
timestamp 1698431365
transform 1 0 7504 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_90
timestamp 1698431365
transform 1 0 11424 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_113
timestamp 1698431365
transform 1 0 14000 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_117
timestamp 1698431365
transform 1 0 14448 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_133
timestamp 1698431365
transform 1 0 16240 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_141
timestamp 1698431365
transform 1 0 17136 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_145
timestamp 1698431365
transform 1 0 17584 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_177
timestamp 1698431365
transform 1 0 21168 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_181
timestamp 1698431365
transform 1 0 21616 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_189
timestamp 1698431365
transform 1 0 22512 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_224
timestamp 1698431365
transform 1 0 26432 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_232
timestamp 1698431365
transform 1 0 27328 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_236
timestamp 1698431365
transform 1 0 27776 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_238
timestamp 1698431365
transform 1 0 28000 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_259
timestamp 1698431365
transform 1 0 30352 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_269
timestamp 1698431365
transform 1 0 31472 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_299
timestamp 1698431365
transform 1 0 34832 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_303
timestamp 1698431365
transform 1 0 35280 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_309
timestamp 1698431365
transform 1 0 35952 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_313
timestamp 1698431365
transform 1 0 36400 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_321
timestamp 1698431365
transform 1 0 37296 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_325
timestamp 1698431365
transform 1 0 37744 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_349
timestamp 1698431365
transform 1 0 40432 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_379
timestamp 1698431365
transform 1 0 43792 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_2
timestamp 1698431365
transform 1 0 1568 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_10
timestamp 1698431365
transform 1 0 2464 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_38
timestamp 1698431365
transform 1 0 5600 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_40
timestamp 1698431365
transform 1 0 5824 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_72
timestamp 1698431365
transform 1 0 9408 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_76
timestamp 1698431365
transform 1 0 9856 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_90
timestamp 1698431365
transform 1 0 11424 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_94
timestamp 1698431365
transform 1 0 11872 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_98
timestamp 1698431365
transform 1 0 12320 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_102
timestamp 1698431365
transform 1 0 12768 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_104
timestamp 1698431365
transform 1 0 12992 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_107
timestamp 1698431365
transform 1 0 13328 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_111
timestamp 1698431365
transform 1 0 13776 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_115
timestamp 1698431365
transform 1 0 14224 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_119
timestamp 1698431365
transform 1 0 14672 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_121
timestamp 1698431365
transform 1 0 14896 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_132
timestamp 1698431365
transform 1 0 16128 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_142
timestamp 1698431365
transform 1 0 17248 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_146
timestamp 1698431365
transform 1 0 17696 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_148
timestamp 1698431365
transform 1 0 17920 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_165
timestamp 1698431365
transform 1 0 19824 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_169
timestamp 1698431365
transform 1 0 20272 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_185
timestamp 1698431365
transform 1 0 22064 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_195
timestamp 1698431365
transform 1 0 23184 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_199
timestamp 1698431365
transform 1 0 23632 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_206
timestamp 1698431365
transform 1 0 24416 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_212
timestamp 1698431365
transform 1 0 25088 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_220
timestamp 1698431365
transform 1 0 25984 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_261
timestamp 1698431365
transform 1 0 30576 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_276
timestamp 1698431365
transform 1 0 32256 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_282
timestamp 1698431365
transform 1 0 32928 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_284
timestamp 1698431365
transform 1 0 33152 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_287
timestamp 1698431365
transform 1 0 33488 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_291
timestamp 1698431365
transform 1 0 33936 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_295
timestamp 1698431365
transform 1 0 34384 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_299
timestamp 1698431365
transform 1 0 34832 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_311
timestamp 1698431365
transform 1 0 36176 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_360
timestamp 1698431365
transform 1 0 41664 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_408
timestamp 1698431365
transform 1 0 47040 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_418
timestamp 1698431365
transform 1 0 48160 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_45
timestamp 1698431365
transform 1 0 6384 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_49
timestamp 1698431365
transform 1 0 6832 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_65
timestamp 1698431365
transform 1 0 8624 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_92
timestamp 1698431365
transform 1 0 11648 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_100
timestamp 1698431365
transform 1 0 12544 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_102
timestamp 1698431365
transform 1 0 12768 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_148
timestamp 1698431365
transform 1 0 17920 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_152
timestamp 1698431365
transform 1 0 18368 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_156
timestamp 1698431365
transform 1 0 18816 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_158
timestamp 1698431365
transform 1 0 19040 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_161
timestamp 1698431365
transform 1 0 19376 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_170
timestamp 1698431365
transform 1 0 20384 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_174
timestamp 1698431365
transform 1 0 20832 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_214
timestamp 1698431365
transform 1 0 25312 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_218
timestamp 1698431365
transform 1 0 25760 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_240
timestamp 1698431365
transform 1 0 28224 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_242
timestamp 1698431365
transform 1 0 28448 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_247
timestamp 1698431365
transform 1 0 29008 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_291
timestamp 1698431365
transform 1 0 33936 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_317
timestamp 1698431365
transform 1 0 36848 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_319
timestamp 1698431365
transform 1 0 37072 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_365
timestamp 1698431365
transform 1 0 42224 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_2
timestamp 1698431365
transform 1 0 1568 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_18
timestamp 1698431365
transform 1 0 3360 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_26
timestamp 1698431365
transform 1 0 4256 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_37
timestamp 1698431365
transform 1 0 5488 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_67
timestamp 1698431365
transform 1 0 8848 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_69
timestamp 1698431365
transform 1 0 9072 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_72
timestamp 1698431365
transform 1 0 9408 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_87
timestamp 1698431365
transform 1 0 11088 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_105
timestamp 1698431365
transform 1 0 13104 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_138
timestamp 1698431365
transform 1 0 16800 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_142
timestamp 1698431365
transform 1 0 17248 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_146
timestamp 1698431365
transform 1 0 17696 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_153
timestamp 1698431365
transform 1 0 18480 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_191
timestamp 1698431365
transform 1 0 22736 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_212
timestamp 1698431365
transform 1 0 25088 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_216
timestamp 1698431365
transform 1 0 25536 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_220
timestamp 1698431365
transform 1 0 25984 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_223
timestamp 1698431365
transform 1 0 26320 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_244
timestamp 1698431365
transform 1 0 28672 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_273
timestamp 1698431365
transform 1 0 31920 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_277
timestamp 1698431365
transform 1 0 32368 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_279
timestamp 1698431365
transform 1 0 32592 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_282
timestamp 1698431365
transform 1 0 32928 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_284
timestamp 1698431365
transform 1 0 33152 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_311
timestamp 1698431365
transform 1 0 36176 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_313
timestamp 1698431365
transform 1 0 36400 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_367
timestamp 1698431365
transform 1 0 42448 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_371
timestamp 1698431365
transform 1 0 42896 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_418
timestamp 1698431365
transform 1 0 48160 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_31
timestamp 1698431365
transform 1 0 4816 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_37
timestamp 1698431365
transform 1 0 5488 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_45
timestamp 1698431365
transform 1 0 6384 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_49
timestamp 1698431365
transform 1 0 6832 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_87
timestamp 1698431365
transform 1 0 11088 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_107
timestamp 1698431365
transform 1 0 13328 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_191
timestamp 1698431365
transform 1 0 22736 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_213
timestamp 1698431365
transform 1 0 25200 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_215
timestamp 1698431365
transform 1 0 25424 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_235
timestamp 1698431365
transform 1 0 27664 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_239
timestamp 1698431365
transform 1 0 28112 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_247
timestamp 1698431365
transform 1 0 29008 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_255
timestamp 1698431365
transform 1 0 29904 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_269
timestamp 1698431365
transform 1 0 31472 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_285
timestamp 1698431365
transform 1 0 33264 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_297
timestamp 1698431365
transform 1 0 34608 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_299
timestamp 1698431365
transform 1 0 34832 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_314
timestamp 1698431365
transform 1 0 36512 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_317
timestamp 1698431365
transform 1 0 36848 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_387
timestamp 1698431365
transform 1 0 44688 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_2
timestamp 1698431365
transform 1 0 1568 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_18
timestamp 1698431365
transform 1 0 3360 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_26
timestamp 1698431365
transform 1 0 4256 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_28
timestamp 1698431365
transform 1 0 4480 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_43
timestamp 1698431365
transform 1 0 6160 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_57
timestamp 1698431365
transform 1 0 7728 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_65
timestamp 1698431365
transform 1 0 8624 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_69
timestamp 1698431365
transform 1 0 9072 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_76
timestamp 1698431365
transform 1 0 9856 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_78
timestamp 1698431365
transform 1 0 10080 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_81
timestamp 1698431365
transform 1 0 10416 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_127
timestamp 1698431365
transform 1 0 15568 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_131
timestamp 1698431365
transform 1 0 16016 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_138
timestamp 1698431365
transform 1 0 16800 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_148
timestamp 1698431365
transform 1 0 17920 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_164
timestamp 1698431365
transform 1 0 19712 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_198
timestamp 1698431365
transform 1 0 23520 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_200
timestamp 1698431365
transform 1 0 23744 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_212
timestamp 1698431365
transform 1 0 25088 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_216
timestamp 1698431365
transform 1 0 25536 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_238
timestamp 1698431365
transform 1 0 28000 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_242
timestamp 1698431365
transform 1 0 28448 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_244
timestamp 1698431365
transform 1 0 28672 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_247
timestamp 1698431365
transform 1 0 29008 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_251
timestamp 1698431365
transform 1 0 29456 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_253
timestamp 1698431365
transform 1 0 29680 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_256
timestamp 1698431365
transform 1 0 30016 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_264
timestamp 1698431365
transform 1 0 30912 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_275
timestamp 1698431365
transform 1 0 32144 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_279
timestamp 1698431365
transform 1 0 32592 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_288
timestamp 1698431365
transform 1 0 33600 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_310
timestamp 1698431365
transform 1 0 36064 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_319
timestamp 1698431365
transform 1 0 37072 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_321
timestamp 1698431365
transform 1 0 37296 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_329
timestamp 1698431365
transform 1 0 38192 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_331
timestamp 1698431365
transform 1 0 38416 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_352
timestamp 1698431365
transform 1 0 40768 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_354
timestamp 1698431365
transform 1 0 40992 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_364
timestamp 1698431365
transform 1 0 42112 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_368
timestamp 1698431365
transform 1 0 42560 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_372
timestamp 1698431365
transform 1 0 43008 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_374
timestamp 1698431365
transform 1 0 43232 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_418
timestamp 1698431365
transform 1 0 48160 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_31
timestamp 1698431365
transform 1 0 4816 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_37
timestamp 1698431365
transform 1 0 5488 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_41
timestamp 1698431365
transform 1 0 5936 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_45
timestamp 1698431365
transform 1 0 6384 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_49
timestamp 1698431365
transform 1 0 6832 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_63
timestamp 1698431365
transform 1 0 8400 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_71
timestamp 1698431365
transform 1 0 9296 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_79
timestamp 1698431365
transform 1 0 10192 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_87
timestamp 1698431365
transform 1 0 11088 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_91
timestamp 1698431365
transform 1 0 11536 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_133
timestamp 1698431365
transform 1 0 16240 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_137
timestamp 1698431365
transform 1 0 16688 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_144
timestamp 1698431365
transform 1 0 17472 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_152
timestamp 1698431365
transform 1 0 18368 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_154
timestamp 1698431365
transform 1 0 18592 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_170
timestamp 1698431365
transform 1 0 20384 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_172
timestamp 1698431365
transform 1 0 20608 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_197
timestamp 1698431365
transform 1 0 23408 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_213
timestamp 1698431365
transform 1 0 25200 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_215
timestamp 1698431365
transform 1 0 25424 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_222
timestamp 1698431365
transform 1 0 26208 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_230
timestamp 1698431365
transform 1 0 27104 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_234
timestamp 1698431365
transform 1 0 27552 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_236
timestamp 1698431365
transform 1 0 27776 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_261
timestamp 1698431365
transform 1 0 30576 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_275
timestamp 1698431365
transform 1 0 32144 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_283
timestamp 1698431365
transform 1 0 33040 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_287
timestamp 1698431365
transform 1 0 33488 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_289
timestamp 1698431365
transform 1 0 33712 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_312
timestamp 1698431365
transform 1 0 36288 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_314
timestamp 1698431365
transform 1 0 36512 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_343
timestamp 1698431365
transform 1 0 39760 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_370
timestamp 1698431365
transform 1 0 42784 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_380
timestamp 1698431365
transform 1 0 43904 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_382
timestamp 1698431365
transform 1 0 44128 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_405
timestamp 1698431365
transform 1 0 46704 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_417
timestamp 1698431365
transform 1 0 48048 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_419
timestamp 1698431365
transform 1 0 48272 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_2
timestamp 1698431365
transform 1 0 1568 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_10
timestamp 1698431365
transform 1 0 2464 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_12
timestamp 1698431365
transform 1 0 2688 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_36
timestamp 1698431365
transform 1 0 5376 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_44
timestamp 1698431365
transform 1 0 6272 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_46
timestamp 1698431365
transform 1 0 6496 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_49
timestamp 1698431365
transform 1 0 6832 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_51
timestamp 1698431365
transform 1 0 7056 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_62
timestamp 1698431365
transform 1 0 8288 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_66
timestamp 1698431365
transform 1 0 8736 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_78
timestamp 1698431365
transform 1 0 10080 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_119
timestamp 1698431365
transform 1 0 14672 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_123
timestamp 1698431365
transform 1 0 15120 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_127
timestamp 1698431365
transform 1 0 15568 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_138
timestamp 1698431365
transform 1 0 16800 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_150
timestamp 1698431365
transform 1 0 18144 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_183
timestamp 1698431365
transform 1 0 21840 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_185
timestamp 1698431365
transform 1 0 22064 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_202
timestamp 1698431365
transform 1 0 23968 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_206
timestamp 1698431365
transform 1 0 24416 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_218
timestamp 1698431365
transform 1 0 25760 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_230
timestamp 1698431365
transform 1 0 27104 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_262
timestamp 1698431365
transform 1 0 30688 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_275
timestamp 1698431365
transform 1 0 32144 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_279
timestamp 1698431365
transform 1 0 32592 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_307
timestamp 1698431365
transform 1 0 35728 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_309
timestamp 1698431365
transform 1 0 35952 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_331
timestamp 1698431365
transform 1 0 38416 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_349
timestamp 1698431365
transform 1 0 40432 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_392
timestamp 1698431365
transform 1 0 45248 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_415
timestamp 1698431365
transform 1 0 47824 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_419
timestamp 1698431365
transform 1 0 48272 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_28
timestamp 1698431365
transform 1 0 4480 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_94
timestamp 1698431365
transform 1 0 11872 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_96
timestamp 1698431365
transform 1 0 12096 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_107
timestamp 1698431365
transform 1 0 13328 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_140
timestamp 1698431365
transform 1 0 17024 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_142
timestamp 1698431365
transform 1 0 17248 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_149
timestamp 1698431365
transform 1 0 18032 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_153
timestamp 1698431365
transform 1 0 18480 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_155
timestamp 1698431365
transform 1 0 18704 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_170
timestamp 1698431365
transform 1 0 20384 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_174
timestamp 1698431365
transform 1 0 20832 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_177
timestamp 1698431365
transform 1 0 21168 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_187
timestamp 1698431365
transform 1 0 22288 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_191
timestamp 1698431365
transform 1 0 22736 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_207
timestamp 1698431365
transform 1 0 24528 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_215
timestamp 1698431365
transform 1 0 25424 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_247
timestamp 1698431365
transform 1 0 29008 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_260
timestamp 1698431365
transform 1 0 30464 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_262
timestamp 1698431365
transform 1 0 30688 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_265
timestamp 1698431365
transform 1 0 31024 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_269
timestamp 1698431365
transform 1 0 31472 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_284
timestamp 1698431365
transform 1 0 33152 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_292
timestamp 1698431365
transform 1 0 34048 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_311
timestamp 1698431365
transform 1 0 36176 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_372
timestamp 1698431365
transform 1 0 43008 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_374
timestamp 1698431365
transform 1 0 43232 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_387
timestamp 1698431365
transform 1 0 44688 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_41
timestamp 1698431365
transform 1 0 5936 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_45
timestamp 1698431365
transform 1 0 6384 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_49
timestamp 1698431365
transform 1 0 6832 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_62
timestamp 1698431365
transform 1 0 8288 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_66
timestamp 1698431365
transform 1 0 8736 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_72
timestamp 1698431365
transform 1 0 9408 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_76
timestamp 1698431365
transform 1 0 9856 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_78
timestamp 1698431365
transform 1 0 10080 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_81
timestamp 1698431365
transform 1 0 10416 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_112
timestamp 1698431365
transform 1 0 13888 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_122
timestamp 1698431365
transform 1 0 15008 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_138
timestamp 1698431365
transform 1 0 16800 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_142
timestamp 1698431365
transform 1 0 17248 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_146
timestamp 1698431365
transform 1 0 17696 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_150
timestamp 1698431365
transform 1 0 18144 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_167
timestamp 1698431365
transform 1 0 20048 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_171
timestamp 1698431365
transform 1 0 20496 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_173
timestamp 1698431365
transform 1 0 20720 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_207
timestamp 1698431365
transform 1 0 24528 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_209
timestamp 1698431365
transform 1 0 24752 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_221
timestamp 1698431365
transform 1 0 26096 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_236
timestamp 1698431365
transform 1 0 27776 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_238
timestamp 1698431365
transform 1 0 28000 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_244
timestamp 1698431365
transform 1 0 28672 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_263
timestamp 1698431365
transform 1 0 30800 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_279
timestamp 1698431365
transform 1 0 32592 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_308
timestamp 1698431365
transform 1 0 35840 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_338
timestamp 1698431365
transform 1 0 39200 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_352
timestamp 1698431365
transform 1 0 40768 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_354
timestamp 1698431365
transform 1 0 40992 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_372
timestamp 1698431365
transform 1 0 43008 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_407
timestamp 1698431365
transform 1 0 46928 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_2
timestamp 1698431365
transform 1 0 1568 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_8
timestamp 1698431365
transform 1 0 2240 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_12
timestamp 1698431365
transform 1 0 2688 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_16
timestamp 1698431365
transform 1 0 3136 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_34
timestamp 1698431365
transform 1 0 5152 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_37
timestamp 1698431365
transform 1 0 5488 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_41
timestamp 1698431365
transform 1 0 5936 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_45
timestamp 1698431365
transform 1 0 6384 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_49
timestamp 1698431365
transform 1 0 6832 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_52
timestamp 1698431365
transform 1 0 7168 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_56
timestamp 1698431365
transform 1 0 7616 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_67
timestamp 1698431365
transform 1 0 8848 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_73
timestamp 1698431365
transform 1 0 9520 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_91
timestamp 1698431365
transform 1 0 11536 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_95
timestamp 1698431365
transform 1 0 11984 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_99
timestamp 1698431365
transform 1 0 12432 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_107
timestamp 1698431365
transform 1 0 13328 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_126
timestamp 1698431365
transform 1 0 15456 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_130
timestamp 1698431365
transform 1 0 15904 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_183
timestamp 1698431365
transform 1 0 21840 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_187
timestamp 1698431365
transform 1 0 22288 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_218
timestamp 1698431365
transform 1 0 25760 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_230
timestamp 1698431365
transform 1 0 27104 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_238
timestamp 1698431365
transform 1 0 28000 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_242
timestamp 1698431365
transform 1 0 28448 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_268
timestamp 1698431365
transform 1 0 31360 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_270
timestamp 1698431365
transform 1 0 31584 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_306
timestamp 1698431365
transform 1 0 35616 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_317
timestamp 1698431365
transform 1 0 36848 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_319
timestamp 1698431365
transform 1 0 37072 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_369
timestamp 1698431365
transform 1 0 42672 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_373
timestamp 1698431365
transform 1 0 43120 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_2
timestamp 1698431365
transform 1 0 1568 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_8
timestamp 1698431365
transform 1 0 2240 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_12
timestamp 1698431365
transform 1 0 2688 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_15
timestamp 1698431365
transform 1 0 3024 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_80
timestamp 1698431365
transform 1 0 10304 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_119
timestamp 1698431365
transform 1 0 14672 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_121
timestamp 1698431365
transform 1 0 14896 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_142
timestamp 1698431365
transform 1 0 17248 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_150
timestamp 1698431365
transform 1 0 18144 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_157
timestamp 1698431365
transform 1 0 18928 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_165
timestamp 1698431365
transform 1 0 19824 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_167
timestamp 1698431365
transform 1 0 20048 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_183
timestamp 1698431365
transform 1 0 21840 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_199
timestamp 1698431365
transform 1 0 23632 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_207
timestamp 1698431365
transform 1 0 24528 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_209
timestamp 1698431365
transform 1 0 24752 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_212
timestamp 1698431365
transform 1 0 25088 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_248
timestamp 1698431365
transform 1 0 29120 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_252
timestamp 1698431365
transform 1 0 29568 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_254
timestamp 1698431365
transform 1 0 29792 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_260
timestamp 1698431365
transform 1 0 30464 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_264
timestamp 1698431365
transform 1 0 30912 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_268
timestamp 1698431365
transform 1 0 31360 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_277
timestamp 1698431365
transform 1 0 32368 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_279
timestamp 1698431365
transform 1 0 32592 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_282
timestamp 1698431365
transform 1 0 32928 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_286
timestamp 1698431365
transform 1 0 33376 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_294
timestamp 1698431365
transform 1 0 34272 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_386
timestamp 1698431365
transform 1 0 44576 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_388
timestamp 1698431365
transform 1 0 44800 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_31
timestamp 1698431365
transform 1 0 4816 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_37
timestamp 1698431365
transform 1 0 5488 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_39
timestamp 1698431365
transform 1 0 5712 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_63
timestamp 1698431365
transform 1 0 8400 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_72
timestamp 1698431365
transform 1 0 9408 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_74
timestamp 1698431365
transform 1 0 9632 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_77
timestamp 1698431365
transform 1 0 9968 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_100
timestamp 1698431365
transform 1 0 12544 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_104
timestamp 1698431365
transform 1 0 12992 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_127
timestamp 1698431365
transform 1 0 15568 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_129
timestamp 1698431365
transform 1 0 15792 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_139
timestamp 1698431365
transform 1 0 16912 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_143
timestamp 1698431365
transform 1 0 17360 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_177
timestamp 1698431365
transform 1 0 21168 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_186
timestamp 1698431365
transform 1 0 22176 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_190
timestamp 1698431365
transform 1 0 22624 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_205
timestamp 1698431365
transform 1 0 24304 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_217
timestamp 1698431365
transform 1 0 25648 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_227
timestamp 1698431365
transform 1 0 26768 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_235
timestamp 1698431365
transform 1 0 27664 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_243
timestamp 1698431365
transform 1 0 28560 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_247
timestamp 1698431365
transform 1 0 29008 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_255
timestamp 1698431365
transform 1 0 29904 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_259
timestamp 1698431365
transform 1 0 30352 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_311
timestamp 1698431365
transform 1 0 36176 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_317
timestamp 1698431365
transform 1 0 36848 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_327
timestamp 1698431365
transform 1 0 37968 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_358
timestamp 1698431365
transform 1 0 41440 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_383
timestamp 1698431365
transform 1 0 44240 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_387
timestamp 1698431365
transform 1 0 44688 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_31
timestamp 1698431365
transform 1 0 4816 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_35
timestamp 1698431365
transform 1 0 5264 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_47
timestamp 1698431365
transform 1 0 6608 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_67
timestamp 1698431365
transform 1 0 8848 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_69
timestamp 1698431365
transform 1 0 9072 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_72
timestamp 1698431365
transform 1 0 9408 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_76
timestamp 1698431365
transform 1 0 9856 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_124
timestamp 1698431365
transform 1 0 15232 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_128
timestamp 1698431365
transform 1 0 15680 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_132
timestamp 1698431365
transform 1 0 16128 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_136
timestamp 1698431365
transform 1 0 16576 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_177
timestamp 1698431365
transform 1 0 21168 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_202
timestamp 1698431365
transform 1 0 23968 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_212
timestamp 1698431365
transform 1 0 25088 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_228
timestamp 1698431365
transform 1 0 26880 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_232
timestamp 1698431365
transform 1 0 27328 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_234
timestamp 1698431365
transform 1 0 27552 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_240
timestamp 1698431365
transform 1 0 28224 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_258
timestamp 1698431365
transform 1 0 30240 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_278
timestamp 1698431365
transform 1 0 32480 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_308
timestamp 1698431365
transform 1 0 35840 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_316
timestamp 1698431365
transform 1 0 36736 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_348
timestamp 1698431365
transform 1 0 40320 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_372
timestamp 1698431365
transform 1 0 43008 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_402
timestamp 1698431365
transform 1 0 46368 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_404
timestamp 1698431365
transform 1 0 46592 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_31
timestamp 1698431365
transform 1 0 4816 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_37
timestamp 1698431365
transform 1 0 5488 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_50
timestamp 1698431365
transform 1 0 6944 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_62
timestamp 1698431365
transform 1 0 8288 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_64
timestamp 1698431365
transform 1 0 8512 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_82
timestamp 1698431365
transform 1 0 10528 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_86
timestamp 1698431365
transform 1 0 10976 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_88
timestamp 1698431365
transform 1 0 11200 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_91
timestamp 1698431365
transform 1 0 11536 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_95
timestamp 1698431365
transform 1 0 11984 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_99
timestamp 1698431365
transform 1 0 12432 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_115
timestamp 1698431365
transform 1 0 14224 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_150
timestamp 1698431365
transform 1 0 18144 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_160
timestamp 1698431365
transform 1 0 19264 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_168
timestamp 1698431365
transform 1 0 20160 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_172
timestamp 1698431365
transform 1 0 20608 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_174
timestamp 1698431365
transform 1 0 20832 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_177
timestamp 1698431365
transform 1 0 21168 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_181
timestamp 1698431365
transform 1 0 21616 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_187
timestamp 1698431365
transform 1 0 22288 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_201
timestamp 1698431365
transform 1 0 23856 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_205
timestamp 1698431365
transform 1 0 24304 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_209
timestamp 1698431365
transform 1 0 24752 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_211
timestamp 1698431365
transform 1 0 24976 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_241
timestamp 1698431365
transform 1 0 28336 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_276
timestamp 1698431365
transform 1 0 32256 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_282
timestamp 1698431365
transform 1 0 32928 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_296
timestamp 1698431365
transform 1 0 34496 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_312
timestamp 1698431365
transform 1 0 36288 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_314
timestamp 1698431365
transform 1 0 36512 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_317
timestamp 1698431365
transform 1 0 36848 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_321
timestamp 1698431365
transform 1 0 37296 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_325
timestamp 1698431365
transform 1 0 37744 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_380
timestamp 1698431365
transform 1 0 43904 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_382
timestamp 1698431365
transform 1 0 44128 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_387
timestamp 1698431365
transform 1 0 44688 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_8
timestamp 1698431365
transform 1 0 2240 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_12
timestamp 1698431365
transform 1 0 2688 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_16
timestamp 1698431365
transform 1 0 3136 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_20
timestamp 1698431365
transform 1 0 3584 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_22
timestamp 1698431365
transform 1 0 3808 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_25
timestamp 1698431365
transform 1 0 4144 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_58
timestamp 1698431365
transform 1 0 7840 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_109
timestamp 1698431365
transform 1 0 13552 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_119
timestamp 1698431365
transform 1 0 14672 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_123
timestamp 1698431365
transform 1 0 15120 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_129
timestamp 1698431365
transform 1 0 15792 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_133
timestamp 1698431365
transform 1 0 16240 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_142
timestamp 1698431365
transform 1 0 17248 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_146
timestamp 1698431365
transform 1 0 17696 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_177
timestamp 1698431365
transform 1 0 21168 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_185
timestamp 1698431365
transform 1 0 22064 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_209
timestamp 1698431365
transform 1 0 24752 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_212
timestamp 1698431365
transform 1 0 25088 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_237
timestamp 1698431365
transform 1 0 27888 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_245
timestamp 1698431365
transform 1 0 28784 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_255
timestamp 1698431365
transform 1 0 29904 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_276
timestamp 1698431365
transform 1 0 32256 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_282
timestamp 1698431365
transform 1 0 32928 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_298
timestamp 1698431365
transform 1 0 34720 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_315
timestamp 1698431365
transform 1 0 36624 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_323
timestamp 1698431365
transform 1 0 37520 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_347
timestamp 1698431365
transform 1 0 40208 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_349
timestamp 1698431365
transform 1 0 40432 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_358
timestamp 1698431365
transform 1 0 41440 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_368
timestamp 1698431365
transform 1 0 42560 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_398
timestamp 1698431365
transform 1 0 45920 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_400
timestamp 1698431365
transform 1 0 46144 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_416
timestamp 1698431365
transform 1 0 47936 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_31
timestamp 1698431365
transform 1 0 4816 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_37
timestamp 1698431365
transform 1 0 5488 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_43
timestamp 1698431365
transform 1 0 6160 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_84
timestamp 1698431365
transform 1 0 10752 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_94
timestamp 1698431365
transform 1 0 11872 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_98
timestamp 1698431365
transform 1 0 12320 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_101
timestamp 1698431365
transform 1 0 12656 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_153
timestamp 1698431365
transform 1 0 18480 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_177
timestamp 1698431365
transform 1 0 21168 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_185
timestamp 1698431365
transform 1 0 22064 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_255
timestamp 1698431365
transform 1 0 29904 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_291
timestamp 1698431365
transform 1 0 33936 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_299
timestamp 1698431365
transform 1 0 34832 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_303
timestamp 1698431365
transform 1 0 35280 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_311
timestamp 1698431365
transform 1 0 36176 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_337
timestamp 1698431365
transform 1 0 39088 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_339
timestamp 1698431365
transform 1 0 39312 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_363
timestamp 1698431365
transform 1 0 42000 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_367
timestamp 1698431365
transform 1 0 42448 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_382
timestamp 1698431365
transform 1 0 44128 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_384
timestamp 1698431365
transform 1 0 44352 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_387
timestamp 1698431365
transform 1 0 44688 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_16
timestamp 1698431365
transform 1 0 3136 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_20
timestamp 1698431365
transform 1 0 3584 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_23
timestamp 1698431365
transform 1 0 3920 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_27
timestamp 1698431365
transform 1 0 4368 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_31
timestamp 1698431365
transform 1 0 4816 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_35
timestamp 1698431365
transform 1 0 5264 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_39
timestamp 1698431365
transform 1 0 5712 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_118
timestamp 1698431365
transform 1 0 14560 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_120
timestamp 1698431365
transform 1 0 14784 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_123
timestamp 1698431365
transform 1 0 15120 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_127
timestamp 1698431365
transform 1 0 15568 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_129
timestamp 1698431365
transform 1 0 15792 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_142
timestamp 1698431365
transform 1 0 17248 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_152
timestamp 1698431365
transform 1 0 18368 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_156
timestamp 1698431365
transform 1 0 18816 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_159
timestamp 1698431365
transform 1 0 19152 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_181
timestamp 1698431365
transform 1 0 21616 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_185
timestamp 1698431365
transform 1 0 22064 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_189
timestamp 1698431365
transform 1 0 22512 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_191
timestamp 1698431365
transform 1 0 22736 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_198
timestamp 1698431365
transform 1 0 23520 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_206
timestamp 1698431365
transform 1 0 24416 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_270
timestamp 1698431365
transform 1 0 31584 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_278
timestamp 1698431365
transform 1 0 32480 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_282
timestamp 1698431365
transform 1 0 32928 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_290
timestamp 1698431365
transform 1 0 33824 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_309
timestamp 1698431365
transform 1 0 35952 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_325
timestamp 1698431365
transform 1 0 37744 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_329
timestamp 1698431365
transform 1 0 38192 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_340
timestamp 1698431365
transform 1 0 39424 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_344
timestamp 1698431365
transform 1 0 39872 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_346
timestamp 1698431365
transform 1 0 40096 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_349
timestamp 1698431365
transform 1 0 40432 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_352
timestamp 1698431365
transform 1 0 40768 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_356
timestamp 1698431365
transform 1 0 41216 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_360
timestamp 1698431365
transform 1 0 41664 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_362
timestamp 1698431365
transform 1 0 41888 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_377
timestamp 1698431365
transform 1 0 43568 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_381
timestamp 1698431365
transform 1 0 44016 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_31
timestamp 1698431365
transform 1 0 4816 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_37
timestamp 1698431365
transform 1 0 5488 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_39
timestamp 1698431365
transform 1 0 5712 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_73
timestamp 1698431365
transform 1 0 9520 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_111
timestamp 1698431365
transform 1 0 13776 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_113
timestamp 1698431365
transform 1 0 14000 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_143
timestamp 1698431365
transform 1 0 17360 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_159
timestamp 1698431365
transform 1 0 19152 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_177
timestamp 1698431365
transform 1 0 21168 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_181
timestamp 1698431365
transform 1 0 21616 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_185
timestamp 1698431365
transform 1 0 22064 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_189
timestamp 1698431365
transform 1 0 22512 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_193
timestamp 1698431365
transform 1 0 22960 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_229
timestamp 1698431365
transform 1 0 26992 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_247
timestamp 1698431365
transform 1 0 29008 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_277
timestamp 1698431365
transform 1 0 32368 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_285
timestamp 1698431365
transform 1 0 33264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_287
timestamp 1698431365
transform 1 0 33488 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_294
timestamp 1698431365
transform 1 0 34272 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_298
timestamp 1698431365
transform 1 0 34720 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_308
timestamp 1698431365
transform 1 0 35840 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_312
timestamp 1698431365
transform 1 0 36288 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_314
timestamp 1698431365
transform 1 0 36512 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_317
timestamp 1698431365
transform 1 0 36848 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_335
timestamp 1698431365
transform 1 0 38864 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_337
timestamp 1698431365
transform 1 0 39088 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_380
timestamp 1698431365
transform 1 0 43904 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_384
timestamp 1698431365
transform 1 0 44352 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_387
timestamp 1698431365
transform 1 0 44688 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_2
timestamp 1698431365
transform 1 0 1568 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_35
timestamp 1698431365
transform 1 0 5264 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_62
timestamp 1698431365
transform 1 0 8288 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_86
timestamp 1698431365
transform 1 0 10976 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_118
timestamp 1698431365
transform 1 0 14560 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_135
timestamp 1698431365
transform 1 0 16464 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_137
timestamp 1698431365
transform 1 0 16688 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_142
timestamp 1698431365
transform 1 0 17248 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_155
timestamp 1698431365
transform 1 0 18704 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_157
timestamp 1698431365
transform 1 0 18928 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_193
timestamp 1698431365
transform 1 0 22960 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_212
timestamp 1698431365
transform 1 0 25088 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_220
timestamp 1698431365
transform 1 0 25984 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_239
timestamp 1698431365
transform 1 0 28112 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_271
timestamp 1698431365
transform 1 0 31696 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_279
timestamp 1698431365
transform 1 0 32592 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_348
timestamp 1698431365
transform 1 0 40320 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_360
timestamp 1698431365
transform 1 0 41664 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_390
timestamp 1698431365
transform 1 0 45024 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_10
timestamp 1698431365
transform 1 0 2464 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_26
timestamp 1698431365
transform 1 0 4256 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_55
timestamp 1698431365
transform 1 0 7504 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_76
timestamp 1698431365
transform 1 0 9856 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_78
timestamp 1698431365
transform 1 0 10080 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_119
timestamp 1698431365
transform 1 0 14672 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_121
timestamp 1698431365
transform 1 0 14896 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_132
timestamp 1698431365
transform 1 0 16128 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_177
timestamp 1698431365
transform 1 0 21168 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_209
timestamp 1698431365
transform 1 0 24752 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_213
timestamp 1698431365
transform 1 0 25200 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_215
timestamp 1698431365
transform 1 0 25424 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_247
timestamp 1698431365
transform 1 0 29008 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_255
timestamp 1698431365
transform 1 0 29904 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_278
timestamp 1698431365
transform 1 0 32480 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_300
timestamp 1698431365
transform 1 0 34944 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_308
timestamp 1698431365
transform 1 0 35840 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_312
timestamp 1698431365
transform 1 0 36288 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_314
timestamp 1698431365
transform 1 0 36512 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_317
timestamp 1698431365
transform 1 0 36848 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_321
timestamp 1698431365
transform 1 0 37296 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_323
timestamp 1698431365
transform 1 0 37520 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_332
timestamp 1698431365
transform 1 0 38528 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_340
timestamp 1698431365
transform 1 0 39424 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_347
timestamp 1698431365
transform 1 0 40208 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_387
timestamp 1698431365
transform 1 0 44688 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_39
timestamp 1698431365
transform 1 0 5712 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_41
timestamp 1698431365
transform 1 0 5936 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_54
timestamp 1698431365
transform 1 0 7392 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_58
timestamp 1698431365
transform 1 0 7840 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_86
timestamp 1698431365
transform 1 0 10976 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_139
timestamp 1698431365
transform 1 0 16912 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_142
timestamp 1698431365
transform 1 0 17248 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_149
timestamp 1698431365
transform 1 0 18032 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_195
timestamp 1698431365
transform 1 0 23184 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_199
timestamp 1698431365
transform 1 0 23632 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_209
timestamp 1698431365
transform 1 0 24752 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_212
timestamp 1698431365
transform 1 0 25088 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_220
timestamp 1698431365
transform 1 0 25984 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_222
timestamp 1698431365
transform 1 0 26208 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_235
timestamp 1698431365
transform 1 0 27664 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_243
timestamp 1698431365
transform 1 0 28560 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_247
timestamp 1698431365
transform 1 0 29008 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_249
timestamp 1698431365
transform 1 0 29232 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_279
timestamp 1698431365
transform 1 0 32592 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_282
timestamp 1698431365
transform 1 0 32928 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_286
timestamp 1698431365
transform 1 0 33376 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_316
timestamp 1698431365
transform 1 0 36736 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_320
timestamp 1698431365
transform 1 0 37184 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_352
timestamp 1698431365
transform 1 0 40768 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_354
timestamp 1698431365
transform 1 0 40992 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_361
timestamp 1698431365
transform 1 0 41776 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_396
timestamp 1698431365
transform 1 0 45696 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_398
timestamp 1698431365
transform 1 0 45920 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_416
timestamp 1698431365
transform 1 0 47936 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_2
timestamp 1698431365
transform 1 0 1568 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_20
timestamp 1698431365
transform 1 0 3584 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_41
timestamp 1698431365
transform 1 0 5936 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_52
timestamp 1698431365
transform 1 0 7168 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_54
timestamp 1698431365
transform 1 0 7392 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_63
timestamp 1698431365
transform 1 0 8400 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_84
timestamp 1698431365
transform 1 0 10752 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_86
timestamp 1698431365
transform 1 0 10976 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_133
timestamp 1698431365
transform 1 0 16240 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_135
timestamp 1698431365
transform 1 0 16464 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_150
timestamp 1698431365
transform 1 0 18144 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_159
timestamp 1698431365
transform 1 0 19152 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_214
timestamp 1698431365
transform 1 0 25312 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_216
timestamp 1698431365
transform 1 0 25536 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_234
timestamp 1698431365
transform 1 0 27552 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_242
timestamp 1698431365
transform 1 0 28448 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_244
timestamp 1698431365
transform 1 0 28672 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_255
timestamp 1698431365
transform 1 0 29904 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_257
timestamp 1698431365
transform 1 0 30128 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_275
timestamp 1698431365
transform 1 0 32144 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_279
timestamp 1698431365
transform 1 0 32592 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_281
timestamp 1698431365
transform 1 0 32816 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_288
timestamp 1698431365
transform 1 0 33600 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_296
timestamp 1698431365
transform 1 0 34496 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_298
timestamp 1698431365
transform 1 0 34720 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_314
timestamp 1698431365
transform 1 0 36512 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_317
timestamp 1698431365
transform 1 0 36848 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_321
timestamp 1698431365
transform 1 0 37296 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_328
timestamp 1698431365
transform 1 0 38080 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_336
timestamp 1698431365
transform 1 0 38976 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_344
timestamp 1698431365
transform 1 0 39872 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_348
timestamp 1698431365
transform 1 0 40320 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_350
timestamp 1698431365
transform 1 0 40544 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_368
timestamp 1698431365
transform 1 0 42560 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_393
timestamp 1698431365
transform 1 0 45360 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_69
timestamp 1698431365
transform 1 0 9072 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_96
timestamp 1698431365
transform 1 0 12096 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_164
timestamp 1698431365
transform 1 0 19712 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_166
timestamp 1698431365
transform 1 0 19936 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_186
timestamp 1698431365
transform 1 0 22176 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_212
timestamp 1698431365
transform 1 0 25088 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_220
timestamp 1698431365
transform 1 0 25984 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_222
timestamp 1698431365
transform 1 0 26208 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_236
timestamp 1698431365
transform 1 0 27776 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_269
timestamp 1698431365
transform 1 0 31472 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_277
timestamp 1698431365
transform 1 0 32368 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_279
timestamp 1698431365
transform 1 0 32592 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_311
timestamp 1698431365
transform 1 0 36176 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_319
timestamp 1698431365
transform 1 0 37072 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_342
timestamp 1698431365
transform 1 0 39648 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_346
timestamp 1698431365
transform 1 0 40096 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_381
timestamp 1698431365
transform 1 0 44016 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_385
timestamp 1698431365
transform 1 0 44464 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_387
timestamp 1698431365
transform 1 0 44688 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_28
timestamp 1698431365
transform 1 0 4480 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_32
timestamp 1698431365
transform 1 0 4928 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_76
timestamp 1698431365
transform 1 0 9856 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_90
timestamp 1698431365
transform 1 0 11424 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_98
timestamp 1698431365
transform 1 0 12320 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_139
timestamp 1698431365
transform 1 0 16912 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_177
timestamp 1698431365
transform 1 0 21168 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_205
timestamp 1698431365
transform 1 0 24304 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_34_209
timestamp 1698431365
transform 1 0 24752 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_225
timestamp 1698431365
transform 1 0 26544 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_231
timestamp 1698431365
transform 1 0 27216 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_239
timestamp 1698431365
transform 1 0 28112 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_243
timestamp 1698431365
transform 1 0 28560 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_247
timestamp 1698431365
transform 1 0 29008 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_259
timestamp 1698431365
transform 1 0 30352 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_291
timestamp 1698431365
transform 1 0 33936 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_309
timestamp 1698431365
transform 1 0 35952 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_313
timestamp 1698431365
transform 1 0 36400 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_346
timestamp 1698431365
transform 1 0 40096 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_354
timestamp 1698431365
transform 1 0 40992 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_34_361
timestamp 1698431365
transform 1 0 41776 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_377
timestamp 1698431365
transform 1 0 43568 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_387
timestamp 1698431365
transform 1 0 44688 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_37
timestamp 1698431365
transform 1 0 5488 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_65
timestamp 1698431365
transform 1 0 8624 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_69
timestamp 1698431365
transform 1 0 9072 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_81
timestamp 1698431365
transform 1 0 10416 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_85
timestamp 1698431365
transform 1 0 10864 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_107
timestamp 1698431365
transform 1 0 13328 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_121
timestamp 1698431365
transform 1 0 14896 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_123
timestamp 1698431365
transform 1 0 15120 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_142
timestamp 1698431365
transform 1 0 17248 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_144
timestamp 1698431365
transform 1 0 17472 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_195
timestamp 1698431365
transform 1 0 23184 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_241
timestamp 1698431365
transform 1 0 28336 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_255
timestamp 1698431365
transform 1 0 29904 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_259
timestamp 1698431365
transform 1 0 30352 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_275
timestamp 1698431365
transform 1 0 32144 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_279
timestamp 1698431365
transform 1 0 32592 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_282
timestamp 1698431365
transform 1 0 32928 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_284
timestamp 1698431365
transform 1 0 33152 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_291
timestamp 1698431365
transform 1 0 33936 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_336
timestamp 1698431365
transform 1 0 38976 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_352
timestamp 1698431365
transform 1 0 40768 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_368
timestamp 1698431365
transform 1 0 42560 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_419
timestamp 1698431365
transform 1 0 48272 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_10
timestamp 1698431365
transform 1 0 2464 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_12
timestamp 1698431365
transform 1 0 2688 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_33
timestamp 1698431365
transform 1 0 5040 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_37
timestamp 1698431365
transform 1 0 5488 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_39
timestamp 1698431365
transform 1 0 5712 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_42
timestamp 1698431365
transform 1 0 6048 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_53
timestamp 1698431365
transform 1 0 7280 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_57
timestamp 1698431365
transform 1 0 7728 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_59
timestamp 1698431365
transform 1 0 7952 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_107
timestamp 1698431365
transform 1 0 13328 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_177
timestamp 1698431365
transform 1 0 21168 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_181
timestamp 1698431365
transform 1 0 21616 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_183
timestamp 1698431365
transform 1 0 21840 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_198
timestamp 1698431365
transform 1 0 23520 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_239
timestamp 1698431365
transform 1 0 28112 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_243
timestamp 1698431365
transform 1 0 28560 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_305
timestamp 1698431365
transform 1 0 35504 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_313
timestamp 1698431365
transform 1 0 36400 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_317
timestamp 1698431365
transform 1 0 36848 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_319
timestamp 1698431365
transform 1 0 37072 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_366
timestamp 1698431365
transform 1 0 42336 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_393
timestamp 1698431365
transform 1 0 45360 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_10
timestamp 1698431365
transform 1 0 2464 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_31
timestamp 1698431365
transform 1 0 4816 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_35
timestamp 1698431365
transform 1 0 5264 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_47
timestamp 1698431365
transform 1 0 6608 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_51
timestamp 1698431365
transform 1 0 7056 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_63
timestamp 1698431365
transform 1 0 8400 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_67
timestamp 1698431365
transform 1 0 8848 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_72
timestamp 1698431365
transform 1 0 9408 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_125
timestamp 1698431365
transform 1 0 15344 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_139
timestamp 1698431365
transform 1 0 16912 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_146
timestamp 1698431365
transform 1 0 17696 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_150
timestamp 1698431365
transform 1 0 18144 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_154
timestamp 1698431365
transform 1 0 18592 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_156
timestamp 1698431365
transform 1 0 18816 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_159
timestamp 1698431365
transform 1 0 19152 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_165
timestamp 1698431365
transform 1 0 19824 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_169
timestamp 1698431365
transform 1 0 20272 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_173
timestamp 1698431365
transform 1 0 20720 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_176
timestamp 1698431365
transform 1 0 21056 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_180
timestamp 1698431365
transform 1 0 21504 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_187
timestamp 1698431365
transform 1 0 22288 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_189
timestamp 1698431365
transform 1 0 22512 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_205
timestamp 1698431365
transform 1 0 24304 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_209
timestamp 1698431365
transform 1 0 24752 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_212
timestamp 1698431365
transform 1 0 25088 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_220
timestamp 1698431365
transform 1 0 25984 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_37_227
timestamp 1698431365
transform 1 0 26768 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_243
timestamp 1698431365
transform 1 0 28560 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_247
timestamp 1698431365
transform 1 0 29008 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_249
timestamp 1698431365
transform 1 0 29232 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_256
timestamp 1698431365
transform 1 0 30016 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_279
timestamp 1698431365
transform 1 0 32592 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_37_282
timestamp 1698431365
transform 1 0 32928 0 -1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_314
timestamp 1698431365
transform 1 0 36512 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_316
timestamp 1698431365
transform 1 0 36736 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_323
timestamp 1698431365
transform 1 0 37520 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_327
timestamp 1698431365
transform 1 0 37968 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_352
timestamp 1698431365
transform 1 0 40768 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_8
timestamp 1698431365
transform 1 0 2240 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_10
timestamp 1698431365
transform 1 0 2464 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_33
timestamp 1698431365
transform 1 0 5040 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_37
timestamp 1698431365
transform 1 0 5488 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_39
timestamp 1698431365
transform 1 0 5712 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_107
timestamp 1698431365
transform 1 0 13328 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_109
timestamp 1698431365
transform 1 0 13552 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_130
timestamp 1698431365
transform 1 0 15904 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_189
timestamp 1698431365
transform 1 0 22512 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_191
timestamp 1698431365
transform 1 0 22736 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_208
timestamp 1698431365
transform 1 0 24640 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_212
timestamp 1698431365
transform 1 0 25088 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_216
timestamp 1698431365
transform 1 0 25536 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_218
timestamp 1698431365
transform 1 0 25760 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_38_225
timestamp 1698431365
transform 1 0 26544 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_241
timestamp 1698431365
transform 1 0 28336 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_284
timestamp 1698431365
transform 1 0 33152 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_288
timestamp 1698431365
transform 1 0 33600 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_296
timestamp 1698431365
transform 1 0 34496 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_312
timestamp 1698431365
transform 1 0 36288 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_314
timestamp 1698431365
transform 1 0 36512 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_317
timestamp 1698431365
transform 1 0 36848 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_319
timestamp 1698431365
transform 1 0 37072 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_354
timestamp 1698431365
transform 1 0 40992 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_358
timestamp 1698431365
transform 1 0 41440 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_387
timestamp 1698431365
transform 1 0 44688 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_16
timestamp 1698431365
transform 1 0 3136 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_27
timestamp 1698431365
transform 1 0 4368 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_51
timestamp 1698431365
transform 1 0 7056 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_55
timestamp 1698431365
transform 1 0 7504 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_64
timestamp 1698431365
transform 1 0 8512 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_85
timestamp 1698431365
transform 1 0 10864 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_198
timestamp 1698431365
transform 1 0 23520 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_279
timestamp 1698431365
transform 1 0 32592 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_319
timestamp 1698431365
transform 1 0 37072 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_349
timestamp 1698431365
transform 1 0 40432 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_389
timestamp 1698431365
transform 1 0 44912 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_393
timestamp 1698431365
transform 1 0 45360 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_25
timestamp 1698431365
transform 1 0 4144 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_31
timestamp 1698431365
transform 1 0 4816 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_45
timestamp 1698431365
transform 1 0 6384 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_63
timestamp 1698431365
transform 1 0 8400 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_76
timestamp 1698431365
transform 1 0 9856 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_107
timestamp 1698431365
transform 1 0 13328 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_138
timestamp 1698431365
transform 1 0 16800 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_140
timestamp 1698431365
transform 1 0 17024 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_173
timestamp 1698431365
transform 1 0 20720 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_187
timestamp 1698431365
transform 1 0 22288 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_201
timestamp 1698431365
transform 1 0 23856 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_205
timestamp 1698431365
transform 1 0 24304 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_212
timestamp 1698431365
transform 1 0 25088 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_216
timestamp 1698431365
transform 1 0 25536 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_218
timestamp 1698431365
transform 1 0 25760 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_230
timestamp 1698431365
transform 1 0 27104 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_238
timestamp 1698431365
transform 1 0 28000 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_242
timestamp 1698431365
transform 1 0 28448 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_244
timestamp 1698431365
transform 1 0 28672 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_291
timestamp 1698431365
transform 1 0 33936 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_301
timestamp 1698431365
transform 1 0 35056 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_309
timestamp 1698431365
transform 1 0 35952 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_313
timestamp 1698431365
transform 1 0 36400 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_317
timestamp 1698431365
transform 1 0 36848 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_347
timestamp 1698431365
transform 1 0 40208 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_351
timestamp 1698431365
transform 1 0 40656 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_383
timestamp 1698431365
transform 1 0 44240 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_387
timestamp 1698431365
transform 1 0 44688 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_2
timestamp 1698431365
transform 1 0 1568 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_4
timestamp 1698431365
transform 1 0 1792 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_34
timestamp 1698431365
transform 1 0 5152 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_36
timestamp 1698431365
transform 1 0 5376 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_52
timestamp 1698431365
transform 1 0 7168 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_72
timestamp 1698431365
transform 1 0 9408 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_81
timestamp 1698431365
transform 1 0 10416 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_87
timestamp 1698431365
transform 1 0 11088 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_142
timestamp 1698431365
transform 1 0 17248 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_208
timestamp 1698431365
transform 1 0 24640 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_212
timestamp 1698431365
transform 1 0 25088 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_216
timestamp 1698431365
transform 1 0 25536 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_282
timestamp 1698431365
transform 1 0 32928 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_286
timestamp 1698431365
transform 1 0 33376 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_294
timestamp 1698431365
transform 1 0 34272 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_310
timestamp 1698431365
transform 1 0 36064 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_318
timestamp 1698431365
transform 1 0 36960 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_322
timestamp 1698431365
transform 1 0 37408 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_339
timestamp 1698431365
transform 1 0 39312 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_343
timestamp 1698431365
transform 1 0 39760 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_345
timestamp 1698431365
transform 1 0 39984 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_348
timestamp 1698431365
transform 1 0 40320 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_352
timestamp 1698431365
transform 1 0 40768 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_358
timestamp 1698431365
transform 1 0 41440 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_417
timestamp 1698431365
transform 1 0 48048 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_419
timestamp 1698431365
transform 1 0 48272 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_31
timestamp 1698431365
transform 1 0 4816 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_60
timestamp 1698431365
transform 1 0 8064 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_62
timestamp 1698431365
transform 1 0 8288 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_65
timestamp 1698431365
transform 1 0 8624 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_69
timestamp 1698431365
transform 1 0 9072 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_93
timestamp 1698431365
transform 1 0 11760 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_97
timestamp 1698431365
transform 1 0 12208 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_107
timestamp 1698431365
transform 1 0 13328 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_177
timestamp 1698431365
transform 1 0 21168 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_199
timestamp 1698431365
transform 1 0 23632 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_236
timestamp 1698431365
transform 1 0 27776 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_240
timestamp 1698431365
transform 1 0 28224 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_244
timestamp 1698431365
transform 1 0 28672 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_247
timestamp 1698431365
transform 1 0 29008 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_314
timestamp 1698431365
transform 1 0 36512 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_346
timestamp 1698431365
transform 1 0 40096 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_353
timestamp 1698431365
transform 1 0 40880 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_393
timestamp 1698431365
transform 1 0 45360 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_8
timestamp 1698431365
transform 1 0 2240 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_12
timestamp 1698431365
transform 1 0 2688 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_16
timestamp 1698431365
transform 1 0 3136 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_39
timestamp 1698431365
transform 1 0 5712 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_48
timestamp 1698431365
transform 1 0 6720 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_56
timestamp 1698431365
transform 1 0 7616 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_58
timestamp 1698431365
transform 1 0 7840 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_72
timestamp 1698431365
transform 1 0 9408 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_74
timestamp 1698431365
transform 1 0 9632 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_132
timestamp 1698431365
transform 1 0 16128 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_139
timestamp 1698431365
transform 1 0 16912 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_142
timestamp 1698431365
transform 1 0 17248 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_148
timestamp 1698431365
transform 1 0 17920 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_152
timestamp 1698431365
transform 1 0 18368 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_156
timestamp 1698431365
transform 1 0 18816 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_207
timestamp 1698431365
transform 1 0 24528 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_209
timestamp 1698431365
transform 1 0 24752 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_43_212
timestamp 1698431365
transform 1 0 25088 0 -1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_244
timestamp 1698431365
transform 1 0 28672 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_246
timestamp 1698431365
transform 1 0 28896 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_253
timestamp 1698431365
transform 1 0 29680 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_261
timestamp 1698431365
transform 1 0 30576 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_278
timestamp 1698431365
transform 1 0 32480 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_282
timestamp 1698431365
transform 1 0 32928 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_298
timestamp 1698431365
transform 1 0 34720 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_302
timestamp 1698431365
transform 1 0 35168 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_309
timestamp 1698431365
transform 1 0 35952 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_313
timestamp 1698431365
transform 1 0 36400 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_327
timestamp 1698431365
transform 1 0 37968 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_335
timestamp 1698431365
transform 1 0 38864 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_339
timestamp 1698431365
transform 1 0 39312 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_342
timestamp 1698431365
transform 1 0 39648 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_346
timestamp 1698431365
transform 1 0 40096 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_352
timestamp 1698431365
transform 1 0 40768 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_391
timestamp 1698431365
transform 1 0 45136 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_393
timestamp 1698431365
transform 1 0 45360 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_33
timestamp 1698431365
transform 1 0 5040 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_37
timestamp 1698431365
transform 1 0 5488 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_39
timestamp 1698431365
transform 1 0 5712 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_69
timestamp 1698431365
transform 1 0 9072 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_107
timestamp 1698431365
transform 1 0 13328 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_141
timestamp 1698431365
transform 1 0 17136 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_151
timestamp 1698431365
transform 1 0 18256 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_158
timestamp 1698431365
transform 1 0 19040 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_160
timestamp 1698431365
transform 1 0 19264 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_163
timestamp 1698431365
transform 1 0 19600 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_174
timestamp 1698431365
transform 1 0 20832 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_185
timestamp 1698431365
transform 1 0 22064 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_194
timestamp 1698431365
transform 1 0 23072 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_198
timestamp 1698431365
transform 1 0 23520 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_201
timestamp 1698431365
transform 1 0 23856 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_205
timestamp 1698431365
transform 1 0 24304 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_44_209
timestamp 1698431365
transform 1 0 24752 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_225
timestamp 1698431365
transform 1 0 26544 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_229
timestamp 1698431365
transform 1 0 26992 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_237
timestamp 1698431365
transform 1 0 27888 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_247
timestamp 1698431365
transform 1 0 29008 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_277
timestamp 1698431365
transform 1 0 32368 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_281
timestamp 1698431365
transform 1 0 32816 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_289
timestamp 1698431365
transform 1 0 33712 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_293
timestamp 1698431365
transform 1 0 34160 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_302
timestamp 1698431365
transform 1 0 35168 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_306
timestamp 1698431365
transform 1 0 35616 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_308
timestamp 1698431365
transform 1 0 35840 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_317
timestamp 1698431365
transform 1 0 36848 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_333
timestamp 1698431365
transform 1 0 38640 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_366
timestamp 1698431365
transform 1 0 42336 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_387
timestamp 1698431365
transform 1 0 44688 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_52
timestamp 1698431365
transform 1 0 7168 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_61
timestamp 1698431365
transform 1 0 8176 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_63
timestamp 1698431365
transform 1 0 8400 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_66
timestamp 1698431365
transform 1 0 8736 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_72
timestamp 1698431365
transform 1 0 9408 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_76
timestamp 1698431365
transform 1 0 9856 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_79
timestamp 1698431365
transform 1 0 10192 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_83
timestamp 1698431365
transform 1 0 10640 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_87
timestamp 1698431365
transform 1 0 11088 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_114
timestamp 1698431365
transform 1 0 14112 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_116
timestamp 1698431365
transform 1 0 14336 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_129
timestamp 1698431365
transform 1 0 15792 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_133
timestamp 1698431365
transform 1 0 16240 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_137
timestamp 1698431365
transform 1 0 16688 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_142
timestamp 1698431365
transform 1 0 17248 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_173
timestamp 1698431365
transform 1 0 20720 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_175
timestamp 1698431365
transform 1 0 20944 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_186
timestamp 1698431365
transform 1 0 22176 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_188
timestamp 1698431365
transform 1 0 22400 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_201
timestamp 1698431365
transform 1 0 23856 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_205
timestamp 1698431365
transform 1 0 24304 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_209
timestamp 1698431365
transform 1 0 24752 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_218
timestamp 1698431365
transform 1 0 25760 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_270
timestamp 1698431365
transform 1 0 31584 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_274
timestamp 1698431365
transform 1 0 32032 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_278
timestamp 1698431365
transform 1 0 32480 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_288
timestamp 1698431365
transform 1 0 33600 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_305
timestamp 1698431365
transform 1 0 35504 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_358
timestamp 1698431365
transform 1 0 41440 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_362
timestamp 1698431365
transform 1 0 41888 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_395
timestamp 1698431365
transform 1 0 45584 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_418
timestamp 1698431365
transform 1 0 48160 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_29
timestamp 1698431365
transform 1 0 4592 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_33
timestamp 1698431365
transform 1 0 5040 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_37
timestamp 1698431365
transform 1 0 5488 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_39
timestamp 1698431365
transform 1 0 5712 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_46
timestamp 1698431365
transform 1 0 6496 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_48
timestamp 1698431365
transform 1 0 6720 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_100
timestamp 1698431365
transform 1 0 12544 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_102
timestamp 1698431365
transform 1 0 12768 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_121
timestamp 1698431365
transform 1 0 14896 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_125
timestamp 1698431365
transform 1 0 15344 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_143
timestamp 1698431365
transform 1 0 17360 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_147
timestamp 1698431365
transform 1 0 17808 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_172
timestamp 1698431365
transform 1 0 20608 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_174
timestamp 1698431365
transform 1 0 20832 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_177
timestamp 1698431365
transform 1 0 21168 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_181
timestamp 1698431365
transform 1 0 21616 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_183
timestamp 1698431365
transform 1 0 21840 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_229
timestamp 1698431365
transform 1 0 26992 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_233
timestamp 1698431365
transform 1 0 27440 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_241
timestamp 1698431365
transform 1 0 28336 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_247
timestamp 1698431365
transform 1 0 29008 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_46_251
timestamp 1698431365
transform 1 0 29456 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_267
timestamp 1698431365
transform 1 0 31248 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_269
timestamp 1698431365
transform 1 0 31472 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_307
timestamp 1698431365
transform 1 0 35728 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_311
timestamp 1698431365
transform 1 0 36176 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_317
timestamp 1698431365
transform 1 0 36848 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_365
timestamp 1698431365
transform 1 0 42224 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_369
timestamp 1698431365
transform 1 0 42672 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_387
timestamp 1698431365
transform 1 0 44688 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_37
timestamp 1698431365
transform 1 0 5488 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_39
timestamp 1698431365
transform 1 0 5712 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_68
timestamp 1698431365
transform 1 0 8960 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_128
timestamp 1698431365
transform 1 0 15680 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_142
timestamp 1698431365
transform 1 0 17248 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_146
timestamp 1698431365
transform 1 0 17696 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_162
timestamp 1698431365
transform 1 0 19488 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_177
timestamp 1698431365
transform 1 0 21168 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_185
timestamp 1698431365
transform 1 0 22064 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_200
timestamp 1698431365
transform 1 0 23744 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_208
timestamp 1698431365
transform 1 0 24640 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_212
timestamp 1698431365
transform 1 0 25088 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_216
timestamp 1698431365
transform 1 0 25536 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_232
timestamp 1698431365
transform 1 0 27328 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_236
timestamp 1698431365
transform 1 0 27776 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_253
timestamp 1698431365
transform 1 0 29680 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_257
timestamp 1698431365
transform 1 0 30128 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_261
timestamp 1698431365
transform 1 0 30576 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_277
timestamp 1698431365
transform 1 0 32368 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_279
timestamp 1698431365
transform 1 0 32592 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_298
timestamp 1698431365
transform 1 0 34720 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_308
timestamp 1698431365
transform 1 0 35840 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_343
timestamp 1698431365
transform 1 0 39760 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_347
timestamp 1698431365
transform 1 0 40208 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_349
timestamp 1698431365
transform 1 0 40432 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_382
timestamp 1698431365
transform 1 0 44128 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_2
timestamp 1698431365
transform 1 0 1568 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_107
timestamp 1698431365
transform 1 0 13328 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_126
timestamp 1698431365
transform 1 0 15456 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_145
timestamp 1698431365
transform 1 0 17584 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_149
timestamp 1698431365
transform 1 0 18032 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_158
timestamp 1698431365
transform 1 0 19040 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_160
timestamp 1698431365
transform 1 0 19264 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_172
timestamp 1698431365
transform 1 0 20608 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_174
timestamp 1698431365
transform 1 0 20832 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_185
timestamp 1698431365
transform 1 0 22064 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_48_195
timestamp 1698431365
transform 1 0 23184 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_205
timestamp 1698431365
transform 1 0 24304 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_209
timestamp 1698431365
transform 1 0 24752 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_212
timestamp 1698431365
transform 1 0 25088 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_247
timestamp 1698431365
transform 1 0 29008 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_278
timestamp 1698431365
transform 1 0 32480 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_282
timestamp 1698431365
transform 1 0 32928 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_307
timestamp 1698431365
transform 1 0 35728 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_317
timestamp 1698431365
transform 1 0 36848 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_348
timestamp 1698431365
transform 1 0 40320 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_371
timestamp 1698431365
transform 1 0 42896 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_378
timestamp 1698431365
transform 1 0 43680 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_382
timestamp 1698431365
transform 1 0 44128 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_384
timestamp 1698431365
transform 1 0 44352 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_387
timestamp 1698431365
transform 1 0 44688 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_10
timestamp 1698431365
transform 1 0 2464 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_14
timestamp 1698431365
transform 1 0 2912 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_17
timestamp 1698431365
transform 1 0 3248 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_23
timestamp 1698431365
transform 1 0 3920 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_72
timestamp 1698431365
transform 1 0 9408 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_76
timestamp 1698431365
transform 1 0 9856 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_97
timestamp 1698431365
transform 1 0 12208 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_114
timestamp 1698431365
transform 1 0 14112 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_139
timestamp 1698431365
transform 1 0 16912 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_209
timestamp 1698431365
transform 1 0 24752 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_227
timestamp 1698431365
transform 1 0 26768 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_237
timestamp 1698431365
transform 1 0 27888 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_247
timestamp 1698431365
transform 1 0 29008 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_255
timestamp 1698431365
transform 1 0 29904 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_264
timestamp 1698431365
transform 1 0 30912 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_272
timestamp 1698431365
transform 1 0 31808 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_276
timestamp 1698431365
transform 1 0 32256 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_340
timestamp 1698431365
transform 1 0 39424 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_344
timestamp 1698431365
transform 1 0 39872 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_348
timestamp 1698431365
transform 1 0 40320 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_352
timestamp 1698431365
transform 1 0 40768 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_356
timestamp 1698431365
transform 1 0 41216 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_2
timestamp 1698431365
transform 1 0 1568 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_6
timestamp 1698431365
transform 1 0 2016 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_12
timestamp 1698431365
transform 1 0 2688 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_16
timestamp 1698431365
transform 1 0 3136 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_20
timestamp 1698431365
transform 1 0 3584 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_22
timestamp 1698431365
transform 1 0 3808 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_25
timestamp 1698431365
transform 1 0 4144 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_29
timestamp 1698431365
transform 1 0 4592 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_33
timestamp 1698431365
transform 1 0 5040 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_107
timestamp 1698431365
transform 1 0 13328 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_124
timestamp 1698431365
transform 1 0 15232 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_126
timestamp 1698431365
transform 1 0 15456 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_172
timestamp 1698431365
transform 1 0 20608 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_174
timestamp 1698431365
transform 1 0 20832 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_50_177
timestamp 1698431365
transform 1 0 21168 0 1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_193
timestamp 1698431365
transform 1 0 22960 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_223
timestamp 1698431365
transform 1 0 26320 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_227
timestamp 1698431365
transform 1 0 26768 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_234
timestamp 1698431365
transform 1 0 27552 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_242
timestamp 1698431365
transform 1 0 28448 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_244
timestamp 1698431365
transform 1 0 28672 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_262
timestamp 1698431365
transform 1 0 30688 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_264
timestamp 1698431365
transform 1 0 30912 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_306
timestamp 1698431365
transform 1 0 35616 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_308
timestamp 1698431365
transform 1 0 35840 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_384
timestamp 1698431365
transform 1 0 44352 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_387
timestamp 1698431365
transform 1 0 44688 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_389
timestamp 1698431365
transform 1 0 44912 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_2
timestamp 1698431365
transform 1 0 1568 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_6
timestamp 1698431365
transform 1 0 2016 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_51_10
timestamp 1698431365
transform 1 0 2464 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_18
timestamp 1698431365
transform 1 0 3360 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_22
timestamp 1698431365
transform 1 0 3808 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_25
timestamp 1698431365
transform 1 0 4144 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_29
timestamp 1698431365
transform 1 0 4592 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_33
timestamp 1698431365
transform 1 0 5040 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_37
timestamp 1698431365
transform 1 0 5488 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_96
timestamp 1698431365
transform 1 0 12096 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_137
timestamp 1698431365
transform 1 0 16688 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_139
timestamp 1698431365
transform 1 0 16912 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_142
timestamp 1698431365
transform 1 0 17248 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_146
timestamp 1698431365
transform 1 0 17696 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_161
timestamp 1698431365
transform 1 0 19376 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_163
timestamp 1698431365
transform 1 0 19600 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_166
timestamp 1698431365
transform 1 0 19936 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_170
timestamp 1698431365
transform 1 0 20384 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_174
timestamp 1698431365
transform 1 0 20832 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_212
timestamp 1698431365
transform 1 0 25088 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_216
timestamp 1698431365
transform 1 0 25536 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_246
timestamp 1698431365
transform 1 0 28896 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_250
timestamp 1698431365
transform 1 0 29344 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_349
timestamp 1698431365
transform 1 0 40432 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_358
timestamp 1698431365
transform 1 0 41440 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_389
timestamp 1698431365
transform 1 0 44912 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_52_2
timestamp 1698431365
transform 1 0 1568 0 1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_52_18
timestamp 1698431365
transform 1 0 3360 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_26
timestamp 1698431365
transform 1 0 4256 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_30
timestamp 1698431365
transform 1 0 4704 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_33
timestamp 1698431365
transform 1 0 5040 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_37
timestamp 1698431365
transform 1 0 5488 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_41
timestamp 1698431365
transform 1 0 5936 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_43
timestamp 1698431365
transform 1 0 6160 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_46
timestamp 1698431365
transform 1 0 6496 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_50
timestamp 1698431365
transform 1 0 6944 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_59
timestamp 1698431365
transform 1 0 7952 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_107
timestamp 1698431365
transform 1 0 13328 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_111
timestamp 1698431365
transform 1 0 13776 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_113
timestamp 1698431365
transform 1 0 14000 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_121
timestamp 1698431365
transform 1 0 14896 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_127
timestamp 1698431365
transform 1 0 15568 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_131
timestamp 1698431365
transform 1 0 16016 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_137
timestamp 1698431365
transform 1 0 16688 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_141
timestamp 1698431365
transform 1 0 17136 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_174
timestamp 1698431365
transform 1 0 20832 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_177
timestamp 1698431365
transform 1 0 21168 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_222
timestamp 1698431365
transform 1 0 26208 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_226
timestamp 1698431365
transform 1 0 26656 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_247
timestamp 1698431365
transform 1 0 29008 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_251
timestamp 1698431365
transform 1 0 29456 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_312
timestamp 1698431365
transform 1 0 36288 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_314
timestamp 1698431365
transform 1 0 36512 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_317
timestamp 1698431365
transform 1 0 36848 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_321
timestamp 1698431365
transform 1 0 37296 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_323
timestamp 1698431365
transform 1 0 37520 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_402
timestamp 1698431365
transform 1 0 46368 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_419
timestamp 1698431365
transform 1 0 48272 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_53_2
timestamp 1698431365
transform 1 0 1568 0 -1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_53_34
timestamp 1698431365
transform 1 0 5152 0 -1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_50
timestamp 1698431365
transform 1 0 6944 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_56
timestamp 1698431365
transform 1 0 7616 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_58
timestamp 1698431365
transform 1 0 7840 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_61
timestamp 1698431365
transform 1 0 8176 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_65
timestamp 1698431365
transform 1 0 8624 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_67
timestamp 1698431365
transform 1 0 8848 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_72
timestamp 1698431365
transform 1 0 9408 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_76
timestamp 1698431365
transform 1 0 9856 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_142
timestamp 1698431365
transform 1 0 17248 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_209
timestamp 1698431365
transform 1 0 24752 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_262
timestamp 1698431365
transform 1 0 30688 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_264
timestamp 1698431365
transform 1 0 30912 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_282
timestamp 1698431365
transform 1 0 32928 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_286
timestamp 1698431365
transform 1 0 33376 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_288
timestamp 1698431365
transform 1 0 33600 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_347
timestamp 1698431365
transform 1 0 40208 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_349
timestamp 1698431365
transform 1 0 40432 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_352
timestamp 1698431365
transform 1 0 40768 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_356
timestamp 1698431365
transform 1 0 41216 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_415
timestamp 1698431365
transform 1 0 47824 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_54_6
timestamp 1698431365
transform 1 0 2016 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_22
timestamp 1698431365
transform 1 0 3808 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_30
timestamp 1698431365
transform 1 0 4704 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_54_36
timestamp 1698431365
transform 1 0 5376 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_52
timestamp 1698431365
transform 1 0 7168 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_56
timestamp 1698431365
transform 1 0 7616 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_58
timestamp 1698431365
transform 1 0 7840 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_61
timestamp 1698431365
transform 1 0 8176 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_65
timestamp 1698431365
transform 1 0 8624 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_67
timestamp 1698431365
transform 1 0 8848 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_70
timestamp 1698431365
transform 1 0 9184 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_74
timestamp 1698431365
transform 1 0 9632 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_84
timestamp 1698431365
transform 1 0 10752 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_88
timestamp 1698431365
transform 1 0 11200 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_90
timestamp 1698431365
transform 1 0 11424 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_93
timestamp 1698431365
transform 1 0 11760 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_97
timestamp 1698431365
transform 1 0 12208 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_101
timestamp 1698431365
transform 1 0 12656 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_104
timestamp 1698431365
transform 1 0 12992 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_106
timestamp 1698431365
transform 1 0 13216 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_115
timestamp 1698431365
transform 1 0 14224 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_119
timestamp 1698431365
transform 1 0 14672 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_127
timestamp 1698431365
transform 1 0 15568 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_131
timestamp 1698431365
transform 1 0 16016 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_135
timestamp 1698431365
transform 1 0 16464 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_138
timestamp 1698431365
transform 1 0 16800 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_142
timestamp 1698431365
transform 1 0 17248 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_144
timestamp 1698431365
transform 1 0 17472 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_147
timestamp 1698431365
transform 1 0 17808 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_157
timestamp 1698431365
transform 1 0 18928 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_159
timestamp 1698431365
transform 1 0 19152 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_172
timestamp 1698431365
transform 1 0 20608 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_176
timestamp 1698431365
transform 1 0 21056 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_402
timestamp 1698431365
transform 1 0 46368 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_410
timestamp 1698431365
transform 1 0 47264 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold1 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 39648 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  hold2
timestamp 1698431365
transform -1 0 27888 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input1
timestamp 1698431365
transform 1 0 1568 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input2
timestamp 1698431365
transform -1 0 14224 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input3
timestamp 1698431365
transform 1 0 1568 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input4
timestamp 1698431365
transform 1 0 1568 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input5
timestamp 1698431365
transform 1 0 1568 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input6
timestamp 1698431365
transform 1 0 1568 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input7
timestamp 1698431365
transform 1 0 1568 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input8
timestamp 1698431365
transform 1 0 2464 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input9
timestamp 1698431365
transform -1 0 5040 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input10
timestamp 1698431365
transform 1 0 1568 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input11
timestamp 1698431365
transform 1 0 2240 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input12
timestamp 1698431365
transform 1 0 1568 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input13
timestamp 1698431365
transform 1 0 1568 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input14
timestamp 1698431365
transform 1 0 2464 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input15
timestamp 1698431365
transform 1 0 1568 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input16
timestamp 1698431365
transform 1 0 1568 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input17
timestamp 1698431365
transform 1 0 2912 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input18
timestamp 1698431365
transform 1 0 1568 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input19
timestamp 1698431365
transform 1 0 3136 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input20
timestamp 1698431365
transform -1 0 24752 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input21
timestamp 1698431365
transform 1 0 18256 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input22
timestamp 1698431365
transform -1 0 20384 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input23
timestamp 1698431365
transform 1 0 1568 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input24
timestamp 1698431365
transform -1 0 15568 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input25
timestamp 1698431365
transform -1 0 36512 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input26
timestamp 1698431365
transform -1 0 48160 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input27
timestamp 1698431365
transform 1 0 47712 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input28
timestamp 1698431365
transform -1 0 9856 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input29
timestamp 1698431365
transform -1 0 13104 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input30
timestamp 1698431365
transform -1 0 12880 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input31
timestamp 1698431365
transform -1 0 13664 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input32
timestamp 1698431365
transform -1 0 23632 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input33
timestamp 1698431365
transform -1 0 7504 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input34
timestamp 1698431365
transform -1 0 8176 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input35
timestamp 1698431365
transform 1 0 16800 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input36
timestamp 1698431365
transform 1 0 24416 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input37
timestamp 1698431365
transform 1 0 23632 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input38
timestamp 1698431365
transform 1 0 32032 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input39
timestamp 1698431365
transform 1 0 36848 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input40
timestamp 1698431365
transform -1 0 35168 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input41
timestamp 1698431365
transform -1 0 47936 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input42
timestamp 1698431365
transform -1 0 47040 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input43
timestamp 1698431365
transform 1 0 31024 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input44
timestamp 1698431365
transform -1 0 48272 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input45
timestamp 1698431365
transform 1 0 8288 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input46
timestamp 1698431365
transform 1 0 22960 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input47
timestamp 1698431365
transform -1 0 45472 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input48
timestamp 1698431365
transform -1 0 42560 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input49
timestamp 1698431365
transform -1 0 48384 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input50
timestamp 1698431365
transform -1 0 47712 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input51
timestamp 1698431365
transform -1 0 19936 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input52
timestamp 1698431365
transform 1 0 2240 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output53 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 45472 0 -1 26656
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output54
timestamp 1698431365
transform 1 0 45472 0 -1 7840
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output55
timestamp 1698431365
transform -1 0 48384 0 1 9408
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output56
timestamp 1698431365
transform 1 0 9856 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output57
timestamp 1698431365
transform -1 0 17024 0 -1 6272
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output58
timestamp 1698431365
transform 1 0 13552 0 1 6272
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output59
timestamp 1698431365
transform 1 0 13664 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output60
timestamp 1698431365
transform 1 0 45472 0 1 23520
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output61
timestamp 1698431365
transform -1 0 4480 0 1 17248
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output62
timestamp 1698431365
transform 1 0 9520 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output63
timestamp 1698431365
transform 1 0 17472 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output64
timestamp 1698431365
transform 1 0 45472 0 1 20384
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output65
timestamp 1698431365
transform 1 0 25088 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output66
timestamp 1698431365
transform 1 0 45472 0 1 18816
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output67
timestamp 1698431365
transform -1 0 39424 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output68
timestamp 1698431365
transform 1 0 40768 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output69
timestamp 1698431365
transform 1 0 43680 0 -1 6272
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output70
timestamp 1698431365
transform 1 0 44688 0 1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output71
timestamp 1698431365
transform 1 0 40432 0 1 6272
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output72
timestamp 1698431365
transform 1 0 40768 0 -1 6272
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output73
timestamp 1698431365
transform 1 0 45472 0 1 7840
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output74
timestamp 1698431365
transform 1 0 45472 0 -1 9408
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output75
timestamp 1698431365
transform 1 0 43456 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output76
timestamp 1698431365
transform 1 0 39648 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output77
timestamp 1698431365
transform 1 0 32704 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output78
timestamp 1698431365
transform 1 0 20944 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output79
timestamp 1698431365
transform 1 0 28224 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output80
timestamp 1698431365
transform 1 0 29792 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output81
timestamp 1698431365
transform 1 0 21952 0 -1 43904
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output82
timestamp 1698431365
transform 1 0 43456 0 1 45472
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output83
timestamp 1698431365
transform -1 0 42672 0 1 42336
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output84
timestamp 1698431365
transform 1 0 45472 0 1 40768
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output85
timestamp 1698431365
transform 1 0 45472 0 -1 40768
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output86
timestamp 1698431365
transform 1 0 39648 0 1 45472
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output87
timestamp 1698431365
transform 1 0 40880 0 1 43904
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output88
timestamp 1698431365
transform 1 0 35840 0 -1 43904
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output89
timestamp 1698431365
transform -1 0 39760 0 1 42336
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output90
timestamp 1698431365
transform 1 0 45472 0 -1 43904
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output91
timestamp 1698431365
transform 1 0 44912 0 -1 45472
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output92
timestamp 1698431365
transform 1 0 28224 0 1 45472
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output93
timestamp 1698431365
transform -1 0 48384 0 1 42336
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output94
timestamp 1698431365
transform -1 0 44800 0 -1 36064
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output95
timestamp 1698431365
transform 1 0 32032 0 1 45472
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output96
timestamp 1698431365
transform 1 0 33376 0 1 43904
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output97
timestamp 1698431365
transform 1 0 35840 0 1 45472
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output98
timestamp 1698431365
transform 1 0 32928 0 -1 43904
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output99
timestamp 1698431365
transform 1 0 45472 0 1 36064
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output100
timestamp 1698431365
transform 1 0 41552 0 1 32928
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output101
timestamp 1698431365
transform 1 0 45472 0 1 34496
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output102
timestamp 1698431365
transform 1 0 45472 0 -1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output103
timestamp 1698431365
transform 1 0 45472 0 -1 32928
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output104
timestamp 1698431365
transform 1 0 31024 0 1 42336
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output105
timestamp 1698431365
transform 1 0 42560 0 -1 32928
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output106
timestamp 1698431365
transform 1 0 45472 0 1 31360
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output107
timestamp 1698431365
transform -1 0 48384 0 -1 25088
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output108
timestamp 1698431365
transform -1 0 48384 0 -1 34496
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output109
timestamp 1698431365
transform 1 0 45472 0 1 28224
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output110
timestamp 1698431365
transform 1 0 45472 0 -1 29792
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output111
timestamp 1698431365
transform -1 0 24192 0 1 45472
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output112
timestamp 1698431365
transform 1 0 25088 0 1 45472
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output113
timestamp 1698431365
transform -1 0 4480 0 1 29792
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_55 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698431365
transform -1 0 48608 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_56
timestamp 1698431365
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698431365
transform -1 0 48608 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_57
timestamp 1698431365
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698431365
transform -1 0 48608 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_58
timestamp 1698431365
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698431365
transform -1 0 48608 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_59
timestamp 1698431365
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698431365
transform -1 0 48608 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_60
timestamp 1698431365
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698431365
transform -1 0 48608 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_61
timestamp 1698431365
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698431365
transform -1 0 48608 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_62
timestamp 1698431365
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698431365
transform -1 0 48608 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_63
timestamp 1698431365
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698431365
transform -1 0 48608 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_64
timestamp 1698431365
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698431365
transform -1 0 48608 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_65
timestamp 1698431365
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698431365
transform -1 0 48608 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_66
timestamp 1698431365
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698431365
transform -1 0 48608 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_67
timestamp 1698431365
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698431365
transform -1 0 48608 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_68
timestamp 1698431365
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698431365
transform -1 0 48608 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_69
timestamp 1698431365
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698431365
transform -1 0 48608 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_70
timestamp 1698431365
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698431365
transform -1 0 48608 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_71
timestamp 1698431365
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698431365
transform -1 0 48608 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_72
timestamp 1698431365
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698431365
transform -1 0 48608 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_73
timestamp 1698431365
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698431365
transform -1 0 48608 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_74
timestamp 1698431365
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698431365
transform -1 0 48608 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_75
timestamp 1698431365
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698431365
transform -1 0 48608 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_76
timestamp 1698431365
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698431365
transform -1 0 48608 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_77
timestamp 1698431365
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1698431365
transform -1 0 48608 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_78
timestamp 1698431365
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1698431365
transform -1 0 48608 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_79
timestamp 1698431365
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1698431365
transform -1 0 48608 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_80
timestamp 1698431365
transform 1 0 1344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1698431365
transform -1 0 48608 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_81
timestamp 1698431365
transform 1 0 1344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1698431365
transform -1 0 48608 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_82
timestamp 1698431365
transform 1 0 1344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1698431365
transform -1 0 48608 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_83
timestamp 1698431365
transform 1 0 1344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1698431365
transform -1 0 48608 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_84
timestamp 1698431365
transform 1 0 1344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1698431365
transform -1 0 48608 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Left_85
timestamp 1698431365
transform 1 0 1344 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1698431365
transform -1 0 48608 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Left_86
timestamp 1698431365
transform 1 0 1344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1698431365
transform -1 0 48608 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Left_87
timestamp 1698431365
transform 1 0 1344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1698431365
transform -1 0 48608 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Left_88
timestamp 1698431365
transform 1 0 1344 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1698431365
transform -1 0 48608 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Left_89
timestamp 1698431365
transform 1 0 1344 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1698431365
transform -1 0 48608 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Left_90
timestamp 1698431365
transform 1 0 1344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Right_35
timestamp 1698431365
transform -1 0 48608 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Left_91
timestamp 1698431365
transform 1 0 1344 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Right_36
timestamp 1698431365
transform -1 0 48608 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Left_92
timestamp 1698431365
transform 1 0 1344 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Right_37
timestamp 1698431365
transform -1 0 48608 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Left_93
timestamp 1698431365
transform 1 0 1344 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Right_38
timestamp 1698431365
transform -1 0 48608 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Left_94
timestamp 1698431365
transform 1 0 1344 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Right_39
timestamp 1698431365
transform -1 0 48608 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Left_95
timestamp 1698431365
transform 1 0 1344 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Right_40
timestamp 1698431365
transform -1 0 48608 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Left_96
timestamp 1698431365
transform 1 0 1344 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Right_41
timestamp 1698431365
transform -1 0 48608 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Left_97
timestamp 1698431365
transform 1 0 1344 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Right_42
timestamp 1698431365
transform -1 0 48608 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Left_98
timestamp 1698431365
transform 1 0 1344 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Right_43
timestamp 1698431365
transform -1 0 48608 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Left_99
timestamp 1698431365
transform 1 0 1344 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Right_44
timestamp 1698431365
transform -1 0 48608 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_45_Left_100
timestamp 1698431365
transform 1 0 1344 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_45_Right_45
timestamp 1698431365
transform -1 0 48608 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_46_Left_101
timestamp 1698431365
transform 1 0 1344 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_46_Right_46
timestamp 1698431365
transform -1 0 48608 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_47_Left_102
timestamp 1698431365
transform 1 0 1344 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_47_Right_47
timestamp 1698431365
transform -1 0 48608 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_48_Left_103
timestamp 1698431365
transform 1 0 1344 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_48_Right_48
timestamp 1698431365
transform -1 0 48608 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_49_Left_104
timestamp 1698431365
transform 1 0 1344 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_49_Right_49
timestamp 1698431365
transform -1 0 48608 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_50_Left_105
timestamp 1698431365
transform 1 0 1344 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_50_Right_50
timestamp 1698431365
transform -1 0 48608 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_51_Left_106
timestamp 1698431365
transform 1 0 1344 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_51_Right_51
timestamp 1698431365
transform -1 0 48608 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_52_Left_107
timestamp 1698431365
transform 1 0 1344 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_52_Right_52
timestamp 1698431365
transform -1 0 48608 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_53_Left_108
timestamp 1698431365
transform 1 0 1344 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_53_Right_53
timestamp 1698431365
transform -1 0 48608 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_54_Left_109
timestamp 1698431365
transform 1 0 1344 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_54_Right_54
timestamp 1698431365
transform -1 0 48608 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  spimemio_114 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 47936 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  spimemio_115
timestamp 1698431365
transform -1 0 2016 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  spimemio_116
timestamp 1698431365
transform -1 0 2016 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  spimemio_117
timestamp 1698431365
transform -1 0 2464 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  spimemio_118
timestamp 1698431365
transform 1 0 47488 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  spimemio_119
timestamp 1698431365
transform -1 0 2016 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  spimemio_120
timestamp 1698431365
transform 1 0 44016 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  spimemio_121
timestamp 1698431365
transform 1 0 47936 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  spimemio_122
timestamp 1698431365
transform 1 0 46592 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  spimemio_123
timestamp 1698431365
transform 1 0 47936 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  spimemio_124
timestamp 1698431365
transform 1 0 42224 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  spimemio_125
timestamp 1698431365
transform 1 0 45024 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  spimemio_126
timestamp 1698431365
transform 1 0 47936 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  spimemio_127
timestamp 1698431365
transform -1 0 2016 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  spimemio_128
timestamp 1698431365
transform 1 0 45024 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  spimemio_129
timestamp 1698431365
transform -1 0 2016 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_110 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5152 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_111
timestamp 1698431365
transform 1 0 8960 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_112
timestamp 1698431365
transform 1 0 12768 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_113
timestamp 1698431365
transform 1 0 16576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_114
timestamp 1698431365
transform 1 0 20384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_115
timestamp 1698431365
transform 1 0 24192 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_116
timestamp 1698431365
transform 1 0 28000 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_117
timestamp 1698431365
transform 1 0 31808 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_118
timestamp 1698431365
transform 1 0 35616 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_119
timestamp 1698431365
transform 1 0 39424 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_120
timestamp 1698431365
transform 1 0 43232 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_121
timestamp 1698431365
transform 1 0 47040 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_122
timestamp 1698431365
transform 1 0 9184 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_123
timestamp 1698431365
transform 1 0 17024 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_124
timestamp 1698431365
transform 1 0 24864 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_125
timestamp 1698431365
transform 1 0 32704 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_126
timestamp 1698431365
transform 1 0 40544 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_127
timestamp 1698431365
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_128
timestamp 1698431365
transform 1 0 13104 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_129
timestamp 1698431365
transform 1 0 20944 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_130
timestamp 1698431365
transform 1 0 28784 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_131
timestamp 1698431365
transform 1 0 36624 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_132
timestamp 1698431365
transform 1 0 44464 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_133
timestamp 1698431365
transform 1 0 9184 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_134
timestamp 1698431365
transform 1 0 17024 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_135
timestamp 1698431365
transform 1 0 24864 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_136
timestamp 1698431365
transform 1 0 32704 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_137
timestamp 1698431365
transform 1 0 40544 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_138
timestamp 1698431365
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_139
timestamp 1698431365
transform 1 0 13104 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_140
timestamp 1698431365
transform 1 0 20944 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_141
timestamp 1698431365
transform 1 0 28784 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_142
timestamp 1698431365
transform 1 0 36624 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_143
timestamp 1698431365
transform 1 0 44464 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_144
timestamp 1698431365
transform 1 0 9184 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_145
timestamp 1698431365
transform 1 0 17024 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_146
timestamp 1698431365
transform 1 0 24864 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_147
timestamp 1698431365
transform 1 0 32704 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_148
timestamp 1698431365
transform 1 0 40544 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_149
timestamp 1698431365
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_150
timestamp 1698431365
transform 1 0 13104 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_151
timestamp 1698431365
transform 1 0 20944 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_152
timestamp 1698431365
transform 1 0 28784 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_153
timestamp 1698431365
transform 1 0 36624 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_154
timestamp 1698431365
transform 1 0 44464 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_155
timestamp 1698431365
transform 1 0 9184 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_156
timestamp 1698431365
transform 1 0 17024 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_157
timestamp 1698431365
transform 1 0 24864 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_158
timestamp 1698431365
transform 1 0 32704 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_159
timestamp 1698431365
transform 1 0 40544 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_160
timestamp 1698431365
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_161
timestamp 1698431365
transform 1 0 13104 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_162
timestamp 1698431365
transform 1 0 20944 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_163
timestamp 1698431365
transform 1 0 28784 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_164
timestamp 1698431365
transform 1 0 36624 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_165
timestamp 1698431365
transform 1 0 44464 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_166
timestamp 1698431365
transform 1 0 9184 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_167
timestamp 1698431365
transform 1 0 17024 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_168
timestamp 1698431365
transform 1 0 24864 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_169
timestamp 1698431365
transform 1 0 32704 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_170
timestamp 1698431365
transform 1 0 40544 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_171
timestamp 1698431365
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_172
timestamp 1698431365
transform 1 0 13104 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_173
timestamp 1698431365
transform 1 0 20944 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_174
timestamp 1698431365
transform 1 0 28784 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_175
timestamp 1698431365
transform 1 0 36624 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_176
timestamp 1698431365
transform 1 0 44464 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_177
timestamp 1698431365
transform 1 0 9184 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_178
timestamp 1698431365
transform 1 0 17024 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_179
timestamp 1698431365
transform 1 0 24864 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_180
timestamp 1698431365
transform 1 0 32704 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_181
timestamp 1698431365
transform 1 0 40544 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_182
timestamp 1698431365
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_183
timestamp 1698431365
transform 1 0 13104 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_184
timestamp 1698431365
transform 1 0 20944 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_185
timestamp 1698431365
transform 1 0 28784 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_186
timestamp 1698431365
transform 1 0 36624 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_187
timestamp 1698431365
transform 1 0 44464 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_188
timestamp 1698431365
transform 1 0 9184 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_189
timestamp 1698431365
transform 1 0 17024 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_190
timestamp 1698431365
transform 1 0 24864 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_191
timestamp 1698431365
transform 1 0 32704 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_192
timestamp 1698431365
transform 1 0 40544 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_193
timestamp 1698431365
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_194
timestamp 1698431365
transform 1 0 13104 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_195
timestamp 1698431365
transform 1 0 20944 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_196
timestamp 1698431365
transform 1 0 28784 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_197
timestamp 1698431365
transform 1 0 36624 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_198
timestamp 1698431365
transform 1 0 44464 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_199
timestamp 1698431365
transform 1 0 9184 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_200
timestamp 1698431365
transform 1 0 17024 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_201
timestamp 1698431365
transform 1 0 24864 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_202
timestamp 1698431365
transform 1 0 32704 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_203
timestamp 1698431365
transform 1 0 40544 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_204
timestamp 1698431365
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_205
timestamp 1698431365
transform 1 0 13104 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_206
timestamp 1698431365
transform 1 0 20944 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_207
timestamp 1698431365
transform 1 0 28784 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_208
timestamp 1698431365
transform 1 0 36624 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_209
timestamp 1698431365
transform 1 0 44464 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_210
timestamp 1698431365
transform 1 0 9184 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_211
timestamp 1698431365
transform 1 0 17024 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_212
timestamp 1698431365
transform 1 0 24864 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_213
timestamp 1698431365
transform 1 0 32704 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_214
timestamp 1698431365
transform 1 0 40544 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_215
timestamp 1698431365
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_216
timestamp 1698431365
transform 1 0 13104 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_217
timestamp 1698431365
transform 1 0 20944 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_218
timestamp 1698431365
transform 1 0 28784 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_219
timestamp 1698431365
transform 1 0 36624 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_220
timestamp 1698431365
transform 1 0 44464 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_221
timestamp 1698431365
transform 1 0 9184 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_222
timestamp 1698431365
transform 1 0 17024 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_223
timestamp 1698431365
transform 1 0 24864 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_224
timestamp 1698431365
transform 1 0 32704 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_225
timestamp 1698431365
transform 1 0 40544 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_226
timestamp 1698431365
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_227
timestamp 1698431365
transform 1 0 13104 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_228
timestamp 1698431365
transform 1 0 20944 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_229
timestamp 1698431365
transform 1 0 28784 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_230
timestamp 1698431365
transform 1 0 36624 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_231
timestamp 1698431365
transform 1 0 44464 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_232
timestamp 1698431365
transform 1 0 9184 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_233
timestamp 1698431365
transform 1 0 17024 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_234
timestamp 1698431365
transform 1 0 24864 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_235
timestamp 1698431365
transform 1 0 32704 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_236
timestamp 1698431365
transform 1 0 40544 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_237
timestamp 1698431365
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_238
timestamp 1698431365
transform 1 0 13104 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_239
timestamp 1698431365
transform 1 0 20944 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_240
timestamp 1698431365
transform 1 0 28784 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_241
timestamp 1698431365
transform 1 0 36624 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_242
timestamp 1698431365
transform 1 0 44464 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_243
timestamp 1698431365
transform 1 0 9184 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_244
timestamp 1698431365
transform 1 0 17024 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_245
timestamp 1698431365
transform 1 0 24864 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_246
timestamp 1698431365
transform 1 0 32704 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_247
timestamp 1698431365
transform 1 0 40544 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_248
timestamp 1698431365
transform 1 0 5264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_249
timestamp 1698431365
transform 1 0 13104 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_250
timestamp 1698431365
transform 1 0 20944 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_251
timestamp 1698431365
transform 1 0 28784 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_252
timestamp 1698431365
transform 1 0 36624 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_253
timestamp 1698431365
transform 1 0 44464 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_254
timestamp 1698431365
transform 1 0 9184 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_255
timestamp 1698431365
transform 1 0 17024 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_256
timestamp 1698431365
transform 1 0 24864 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_257
timestamp 1698431365
transform 1 0 32704 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_258
timestamp 1698431365
transform 1 0 40544 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_259
timestamp 1698431365
transform 1 0 5264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_260
timestamp 1698431365
transform 1 0 13104 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_261
timestamp 1698431365
transform 1 0 20944 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_262
timestamp 1698431365
transform 1 0 28784 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_263
timestamp 1698431365
transform 1 0 36624 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_264
timestamp 1698431365
transform 1 0 44464 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_265
timestamp 1698431365
transform 1 0 9184 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_266
timestamp 1698431365
transform 1 0 17024 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_267
timestamp 1698431365
transform 1 0 24864 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_268
timestamp 1698431365
transform 1 0 32704 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_269
timestamp 1698431365
transform 1 0 40544 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_270
timestamp 1698431365
transform 1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_271
timestamp 1698431365
transform 1 0 13104 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_272
timestamp 1698431365
transform 1 0 20944 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_273
timestamp 1698431365
transform 1 0 28784 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_274
timestamp 1698431365
transform 1 0 36624 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_275
timestamp 1698431365
transform 1 0 44464 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_276
timestamp 1698431365
transform 1 0 9184 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_277
timestamp 1698431365
transform 1 0 17024 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_278
timestamp 1698431365
transform 1 0 24864 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_279
timestamp 1698431365
transform 1 0 32704 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_280
timestamp 1698431365
transform 1 0 40544 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_281
timestamp 1698431365
transform 1 0 5264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_282
timestamp 1698431365
transform 1 0 13104 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_283
timestamp 1698431365
transform 1 0 20944 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_284
timestamp 1698431365
transform 1 0 28784 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_285
timestamp 1698431365
transform 1 0 36624 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_286
timestamp 1698431365
transform 1 0 44464 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_287
timestamp 1698431365
transform 1 0 9184 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_288
timestamp 1698431365
transform 1 0 17024 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_289
timestamp 1698431365
transform 1 0 24864 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_290
timestamp 1698431365
transform 1 0 32704 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_291
timestamp 1698431365
transform 1 0 40544 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_292
timestamp 1698431365
transform 1 0 5264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_293
timestamp 1698431365
transform 1 0 13104 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_294
timestamp 1698431365
transform 1 0 20944 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_295
timestamp 1698431365
transform 1 0 28784 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_296
timestamp 1698431365
transform 1 0 36624 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_297
timestamp 1698431365
transform 1 0 44464 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_298
timestamp 1698431365
transform 1 0 9184 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_299
timestamp 1698431365
transform 1 0 17024 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_300
timestamp 1698431365
transform 1 0 24864 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_301
timestamp 1698431365
transform 1 0 32704 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_302
timestamp 1698431365
transform 1 0 40544 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_303
timestamp 1698431365
transform 1 0 5264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_304
timestamp 1698431365
transform 1 0 13104 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_305
timestamp 1698431365
transform 1 0 20944 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_306
timestamp 1698431365
transform 1 0 28784 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_307
timestamp 1698431365
transform 1 0 36624 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_308
timestamp 1698431365
transform 1 0 44464 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_309
timestamp 1698431365
transform 1 0 9184 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_310
timestamp 1698431365
transform 1 0 17024 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_311
timestamp 1698431365
transform 1 0 24864 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_312
timestamp 1698431365
transform 1 0 32704 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_313
timestamp 1698431365
transform 1 0 40544 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_314
timestamp 1698431365
transform 1 0 5264 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_315
timestamp 1698431365
transform 1 0 13104 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_316
timestamp 1698431365
transform 1 0 20944 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_317
timestamp 1698431365
transform 1 0 28784 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_318
timestamp 1698431365
transform 1 0 36624 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_319
timestamp 1698431365
transform 1 0 44464 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_320
timestamp 1698431365
transform 1 0 9184 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_321
timestamp 1698431365
transform 1 0 17024 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_322
timestamp 1698431365
transform 1 0 24864 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_323
timestamp 1698431365
transform 1 0 32704 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_324
timestamp 1698431365
transform 1 0 40544 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_325
timestamp 1698431365
transform 1 0 5264 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_326
timestamp 1698431365
transform 1 0 13104 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_327
timestamp 1698431365
transform 1 0 20944 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_328
timestamp 1698431365
transform 1 0 28784 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_329
timestamp 1698431365
transform 1 0 36624 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_330
timestamp 1698431365
transform 1 0 44464 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_331
timestamp 1698431365
transform 1 0 9184 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_332
timestamp 1698431365
transform 1 0 17024 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_333
timestamp 1698431365
transform 1 0 24864 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_334
timestamp 1698431365
transform 1 0 32704 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_335
timestamp 1698431365
transform 1 0 40544 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_336
timestamp 1698431365
transform 1 0 5264 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_337
timestamp 1698431365
transform 1 0 13104 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_338
timestamp 1698431365
transform 1 0 20944 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_339
timestamp 1698431365
transform 1 0 28784 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_340
timestamp 1698431365
transform 1 0 36624 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_341
timestamp 1698431365
transform 1 0 44464 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_342
timestamp 1698431365
transform 1 0 9184 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_343
timestamp 1698431365
transform 1 0 17024 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_344
timestamp 1698431365
transform 1 0 24864 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_345
timestamp 1698431365
transform 1 0 32704 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_346
timestamp 1698431365
transform 1 0 40544 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_347
timestamp 1698431365
transform 1 0 5264 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_348
timestamp 1698431365
transform 1 0 13104 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_349
timestamp 1698431365
transform 1 0 20944 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_350
timestamp 1698431365
transform 1 0 28784 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_351
timestamp 1698431365
transform 1 0 36624 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_352
timestamp 1698431365
transform 1 0 44464 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_353
timestamp 1698431365
transform 1 0 9184 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_354
timestamp 1698431365
transform 1 0 17024 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_355
timestamp 1698431365
transform 1 0 24864 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_356
timestamp 1698431365
transform 1 0 32704 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_357
timestamp 1698431365
transform 1 0 40544 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_358
timestamp 1698431365
transform 1 0 5264 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_359
timestamp 1698431365
transform 1 0 13104 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_360
timestamp 1698431365
transform 1 0 20944 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_361
timestamp 1698431365
transform 1 0 28784 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_362
timestamp 1698431365
transform 1 0 36624 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_363
timestamp 1698431365
transform 1 0 44464 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_364
timestamp 1698431365
transform 1 0 9184 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_365
timestamp 1698431365
transform 1 0 17024 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_366
timestamp 1698431365
transform 1 0 24864 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_367
timestamp 1698431365
transform 1 0 32704 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_368
timestamp 1698431365
transform 1 0 40544 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_369
timestamp 1698431365
transform 1 0 5264 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_370
timestamp 1698431365
transform 1 0 13104 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_371
timestamp 1698431365
transform 1 0 20944 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_372
timestamp 1698431365
transform 1 0 28784 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_373
timestamp 1698431365
transform 1 0 36624 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_374
timestamp 1698431365
transform 1 0 44464 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_375
timestamp 1698431365
transform 1 0 9184 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_376
timestamp 1698431365
transform 1 0 17024 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_377
timestamp 1698431365
transform 1 0 24864 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_378
timestamp 1698431365
transform 1 0 32704 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_379
timestamp 1698431365
transform 1 0 40544 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_380
timestamp 1698431365
transform 1 0 5264 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_381
timestamp 1698431365
transform 1 0 13104 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_382
timestamp 1698431365
transform 1 0 20944 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_383
timestamp 1698431365
transform 1 0 28784 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_384
timestamp 1698431365
transform 1 0 36624 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_385
timestamp 1698431365
transform 1 0 44464 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_386
timestamp 1698431365
transform 1 0 9184 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_387
timestamp 1698431365
transform 1 0 17024 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_388
timestamp 1698431365
transform 1 0 24864 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_389
timestamp 1698431365
transform 1 0 32704 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_390
timestamp 1698431365
transform 1 0 40544 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_391
timestamp 1698431365
transform 1 0 5264 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_392
timestamp 1698431365
transform 1 0 13104 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_393
timestamp 1698431365
transform 1 0 20944 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_394
timestamp 1698431365
transform 1 0 28784 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_395
timestamp 1698431365
transform 1 0 36624 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_396
timestamp 1698431365
transform 1 0 44464 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_397
timestamp 1698431365
transform 1 0 9184 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_398
timestamp 1698431365
transform 1 0 17024 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_399
timestamp 1698431365
transform 1 0 24864 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_400
timestamp 1698431365
transform 1 0 32704 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_401
timestamp 1698431365
transform 1 0 40544 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_402
timestamp 1698431365
transform 1 0 5264 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_403
timestamp 1698431365
transform 1 0 13104 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_404
timestamp 1698431365
transform 1 0 20944 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_405
timestamp 1698431365
transform 1 0 28784 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_406
timestamp 1698431365
transform 1 0 36624 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_407
timestamp 1698431365
transform 1 0 44464 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_408
timestamp 1698431365
transform 1 0 9184 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_409
timestamp 1698431365
transform 1 0 17024 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_410
timestamp 1698431365
transform 1 0 24864 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_411
timestamp 1698431365
transform 1 0 32704 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_412
timestamp 1698431365
transform 1 0 40544 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_413
timestamp 1698431365
transform 1 0 5152 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_414
timestamp 1698431365
transform 1 0 8960 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_415
timestamp 1698431365
transform 1 0 12768 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_416
timestamp 1698431365
transform 1 0 16576 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_417
timestamp 1698431365
transform 1 0 20384 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_418
timestamp 1698431365
transform 1 0 24192 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_419
timestamp 1698431365
transform 1 0 28000 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_420
timestamp 1698431365
transform 1 0 31808 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_421
timestamp 1698431365
transform 1 0 35616 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_422
timestamp 1698431365
transform 1 0 39424 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_423
timestamp 1698431365
transform 1 0 43232 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_424
timestamp 1698431365
transform 1 0 47040 0 1 45472
box -86 -86 310 870
<< labels >>
flabel metal3 s 0 25536 800 25648 0 FreeSans 448 0 0 0 addr[0]
port 0 nsew signal input
flabel metal2 s 13440 49200 13552 50000 0 FreeSans 448 90 0 0 addr[10]
port 1 nsew signal input
flabel metal3 s 0 40320 800 40432 0 FreeSans 448 0 0 0 addr[11]
port 2 nsew signal input
flabel metal3 s 0 35616 800 35728 0 FreeSans 448 0 0 0 addr[12]
port 3 nsew signal input
flabel metal3 s 0 32256 800 32368 0 FreeSans 448 0 0 0 addr[13]
port 4 nsew signal input
flabel metal3 s 0 30912 800 31024 0 FreeSans 448 0 0 0 addr[14]
port 5 nsew signal input
flabel metal3 s 0 38304 800 38416 0 FreeSans 448 0 0 0 addr[15]
port 6 nsew signal input
flabel metal3 s 0 39648 800 39760 0 FreeSans 448 0 0 0 addr[16]
port 7 nsew signal input
flabel metal3 s 0 32928 800 33040 0 FreeSans 448 0 0 0 addr[17]
port 8 nsew signal input
flabel metal3 s 0 34944 800 35056 0 FreeSans 448 0 0 0 addr[18]
port 9 nsew signal input
flabel metal3 s 0 24864 800 24976 0 FreeSans 448 0 0 0 addr[19]
port 10 nsew signal input
flabel metal3 s 0 23520 800 23632 0 FreeSans 448 0 0 0 addr[1]
port 11 nsew signal input
flabel metal3 s 0 28224 800 28336 0 FreeSans 448 0 0 0 addr[20]
port 12 nsew signal input
flabel metal3 s 0 33600 800 33712 0 FreeSans 448 0 0 0 addr[21]
port 13 nsew signal input
flabel metal3 s 0 31584 800 31696 0 FreeSans 448 0 0 0 addr[22]
port 14 nsew signal input
flabel metal3 s 0 30240 800 30352 0 FreeSans 448 0 0 0 addr[23]
port 15 nsew signal input
flabel metal3 s 0 28896 800 29008 0 FreeSans 448 0 0 0 addr[2]
port 16 nsew signal input
flabel metal3 s 0 26208 800 26320 0 FreeSans 448 0 0 0 addr[3]
port 17 nsew signal input
flabel metal3 s 0 27552 800 27664 0 FreeSans 448 0 0 0 addr[4]
port 18 nsew signal input
flabel metal2 s 22848 49200 22960 50000 0 FreeSans 448 90 0 0 addr[5]
port 19 nsew signal input
flabel metal2 s 18144 49200 18256 50000 0 FreeSans 448 90 0 0 addr[6]
port 20 nsew signal input
flabel metal2 s 20160 49200 20272 50000 0 FreeSans 448 90 0 0 addr[7]
port 21 nsew signal input
flabel metal3 s 0 37632 800 37744 0 FreeSans 448 0 0 0 addr[8]
port 22 nsew signal input
flabel metal2 s 14784 49200 14896 50000 0 FreeSans 448 90 0 0 addr[9]
port 23 nsew signal input
flabel metal2 s 33600 0 33712 800 0 FreeSans 448 90 0 0 cfgreg_di[0]
port 24 nsew signal input
flabel metal2 s 43680 0 43792 800 0 FreeSans 448 90 0 0 cfgreg_di[10]
port 25 nsew signal input
flabel metal2 s 45024 0 45136 800 0 FreeSans 448 90 0 0 cfgreg_di[11]
port 26 nsew signal input
flabel metal2 s 3360 0 3472 800 0 FreeSans 448 90 0 0 cfgreg_di[12]
port 27 nsew signal input
flabel metal2 s 2016 0 2128 800 0 FreeSans 448 90 0 0 cfgreg_di[13]
port 28 nsew signal input
flabel metal2 s 2688 0 2800 800 0 FreeSans 448 90 0 0 cfgreg_di[14]
port 29 nsew signal input
flabel metal2 s 20160 0 20272 800 0 FreeSans 448 90 0 0 cfgreg_di[15]
port 30 nsew signal input
flabel metal2 s 10752 0 10864 800 0 FreeSans 448 90 0 0 cfgreg_di[16]
port 31 nsew signal input
flabel metal2 s 12768 0 12880 800 0 FreeSans 448 90 0 0 cfgreg_di[17]
port 32 nsew signal input
flabel metal2 s 12096 0 12208 800 0 FreeSans 448 90 0 0 cfgreg_di[18]
port 33 nsew signal input
flabel metal2 s 14112 0 14224 800 0 FreeSans 448 90 0 0 cfgreg_di[19]
port 34 nsew signal input
flabel metal2 s 22176 0 22288 800 0 FreeSans 448 90 0 0 cfgreg_di[1]
port 35 nsew signal input
flabel metal2 s 6720 0 6832 800 0 FreeSans 448 90 0 0 cfgreg_di[20]
port 36 nsew signal input
flabel metal2 s 7392 0 7504 800 0 FreeSans 448 90 0 0 cfgreg_di[21]
port 37 nsew signal input
flabel metal2 s 16800 0 16912 800 0 FreeSans 448 90 0 0 cfgreg_di[22]
port 38 nsew signal input
flabel metal2 s 4032 0 4144 800 0 FreeSans 448 90 0 0 cfgreg_di[23]
port 39 nsew signal input
flabel metal2 s 4704 0 4816 800 0 FreeSans 448 90 0 0 cfgreg_di[24]
port 40 nsew signal input
flabel metal2 s 5376 0 5488 800 0 FreeSans 448 90 0 0 cfgreg_di[25]
port 41 nsew signal input
flabel metal2 s 6048 0 6160 800 0 FreeSans 448 90 0 0 cfgreg_di[26]
port 42 nsew signal input
flabel metal2 s 18144 0 18256 800 0 FreeSans 448 90 0 0 cfgreg_di[27]
port 43 nsew signal input
flabel metal2 s 8064 0 8176 800 0 FreeSans 448 90 0 0 cfgreg_di[28]
port 44 nsew signal input
flabel metal2 s 672 0 784 800 0 FreeSans 448 90 0 0 cfgreg_di[29]
port 45 nsew signal input
flabel metal2 s 24864 0 24976 800 0 FreeSans 448 90 0 0 cfgreg_di[2]
port 46 nsew signal input
flabel metal2 s 19488 0 19600 800 0 FreeSans 448 90 0 0 cfgreg_di[30]
port 47 nsew signal input
flabel metal2 s 23520 0 23632 800 0 FreeSans 448 90 0 0 cfgreg_di[31]
port 48 nsew signal input
flabel metal2 s 30240 0 30352 800 0 FreeSans 448 90 0 0 cfgreg_di[3]
port 49 nsew signal input
flabel metal2 s 35616 0 35728 800 0 FreeSans 448 90 0 0 cfgreg_di[4]
port 50 nsew signal input
flabel metal2 s 31584 0 31696 800 0 FreeSans 448 90 0 0 cfgreg_di[5]
port 51 nsew signal input
flabel metal2 s 8736 0 8848 800 0 FreeSans 448 90 0 0 cfgreg_di[6]
port 52 nsew signal input
flabel metal2 s 1344 0 1456 800 0 FreeSans 448 90 0 0 cfgreg_di[7]
port 53 nsew signal input
flabel metal2 s 43008 0 43120 800 0 FreeSans 448 90 0 0 cfgreg_di[8]
port 54 nsew signal input
flabel metal2 s 42336 0 42448 800 0 FreeSans 448 90 0 0 cfgreg_di[9]
port 55 nsew signal input
flabel metal3 s 49200 25536 50000 25648 0 FreeSans 448 0 0 0 cfgreg_do[0]
port 56 nsew signal tristate
flabel metal3 s 49200 7392 50000 7504 0 FreeSans 448 0 0 0 cfgreg_do[10]
port 57 nsew signal tristate
flabel metal3 s 49200 9408 50000 9520 0 FreeSans 448 0 0 0 cfgreg_do[11]
port 58 nsew signal tristate
flabel metal3 s 0 5376 800 5488 0 FreeSans 448 0 0 0 cfgreg_do[12]
port 59 nsew signal tristate
flabel metal3 s 0 2688 800 2800 0 FreeSans 448 0 0 0 cfgreg_do[13]
port 60 nsew signal tristate
flabel metal3 s 49200 44352 50000 44464 0 FreeSans 448 0 0 0 cfgreg_do[14]
port 61 nsew signal tristate
flabel metal3 s 0 4032 800 4144 0 FreeSans 448 0 0 0 cfgreg_do[15]
port 62 nsew signal tristate
flabel metal2 s 11424 0 11536 800 0 FreeSans 448 90 0 0 cfgreg_do[16]
port 63 nsew signal tristate
flabel metal2 s 14784 0 14896 800 0 FreeSans 448 90 0 0 cfgreg_do[17]
port 64 nsew signal tristate
flabel metal2 s 13440 0 13552 800 0 FreeSans 448 90 0 0 cfgreg_do[18]
port 65 nsew signal tristate
flabel metal2 s 16128 0 16240 800 0 FreeSans 448 90 0 0 cfgreg_do[19]
port 66 nsew signal tristate
flabel metal3 s 49200 23520 50000 23632 0 FreeSans 448 0 0 0 cfgreg_do[1]
port 67 nsew signal tristate
flabel metal3 s 0 17472 800 17584 0 FreeSans 448 0 0 0 cfgreg_do[20]
port 68 nsew signal tristate
flabel metal2 s 9408 0 9520 800 0 FreeSans 448 90 0 0 cfgreg_do[21]
port 69 nsew signal tristate
flabel metal2 s 17472 0 17584 800 0 FreeSans 448 90 0 0 cfgreg_do[22]
port 70 nsew signal tristate
flabel metal3 s 49200 4704 50000 4816 0 FreeSans 448 0 0 0 cfgreg_do[23]
port 71 nsew signal tristate
flabel metal3 s 49200 43680 50000 43792 0 FreeSans 448 0 0 0 cfgreg_do[24]
port 72 nsew signal tristate
flabel metal3 s 49200 45024 50000 45136 0 FreeSans 448 0 0 0 cfgreg_do[25]
port 73 nsew signal tristate
flabel metal3 s 49200 4032 50000 4144 0 FreeSans 448 0 0 0 cfgreg_do[26]
port 74 nsew signal tristate
flabel metal3 s 49200 3360 50000 3472 0 FreeSans 448 0 0 0 cfgreg_do[27]
port 75 nsew signal tristate
flabel metal3 s 49200 46368 50000 46480 0 FreeSans 448 0 0 0 cfgreg_do[28]
port 76 nsew signal tristate
flabel metal3 s 49200 43008 50000 43120 0 FreeSans 448 0 0 0 cfgreg_do[29]
port 77 nsew signal tristate
flabel metal3 s 49200 22176 50000 22288 0 FreeSans 448 0 0 0 cfgreg_do[2]
port 78 nsew signal tristate
flabel metal3 s 0 3360 800 3472 0 FreeSans 448 0 0 0 cfgreg_do[30]
port 79 nsew signal tristate
flabel metal2 s 26880 0 26992 800 0 FreeSans 448 90 0 0 cfgreg_do[31]
port 80 nsew signal tristate
flabel metal3 s 49200 20160 50000 20272 0 FreeSans 448 0 0 0 cfgreg_do[3]
port 81 nsew signal tristate
flabel metal2 s 36960 0 37072 800 0 FreeSans 448 90 0 0 cfgreg_do[4]
port 82 nsew signal tristate
flabel metal2 s 38304 0 38416 800 0 FreeSans 448 90 0 0 cfgreg_do[5]
port 83 nsew signal tristate
flabel metal3 s 49200 42336 50000 42448 0 FreeSans 448 0 0 0 cfgreg_do[6]
port 84 nsew signal tristate
flabel metal3 s 0 45024 800 45136 0 FreeSans 448 0 0 0 cfgreg_do[7]
port 85 nsew signal tristate
flabel metal2 s 40992 0 41104 800 0 FreeSans 448 90 0 0 cfgreg_do[8]
port 86 nsew signal tristate
flabel metal2 s 41664 0 41776 800 0 FreeSans 448 90 0 0 cfgreg_do[9]
port 87 nsew signal tristate
flabel metal2 s 30912 0 31024 800 0 FreeSans 448 90 0 0 cfgreg_we[0]
port 88 nsew signal input
flabel metal2 s 44352 0 44464 800 0 FreeSans 448 90 0 0 cfgreg_we[1]
port 89 nsew signal input
flabel metal2 s 10080 0 10192 800 0 FreeSans 448 90 0 0 cfgreg_we[2]
port 90 nsew signal input
flabel metal2 s 22848 0 22960 800 0 FreeSans 448 90 0 0 cfgreg_we[3]
port 91 nsew signal input
flabel metal3 s 0 44352 800 44464 0 FreeSans 448 0 0 0 clk
port 92 nsew signal input
flabel metal2 s 0 0 112 800 0 FreeSans 448 90 0 0 flash_in[0]
port 93 nsew signal input
flabel metal2 s 15456 0 15568 800 0 FreeSans 448 90 0 0 flash_in[1]
port 94 nsew signal input
flabel metal3 s 49200 24864 50000 24976 0 FreeSans 448 0 0 0 flash_in[2]
port 95 nsew signal input
flabel metal3 s 49200 24192 50000 24304 0 FreeSans 448 0 0 0 flash_in[3]
port 96 nsew signal input
flabel metal3 s 49200 21504 50000 21616 0 FreeSans 448 0 0 0 flash_in[4]
port 97 nsew signal input
flabel metal3 s 49200 20832 50000 20944 0 FreeSans 448 0 0 0 flash_in[5]
port 98 nsew signal input
flabel metal3 s 49200 45696 50000 45808 0 FreeSans 448 0 0 0 flash_oeb[0]
port 99 nsew signal tristate
flabel metal3 s 0 4704 800 4816 0 FreeSans 448 0 0 0 flash_oeb[1]
port 100 nsew signal tristate
flabel metal2 s 40320 0 40432 800 0 FreeSans 448 90 0 0 flash_oeb[2]
port 101 nsew signal tristate
flabel metal2 s 39648 0 39760 800 0 FreeSans 448 90 0 0 flash_oeb[3]
port 102 nsew signal tristate
flabel metal3 s 49200 8064 50000 8176 0 FreeSans 448 0 0 0 flash_oeb[4]
port 103 nsew signal tristate
flabel metal3 s 49200 8736 50000 8848 0 FreeSans 448 0 0 0 flash_oeb[5]
port 104 nsew signal tristate
flabel metal2 s 38976 0 39088 800 0 FreeSans 448 90 0 0 flash_out[0]
port 105 nsew signal tristate
flabel metal2 s 37632 0 37744 800 0 FreeSans 448 90 0 0 flash_out[1]
port 106 nsew signal tristate
flabel metal2 s 32928 0 33040 800 0 FreeSans 448 90 0 0 flash_out[2]
port 107 nsew signal tristate
flabel metal2 s 20832 0 20944 800 0 FreeSans 448 90 0 0 flash_out[3]
port 108 nsew signal tristate
flabel metal2 s 26208 0 26320 800 0 FreeSans 448 90 0 0 flash_out[4]
port 109 nsew signal tristate
flabel metal2 s 29568 0 29680 800 0 FreeSans 448 90 0 0 flash_out[5]
port 110 nsew signal tristate
flabel metal2 s 23520 49200 23632 50000 0 FreeSans 448 90 0 0 rdata[0]
port 111 nsew signal tristate
flabel metal2 s 38304 49200 38416 50000 0 FreeSans 448 90 0 0 rdata[10]
port 112 nsew signal tristate
flabel metal2 s 39648 49200 39760 50000 0 FreeSans 448 90 0 0 rdata[11]
port 113 nsew signal tristate
flabel metal3 s 49200 39648 50000 39760 0 FreeSans 448 0 0 0 rdata[12]
port 114 nsew signal tristate
flabel metal3 s 49200 38976 50000 39088 0 FreeSans 448 0 0 0 rdata[13]
port 115 nsew signal tristate
flabel metal2 s 34944 49200 35056 50000 0 FreeSans 448 90 0 0 rdata[14]
port 116 nsew signal tristate
flabel metal2 s 37632 49200 37744 50000 0 FreeSans 448 90 0 0 rdata[15]
port 117 nsew signal tristate
flabel metal2 s 33600 49200 33712 50000 0 FreeSans 448 90 0 0 rdata[16]
port 118 nsew signal tristate
flabel metal2 s 36288 49200 36400 50000 0 FreeSans 448 90 0 0 rdata[17]
port 119 nsew signal tristate
flabel metal3 s 49200 41664 50000 41776 0 FreeSans 448 0 0 0 rdata[18]
port 120 nsew signal tristate
flabel metal2 s 44352 49200 44464 50000 0 FreeSans 448 90 0 0 rdata[19]
port 121 nsew signal tristate
flabel metal2 s 26208 49200 26320 50000 0 FreeSans 448 90 0 0 rdata[1]
port 122 nsew signal tristate
flabel metal3 s 49200 40320 50000 40432 0 FreeSans 448 0 0 0 rdata[20]
port 123 nsew signal tristate
flabel metal3 s 49200 34944 50000 35056 0 FreeSans 448 0 0 0 rdata[21]
port 124 nsew signal tristate
flabel metal2 s 30240 49200 30352 50000 0 FreeSans 448 90 0 0 rdata[22]
port 125 nsew signal tristate
flabel metal2 s 31584 49200 31696 50000 0 FreeSans 448 90 0 0 rdata[23]
port 126 nsew signal tristate
flabel metal2 s 32928 49200 33040 50000 0 FreeSans 448 90 0 0 rdata[24]
port 127 nsew signal tristate
flabel metal2 s 32256 49200 32368 50000 0 FreeSans 448 90 0 0 rdata[25]
port 128 nsew signal tristate
flabel metal3 s 49200 33600 50000 33712 0 FreeSans 448 0 0 0 rdata[26]
port 129 nsew signal tristate
flabel metal3 s 49200 32256 50000 32368 0 FreeSans 448 0 0 0 rdata[27]
port 130 nsew signal tristate
flabel metal3 s 49200 31584 50000 31696 0 FreeSans 448 0 0 0 rdata[28]
port 131 nsew signal tristate
flabel metal3 s 49200 34272 50000 34384 0 FreeSans 448 0 0 0 rdata[29]
port 132 nsew signal tristate
flabel metal3 s 49200 29568 50000 29680 0 FreeSans 448 0 0 0 rdata[2]
port 133 nsew signal tristate
flabel metal2 s 30912 49200 31024 50000 0 FreeSans 448 90 0 0 rdata[30]
port 134 nsew signal tristate
flabel metal3 s 49200 30912 50000 31024 0 FreeSans 448 0 0 0 rdata[31]
port 135 nsew signal tristate
flabel metal3 s 49200 28896 50000 29008 0 FreeSans 448 0 0 0 rdata[3]
port 136 nsew signal tristate
flabel metal3 s 49200 22848 50000 22960 0 FreeSans 448 0 0 0 rdata[4]
port 137 nsew signal tristate
flabel metal3 s 49200 30240 50000 30352 0 FreeSans 448 0 0 0 rdata[5]
port 138 nsew signal tristate
flabel metal3 s 49200 27552 50000 27664 0 FreeSans 448 0 0 0 rdata[6]
port 139 nsew signal tristate
flabel metal3 s 49200 28224 50000 28336 0 FreeSans 448 0 0 0 rdata[7]
port 140 nsew signal tristate
flabel metal2 s 25536 49200 25648 50000 0 FreeSans 448 90 0 0 rdata[8]
port 141 nsew signal tristate
flabel metal2 s 26880 49200 26992 50000 0 FreeSans 448 90 0 0 rdata[9]
port 142 nsew signal tristate
flabel metal3 s 0 29568 800 29680 0 FreeSans 448 0 0 0 ready
port 143 nsew signal tristate
flabel metal2 s 18816 0 18928 800 0 FreeSans 448 90 0 0 resetn
port 144 nsew signal input
flabel metal3 s 0 26880 800 26992 0 FreeSans 448 0 0 0 valid
port 145 nsew signal input
flabel metal4 s 4448 3076 4768 46316 0 FreeSans 1280 90 0 0 vdd
port 146 nsew power bidirectional
flabel metal4 s 35168 3076 35488 46316 0 FreeSans 1280 90 0 0 vdd
port 146 nsew power bidirectional
flabel metal4 s 19808 3076 20128 46316 0 FreeSans 1280 90 0 0 vss
port 147 nsew ground bidirectional
rlabel metal1 24976 46256 24976 46256 0 vdd
rlabel metal1 24976 45472 24976 45472 0 vss
rlabel metal2 2520 14896 2520 14896 0 _0000_
rlabel metal3 4088 18984 4088 18984 0 _0001_
rlabel metal2 2520 11760 2520 11760 0 _0002_
rlabel metal2 7000 15148 7000 15148 0 _0003_
rlabel metal2 13272 15624 13272 15624 0 _0004_
rlabel metal2 2520 20664 2520 20664 0 _0005_
rlabel metal2 13832 11088 13832 11088 0 _0006_
rlabel metal3 3864 18312 3864 18312 0 _0007_
rlabel metal2 3920 9912 3920 9912 0 _0008_
rlabel metal2 8008 15484 8008 15484 0 _0009_
rlabel metal2 3864 16240 3864 16240 0 _0010_
rlabel metal2 2520 13328 2520 13328 0 _0011_
rlabel metal2 7504 15848 7504 15848 0 _0012_
rlabel metal2 29064 45248 29064 45248 0 _0013_
rlabel metal2 27384 38304 27384 38304 0 _0014_
rlabel metal2 37464 40712 37464 40712 0 _0015_
rlabel metal2 38584 43904 38584 43904 0 _0016_
rlabel metal2 44856 36736 44856 36736 0 _0017_
rlabel metal2 40320 36344 40320 36344 0 _0018_
rlabel metal2 33768 36120 33768 36120 0 _0019_
rlabel metal2 37800 36960 37800 36960 0 _0020_
rlabel metal3 23856 18424 23856 18424 0 _0021_
rlabel metal2 31304 42784 31304 42784 0 _0022_
rlabel metal2 33880 41440 33880 41440 0 _0023_
rlabel metal3 42392 40936 42392 40936 0 _0024_
rlabel metal2 43960 43848 43960 43848 0 _0025_
rlabel metal2 41720 37688 41720 37688 0 _0026_
rlabel metal3 45696 33432 45696 33432 0 _0027_
rlabel metal2 32088 34552 32088 34552 0 _0028_
rlabel metal2 36120 34440 36120 34440 0 _0029_
rlabel metal2 26600 17248 26600 17248 0 _0030_
rlabel metal2 29624 22008 29624 22008 0 _0031_
rlabel metal3 31752 20888 31752 20888 0 _0032_
rlabel metal2 31584 23800 31584 23800 0 _0033_
rlabel metal3 30520 24920 30520 24920 0 _0034_
rlabel metal2 26264 22008 26264 22008 0 _0035_
rlabel metal2 26488 19600 26488 19600 0 _0036_
rlabel metal3 45528 12824 45528 12824 0 _0037_
rlabel metal2 38920 9296 38920 9296 0 _0038_
rlabel metal2 21448 44352 21448 44352 0 _0039_
rlabel metal2 24248 42392 24248 42392 0 _0040_
rlabel metal2 37800 29848 37800 29848 0 _0041_
rlabel metal3 44856 28504 44856 28504 0 _0042_
rlabel metal2 45304 21448 45304 21448 0 _0043_
rlabel metal2 46088 30688 46088 30688 0 _0044_
rlabel metal2 30296 27328 30296 27328 0 _0045_
rlabel metal2 34440 27328 34440 27328 0 _0046_
rlabel metal2 25256 45024 25256 45024 0 _0047_
rlabel metal2 25256 39256 25256 39256 0 _0048_
rlabel metal2 37016 41944 37016 41944 0 _0049_
rlabel metal2 37912 45416 37912 45416 0 _0050_
rlabel metal2 43288 39928 43288 39928 0 _0051_
rlabel metal2 40936 39256 40936 39256 0 _0052_
rlabel metal2 33096 39256 33096 39256 0 _0053_
rlabel metal2 36456 38304 36456 38304 0 _0054_
rlabel metal2 31080 45024 31080 45024 0 _0055_
rlabel metal2 34664 45416 34664 45416 0 _0056_
rlabel metal2 45304 41440 45304 41440 0 _0057_
rlabel metal2 42616 45416 42616 45416 0 _0058_
rlabel metal3 45696 39704 45696 39704 0 _0059_
rlabel metal2 45752 37212 45752 37212 0 _0060_
rlabel metal2 28728 36568 28728 36568 0 _0061_
rlabel metal2 29960 33824 29960 33824 0 _0062_
rlabel metal2 30296 41272 30296 41272 0 _0063_
rlabel metal2 30072 38528 30072 38528 0 _0064_
rlabel metal3 39312 33096 39312 33096 0 _0065_
rlabel metal2 39928 31864 39928 31864 0 _0066_
rlabel metal2 44968 31304 44968 31304 0 _0067_
rlabel metal2 41720 34440 41720 34440 0 _0068_
rlabel metal2 29960 31892 29960 31892 0 _0069_
rlabel metal2 33432 31416 33432 31416 0 _0070_
rlabel metal3 13552 16296 13552 16296 0 _0071_
rlabel metal3 14672 9688 14672 9688 0 _0072_
rlabel metal3 14728 9240 14728 9240 0 _0073_
rlabel metal2 13888 8904 13888 8904 0 _0074_
rlabel metal2 27832 10192 27832 10192 0 _0075_
rlabel metal2 18648 19712 18648 19712 0 _0076_
rlabel metal2 19544 17192 19544 17192 0 _0077_
rlabel metal2 17976 14168 17976 14168 0 _0078_
rlabel metal2 21784 18760 21784 18760 0 _0079_
rlabel metal2 26824 24640 26824 24640 0 _0080_
rlabel metal2 27160 27552 27160 27552 0 _0081_
rlabel metal2 23240 24416 23240 24416 0 _0082_
rlabel metal2 24024 26208 24024 26208 0 _0083_
rlabel metal2 15624 12600 15624 12600 0 _0084_
rlabel metal2 14728 18032 14728 18032 0 _0085_
rlabel metal2 18648 11928 18648 11928 0 _0086_
rlabel metal2 27048 43008 27048 43008 0 _0087_
rlabel metal2 27776 41272 27776 41272 0 _0088_
rlabel metal2 36680 31500 36680 31500 0 _0089_
rlabel metal2 41720 29736 41720 29736 0 _0090_
rlabel metal2 44632 25144 44632 25144 0 _0091_
rlabel metal3 45696 27160 45696 27160 0 _0092_
rlabel metal2 29176 30296 29176 30296 0 _0093_
rlabel metal2 33432 28896 33432 28896 0 _0094_
rlabel metal3 13384 21672 13384 21672 0 _0095_
rlabel metal2 2520 22512 2520 22512 0 _0096_
rlabel metal2 6440 22736 6440 22736 0 _0097_
rlabel metal2 23240 7448 23240 7448 0 _0098_
rlabel metal2 16968 5432 16968 5432 0 _0099_
rlabel metal2 7224 7000 7224 7000 0 _0100_
rlabel metal2 6272 4424 6272 4424 0 _0101_
rlabel metal2 6664 4256 6664 4256 0 _0102_
rlabel metal3 11368 4200 11368 4200 0 _0103_
rlabel metal2 11592 7112 11592 7112 0 _0104_
rlabel metal2 14504 6272 14504 6272 0 _0105_
rlabel metal2 40152 5432 40152 5432 0 _0106_
rlabel metal2 42168 7616 42168 7616 0 _0107_
rlabel metal2 45864 6664 45864 6664 0 _0108_
rlabel metal3 44128 4424 44128 4424 0 _0109_
rlabel metal2 36512 5992 36512 5992 0 _0110_
rlabel metal2 38752 4424 38752 4424 0 _0111_
rlabel metal2 32648 5432 32648 5432 0 _0112_
rlabel metal2 19488 4424 19488 4424 0 _0113_
rlabel metal2 24248 5432 24248 5432 0 _0114_
rlabel metal2 27496 4480 27496 4480 0 _0115_
rlabel metal2 22792 6160 22792 6160 0 _0116_
rlabel metal2 41496 11032 41496 11032 0 _0117_
rlabel metal2 33768 25760 33768 25760 0 _0118_
rlabel metal2 35336 20272 35336 20272 0 _0119_
rlabel metal2 39144 21392 39144 21392 0 _0120_
rlabel metal2 45416 21728 45416 21728 0 _0121_
rlabel metal2 43624 23352 43624 23352 0 _0122_
rlabel metal2 43400 25424 43400 25424 0 _0123_
rlabel metal2 38472 25704 38472 25704 0 _0124_
rlabel metal2 38248 27104 38248 27104 0 _0125_
rlabel metal2 31528 9968 31528 9968 0 _0126_
rlabel metal2 32536 11536 32536 11536 0 _0127_
rlabel metal2 24136 11760 24136 11760 0 _0128_
rlabel metal3 25480 10696 25480 10696 0 _0129_
rlabel metal2 22680 12432 22680 12432 0 _0130_
rlabel metal2 23240 10080 23240 10080 0 _0131_
rlabel metal2 46088 17304 46088 17304 0 _0132_
rlabel metal3 46480 16744 46480 16744 0 _0133_
rlabel metal2 2520 8792 2520 8792 0 _0134_
rlabel metal2 4088 8400 4088 8400 0 _0135_
rlabel metal2 6888 9184 6888 9184 0 _0136_
rlabel metal2 45640 11032 45640 11032 0 _0137_
rlabel metal2 41608 9464 41608 9464 0 _0138_
rlabel metal2 33880 10920 33880 10920 0 _0139_
rlabel metal2 31584 13048 31584 13048 0 _0140_
rlabel metal2 19992 26432 19992 26432 0 _0141_
rlabel metal2 18872 23464 18872 23464 0 _0142_
rlabel metal2 24808 30912 24808 30912 0 _0143_
rlabel metal3 23072 31752 23072 31752 0 _0144_
rlabel metal3 25144 33992 25144 33992 0 _0145_
rlabel metal2 24584 36120 24584 36120 0 _0146_
rlabel metal2 19096 43064 19096 43064 0 _0147_
rlabel metal2 21672 38808 21672 38808 0 _0148_
rlabel metal2 18424 43120 18424 43120 0 _0149_
rlabel metal2 17304 41944 17304 41944 0 _0150_
rlabel metal2 13720 43120 13720 43120 0 _0151_
rlabel metal2 13888 41944 13888 41944 0 _0152_
rlabel metal3 10528 43624 10528 43624 0 _0153_
rlabel metal3 6944 36568 6944 36568 0 _0154_
rlabel metal2 2968 40600 2968 40600 0 _0155_
rlabel metal2 3752 39648 3752 39648 0 _0156_
rlabel metal2 2520 38668 2520 38668 0 _0157_
rlabel metal2 2408 36120 2408 36120 0 _0158_
rlabel metal2 2576 24024 2576 24024 0 _0159_
rlabel metal3 15848 25592 15848 25592 0 _0160_
rlabel metal2 2520 26152 2520 26152 0 _0161_
rlabel metal2 15624 43680 15624 43680 0 _0162_
rlabel metal3 3808 27720 3808 27720 0 _0163_
rlabel metal2 6888 43680 6888 43680 0 _0164_
rlabel metal2 46536 19264 46536 19264 0 _0165_
rlabel metal2 31584 37352 31584 37352 0 _0166_
rlabel metal2 31304 36344 31304 36344 0 _0167_
rlabel metal2 31192 33040 31192 33040 0 _0168_
rlabel metal2 30968 41272 30968 41272 0 _0169_
rlabel metal2 31136 37464 31136 37464 0 _0170_
rlabel metal2 44072 34888 44072 34888 0 _0171_
rlabel metal2 40264 33040 40264 33040 0 _0172_
rlabel metal3 39816 31192 39816 31192 0 _0173_
rlabel metal2 44520 31640 44520 31640 0 _0174_
rlabel metal3 42000 34888 42000 34888 0 _0175_
rlabel metal3 30884 31080 30884 31080 0 _0176_
rlabel metal3 30184 31192 30184 31192 0 _0177_
rlabel metal2 34048 30968 34048 30968 0 _0178_
rlabel metal3 8792 16968 8792 16968 0 _0179_
rlabel metal2 8736 20552 8736 20552 0 _0180_
rlabel metal3 4480 9016 4480 9016 0 _0181_
rlabel metal2 15176 8372 15176 8372 0 _0182_
rlabel metal2 10248 13608 10248 13608 0 _0183_
rlabel metal2 10472 13664 10472 13664 0 _0184_
rlabel metal3 7336 12712 7336 12712 0 _0185_
rlabel metal2 9800 11648 9800 11648 0 _0186_
rlabel metal2 10472 10192 10472 10192 0 _0187_
rlabel metal2 10360 10640 10360 10640 0 _0188_
rlabel metal2 11200 9688 11200 9688 0 _0189_
rlabel metal2 15176 8792 15176 8792 0 _0190_
rlabel metal2 16296 9016 16296 9016 0 _0191_
rlabel metal2 16408 8008 16408 8008 0 _0192_
rlabel metal2 6664 7896 6664 7896 0 _0193_
rlabel metal2 13720 9016 13720 9016 0 _0194_
rlabel metal2 28056 8792 28056 8792 0 _0195_
rlabel metal3 30352 10584 30352 10584 0 _0196_
rlabel metal2 29064 9912 29064 9912 0 _0197_
rlabel metal2 31528 11956 31528 11956 0 _0198_
rlabel metal3 13496 13944 13496 13944 0 _0199_
rlabel metal2 16688 23128 16688 23128 0 _0200_
rlabel metal2 18200 24976 18200 24976 0 _0201_
rlabel metal2 18984 22736 18984 22736 0 _0202_
rlabel metal2 15400 20384 15400 20384 0 _0203_
rlabel metal2 13720 19040 13720 19040 0 _0204_
rlabel metal2 12264 22848 12264 22848 0 _0205_
rlabel metal3 13104 23688 13104 23688 0 _0206_
rlabel metal2 12040 25088 12040 25088 0 _0207_
rlabel metal2 10920 21728 10920 21728 0 _0208_
rlabel metal2 13328 24920 13328 24920 0 _0209_
rlabel metal2 18984 19264 18984 19264 0 _0210_
rlabel metal3 20944 17640 20944 17640 0 _0211_
rlabel metal2 19656 19264 19656 19264 0 _0212_
rlabel metal2 18704 18648 18704 18648 0 _0213_
rlabel metal3 14112 23128 14112 23128 0 _0214_
rlabel metal2 11816 20328 11816 20328 0 _0215_
rlabel metal3 12768 19992 12768 19992 0 _0216_
rlabel metal2 14056 19936 14056 19936 0 _0217_
rlabel metal2 17416 19264 17416 19264 0 _0218_
rlabel metal2 16184 24136 16184 24136 0 _0219_
rlabel metal2 16520 19880 16520 19880 0 _0220_
rlabel metal2 17304 19264 17304 19264 0 _0221_
rlabel metal2 19320 16744 19320 16744 0 _0222_
rlabel metal2 18984 16912 18984 16912 0 _0223_
rlabel metal3 14784 14280 14784 14280 0 _0224_
rlabel metal3 16072 19880 16072 19880 0 _0225_
rlabel metal2 16128 20216 16128 20216 0 _0226_
rlabel metal3 17808 15176 17808 15176 0 _0227_
rlabel metal2 18312 14448 18312 14448 0 _0228_
rlabel metal2 10808 24192 10808 24192 0 _0229_
rlabel metal2 14168 19768 14168 19768 0 _0230_
rlabel metal2 14504 19208 14504 19208 0 _0231_
rlabel metal3 20776 19712 20776 19712 0 _0232_
rlabel metal3 20888 19208 20888 19208 0 _0233_
rlabel metal2 15176 20272 15176 20272 0 _0234_
rlabel metal3 17192 23800 17192 23800 0 _0235_
rlabel metal2 16408 24304 16408 24304 0 _0236_
rlabel metal2 15400 12544 15400 12544 0 _0237_
rlabel metal2 16184 23520 16184 23520 0 _0238_
rlabel metal3 16184 23968 16184 23968 0 _0239_
rlabel metal2 26824 23240 26824 23240 0 _0240_
rlabel metal2 24472 26320 24472 26320 0 _0241_
rlabel metal2 26488 24360 26488 24360 0 _0242_
rlabel metal2 18256 23464 18256 23464 0 _0243_
rlabel metal2 12488 25984 12488 25984 0 _0244_
rlabel metal2 18480 26824 18480 26824 0 _0245_
rlabel metal3 22736 26040 22736 26040 0 _0246_
rlabel metal2 26712 27160 26712 27160 0 _0247_
rlabel metal2 18088 24304 18088 24304 0 _0248_
rlabel metal2 17864 23576 17864 23576 0 _0249_
rlabel metal3 21056 22904 21056 22904 0 _0250_
rlabel metal2 23352 24024 23352 24024 0 _0251_
rlabel metal2 18200 25312 18200 25312 0 _0252_
rlabel metal2 17304 25256 17304 25256 0 _0253_
rlabel metal2 23800 25872 23800 25872 0 _0254_
rlabel metal2 23464 26096 23464 26096 0 _0255_
rlabel metal2 15176 12488 15176 12488 0 _0256_
rlabel metal3 16184 12040 16184 12040 0 _0257_
rlabel metal3 15568 18200 15568 18200 0 _0258_
rlabel metal3 19040 12040 19040 12040 0 _0259_
rlabel metal2 26600 28168 26600 28168 0 _0260_
rlabel metal3 28392 29960 28392 29960 0 _0261_
rlabel metal2 29624 28896 29624 28896 0 _0262_
rlabel metal3 28336 42616 28336 42616 0 _0263_
rlabel metal2 28280 40824 28280 40824 0 _0264_
rlabel metal2 37688 32256 37688 32256 0 _0265_
rlabel metal2 41216 28840 41216 28840 0 _0266_
rlabel metal2 31864 29344 31864 29344 0 _0267_
rlabel metal3 45472 23352 45472 23352 0 _0268_
rlabel metal3 46424 28056 46424 28056 0 _0269_
rlabel metal3 30240 28840 30240 28840 0 _0270_
rlabel metal2 33208 29288 33208 29288 0 _0271_
rlabel metal2 13720 22176 13720 22176 0 _0272_
rlabel metal3 12264 22344 12264 22344 0 _0273_
rlabel metal2 17080 29120 17080 29120 0 _0274_
rlabel metal2 16856 26600 16856 26600 0 _0275_
rlabel metal3 7616 23240 7616 23240 0 _0276_
rlabel metal2 18648 39312 18648 39312 0 _0277_
rlabel metal2 16296 43400 16296 43400 0 _0278_
rlabel metal2 10136 22456 10136 22456 0 _0279_
rlabel metal2 7448 22848 7448 22848 0 _0280_
rlabel metal2 19768 43064 19768 43064 0 _0281_
rlabel metal2 6328 21952 6328 21952 0 _0282_
rlabel metal2 19432 5992 19432 5992 0 _0283_
rlabel metal2 25704 4704 25704 4704 0 _0284_
rlabel metal2 17864 4760 17864 4760 0 _0285_
rlabel metal2 23688 6608 23688 6608 0 _0286_
rlabel metal2 15512 4704 15512 4704 0 _0287_
rlabel metal3 19152 5992 19152 5992 0 _0288_
rlabel metal2 17808 5880 17808 5880 0 _0289_
rlabel metal2 17528 4984 17528 4984 0 _0290_
rlabel metal2 18536 5432 18536 5432 0 _0291_
rlabel metal2 7784 5656 7784 5656 0 _0292_
rlabel metal3 7840 5880 7840 5880 0 _0293_
rlabel metal2 8232 5768 8232 5768 0 _0294_
rlabel metal2 7560 6720 7560 6720 0 _0295_
rlabel metal2 6216 3976 6216 3976 0 _0296_
rlabel metal2 7280 4088 7280 4088 0 _0297_
rlabel metal2 6048 5096 6048 5096 0 _0298_
rlabel metal3 12544 5992 12544 5992 0 _0299_
rlabel metal3 12936 6440 12936 6440 0 _0300_
rlabel metal2 8120 5544 8120 5544 0 _0301_
rlabel metal2 11368 5768 11368 5768 0 _0302_
rlabel metal2 6552 4032 6552 4032 0 _0303_
rlabel metal2 8568 4872 8568 4872 0 _0304_
rlabel metal2 13496 5376 13496 5376 0 _0305_
rlabel metal2 8904 4648 8904 4648 0 _0306_
rlabel metal3 18424 6720 18424 6720 0 _0307_
rlabel metal2 13272 5824 13272 5824 0 _0308_
rlabel metal3 12712 6104 12712 6104 0 _0309_
rlabel metal2 12152 6832 12152 6832 0 _0310_
rlabel metal2 15288 6496 15288 6496 0 _0311_
rlabel metal2 14840 5600 14840 5600 0 _0312_
rlabel metal2 42840 4144 42840 4144 0 _0313_
rlabel metal3 22456 6664 22456 6664 0 _0314_
rlabel metal2 40152 4704 40152 4704 0 _0315_
rlabel metal2 40488 4872 40488 4872 0 _0316_
rlabel metal3 41552 7336 41552 7336 0 _0317_
rlabel metal2 44856 6384 44856 6384 0 _0318_
rlabel metal2 43736 7224 43736 7224 0 _0319_
rlabel metal2 43512 7056 43512 7056 0 _0320_
rlabel metal2 43848 5040 43848 5040 0 _0321_
rlabel metal2 44184 5712 44184 5712 0 _0322_
rlabel metal2 45416 9856 45416 9856 0 _0323_
rlabel metal2 47208 5712 47208 5712 0 _0324_
rlabel metal3 42392 3304 42392 3304 0 _0325_
rlabel metal2 38920 5656 38920 5656 0 _0326_
rlabel metal3 44968 8904 44968 8904 0 _0327_
rlabel metal2 30128 4872 30128 4872 0 _0328_
rlabel metal2 25816 4704 25816 4704 0 _0329_
rlabel metal2 33768 6272 33768 6272 0 _0330_
rlabel metal2 35672 5208 35672 5208 0 _0331_
rlabel metal2 36344 5880 36344 5880 0 _0332_
rlabel metal2 24584 4648 24584 4648 0 _0333_
rlabel metal3 35336 5096 35336 5096 0 _0334_
rlabel metal2 35224 5264 35224 5264 0 _0335_
rlabel metal3 37016 5096 37016 5096 0 _0336_
rlabel metal3 34944 5880 34944 5880 0 _0337_
rlabel metal2 33880 4704 33880 4704 0 _0338_
rlabel metal2 35000 5376 35000 5376 0 _0339_
rlabel metal3 22680 5320 22680 5320 0 _0340_
rlabel metal2 22792 4368 22792 4368 0 _0341_
rlabel metal2 20216 4816 20216 4816 0 _0342_
rlabel metal2 24696 4760 24696 4760 0 _0343_
rlabel metal2 24584 4144 24584 4144 0 _0344_
rlabel metal2 25648 4200 25648 4200 0 _0345_
rlabel metal2 33096 4760 33096 4760 0 _0346_
rlabel metal2 29288 5376 29288 5376 0 _0347_
rlabel metal2 28896 5208 28896 5208 0 _0348_
rlabel metal2 22624 6104 22624 6104 0 _0349_
rlabel metal2 22232 5600 22232 5600 0 _0350_
rlabel metal3 39816 22288 39816 22288 0 _0351_
rlabel metal2 35168 23352 35168 23352 0 _0352_
rlabel metal2 35672 16520 35672 16520 0 _0353_
rlabel metal2 37688 22568 37688 22568 0 _0354_
rlabel metal2 38920 23632 38920 23632 0 _0355_
rlabel metal2 34552 25144 34552 25144 0 _0356_
rlabel metal2 35112 21560 35112 21560 0 _0357_
rlabel metal2 34776 21672 34776 21672 0 _0358_
rlabel metal2 42952 24304 42952 24304 0 _0359_
rlabel metal2 43736 20552 43736 20552 0 _0360_
rlabel metal3 38304 21672 38304 21672 0 _0361_
rlabel metal2 38808 22400 38808 22400 0 _0362_
rlabel metal2 39816 25984 39816 25984 0 _0363_
rlabel metal2 39368 22456 39368 22456 0 _0364_
rlabel metal3 41832 24696 41832 24696 0 _0365_
rlabel metal2 42168 20440 42168 20440 0 _0366_
rlabel metal2 43736 21896 43736 21896 0 _0367_
rlabel metal2 43176 22624 43176 22624 0 _0368_
rlabel metal2 41832 22176 41832 22176 0 _0369_
rlabel metal3 41552 22232 41552 22232 0 _0370_
rlabel metal2 42616 23856 42616 23856 0 _0371_
rlabel metal3 39032 26936 39032 26936 0 _0372_
rlabel metal2 43288 23968 43288 23968 0 _0373_
rlabel metal2 40712 24136 40712 24136 0 _0374_
rlabel metal2 43064 25424 43064 25424 0 _0375_
rlabel metal2 43400 24808 43400 24808 0 _0376_
rlabel metal2 41384 25704 41384 25704 0 _0377_
rlabel metal2 38696 25536 38696 25536 0 _0378_
rlabel metal2 38136 25536 38136 25536 0 _0379_
rlabel metal2 39256 24976 39256 24976 0 _0380_
rlabel metal2 39480 25928 39480 25928 0 _0381_
rlabel metal2 40040 26712 40040 26712 0 _0382_
rlabel metal2 23688 16352 23688 16352 0 _0383_
rlabel metal2 30632 10864 30632 10864 0 _0384_
rlabel metal2 31640 10584 31640 10584 0 _0385_
rlabel metal2 31192 12656 31192 12656 0 _0386_
rlabel metal2 30072 11872 30072 11872 0 _0387_
rlabel metal2 26656 14728 26656 14728 0 _0388_
rlabel metal2 26040 14840 26040 14840 0 _0389_
rlabel metal2 27944 15680 27944 15680 0 _0390_
rlabel metal2 23464 15540 23464 15540 0 _0391_
rlabel metal2 24024 12824 24024 12824 0 _0392_
rlabel metal2 25032 13328 25032 13328 0 _0393_
rlabel metal3 25200 15288 25200 15288 0 _0394_
rlabel metal2 24696 13160 24696 13160 0 _0395_
rlabel metal3 24976 14616 24976 14616 0 _0396_
rlabel metal2 23576 14000 23576 14000 0 _0397_
rlabel metal2 23016 12488 23016 12488 0 _0398_
rlabel metal2 27048 14056 27048 14056 0 _0399_
rlabel metal3 25984 14280 25984 14280 0 _0400_
rlabel metal2 24696 14056 24696 14056 0 _0401_
rlabel metal2 43960 18088 43960 18088 0 _0402_
rlabel metal2 44744 18480 44744 18480 0 _0403_
rlabel metal2 47656 17528 47656 17528 0 _0404_
rlabel metal3 46760 16856 46760 16856 0 _0405_
rlabel metal2 45752 17584 45752 17584 0 _0406_
rlabel metal2 45472 16744 45472 16744 0 _0407_
rlabel metal3 41216 14616 41216 14616 0 _0408_
rlabel metal2 42168 16016 42168 16016 0 _0409_
rlabel metal2 38024 16184 38024 16184 0 _0410_
rlabel metal2 39648 18424 39648 18424 0 _0411_
rlabel metal3 40936 18648 40936 18648 0 _0412_
rlabel metal2 41496 15568 41496 15568 0 _0413_
rlabel metal3 42336 15288 42336 15288 0 _0414_
rlabel metal2 9464 10864 9464 10864 0 _0415_
rlabel metal2 9688 10976 9688 10976 0 _0416_
rlabel metal2 6664 10920 6664 10920 0 _0417_
rlabel via2 5208 9128 5208 9128 0 _0418_
rlabel metal2 4200 9688 4200 9688 0 _0419_
rlabel metal2 5320 9296 5320 9296 0 _0420_
rlabel metal2 7896 9912 7896 9912 0 _0421_
rlabel metal2 7448 9688 7448 9688 0 _0422_
rlabel metal3 44184 10584 44184 10584 0 _0423_
rlabel metal2 31136 11368 31136 11368 0 _0424_
rlabel metal2 30632 11312 30632 11312 0 _0425_
rlabel metal2 28896 11144 28896 11144 0 _0426_
rlabel metal2 29512 13440 29512 13440 0 _0427_
rlabel metal2 31136 14392 31136 14392 0 _0428_
rlabel metal3 16800 39592 16800 39592 0 _0429_
rlabel metal2 20328 24472 20328 24472 0 _0430_
rlabel metal2 19376 25368 19376 25368 0 _0431_
rlabel metal2 19320 23800 19320 23800 0 _0432_
rlabel metal2 23128 31808 23128 31808 0 _0433_
rlabel metal2 24416 37240 24416 37240 0 _0434_
rlabel metal2 24528 31192 24528 31192 0 _0435_
rlabel metal3 15736 29512 15736 29512 0 _0436_
rlabel metal2 22456 37800 22456 37800 0 _0437_
rlabel metal2 22120 26992 22120 26992 0 _0438_
rlabel metal3 17640 27832 17640 27832 0 _0439_
rlabel metal2 17808 31192 17808 31192 0 _0440_
rlabel metal2 22344 30184 22344 30184 0 _0441_
rlabel metal3 23128 30296 23128 30296 0 _0442_
rlabel metal2 17416 41552 17416 41552 0 _0443_
rlabel metal2 20776 30352 20776 30352 0 _0444_
rlabel metal3 18424 38808 18424 38808 0 _0445_
rlabel metal3 19712 30184 19712 30184 0 _0446_
rlabel metal2 20664 31024 20664 31024 0 _0447_
rlabel metal2 17864 29288 17864 29288 0 _0448_
rlabel metal2 23016 31920 23016 31920 0 _0449_
rlabel metal4 15848 19432 15848 19432 0 _0450_
rlabel metal3 23520 33320 23520 33320 0 _0451_
rlabel metal2 24248 33432 24248 33432 0 _0452_
rlabel metal2 24864 34104 24864 34104 0 _0453_
rlabel metal2 24136 38668 24136 38668 0 _0454_
rlabel metal2 23016 37520 23016 37520 0 _0455_
rlabel metal3 23912 35896 23912 35896 0 _0456_
rlabel metal2 24248 36400 24248 36400 0 _0457_
rlabel metal3 19040 34664 19040 34664 0 _0458_
rlabel metal2 17304 35140 17304 35140 0 _0459_
rlabel metal2 18536 35000 18536 35000 0 _0460_
rlabel metal2 18816 41272 18816 41272 0 _0461_
rlabel metal3 20720 43512 20720 43512 0 _0462_
rlabel metal2 19432 43064 19432 43064 0 _0463_
rlabel metal2 22120 35672 22120 35672 0 _0464_
rlabel metal2 21392 36232 21392 36232 0 _0465_
rlabel metal2 21224 39032 21224 39032 0 _0466_
rlabel metal3 19264 39480 19264 39480 0 _0467_
rlabel metal2 18424 39116 18424 39116 0 _0468_
rlabel metal2 18928 41048 18928 41048 0 _0469_
rlabel metal2 17640 24024 17640 24024 0 _0470_
rlabel metal2 16464 39816 16464 39816 0 _0471_
rlabel metal2 16520 40992 16520 40992 0 _0472_
rlabel metal2 17640 39760 17640 39760 0 _0473_
rlabel metal2 15680 37352 15680 37352 0 _0474_
rlabel metal2 16072 37632 16072 37632 0 _0475_
rlabel metal2 13664 40600 13664 40600 0 _0476_
rlabel metal2 14336 42728 14336 42728 0 _0477_
rlabel metal3 13216 39816 13216 39816 0 _0478_
rlabel metal2 12488 41328 12488 41328 0 _0479_
rlabel metal2 10248 36008 10248 36008 0 _0480_
rlabel metal3 10640 40488 10640 40488 0 _0481_
rlabel metal2 11928 43624 11928 43624 0 _0482_
rlabel metal2 3304 39648 3304 39648 0 _0483_
rlabel metal2 6104 35476 6104 35476 0 _0484_
rlabel metal2 8008 33992 8008 33992 0 _0485_
rlabel metal2 7728 35000 7728 35000 0 _0486_
rlabel metal2 3192 27776 3192 27776 0 _0487_
rlabel metal3 8008 38136 8008 38136 0 _0488_
rlabel metal2 8232 37072 8232 37072 0 _0489_
rlabel metal3 6552 39144 6552 39144 0 _0490_
rlabel metal2 3976 39592 3976 39592 0 _0491_
rlabel metal2 6664 37744 6664 37744 0 _0492_
rlabel metal2 6104 37632 6104 37632 0 _0493_
rlabel metal3 3808 37464 3808 37464 0 _0494_
rlabel metal2 6552 35672 6552 35672 0 _0495_
rlabel metal2 3304 36848 3304 36848 0 _0496_
rlabel metal2 4312 32536 4312 32536 0 _0497_
rlabel metal2 4760 33040 4760 33040 0 _0498_
rlabel metal2 2968 35280 2968 35280 0 _0499_
rlabel metal2 2184 26544 2184 26544 0 _0500_
rlabel metal2 10696 26600 10696 26600 0 _0501_
rlabel metal3 15260 27048 15260 27048 0 _0502_
rlabel metal2 11704 26600 11704 26600 0 _0503_
rlabel metal2 4648 26488 4648 26488 0 _0504_
rlabel metal3 13104 26264 13104 26264 0 _0505_
rlabel metal2 15512 26376 15512 26376 0 _0506_
rlabel metal2 15176 26712 15176 26712 0 _0507_
rlabel metal2 6328 27216 6328 27216 0 _0508_
rlabel metal2 5208 27104 5208 27104 0 _0509_
rlabel metal2 17248 39816 17248 39816 0 _0510_
rlabel metal2 15736 44576 15736 44576 0 _0511_
rlabel metal2 16520 43792 16520 43792 0 _0512_
rlabel metal2 8232 28896 8232 28896 0 _0513_
rlabel metal2 7112 28616 7112 28616 0 _0514_
rlabel metal2 5656 27944 5656 27944 0 _0515_
rlabel metal2 5320 31192 5320 31192 0 _0516_
rlabel metal2 4536 31864 4536 31864 0 _0517_
rlabel metal2 1456 36568 1456 36568 0 _0518_
rlabel metal2 8008 44296 8008 44296 0 _0519_
rlabel metal2 44240 18312 44240 18312 0 _0520_
rlabel metal3 45864 18312 45864 18312 0 _0521_
rlabel metal2 22232 31192 22232 31192 0 _0522_
rlabel metal2 20608 29624 20608 29624 0 _0523_
rlabel metal2 12824 29344 12824 29344 0 _0524_
rlabel metal2 5320 39704 5320 39704 0 _0525_
rlabel metal2 7336 37632 7336 37632 0 _0526_
rlabel metal2 13272 36568 13272 36568 0 _0527_
rlabel metal2 14504 30184 14504 30184 0 _0528_
rlabel metal2 11368 23352 11368 23352 0 _0529_
rlabel metal3 3416 34328 3416 34328 0 _0530_
rlabel metal2 10248 32480 10248 32480 0 _0531_
rlabel metal2 12376 43064 12376 43064 0 _0532_
rlabel metal3 11144 35784 11144 35784 0 _0533_
rlabel metal2 10752 35448 10752 35448 0 _0534_
rlabel metal2 2576 34328 2576 34328 0 _0535_
rlabel metal2 3136 41832 3136 41832 0 _0536_
rlabel metal2 10584 34160 10584 34160 0 _0537_
rlabel metal2 14168 33992 14168 33992 0 _0538_
rlabel metal2 24696 34216 24696 34216 0 _0539_
rlabel metal2 21784 33432 21784 33432 0 _0540_
rlabel metal2 21000 40320 21000 40320 0 _0541_
rlabel metal2 17528 33208 17528 33208 0 _0542_
rlabel metal3 10024 34888 10024 34888 0 _0543_
rlabel metal2 6944 39592 6944 39592 0 _0544_
rlabel metal2 8904 34776 8904 34776 0 _0545_
rlabel metal2 10360 33600 10360 33600 0 _0546_
rlabel metal2 6328 31192 6328 31192 0 _0547_
rlabel metal2 6440 30576 6440 30576 0 _0548_
rlabel metal2 11144 32704 11144 32704 0 _0549_
rlabel metal2 15512 34832 15512 34832 0 _0550_
rlabel metal2 12264 39144 12264 39144 0 _0551_
rlabel metal2 11592 34048 11592 34048 0 _0552_
rlabel metal2 2408 31024 2408 31024 0 _0553_
rlabel metal2 2744 29008 2744 29008 0 _0554_
rlabel metal2 12824 31696 12824 31696 0 _0555_
rlabel metal2 19320 40208 19320 40208 0 _0556_
rlabel metal3 17808 37912 17808 37912 0 _0557_
rlabel metal3 17752 37744 17752 37744 0 _0558_
rlabel metal2 16856 34384 16856 34384 0 _0559_
rlabel metal2 12488 32480 12488 32480 0 _0560_
rlabel metal2 10808 26376 10808 26376 0 _0561_
rlabel metal2 11928 30576 11928 30576 0 _0562_
rlabel metal2 3808 24920 3808 24920 0 _0563_
rlabel metal2 12152 32424 12152 32424 0 _0564_
rlabel metal2 11928 32592 11928 32592 0 _0565_
rlabel metal3 15624 33152 15624 33152 0 _0566_
rlabel metal2 14840 30296 14840 30296 0 _0567_
rlabel metal2 22792 27888 22792 27888 0 _0568_
rlabel metal2 21336 25312 21336 25312 0 _0569_
rlabel metal2 17752 28336 17752 28336 0 _0570_
rlabel metal3 8680 27832 8680 27832 0 _0571_
rlabel metal2 12992 26488 12992 26488 0 _0572_
rlabel metal2 15904 41944 15904 41944 0 _0573_
rlabel metal2 12096 38024 12096 38024 0 _0574_
rlabel metal2 9128 27104 9128 27104 0 _0575_
rlabel metal2 12488 29064 12488 29064 0 _0576_
rlabel metal2 15512 40544 15512 40544 0 _0577_
rlabel metal2 6272 39816 6272 39816 0 _0578_
rlabel metal3 14000 40376 14000 40376 0 _0579_
rlabel metal4 13048 35000 13048 35000 0 _0580_
rlabel metal2 15176 30464 15176 30464 0 _0581_
rlabel metal2 2856 37968 2856 37968 0 _0582_
rlabel metal3 6328 28840 6328 28840 0 _0583_
rlabel metal2 15512 31304 15512 31304 0 _0584_
rlabel metal2 23352 32480 23352 32480 0 _0585_
rlabel metal2 19432 31416 19432 31416 0 _0586_
rlabel metal2 19656 30744 19656 30744 0 _0587_
rlabel metal2 21672 36568 21672 36568 0 _0588_
rlabel metal2 19712 33432 19712 33432 0 _0589_
rlabel metal3 17080 33992 17080 33992 0 _0590_
rlabel metal2 16184 31248 16184 31248 0 _0591_
rlabel metal3 19936 29624 19936 29624 0 _0592_
rlabel metal2 15624 29400 15624 29400 0 _0593_
rlabel metal2 16408 30408 16408 30408 0 _0594_
rlabel metal3 17976 40376 17976 40376 0 _0595_
rlabel metal3 16128 39032 16128 39032 0 _0596_
rlabel metal2 15960 37352 15960 37352 0 _0597_
rlabel metal2 16576 30968 16576 30968 0 _0598_
rlabel metal2 16744 31472 16744 31472 0 _0599_
rlabel metal3 10920 32536 10920 32536 0 _0600_
rlabel metal2 23016 35056 23016 35056 0 _0601_
rlabel metal4 15400 33320 15400 33320 0 _0602_
rlabel metal3 16184 32424 16184 32424 0 _0603_
rlabel metal3 6608 34328 6608 34328 0 _0604_
rlabel metal2 6608 38808 6608 38808 0 _0605_
rlabel metal2 9912 33376 9912 33376 0 _0606_
rlabel metal2 17752 32536 17752 32536 0 _0607_
rlabel metal2 10136 25648 10136 25648 0 _0608_
rlabel metal2 18536 29680 18536 29680 0 _0609_
rlabel metal2 4536 16744 4536 16744 0 _0610_
rlabel metal2 14280 27272 14280 27272 0 _0611_
rlabel metal2 14728 32032 14728 32032 0 _0612_
rlabel metal3 15372 34216 15372 34216 0 _0613_
rlabel metal3 13496 34888 13496 34888 0 _0614_
rlabel metal3 14616 35000 14616 35000 0 _0615_
rlabel metal2 14896 34104 14896 34104 0 _0616_
rlabel metal2 11480 34384 11480 34384 0 _0617_
rlabel metal3 12936 34104 12936 34104 0 _0618_
rlabel metal2 8904 33600 8904 33600 0 _0619_
rlabel metal2 13608 33992 13608 33992 0 _0620_
rlabel metal3 11872 35336 11872 35336 0 _0621_
rlabel metal2 9352 23800 9352 23800 0 _0622_
rlabel metal2 9184 20776 9184 20776 0 _0623_
rlabel metal3 8400 20776 8400 20776 0 _0624_
rlabel metal2 5880 17640 5880 17640 0 _0625_
rlabel metal2 8064 23352 8064 23352 0 _0626_
rlabel metal3 11480 25592 11480 25592 0 _0627_
rlabel metal2 5880 41664 5880 41664 0 _0628_
rlabel metal2 22736 39592 22736 39592 0 _0629_
rlabel metal3 22344 41104 22344 41104 0 _0630_
rlabel metal2 17528 41944 17528 41944 0 _0631_
rlabel metal2 9352 42280 9352 42280 0 _0632_
rlabel metal2 10136 42448 10136 42448 0 _0633_
rlabel metal2 9800 40880 9800 40880 0 _0634_
rlabel metal2 8456 28280 8456 28280 0 _0635_
rlabel metal2 12936 27328 12936 27328 0 _0636_
rlabel metal2 10584 28896 10584 28896 0 _0637_
rlabel metal2 2632 29064 2632 29064 0 _0638_
rlabel metal3 3052 29512 3052 29512 0 _0639_
rlabel metal2 16856 40040 16856 40040 0 _0640_
rlabel metal2 4984 28840 4984 28840 0 _0641_
rlabel metal3 4984 29400 4984 29400 0 _0642_
rlabel metal3 3164 32648 3164 32648 0 _0643_
rlabel metal2 4872 37464 4872 37464 0 _0644_
rlabel metal2 13272 39480 13272 39480 0 _0645_
rlabel metal2 11592 40824 11592 40824 0 _0646_
rlabel metal2 7728 40152 7728 40152 0 _0647_
rlabel metal2 3248 35448 3248 35448 0 _0648_
rlabel metal2 3416 30632 3416 30632 0 _0649_
rlabel metal2 3528 31808 3528 31808 0 _0650_
rlabel metal2 8680 29120 8680 29120 0 _0651_
rlabel metal3 8120 31752 8120 31752 0 _0652_
rlabel metal2 8232 29904 8232 29904 0 _0653_
rlabel metal3 4704 30856 4704 30856 0 _0654_
rlabel metal2 6328 24192 6328 24192 0 _0655_
rlabel metal3 8176 30184 8176 30184 0 _0656_
rlabel metal2 18312 35616 18312 35616 0 _0657_
rlabel metal2 19376 39704 19376 39704 0 _0658_
rlabel metal2 16576 37240 16576 37240 0 _0659_
rlabel metal2 16184 35588 16184 35588 0 _0660_
rlabel metal2 20664 40320 20664 40320 0 _0661_
rlabel metal2 17080 41440 17080 41440 0 _0662_
rlabel metal2 16072 39648 16072 39648 0 _0663_
rlabel metal2 16072 33880 16072 33880 0 _0664_
rlabel metal2 14616 31192 14616 31192 0 _0665_
rlabel metal2 15624 34944 15624 34944 0 _0666_
rlabel metal2 10136 31304 10136 31304 0 _0667_
rlabel metal2 13720 30296 13720 30296 0 _0668_
rlabel metal2 15736 28280 15736 28280 0 _0669_
rlabel metal2 14056 31136 14056 31136 0 _0670_
rlabel metal2 14504 30912 14504 30912 0 _0671_
rlabel metal2 8176 35112 8176 35112 0 _0672_
rlabel metal2 20328 39200 20328 39200 0 _0673_
rlabel metal3 10080 41944 10080 41944 0 _0674_
rlabel metal2 8848 37240 8848 37240 0 _0675_
rlabel metal2 9912 36064 9912 36064 0 _0676_
rlabel metal2 7560 33936 7560 33936 0 _0677_
rlabel metal2 7728 34664 7728 34664 0 _0678_
rlabel metal2 8120 32928 8120 32928 0 _0679_
rlabel metal2 7896 30968 7896 30968 0 _0680_
rlabel metal2 9072 35448 9072 35448 0 _0681_
rlabel metal2 20552 31584 20552 31584 0 _0682_
rlabel metal3 8736 30744 8736 30744 0 _0683_
rlabel metal2 6552 24192 6552 24192 0 _0684_
rlabel metal2 7224 25872 7224 25872 0 _0685_
rlabel metal2 5600 35000 5600 35000 0 _0686_
rlabel metal2 7112 38864 7112 38864 0 _0687_
rlabel metal2 6104 38668 6104 38668 0 _0688_
rlabel metal2 7448 26488 7448 26488 0 _0689_
rlabel metal3 7672 26824 7672 26824 0 _0690_
rlabel metal2 9912 26096 9912 26096 0 _0691_
rlabel metal2 10136 26208 10136 26208 0 _0692_
rlabel metal2 7784 25424 7784 25424 0 _0693_
rlabel metal2 5656 26544 5656 26544 0 _0694_
rlabel metal2 7896 25144 7896 25144 0 _0695_
rlabel metal2 6776 25760 6776 25760 0 _0696_
rlabel metal2 8904 24808 8904 24808 0 _0697_
rlabel metal3 9800 36344 9800 36344 0 _0698_
rlabel metal2 10584 38136 10584 38136 0 _0699_
rlabel metal3 12880 36680 12880 36680 0 _0700_
rlabel metal2 18760 36624 18760 36624 0 _0701_
rlabel metal2 14056 39060 14056 39060 0 _0702_
rlabel metal2 13944 39060 13944 39060 0 _0703_
rlabel metal2 12824 37688 12824 37688 0 _0704_
rlabel metal2 10696 37520 10696 37520 0 _0705_
rlabel metal2 10360 37632 10360 37632 0 _0706_
rlabel metal2 12040 36568 12040 36568 0 _0707_
rlabel metal3 17304 37016 17304 37016 0 _0708_
rlabel metal2 21112 34048 21112 34048 0 _0709_
rlabel metal2 22120 32312 22120 32312 0 _0710_
rlabel metal2 21336 33824 21336 33824 0 _0711_
rlabel metal2 22792 29064 22792 29064 0 _0712_
rlabel metal2 21896 32368 21896 32368 0 _0713_
rlabel metal2 20776 35280 20776 35280 0 _0714_
rlabel metal2 20216 39536 20216 39536 0 _0715_
rlabel metal2 18480 36456 18480 36456 0 _0716_
rlabel metal3 16856 36344 16856 36344 0 _0717_
rlabel metal2 15064 35952 15064 35952 0 _0718_
rlabel metal2 20216 37632 20216 37632 0 _0719_
rlabel metal2 20384 39592 20384 39592 0 _0720_
rlabel metal2 21896 37464 21896 37464 0 _0721_
rlabel metal2 20776 37296 20776 37296 0 _0722_
rlabel metal2 23464 35672 23464 35672 0 _0723_
rlabel metal2 23240 33824 23240 33824 0 _0724_
rlabel metal2 22680 37240 22680 37240 0 _0725_
rlabel metal2 22232 36008 22232 36008 0 _0726_
rlabel metal2 14728 35840 14728 35840 0 _0727_
rlabel metal2 10024 24472 10024 24472 0 _0728_
rlabel metal2 8008 21840 8008 21840 0 _0729_
rlabel metal2 7224 17752 7224 17752 0 _0730_
rlabel metal2 19992 8372 19992 8372 0 _0731_
rlabel metal2 21168 21560 21168 21560 0 _0732_
rlabel metal2 23016 21952 23016 21952 0 _0733_
rlabel metal2 8680 17584 8680 17584 0 _0734_
rlabel metal2 45192 15596 45192 15596 0 _0735_
rlabel metal3 46648 15288 46648 15288 0 _0736_
rlabel metal2 42168 11872 42168 11872 0 _0737_
rlabel metal2 44184 12824 44184 12824 0 _0738_
rlabel metal2 37240 13608 37240 13608 0 _0739_
rlabel metal2 46312 11424 46312 11424 0 _0740_
rlabel metal2 42504 16072 42504 16072 0 _0741_
rlabel metal2 43960 15512 43960 15512 0 _0742_
rlabel metal2 43960 13160 43960 13160 0 _0743_
rlabel metal2 35336 14672 35336 14672 0 _0744_
rlabel metal3 32312 13720 32312 13720 0 _0745_
rlabel metal2 35560 15204 35560 15204 0 _0746_
rlabel metal2 43176 12824 43176 12824 0 _0747_
rlabel metal2 21896 13384 21896 13384 0 _0748_
rlabel metal2 39704 15344 39704 15344 0 _0749_
rlabel metal3 41272 15848 41272 15848 0 _0750_
rlabel metal2 40488 14000 40488 14000 0 _0751_
rlabel metal2 47096 14280 47096 14280 0 _0752_
rlabel metal2 43064 15064 43064 15064 0 _0753_
rlabel metal2 42168 14056 42168 14056 0 _0754_
rlabel metal3 40824 14336 40824 14336 0 _0755_
rlabel metal2 23016 13552 23016 13552 0 _0756_
rlabel metal2 20104 13384 20104 13384 0 _0757_
rlabel metal2 21280 15848 21280 15848 0 _0758_
rlabel metal2 6608 17080 6608 17080 0 _0759_
rlabel metal2 5768 17248 5768 17248 0 _0760_
rlabel metal2 4816 17528 4816 17528 0 _0761_
rlabel metal2 5656 19880 5656 19880 0 _0762_
rlabel metal3 4928 12152 4928 12152 0 _0763_
rlabel metal2 21840 15960 21840 15960 0 _0764_
rlabel metal2 17304 17360 17304 17360 0 _0765_
rlabel metal2 7448 18704 7448 18704 0 _0766_
rlabel metal2 7504 17080 7504 17080 0 _0767_
rlabel metal2 4984 12992 4984 12992 0 _0768_
rlabel metal3 10472 15512 10472 15512 0 _0769_
rlabel metal3 21616 15624 21616 15624 0 _0770_
rlabel metal2 12712 16688 12712 16688 0 _0771_
rlabel metal2 11368 15344 11368 15344 0 _0772_
rlabel metal3 21560 15400 21560 15400 0 _0773_
rlabel metal2 16856 8008 16856 8008 0 _0774_
rlabel metal2 11816 15680 11816 15680 0 _0775_
rlabel metal2 12264 15792 12264 15792 0 _0776_
rlabel metal2 3752 18928 3752 18928 0 _0777_
rlabel metal2 13664 11256 13664 11256 0 _0778_
rlabel metal2 4648 19432 4648 19432 0 _0779_
rlabel metal2 40208 10808 40208 10808 0 _0780_
rlabel metal2 39928 11928 39928 11928 0 _0781_
rlabel metal3 38360 12152 38360 12152 0 _0782_
rlabel metal2 38808 12208 38808 12208 0 _0783_
rlabel metal2 24248 21728 24248 21728 0 _0784_
rlabel metal3 22624 20776 22624 20776 0 _0785_
rlabel metal2 21448 19376 21448 19376 0 _0786_
rlabel metal3 5376 19880 5376 19880 0 _0787_
rlabel metal2 5152 17080 5152 17080 0 _0788_
rlabel metal3 9352 11256 9352 11256 0 _0789_
rlabel metal2 25256 17360 25256 17360 0 _0790_
rlabel metal2 23240 16912 23240 16912 0 _0791_
rlabel metal2 22232 16016 22232 16016 0 _0792_
rlabel metal2 9576 19208 9576 19208 0 _0793_
rlabel metal3 12264 11144 12264 11144 0 _0794_
rlabel metal2 12824 11424 12824 11424 0 _0795_
rlabel metal2 11312 18536 11312 18536 0 _0796_
rlabel metal2 10808 18312 10808 18312 0 _0797_
rlabel metal2 6104 16856 6104 16856 0 _0798_
rlabel metal2 5096 19320 5096 19320 0 _0799_
rlabel metal2 9016 18200 9016 18200 0 _0800_
rlabel metal2 10024 16128 10024 16128 0 _0801_
rlabel metal2 9352 18536 9352 18536 0 _0802_
rlabel metal3 9072 19992 9072 19992 0 _0803_
rlabel metal2 8344 20104 8344 20104 0 _0804_
rlabel metal2 8792 19544 8792 19544 0 _0805_
rlabel metal2 4928 11368 4928 11368 0 _0806_
rlabel metal2 4312 17192 4312 17192 0 _0807_
rlabel metal2 22568 17360 22568 17360 0 _0808_
rlabel metal3 19936 17528 19936 17528 0 _0809_
rlabel metal2 8960 19208 8960 19208 0 _0810_
rlabel metal2 11368 21224 11368 21224 0 _0811_
rlabel metal3 10416 21448 10416 21448 0 _0812_
rlabel metal2 7952 16744 7952 16744 0 _0813_
rlabel metal3 17080 12152 17080 12152 0 _0814_
rlabel metal3 9856 10472 9856 10472 0 _0815_
rlabel metal2 5320 13272 5320 13272 0 _0816_
rlabel metal2 10416 12152 10416 12152 0 _0817_
rlabel metal3 9128 16184 9128 16184 0 _0818_
rlabel metal3 10136 15960 10136 15960 0 _0819_
rlabel metal2 11256 19712 11256 19712 0 _0820_
rlabel metal2 41720 8904 41720 8904 0 _0821_
rlabel metal2 36456 7168 36456 7168 0 _0822_
rlabel metal2 44184 8792 44184 8792 0 _0823_
rlabel metal2 23128 6608 23128 6608 0 _0824_
rlabel metal2 38304 6664 38304 6664 0 _0825_
rlabel metal2 26152 14056 26152 14056 0 _0826_
rlabel metal2 39816 6160 39816 6160 0 _0827_
rlabel metal2 38472 6440 38472 6440 0 _0828_
rlabel metal2 26600 15204 26600 15204 0 _0829_
rlabel metal2 38920 10696 38920 10696 0 _0830_
rlabel metal2 29624 13944 29624 13944 0 _0831_
rlabel metal2 39312 16856 39312 16856 0 _0832_
rlabel metal2 38808 13552 38808 13552 0 _0833_
rlabel metal2 36456 13384 36456 13384 0 _0834_
rlabel metal2 35168 9576 35168 9576 0 _0835_
rlabel metal2 40488 8288 40488 8288 0 _0836_
rlabel metal2 39256 5880 39256 5880 0 _0837_
rlabel metal2 44688 7448 44688 7448 0 _0838_
rlabel metal2 44744 9072 44744 9072 0 _0839_
rlabel metal2 45248 7672 45248 7672 0 _0840_
rlabel metal2 45080 9016 45080 9016 0 _0841_
rlabel metal2 45080 8512 45080 8512 0 _0842_
rlabel metal3 36232 16072 36232 16072 0 _0843_
rlabel metal2 34664 17248 34664 17248 0 _0844_
rlabel metal2 40936 18704 40936 18704 0 _0845_
rlabel metal3 34216 16856 34216 16856 0 _0846_
rlabel metal2 33488 17080 33488 17080 0 _0847_
rlabel metal2 33208 8512 33208 8512 0 _0848_
rlabel metal2 26040 7840 26040 7840 0 _0849_
rlabel metal2 33320 6384 33320 6384 0 _0850_
rlabel metal3 20608 7560 20608 7560 0 _0851_
rlabel metal2 19432 7728 19432 7728 0 _0852_
rlabel metal2 22232 6384 22232 6384 0 _0853_
rlabel metal2 26264 5768 26264 5768 0 _0854_
rlabel metal3 32592 6776 32592 6776 0 _0855_
rlabel metal2 34216 6664 34216 6664 0 _0856_
rlabel metal2 35560 16744 35560 16744 0 _0857_
rlabel metal2 31584 16184 31584 16184 0 _0858_
rlabel metal2 30072 9072 30072 9072 0 _0859_
rlabel metal2 20888 6552 20888 6552 0 _0860_
rlabel metal3 20216 5880 20216 5880 0 _0861_
rlabel metal2 43288 17024 43288 17024 0 _0862_
rlabel metal3 31528 8232 31528 8232 0 _0863_
rlabel metal2 27496 6664 27496 6664 0 _0864_
rlabel metal2 27720 7056 27720 7056 0 _0865_
rlabel metal3 27216 5880 27216 5880 0 _0866_
rlabel metal2 25816 6048 25816 6048 0 _0867_
rlabel metal2 30856 15064 30856 15064 0 _0868_
rlabel metal2 30184 6496 30184 6496 0 _0869_
rlabel metal2 30408 6720 30408 6720 0 _0870_
rlabel metal2 30072 6048 30072 6048 0 _0871_
rlabel metal2 28952 6048 28952 6048 0 _0872_
rlabel metal2 30296 42672 30296 42672 0 _0873_
rlabel metal2 26936 29120 26936 29120 0 _0874_
rlabel metal2 23016 21112 23016 21112 0 _0875_
rlabel metal2 23744 21000 23744 21000 0 _0876_
rlabel metal3 29512 29512 29512 29512 0 _0877_
rlabel metal3 29848 44072 29848 44072 0 _0878_
rlabel metal2 27384 44800 27384 44800 0 _0879_
rlabel metal2 36344 37128 36344 37128 0 _0880_
rlabel metal2 30408 39256 30408 39256 0 _0881_
rlabel metal2 27720 38360 27720 38360 0 _0882_
rlabel metal2 40376 28616 40376 28616 0 _0883_
rlabel metal2 40040 31304 40040 31304 0 _0884_
rlabel metal3 37576 41160 37576 41160 0 _0885_
rlabel metal2 41328 23128 41328 23128 0 _0886_
rlabel metal2 42280 29792 42280 29792 0 _0887_
rlabel metal2 42952 43232 42952 43232 0 _0888_
rlabel metal2 45024 38136 45024 38136 0 _0889_
rlabel metal3 42840 36456 42840 36456 0 _0890_
rlabel metal2 45080 36400 45080 36400 0 _0891_
rlabel metal3 45304 27944 45304 27944 0 _0892_
rlabel metal2 41048 36344 41048 36344 0 _0893_
rlabel metal2 31640 29792 31640 29792 0 _0894_
rlabel metal2 34384 35672 34384 35672 0 _0895_
rlabel metal2 35448 29680 35448 29680 0 _0896_
rlabel metal2 37800 35896 37800 35896 0 _0897_
rlabel metal2 25592 17136 25592 17136 0 _0898_
rlabel metal2 44856 16128 44856 16128 0 _0899_
rlabel metal2 46424 15736 46424 15736 0 _0900_
rlabel metal3 44016 16856 44016 16856 0 _0901_
rlabel metal2 43736 17360 43736 17360 0 _0902_
rlabel metal2 36680 16968 36680 16968 0 _0903_
rlabel metal2 40040 14224 40040 14224 0 _0904_
rlabel metal2 37800 16800 37800 16800 0 _0905_
rlabel metal2 45080 18928 45080 18928 0 _0906_
rlabel metal2 43512 15680 43512 15680 0 _0907_
rlabel metal2 43400 16352 43400 16352 0 _0908_
rlabel metal2 42280 16576 42280 16576 0 _0909_
rlabel metal2 37912 17808 37912 17808 0 _0910_
rlabel metal2 37128 17920 37128 17920 0 _0911_
rlabel metal2 39144 16296 39144 16296 0 _0912_
rlabel metal2 40600 18536 40600 18536 0 _0913_
rlabel metal2 38136 14896 38136 14896 0 _0914_
rlabel metal2 41272 14224 41272 14224 0 _0915_
rlabel metal2 39256 17584 39256 17584 0 _0916_
rlabel metal2 38696 19152 38696 19152 0 _0917_
rlabel metal2 26600 19656 26600 19656 0 _0918_
rlabel metal3 24976 18312 24976 18312 0 _0919_
rlabel metal3 30184 28504 30184 28504 0 _0920_
rlabel metal2 35224 40992 35224 40992 0 _0921_
rlabel metal2 31640 42280 31640 42280 0 _0922_
rlabel metal2 33656 41104 33656 41104 0 _0923_
rlabel metal2 41160 41160 41160 41160 0 _0924_
rlabel metal2 43848 41384 43848 41384 0 _0925_
rlabel metal2 43736 36512 43736 36512 0 _0926_
rlabel metal2 41496 37520 41496 37520 0 _0927_
rlabel metal2 42280 33768 42280 33768 0 _0928_
rlabel metal2 32424 34440 32424 34440 0 _0929_
rlabel metal2 34832 33544 34832 33544 0 _0930_
rlabel metal3 40152 20104 40152 20104 0 _0931_
rlabel metal3 27048 18256 27048 18256 0 _0932_
rlabel metal2 26376 17304 26376 17304 0 _0933_
rlabel metal2 25928 16408 25928 16408 0 _0934_
rlabel metal2 28952 19264 28952 19264 0 _0935_
rlabel metal2 26936 17136 26936 17136 0 _0936_
rlabel metal2 31192 24696 31192 24696 0 _0937_
rlabel metal2 30296 16464 30296 16464 0 _0938_
rlabel metal2 40264 18256 40264 18256 0 _0939_
rlabel metal3 34328 17528 34328 17528 0 _0940_
rlabel metal2 30072 15904 30072 15904 0 _0941_
rlabel metal2 29736 16128 29736 16128 0 _0942_
rlabel metal2 29232 16184 29232 16184 0 _0943_
rlabel metal2 32088 23352 32088 23352 0 _0944_
rlabel metal3 30352 21560 30352 21560 0 _0945_
rlabel metal2 30520 17192 30520 17192 0 _0946_
rlabel metal2 29848 16800 29848 16800 0 _0947_
rlabel metal2 29512 17976 29512 17976 0 _0948_
rlabel metal2 31864 21448 31864 21448 0 _0949_
rlabel metal2 25480 23352 25480 23352 0 _0950_
rlabel metal2 39928 23464 39928 23464 0 _0951_
rlabel metal2 29960 19264 29960 19264 0 _0952_
rlabel metal2 33544 18368 33544 18368 0 _0953_
rlabel metal2 39984 18424 39984 18424 0 _0954_
rlabel metal3 31752 19208 31752 19208 0 _0955_
rlabel metal3 29960 19320 29960 19320 0 _0956_
rlabel metal3 30184 23352 30184 23352 0 _0957_
rlabel metal2 31696 23240 31696 23240 0 _0958_
rlabel metal2 32312 19656 32312 19656 0 _0959_
rlabel metal2 30800 19208 30800 19208 0 _0960_
rlabel metal2 31304 19264 31304 19264 0 _0961_
rlabel metal4 30968 20720 30968 20720 0 _0962_
rlabel metal2 29288 24360 29288 24360 0 _0963_
rlabel metal2 30632 24528 30632 24528 0 _0964_
rlabel metal2 32200 17416 32200 17416 0 _0965_
rlabel metal2 32536 17752 32536 17752 0 _0966_
rlabel metal2 26040 22848 26040 22848 0 _0967_
rlabel metal2 26040 21784 26040 21784 0 _0968_
rlabel metal3 27272 21560 27272 21560 0 _0969_
rlabel metal2 31528 18760 31528 18760 0 _0970_
rlabel metal2 32200 19656 32200 19656 0 _0971_
rlabel metal2 31976 20440 31976 20440 0 _0972_
rlabel metal2 26264 19208 26264 19208 0 _0973_
rlabel metal2 27048 19488 27048 19488 0 _0974_
rlabel metal2 41608 16240 41608 16240 0 _0975_
rlabel metal3 39704 16968 39704 16968 0 _0976_
rlabel metal2 41384 16408 41384 16408 0 _0977_
rlabel metal3 39200 15512 39200 15512 0 _0978_
rlabel metal2 39144 16800 39144 16800 0 _0979_
rlabel metal2 40376 16184 40376 16184 0 _0980_
rlabel metal2 41160 15904 41160 15904 0 _0981_
rlabel metal4 41496 15232 41496 15232 0 _0982_
rlabel metal2 41048 19600 41048 19600 0 _0983_
rlabel metal2 42056 18032 42056 18032 0 _0984_
rlabel metal2 44968 16016 44968 16016 0 _0985_
rlabel metal2 42168 17808 42168 17808 0 _0986_
rlabel metal2 42112 19208 42112 19208 0 _0987_
rlabel metal2 42448 18312 42448 18312 0 _0988_
rlabel metal3 42224 14504 42224 14504 0 _0989_
rlabel metal2 41608 13160 41608 13160 0 _0990_
rlabel metal2 39816 14168 39816 14168 0 _0991_
rlabel metal2 41720 12936 41720 12936 0 _0992_
rlabel metal2 41496 12992 41496 12992 0 _0993_
rlabel metal2 39144 9352 39144 9352 0 _0994_
rlabel metal3 22736 22232 22736 22232 0 _0995_
rlabel metal2 22680 26572 22680 26572 0 _0996_
rlabel metal2 22456 26544 22456 26544 0 _0997_
rlabel metal2 22120 43792 22120 43792 0 _0998_
rlabel metal2 21672 43792 21672 43792 0 _0999_
rlabel metal2 24584 41888 24584 41888 0 _1000_
rlabel metal2 31640 26992 31640 26992 0 _1001_
rlabel metal2 44072 29232 44072 29232 0 _1002_
rlabel metal2 37912 29400 37912 29400 0 _1003_
rlabel metal2 45080 28672 45080 28672 0 _1004_
rlabel metal2 45080 21056 45080 21056 0 _1005_
rlabel metal2 46648 30968 46648 30968 0 _1006_
rlabel metal2 30856 26936 30856 26936 0 _1007_
rlabel metal2 34776 27720 34776 27720 0 _1008_
rlabel metal3 23016 25928 23016 25928 0 _1009_
rlabel metal2 23464 39984 23464 39984 0 _1010_
rlabel metal3 18200 40600 18200 40600 0 _1011_
rlabel metal2 25368 45528 25368 45528 0 _1012_
rlabel metal2 25592 39536 25592 39536 0 _1013_
rlabel metal2 33992 40208 33992 40208 0 _1014_
rlabel metal2 37800 40768 37800 40768 0 _1015_
rlabel metal3 36736 41384 36736 41384 0 _1016_
rlabel metal3 42112 44520 42112 44520 0 _1017_
rlabel metal2 43064 40432 43064 40432 0 _1018_
rlabel metal2 41160 39480 41160 39480 0 _1019_
rlabel metal2 31976 44464 31976 44464 0 _1020_
rlabel metal3 33768 38808 33768 38808 0 _1021_
rlabel metal2 36232 37968 36232 37968 0 _1022_
rlabel metal2 31360 45304 31360 45304 0 _1023_
rlabel metal2 35448 45304 35448 45304 0 _1024_
rlabel metal2 44632 34384 44632 34384 0 _1025_
rlabel metal2 38136 39200 38136 39200 0 _1026_
rlabel metal2 40264 39704 40264 39704 0 _1027_
rlabel metal3 40768 39816 40768 39816 0 _1028_
rlabel metal2 45080 41272 45080 41272 0 _1029_
rlabel metal2 46536 38808 46536 38808 0 _1030_
rlabel metal2 1736 25256 1736 25256 0 addr[0]
rlabel metal2 13944 46424 13944 46424 0 addr[10]
rlabel metal2 1736 41720 1736 41720 0 addr[11]
rlabel metal2 2912 42504 2912 42504 0 addr[12]
rlabel metal2 1680 34104 1680 34104 0 addr[13]
rlabel metal2 1736 32368 1736 32368 0 addr[14]
rlabel metal2 1736 40488 1736 40488 0 addr[15]
rlabel metal3 2968 39648 2968 39648 0 addr[16]
rlabel metal2 4760 39368 4760 39368 0 addr[17]
rlabel metal2 2464 40600 2464 40600 0 addr[18]
rlabel metal3 1582 24920 1582 24920 0 addr[19]
rlabel metal2 1736 23464 1736 23464 0 addr[1]
rlabel metal2 1736 28840 1736 28840 0 addr[20]
rlabel metal2 2744 34272 2744 34272 0 addr[21]
rlabel metal2 1904 32536 1904 32536 0 addr[22]
rlabel metal2 1736 33152 1736 33152 0 addr[23]
rlabel metal2 3136 26600 3136 26600 0 addr[2]
rlabel metal3 2408 25816 2408 25816 0 addr[3]
rlabel metal2 2184 22344 2184 22344 0 addr[4]
rlabel metal3 23688 45080 23688 45080 0 addr[5]
rlabel metal2 18312 45864 18312 45864 0 addr[6]
rlabel metal2 20160 45864 20160 45864 0 addr[7]
rlabel metal3 1246 37688 1246 37688 0 addr[8]
rlabel metal2 15288 45976 15288 45976 0 addr[9]
rlabel metal2 28728 43176 28728 43176 0 buffer\[0\]
rlabel metal2 39256 41104 39256 41104 0 buffer\[10\]
rlabel metal2 43288 43680 43288 43680 0 buffer\[11\]
rlabel metal2 43904 36680 43904 36680 0 buffer\[12\]
rlabel metal2 42112 38136 42112 38136 0 buffer\[13\]
rlabel metal2 35448 36624 35448 36624 0 buffer\[14\]
rlabel metal2 38248 36792 38248 36792 0 buffer\[15\]
rlabel metal2 32424 44436 32424 44436 0 buffer\[16\]
rlabel metal2 34664 41608 34664 41608 0 buffer\[17\]
rlabel metal2 41832 40880 41832 40880 0 buffer\[18\]
rlabel metal2 37800 39816 37800 39816 0 buffer\[19\]
rlabel metal2 25704 41160 25704 41160 0 buffer\[1\]
rlabel metal2 48216 38080 48216 38080 0 buffer\[20\]
rlabel metal2 48216 32872 48216 32872 0 buffer\[21\]
rlabel metal2 32480 35000 32480 35000 0 buffer\[22\]
rlabel via2 33992 33320 33992 33320 0 buffer\[23\]
rlabel metal3 38416 30856 38416 30856 0 buffer\[2\]
rlabel metal2 43848 29064 43848 29064 0 buffer\[3\]
rlabel metal2 46872 23184 46872 23184 0 buffer\[4\]
rlabel metal2 47320 29288 47320 29288 0 buffer\[5\]
rlabel metal2 31080 27944 31080 27944 0 buffer\[6\]
rlabel metal2 34888 29568 34888 29568 0 buffer\[7\]
rlabel metal2 26936 44744 26936 44744 0 buffer\[8\]
rlabel metal2 29064 38976 29064 38976 0 buffer\[9\]
rlabel metal3 35672 3528 35672 3528 0 cfgreg_di[0]
rlabel metal2 43736 1862 43736 1862 0 cfgreg_di[10]
rlabel metal2 45080 2058 45080 2058 0 cfgreg_di[11]
rlabel metal2 9576 3696 9576 3696 0 cfgreg_di[16]
rlabel metal2 12824 5880 12824 5880 0 cfgreg_di[17]
rlabel metal2 12152 2058 12152 2058 0 cfgreg_di[18]
rlabel metal3 12824 3528 12824 3528 0 cfgreg_di[19]
rlabel metal2 22232 2058 22232 2058 0 cfgreg_di[1]
rlabel metal3 6160 4088 6160 4088 0 cfgreg_di[20]
rlabel metal3 6048 3528 6048 3528 0 cfgreg_di[21]
rlabel metal2 16856 2058 16856 2058 0 cfgreg_di[22]
rlabel metal2 24920 1918 24920 1918 0 cfgreg_di[2]
rlabel metal2 23576 2058 23576 2058 0 cfgreg_di[31]
rlabel metal3 32480 3528 32480 3528 0 cfgreg_di[3]
rlabel metal2 35672 854 35672 854 0 cfgreg_di[4]
rlabel metal2 31640 1246 31640 1246 0 cfgreg_di[5]
rlabel metal2 43064 1974 43064 1974 0 cfgreg_di[8]
rlabel metal2 42392 2058 42392 2058 0 cfgreg_di[9]
rlabel metal2 47992 25816 47992 25816 0 cfgreg_do[0]
rlabel metal2 47992 7392 47992 7392 0 cfgreg_do[10]
rlabel metal3 48258 9464 48258 9464 0 cfgreg_do[11]
rlabel metal2 11480 2058 11480 2058 0 cfgreg_do[16]
rlabel metal2 14840 1806 14840 1806 0 cfgreg_do[17]
rlabel metal2 13496 1974 13496 1974 0 cfgreg_do[18]
rlabel metal2 16184 2198 16184 2198 0 cfgreg_do[19]
rlabel metal2 47992 23800 47992 23800 0 cfgreg_do[1]
rlabel metal3 1358 17528 1358 17528 0 cfgreg_do[20]
rlabel metal3 10080 4088 10080 4088 0 cfgreg_do[21]
rlabel metal3 18088 3640 18088 3640 0 cfgreg_do[22]
rlabel metal2 47992 21616 47992 21616 0 cfgreg_do[2]
rlabel metal2 26936 2086 26936 2086 0 cfgreg_do[31]
rlabel metal2 47992 19768 47992 19768 0 cfgreg_do[3]
rlabel metal2 37016 2198 37016 2198 0 cfgreg_do[4]
rlabel metal2 38360 2478 38360 2478 0 cfgreg_do[5]
rlabel metal3 42952 5656 42952 5656 0 cfgreg_do[8]
rlabel metal3 43792 4872 43792 4872 0 cfgreg_do[9]
rlabel metal3 31080 5992 31080 5992 0 cfgreg_we[0]
rlabel metal2 44576 4088 44576 4088 0 cfgreg_we[1]
rlabel metal2 8456 3584 8456 3584 0 cfgreg_we[2]
rlabel metal2 22904 854 22904 854 0 cfgreg_we[3]
rlabel metal2 24976 24696 24976 24696 0 clk
rlabel metal3 30464 36456 30464 36456 0 clknet_0_clk
rlabel metal2 17528 9296 17528 9296 0 clknet_4_0_0_clk
rlabel metal2 43624 10696 43624 10696 0 clknet_4_10_0_clk
rlabel metal3 42000 26264 42000 26264 0 clknet_4_11_0_clk
rlabel metal2 28560 29400 28560 29400 0 clknet_4_12_0_clk
rlabel metal3 30184 44296 30184 44296 0 clknet_4_13_0_clk
rlabel metal2 45640 30576 45640 30576 0 clknet_4_14_0_clk
rlabel metal2 45080 34552 45080 34552 0 clknet_4_15_0_clk
rlabel metal2 3304 7840 3304 7840 0 clknet_4_1_0_clk
rlabel metal2 24808 6216 24808 6216 0 clknet_4_2_0_clk
rlabel metal2 18592 16856 18592 16856 0 clknet_4_3_0_clk
rlabel metal2 1848 22680 1848 22680 0 clknet_4_4_0_clk
rlabel metal2 17192 45360 17192 45360 0 clknet_4_5_0_clk
rlabel metal2 17528 20384 17528 20384 0 clknet_4_6_0_clk
rlabel metal2 18648 42672 18648 42672 0 clknet_4_7_0_clk
rlabel metal2 34104 16716 34104 16716 0 clknet_4_8_0_clk
rlabel metal2 35224 21392 35224 21392 0 clknet_4_9_0_clk
rlabel metal2 36456 4536 36456 4536 0 config_clk
rlabel metal2 38696 5712 38696 5712 0 config_csb
rlabel metal2 34664 5208 34664 5208 0 config_do\[0\]
rlabel metal2 21616 4200 21616 4200 0 config_do\[1\]
rlabel metal2 26376 5544 26376 5544 0 config_do\[2\]
rlabel metal2 29736 5432 29736 5432 0 config_do\[3\]
rlabel metal2 42280 5544 42280 5544 0 config_oe\[0\]
rlabel metal2 44240 7336 44240 7336 0 config_oe\[1\]
rlabel metal3 46256 8008 46256 8008 0 config_oe\[2\]
rlabel metal2 46984 7840 46984 7840 0 config_oe\[3\]
rlabel metal2 20776 11424 20776 11424 0 din_ddr
rlabel metal2 45192 24416 45192 24416 0 flash_in[2]
rlabel metal2 42392 23352 42392 23352 0 flash_in[3]
rlabel metal2 48272 18424 48272 18424 0 flash_in[4]
rlabel metal2 47544 19656 47544 19656 0 flash_in[5]
rlabel metal3 40992 5096 40992 5096 0 flash_oeb[2]
rlabel metal2 39704 1806 39704 1806 0 flash_oeb[3]
rlabel metal2 47992 8232 47992 8232 0 flash_oeb[4]
rlabel metal3 48650 8792 48650 8792 0 flash_oeb[5]
rlabel metal3 41832 3416 41832 3416 0 flash_out[0]
rlabel metal2 37688 2198 37688 2198 0 flash_out[1]
rlabel metal3 33432 3640 33432 3640 0 flash_out[2]
rlabel metal3 21504 3640 21504 3640 0 flash_out[3]
rlabel metal2 26264 2198 26264 2198 0 flash_out[4]
rlabel metal3 30296 3752 30296 3752 0 flash_out[5]
rlabel metal2 2072 24472 2072 24472 0 net1
rlabel metal2 18312 36848 18312 36848 0 net10
rlabel metal2 42168 31892 42168 31892 0 net100
rlabel metal2 43848 31304 43848 31304 0 net101
rlabel metal2 45864 36232 45864 36232 0 net102
rlabel metal2 40040 30296 40040 30296 0 net103
rlabel metal2 31080 31444 31080 31444 0 net104
rlabel metal2 35336 31752 35336 31752 0 net105
rlabel metal2 45528 28672 45528 28672 0 net106
rlabel metal2 48160 22456 48160 22456 0 net107
rlabel metal2 47992 30688 47992 30688 0 net108
rlabel metal2 45640 27944 45640 27944 0 net109
rlabel metal2 2968 24920 2968 24920 0 net11
rlabel metal3 45640 28784 45640 28784 0 net110
rlabel metal2 23912 45528 23912 45528 0 net111
rlabel metal2 26264 40992 26264 40992 0 net112
rlabel metal2 18312 29848 18312 29848 0 net113
rlabel metal2 48216 42280 48216 42280 0 net114
rlabel metal3 1246 45080 1246 45080 0 net115
rlabel metal3 1246 5432 1246 5432 0 net116
rlabel metal3 1470 2744 1470 2744 0 net117
rlabel metal2 47768 45024 47768 45024 0 net118
rlabel metal3 1246 4088 1246 4088 0 net119
rlabel metal2 2072 23072 2072 23072 0 net12
rlabel metal2 44240 11144 44240 11144 0 net120
rlabel metal2 48272 45640 48272 45640 0 net121
rlabel metal2 46872 45360 46872 45360 0 net122
rlabel metal2 48216 10640 48216 10640 0 net123
rlabel metal2 42504 8792 42504 8792 0 net124
rlabel metal2 45248 43736 45248 43736 0 net125
rlabel metal2 48216 44128 48216 44128 0 net126
rlabel metal2 1736 3360 1736 3360 0 net127
rlabel metal2 45304 43064 45304 43064 0 net128
rlabel metal3 1246 4760 1246 4760 0 net129
rlabel metal2 2296 28896 2296 28896 0 net13
rlabel metal3 37576 10696 37576 10696 0 net130
rlabel metal2 21224 10080 21224 10080 0 net131
rlabel metal3 2968 34552 2968 34552 0 net14
rlabel metal2 11816 23240 11816 23240 0 net15
rlabel metal2 1960 29736 1960 29736 0 net16
rlabel metal2 3416 28672 3416 28672 0 net17
rlabel metal2 2296 27608 2296 27608 0 net18
rlabel metal2 16744 25872 16744 25872 0 net19
rlabel metal2 13440 39592 13440 39592 0 net2
rlabel metal2 24136 38192 24136 38192 0 net20
rlabel metal2 19264 34104 19264 34104 0 net21
rlabel metal2 17696 26376 17696 26376 0 net22
rlabel metal2 17864 39480 17864 39480 0 net23
rlabel metal2 15064 41720 15064 41720 0 net24
rlabel metal2 36008 3696 36008 3696 0 net25
rlabel metal3 47152 4536 47152 4536 0 net26
rlabel metal2 48216 4816 48216 4816 0 net27
rlabel metal2 9352 3584 9352 3584 0 net28
rlabel metal2 8456 4760 8456 4760 0 net29
rlabel metal2 2296 41608 2296 41608 0 net3
rlabel metal2 12320 6104 12320 6104 0 net30
rlabel metal2 13272 3416 13272 3416 0 net31
rlabel metal2 21448 5600 21448 5600 0 net32
rlabel metal3 6552 3416 6552 3416 0 net33
rlabel metal2 7672 3640 7672 3640 0 net34
rlabel metal2 17304 3752 17304 3752 0 net35
rlabel metal2 24920 4312 24920 4312 0 net36
rlabel metal2 24136 5488 24136 5488 0 net37
rlabel metal2 32536 3640 32536 3640 0 net38
rlabel metal2 37352 5040 37352 5040 0 net39
rlabel metal2 2072 37184 2072 37184 0 net4
rlabel metal2 34664 4760 34664 4760 0 net40
rlabel metal2 47432 4200 47432 4200 0 net41
rlabel metal2 46536 4256 46536 4256 0 net42
rlabel metal2 31136 5096 31136 5096 0 net43
rlabel metal2 42728 4256 42728 4256 0 net44
rlabel metal3 9408 5880 9408 5880 0 net45
rlabel metal2 22960 6440 22960 6440 0 net46
rlabel metal2 44968 23912 44968 23912 0 net47
rlabel metal2 42056 23184 42056 23184 0 net48
rlabel metal2 40040 21224 40040 21224 0 net49
rlabel metal2 2296 33432 2296 33432 0 net5
rlabel metal2 43512 19320 43512 19320 0 net50
rlabel metal2 19320 8064 19320 8064 0 net51
rlabel metal2 15288 34944 15288 34944 0 net52
rlabel metal2 45640 26096 45640 26096 0 net53
rlabel metal2 45752 9688 45752 9688 0 net54
rlabel metal2 47880 10080 47880 10080 0 net55
rlabel metal3 12040 13720 12040 13720 0 net56
rlabel metal3 16128 18648 16128 18648 0 net57
rlabel metal2 12656 14280 12656 14280 0 net58
rlabel metal3 17696 20552 17696 20552 0 net59
rlabel metal2 2184 32592 2184 32592 0 net6
rlabel metal2 36008 23856 36008 23856 0 net60
rlabel metal2 3864 17248 3864 17248 0 net61
rlabel metal2 9800 6776 9800 6776 0 net62
rlabel metal2 19096 5264 19096 5264 0 net63
rlabel metal2 45640 21448 45640 21448 0 net64
rlabel metal2 25704 5880 25704 5880 0 net65
rlabel metal3 44688 20104 44688 20104 0 net66
rlabel metal2 38808 6496 38808 6496 0 net67
rlabel metal2 39928 7224 39928 7224 0 net68
rlabel metal3 42056 6440 42056 6440 0 net69
rlabel metal2 2296 39760 2296 39760 0 net7
rlabel metal3 43064 7224 43064 7224 0 net70
rlabel metal3 40376 6552 40376 6552 0 net71
rlabel metal2 40936 7784 40936 7784 0 net72
rlabel metal2 47208 10472 47208 10472 0 net73
rlabel metal3 46928 9016 46928 9016 0 net74
rlabel metal2 39032 7560 39032 7560 0 net75
rlabel metal2 39704 8176 39704 8176 0 net76
rlabel metal2 33320 4368 33320 4368 0 net77
rlabel metal2 20104 5712 20104 5712 0 net78
rlabel metal2 25928 4592 25928 4592 0 net79
rlabel metal3 5824 39480 5824 39480 0 net8
rlabel metal2 29064 5544 29064 5544 0 net80
rlabel metal2 22680 44576 22680 44576 0 net81
rlabel metal2 37576 41664 37576 41664 0 net82
rlabel metal2 42056 43344 42056 43344 0 net83
rlabel via1 45416 38682 45416 38682 0 net84
rlabel metal2 42056 39872 42056 39872 0 net85
rlabel metal2 34888 39928 34888 39928 0 net86
rlabel metal2 37576 38472 37576 38472 0 net87
rlabel metal2 31640 44632 31640 44632 0 net88
rlabel metal2 36792 44240 36792 44240 0 net89
rlabel metal2 3304 34160 3304 34160 0 net9
rlabel metal2 45864 41160 45864 41160 0 net90
rlabel metal2 38360 40712 38360 40712 0 net91
rlabel metal2 28616 45304 28616 45304 0 net92
rlabel metal2 48272 42728 48272 42728 0 net93
rlabel metal2 47880 35616 47880 35616 0 net94
rlabel metal2 30856 35616 30856 35616 0 net95
rlabel metal2 31528 32984 31528 32984 0 net96
rlabel metal2 31304 40768 31304 40768 0 net97
rlabel metal2 31416 37912 31416 37912 0 net98
rlabel metal2 45640 36176 45640 36176 0 net99
rlabel metal3 20328 25368 20328 25368 0 rd_addr\[0\]
rlabel metal2 15288 42784 15288 42784 0 rd_addr\[10\]
rlabel metal3 10976 42728 10976 42728 0 rd_addr\[11\]
rlabel metal2 11704 44072 11704 44072 0 rd_addr\[12\]
rlabel metal2 8568 42504 8568 42504 0 rd_addr\[13\]
rlabel metal2 5096 41160 5096 41160 0 rd_addr\[14\]
rlabel metal2 5096 40544 5096 40544 0 rd_addr\[15\]
rlabel metal2 11928 40824 11928 40824 0 rd_addr\[16\]
rlabel metal3 6440 40600 6440 40600 0 rd_addr\[17\]
rlabel metal2 8232 23688 8232 23688 0 rd_addr\[18\]
rlabel metal3 15848 26992 15848 26992 0 rd_addr\[19\]
rlabel metal2 20664 23408 20664 23408 0 rd_addr\[1\]
rlabel metal2 7000 25928 7000 25928 0 rd_addr\[20\]
rlabel metal2 16408 44240 16408 44240 0 rd_addr\[21\]
rlabel metal3 5152 28616 5152 28616 0 rd_addr\[22\]
rlabel metal2 9016 42168 9016 42168 0 rd_addr\[23\]
rlabel metal2 28168 30688 28168 30688 0 rd_addr\[2\]
rlabel metal2 26600 32200 26600 32200 0 rd_addr\[3\]
rlabel metal2 28168 34384 28168 34384 0 rd_addr\[4\]
rlabel metal2 26936 36288 26936 36288 0 rd_addr\[5\]
rlabel metal2 19992 42784 19992 42784 0 rd_addr\[6\]
rlabel metal2 21000 41888 21000 41888 0 rd_addr\[7\]
rlabel metal2 18648 43680 18648 43680 0 rd_addr\[8\]
rlabel metal3 19096 42056 19096 42056 0 rd_addr\[9\]
rlabel metal3 10864 23016 10864 23016 0 rd_inc
rlabel metal2 15176 22400 15176 22400 0 rd_valid
rlabel metal3 5992 22456 5992 22456 0 rd_wait
rlabel metal2 23576 47810 23576 47810 0 rdata[0]
rlabel metal2 38360 47194 38360 47194 0 rdata[10]
rlabel metal2 40152 44520 40152 44520 0 rdata[11]
rlabel metal2 47880 40488 47880 40488 0 rdata[12]
rlabel metal2 47992 39592 47992 39592 0 rdata[13]
rlabel metal2 35000 47698 35000 47698 0 rdata[14]
rlabel metal2 37688 47250 37688 47250 0 rdata[15]
rlabel metal2 33824 44632 33824 44632 0 rdata[16]
rlabel metal2 36400 46536 36400 46536 0 rdata[17]
rlabel metal2 47992 42504 47992 42504 0 rdata[18]
rlabel metal2 44408 47306 44408 47306 0 rdata[19]
rlabel metal2 26264 47698 26264 47698 0 rdata[1]
rlabel metal3 48146 40376 48146 40376 0 rdata[20]
rlabel metal3 46200 35056 46200 35056 0 rdata[21]
rlabel metal2 30296 47698 30296 47698 0 rdata[22]
rlabel metal2 31752 44800 31752 44800 0 rdata[23]
rlabel metal2 32984 48146 32984 48146 0 rdata[24]
rlabel metal3 33208 43400 33208 43400 0 rdata[25]
rlabel metal2 47432 35000 47432 35000 0 rdata[26]
rlabel metal3 49336 32872 49336 32872 0 rdata[27]
rlabel metal3 48174 31640 48174 31640 0 rdata[28]
rlabel metal2 47992 35672 47992 35672 0 rdata[29]
rlabel metal3 48202 29624 48202 29624 0 rdata[2]
rlabel metal2 30968 46466 30968 46466 0 rdata[30]
rlabel metal3 47306 30968 47306 30968 0 rdata[31]
rlabel metal2 47768 30408 47768 30408 0 rdata[3]
rlabel metal2 46984 23744 46984 23744 0 rdata[4]
rlabel metal3 47810 30296 47810 30296 0 rdata[5]
rlabel metal2 47880 28392 47880 28392 0 rdata[6]
rlabel metal2 47992 28728 47992 28728 0 rdata[7]
rlabel metal2 25592 47306 25592 47306 0 rdata[8]
rlabel metal2 26936 47642 26936 47642 0 rdata[9]
rlabel metal3 1638 29624 1638 29624 0 ready
rlabel metal3 19768 5040 19768 5040 0 resetn
rlabel metal2 19880 6888 19880 6888 0 softreset
rlabel metal2 5992 15148 5992 15148 0 state\[0\]
rlabel metal2 1736 20496 1736 20496 0 state\[10\]
rlabel metal2 5656 12152 5656 12152 0 state\[11\]
rlabel metal2 10696 13944 10696 13944 0 state\[12\]
rlabel metal2 15400 15960 15400 15960 0 state\[1\]
rlabel metal2 10360 21448 10360 21448 0 state\[2\]
rlabel metal3 10080 11368 10080 11368 0 state\[3\]
rlabel metal2 9576 18088 9576 18088 0 state\[4\]
rlabel metal2 5432 13104 5432 13104 0 state\[5\]
rlabel metal2 11256 19096 11256 19096 0 state\[6\]
rlabel metal2 1736 16464 1736 16464 0 state\[7\]
rlabel metal2 4648 12936 4648 12936 0 state\[8\]
rlabel metal2 11256 12600 11256 12600 0 state\[9\]
rlabel metal2 2408 25760 2408 25760 0 valid
rlabel metal2 48160 19880 48160 19880 0 xfer.count\[0\]
rlabel metal2 45976 16912 45976 16912 0 xfer.count\[1\]
rlabel metal2 47880 15484 47880 15484 0 xfer.count\[2\]
rlabel metal2 48216 13104 48216 13104 0 xfer.count\[3\]
rlabel metal3 24752 18648 24752 18648 0 xfer.din_data\[0\]
rlabel metal2 21672 16352 21672 16352 0 xfer.din_data\[1\]
rlabel metal2 19432 15260 19432 15260 0 xfer.din_data\[2\]
rlabel metal2 21560 19208 21560 19208 0 xfer.din_data\[3\]
rlabel metal2 25592 23632 25592 23632 0 xfer.din_data\[4\]
rlabel metal3 28672 26376 28672 26376 0 xfer.din_data\[5\]
rlabel metal3 25032 23128 25032 23128 0 xfer.din_data\[6\]
rlabel metal2 26152 24024 26152 24024 0 xfer.din_data\[7\]
rlabel metal2 17752 12992 17752 12992 0 xfer.din_qspi
rlabel metal2 16856 17304 16856 17304 0 xfer.din_rd
rlabel metal2 4816 8344 4816 8344 0 xfer.din_tag\[0\]
rlabel metal2 6216 7392 6216 7392 0 xfer.din_tag\[1\]
rlabel metal2 9016 8792 9016 8792 0 xfer.din_tag\[2\]
rlabel metal2 19712 9912 19712 9912 0 xfer.din_valid
rlabel metal2 35896 31920 35896 31920 0 xfer.dout_data\[0\]
rlabel metal2 37128 20664 37128 20664 0 xfer.dout_data\[1\]
rlabel metal2 41328 20888 41328 20888 0 xfer.dout_data\[2\]
rlabel metal2 42840 22064 42840 22064 0 xfer.dout_data\[3\]
rlabel metal2 42728 24752 42728 24752 0 xfer.dout_data\[4\]
rlabel metal2 43288 25872 43288 25872 0 xfer.dout_data\[5\]
rlabel metal2 37688 27272 37688 27272 0 xfer.dout_data\[6\]
rlabel metal3 40040 27720 40040 27720 0 xfer.dout_data\[7\]
rlabel metal2 23128 22512 23128 22512 0 xfer.dout_tag\[0\]
rlabel metal2 23464 22120 23464 22120 0 xfer.dout_tag\[1\]
rlabel metal2 23016 15624 23016 15624 0 xfer.dout_tag\[2\]
rlabel metal2 26264 12208 26264 12208 0 xfer.dummy_count\[0\]
rlabel metal2 26152 12432 26152 12432 0 xfer.dummy_count\[1\]
rlabel metal2 23576 14448 23576 14448 0 xfer.dummy_count\[2\]
rlabel metal2 25368 10976 25368 10976 0 xfer.dummy_count\[3\]
rlabel metal2 40264 11368 40264 11368 0 xfer.fetch
rlabel metal2 46872 11424 46872 11424 0 xfer.flash_clk
rlabel metal2 43848 9520 43848 9520 0 xfer.flash_csb
rlabel metal2 33432 7000 33432 7000 0 xfer.flash_io0_do
rlabel metal2 21672 8568 21672 8568 0 xfer.flash_io1_do
rlabel metal2 25480 7112 25480 7112 0 xfer.flash_io2_do
rlabel metal2 29848 7784 29848 7784 0 xfer.flash_io3_do
rlabel metal2 40936 9912 40936 9912 0 xfer.last_fetch
rlabel metal2 25928 18928 25928 18928 0 xfer.obuffer\[0\]
rlabel metal2 30016 18536 30016 18536 0 xfer.obuffer\[1\]
rlabel metal2 30744 22064 30744 22064 0 xfer.obuffer\[2\]
rlabel metal2 32424 20440 32424 20440 0 xfer.obuffer\[3\]
rlabel metal2 32872 17192 32872 17192 0 xfer.obuffer\[4\]
rlabel metal2 30408 24696 30408 24696 0 xfer.obuffer\[5\]
rlabel metal2 27944 22120 27944 22120 0 xfer.obuffer\[6\]
rlabel metal2 28784 20104 28784 20104 0 xfer.obuffer\[7\]
rlabel metal2 20216 12320 20216 12320 0 xfer.resetn
rlabel metal3 38836 11256 38836 11256 0 xfer.xfer_ddr
rlabel metal2 39256 10920 39256 10920 0 xfer.xfer_ddr_q
rlabel metal3 34160 13720 34160 13720 0 xfer.xfer_dspi
rlabel metal2 40040 12600 40040 12600 0 xfer.xfer_qspi
rlabel metal2 33656 9968 33656 9968 0 xfer.xfer_rd
rlabel metal2 16520 10248 16520 10248 0 xfer.xfer_tag\[0\]
rlabel metal2 20272 18648 20272 18648 0 xfer.xfer_tag\[1\]
rlabel metal3 26292 9912 26292 9912 0 xfer.xfer_tag\[2\]
rlabel metal2 32312 6776 32312 6776 0 xfer_io0_90
rlabel metal2 22008 7616 22008 7616 0 xfer_io1_90
rlabel metal2 27832 7448 27832 7448 0 xfer_io2_90
rlabel metal2 31080 7112 31080 7112 0 xfer_io3_90
<< properties >>
string FIXED_BBOX 0 0 50000 50000
<< end >>
